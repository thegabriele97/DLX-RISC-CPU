library ieee;
use ieee.std_logic_1164.all;
use work.myTypes.all;
 
package record_CU is

	-- Control word bits
	type control_word_t is record
		fetch_en            : std_logic; -- F
		fetch_stall         : std_logic; -- S
		pc_en               : std_logic; -- P
		jump_en             : std_logic; -- J
		call                : std_logic; -- L
		ret                 : std_logic; -- E
		rf_rd1_en           : std_logic; -- 1
		rf_rd2_en           : std_logic; -- 2
		sel_cmpb            : std_logic; -- P
		unsigned_id         : std_logic; -- U
		npc_sel             : std_logic; -- N
		hazard_table_wr1    : std_logic; -- H
		id_en               : std_logic; -- D
		ex_en               : std_logic; -- X
		muxa_sel            : std_logic; -- A
		muxb_sel            : std_logic; -- B
		alu_opcode          : alu_op_sig_t; -- -----
		set_cmp             : set_op_sig_t; -- +++
		sel_alu             : std_logic; -- T
		dram_we             : std_logic; -- W
		dram_re             : std_logic; -- R
		data_size           : std_logic_vector(1 downto 0); -- 10
		mem_en              : std_logic; -- M
		wb_mux_sel          : std_logic; -- C
		wb_en               : std_logic; -- K
	end record control_word_t;

	constant RECORD_RTYPE: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        => ALU_ADD,
		set_cmp           => SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_VOID: control_word_t := (
		fetch_en          => '0', 
		fetch_stall       => '0',
		pc_en             => '0',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '0',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        => ALU_ADD,
		set_cmp           => SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_J: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '1',
		pc_en             => '1',
		jump_en           => '1',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '0',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_JAL: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '1',
		pc_en             => '1',
		jump_en           => '1',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_BEQZ: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_BNEZ: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_ADDI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_ADDUI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SUBI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_SUB,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SUBUI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_SUB,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_ANDI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_AND,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_ORI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_OR,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_XORI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_XOR,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_LHI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '0',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '1',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_SLL,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_JR: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '1',
		pc_en             => '1',
		jump_en           => '1',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '1',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_JALR: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '1',
		pc_en             => '1',
		jump_en           => '1',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '1',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '1',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SLLI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_SLL,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_NOP: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '0',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_SRLI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_SRL,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SRAI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_SRA,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SEQI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SNEI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SNE,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SLTI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SLT,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SGTI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SGT,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SLEI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SLE,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SGEI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SGE,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_CALL: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '1',
		pc_en             => '1',
		jump_en           => '1',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_RET: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '1',
		pc_en             => '1',
		jump_en           => '1',
		call              => '0',
		ret               => '1',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '1',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_LB: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '1',
		data_size         => "10",
		mem_en            => '1',
		wb_mux_sel        => '1',
		wb_en             => '1'
	);

	constant RECORD_LH: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '1',
		data_size         => "01",
		mem_en            => '1',
		wb_mux_sel        => '1',
		wb_en             => '1'
	);

	constant RECORD_LW: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '1',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '1',
		wb_en             => '1'
	);

	constant RECORD_LBU: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '1',
		data_size         => "10",
		mem_en            => '1',
		wb_mux_sel        => '1',
		wb_en             => '1'
	);

	constant RECORD_LHU: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '1',
		data_size         => "01",
		mem_en            => '1',
		wb_mux_sel        => '1',
		wb_en             => '1'
	);

	constant RECORD_SB: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '1',
		dram_re           => '0',
		data_size         => "10",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_SH: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '1',
		dram_re           => '0',
		data_size         => "01",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_SW: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '0',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '1',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_BGT: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_BGE: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_BLT: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_BLE: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '1',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '0',
		id_en             => '0',
		ex_en             => '0',
		muxa_sel          => '0',
		muxb_sel          => '0',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '0',
		wb_mux_sel        => '0',
		wb_en             => '0'
	);

	constant RECORD_TICKTMR: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '1',
		unsigned_id       => '0',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SEQ,
		sel_alu           => '0',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SLTUI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SLT,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SGTUI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SGT,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SLEUI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SLE,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

	constant RECORD_SGEUI: control_word_t := (
		fetch_en          => '1', 
		fetch_stall       => '0',
		pc_en             => '1',
		jump_en           => '0',
		call              => '0',
		ret               => '0',
		rf_rd1_en         => '1',
		rf_rd2_en         => '0',
		sel_cmpb          => '0',
		unsigned_id       => '1',
		npc_sel           => '0',
		hazard_table_wr1  => '1',
		id_en             => '1',
		ex_en             => '1',
		muxa_sel          => '0',
		muxb_sel          => '1',
		alu_opcode        =>  ALU_ADD,
		set_cmp           =>  SET_SGE,
		sel_alu           => '1',
		dram_we           => '0',
		dram_re           => '0',
		data_size         => "00",
		mem_en            => '1',
		wb_mux_sel        => '0',
		wb_en             => '1'
	);

end package record_CU;