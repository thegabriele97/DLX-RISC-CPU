
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32.all;

entity mux_N32_M5_0 is

   port( S : in std_logic_vector (4 downto 0);  Q : in std_logic_vector (1023 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end mux_N32_M5_0;

architecture SYN_behav of mux_N32_M5_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705 : std_logic;

begin
   
   U2 : AOI22_X1 port map( A1 => n255, A2 => Q(502), B1 => n254, B2 => Q(566), 
                           ZN => n1);
   U3 : AOI22_X1 port map( A1 => n257, A2 => Q(662), B1 => n256, B2 => Q(470), 
                           ZN => n2);
   U4 : AOI22_X1 port map( A1 => n259, A2 => Q(374), B1 => n258, B2 => Q(310), 
                           ZN => n3);
   U5 : AOI22_X1 port map( A1 => n261, A2 => Q(406), B1 => n260, B2 => Q(278), 
                           ZN => n4);
   U6 : NAND4_X1 port map( A1 => n1, A2 => n2, A3 => n3, A4 => n4, ZN => n5);
   U7 : AOI22_X1 port map( A1 => n263, A2 => Q(342), B1 => n262, B2 => Q(438), 
                           ZN => n6);
   U8 : AOI22_X1 port map( A1 => n265, A2 => Q(246), B1 => n264, B2 => Q(150), 
                           ZN => n7);
   U9 : AOI22_X1 port map( A1 => n267, A2 => Q(86), B1 => n266, B2 => Q(182), 
                           ZN => n8);
   U10 : AOI22_X1 port map( A1 => n269, A2 => Q(214), B1 => n268, B2 => Q(54), 
                           ZN => n9);
   U11 : NAND4_X1 port map( A1 => n6, A2 => n7, A3 => n8, A4 => n9, ZN => n10);
   U12 : AOI22_X1 port map( A1 => n240, A2 => Q(1014), B1 => n239, B2 => Q(950)
                           , ZN => n11);
   U13 : AOI22_X1 port map( A1 => n242, A2 => Q(982), B1 => n241, B2 => Q(918),
                           ZN => n12);
   U14 : AOI222_X1 port map( A1 => n244, A2 => Q(822), B1 => n245, B2 => Q(118)
                           , C1 => n243, C2 => Q(758), ZN => n13);
   U15 : NAND3_X1 port map( A1 => n11, A2 => n12, A3 => n13, ZN => n14);
   U16 : AOI22_X1 port map( A1 => n247, A2 => Q(854), B1 => n246, B2 => Q(726),
                           ZN => n15);
   U17 : AOI22_X1 port map( A1 => n249, A2 => Q(790), B1 => n248, B2 => Q(886),
                           ZN => n16);
   U18 : NAND4_X1 port map( A1 => n495, A2 => n496, A3 => n15, A4 => n16, ZN =>
                           n17);
   U19 : OR4_X1 port map( A1 => n5, A2 => n10, A3 => n14, A4 => n17, ZN => 
                           Y(22));
   U20 : AOI22_X1 port map( A1 => n255, A2 => Q(493), B1 => n254, B2 => Q(557),
                           ZN => n18);
   U21 : AOI22_X1 port map( A1 => n257, A2 => Q(653), B1 => n256, B2 => Q(461),
                           ZN => n19);
   U22 : AOI22_X1 port map( A1 => n259, A2 => Q(365), B1 => n258, B2 => Q(301),
                           ZN => n20);
   U23 : AOI22_X1 port map( A1 => n261, A2 => Q(397), B1 => n260, B2 => Q(269),
                           ZN => n21);
   U24 : NAND4_X1 port map( A1 => n18, A2 => n19, A3 => n20, A4 => n21, ZN => 
                           n22);
   U25 : AOI22_X1 port map( A1 => n263, A2 => Q(333), B1 => n262, B2 => Q(429),
                           ZN => n23);
   U26 : AOI22_X1 port map( A1 => n265, A2 => Q(237), B1 => n264, B2 => Q(141),
                           ZN => n24);
   U27 : AOI22_X1 port map( A1 => n267, A2 => Q(77), B1 => n266, B2 => Q(173), 
                           ZN => n25);
   U28 : AOI22_X1 port map( A1 => n269, A2 => Q(205), B1 => n268, B2 => Q(45), 
                           ZN => n26);
   U29 : NAND4_X1 port map( A1 => n23, A2 => n24, A3 => n25, A4 => n26, ZN => 
                           n27);
   U30 : AOI22_X1 port map( A1 => n240, A2 => Q(1005), B1 => n239, B2 => Q(941)
                           , ZN => n28);
   U31 : AOI22_X1 port map( A1 => n242, A2 => Q(973), B1 => n241, B2 => Q(909),
                           ZN => n29);
   U32 : AOI222_X1 port map( A1 => n244, A2 => Q(813), B1 => n245, B2 => Q(109)
                           , C1 => n243, C2 => Q(749), ZN => n30);
   U33 : NAND3_X1 port map( A1 => n28, A2 => n29, A3 => n30, ZN => n31);
   U34 : AOI22_X1 port map( A1 => n247, A2 => Q(845), B1 => n246, B2 => Q(717),
                           ZN => n32);
   U35 : AOI22_X1 port map( A1 => n249, A2 => Q(781), B1 => n248, B2 => Q(877),
                           ZN => n33);
   U36 : NAND4_X1 port map( A1 => n331, A2 => n332, A3 => n32, A4 => n33, ZN =>
                           n34);
   U37 : OR4_X1 port map( A1 => n22, A2 => n27, A3 => n31, A4 => n34, ZN => 
                           Y(13));
   U38 : AOI22_X1 port map( A1 => n255, A2 => Q(500), B1 => n254, B2 => Q(564),
                           ZN => n35);
   U39 : AOI22_X1 port map( A1 => n257, A2 => Q(660), B1 => n256, B2 => Q(468),
                           ZN => n36);
   U40 : AOI22_X1 port map( A1 => n259, A2 => Q(372), B1 => n258, B2 => Q(308),
                           ZN => n37);
   U41 : AOI22_X1 port map( A1 => n261, A2 => Q(404), B1 => n260, B2 => Q(276),
                           ZN => n38);
   U42 : NAND4_X1 port map( A1 => n35, A2 => n36, A3 => n37, A4 => n38, ZN => 
                           n39);
   U43 : AOI22_X1 port map( A1 => n263, A2 => Q(340), B1 => n262, B2 => Q(436),
                           ZN => n40);
   U44 : AOI22_X1 port map( A1 => n265, A2 => Q(244), B1 => n264, B2 => Q(148),
                           ZN => n41);
   U45 : AOI22_X1 port map( A1 => n267, A2 => Q(84), B1 => n266, B2 => Q(180), 
                           ZN => n42);
   U46 : AOI22_X1 port map( A1 => n269, A2 => Q(212), B1 => n268, B2 => Q(52), 
                           ZN => n43);
   U47 : NAND4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n44);
   U48 : AOI22_X1 port map( A1 => n240, A2 => Q(1012), B1 => n239, B2 => Q(948)
                           , ZN => n45);
   U49 : AOI22_X1 port map( A1 => n242, A2 => Q(980), B1 => n241, B2 => Q(916),
                           ZN => n46);
   U50 : AOI222_X1 port map( A1 => n244, A2 => Q(820), B1 => n245, B2 => Q(116)
                           , C1 => n243, C2 => Q(756), ZN => n47);
   U51 : NAND3_X1 port map( A1 => n45, A2 => n46, A3 => n47, ZN => n48);
   U52 : AOI22_X1 port map( A1 => n247, A2 => Q(852), B1 => n246, B2 => Q(724),
                           ZN => n49);
   U53 : AOI22_X1 port map( A1 => n249, A2 => Q(788), B1 => n248, B2 => Q(884),
                           ZN => n50);
   U54 : NAND4_X1 port map( A1 => n473, A2 => n474, A3 => n49, A4 => n50, ZN =>
                           n51);
   U55 : OR4_X1 port map( A1 => n39, A2 => n44, A3 => n48, A4 => n51, ZN => 
                           Y(20));
   U56 : AOI22_X1 port map( A1 => n255, A2 => Q(489), B1 => n254, B2 => Q(553),
                           ZN => n52);
   U57 : AOI22_X1 port map( A1 => n257, A2 => Q(649), B1 => n256, B2 => Q(457),
                           ZN => n53);
   U58 : AOI22_X1 port map( A1 => n259, A2 => Q(361), B1 => n258, B2 => Q(297),
                           ZN => n54);
   U59 : AOI22_X1 port map( A1 => n261, A2 => Q(393), B1 => n260, B2 => Q(265),
                           ZN => n55);
   U60 : NAND4_X1 port map( A1 => n52, A2 => n53, A3 => n54, A4 => n55, ZN => 
                           n56);
   U61 : AOI22_X1 port map( A1 => n263, A2 => Q(329), B1 => n262, B2 => Q(425),
                           ZN => n57);
   U62 : AOI22_X1 port map( A1 => n265, A2 => Q(233), B1 => n264, B2 => Q(137),
                           ZN => n58);
   U63 : AOI22_X1 port map( A1 => n267, A2 => Q(73), B1 => n266, B2 => Q(169), 
                           ZN => n59);
   U64 : AOI22_X1 port map( A1 => n269, A2 => Q(201), B1 => n268, B2 => Q(41), 
                           ZN => n60);
   U65 : NAND4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           n61);
   U66 : AOI22_X1 port map( A1 => n240, A2 => Q(1001), B1 => n239, B2 => Q(937)
                           , ZN => n62);
   U67 : AOI22_X1 port map( A1 => n242, A2 => Q(969), B1 => n241, B2 => Q(905),
                           ZN => n63);
   U68 : AOI222_X1 port map( A1 => n244, A2 => Q(809), B1 => n245, B2 => Q(105)
                           , C1 => n243, C2 => Q(745), ZN => n64);
   U69 : NAND3_X1 port map( A1 => n62, A2 => n63, A3 => n64, ZN => n65);
   U70 : AOI22_X1 port map( A1 => n247, A2 => Q(841), B1 => n246, B2 => Q(713),
                           ZN => n66);
   U71 : AOI22_X1 port map( A1 => n249, A2 => Q(777), B1 => n248, B2 => Q(873),
                           ZN => n67);
   U72 : NAND4_X1 port map( A1 => n688, A2 => n689, A3 => n66, A4 => n67, ZN =>
                           n68);
   U73 : OR4_X1 port map( A1 => n56, A2 => n61, A3 => n65, A4 => n68, ZN => 
                           Y(9));
   U74 : AOI22_X1 port map( A1 => n255, A2 => Q(491), B1 => n254, B2 => Q(555),
                           ZN => n69);
   U75 : AOI22_X1 port map( A1 => n257, A2 => Q(651), B1 => n256, B2 => Q(459),
                           ZN => n70);
   U76 : AOI22_X1 port map( A1 => n259, A2 => Q(363), B1 => n258, B2 => Q(299),
                           ZN => n71);
   U77 : AOI22_X1 port map( A1 => n261, A2 => Q(395), B1 => n260, B2 => Q(267),
                           ZN => n72);
   U78 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           n73);
   U79 : AOI22_X1 port map( A1 => n263, A2 => Q(331), B1 => n262, B2 => Q(427),
                           ZN => n74);
   U80 : AOI22_X1 port map( A1 => n265, A2 => Q(235), B1 => n264, B2 => Q(139),
                           ZN => n75);
   U81 : AOI22_X1 port map( A1 => n267, A2 => Q(75), B1 => n266, B2 => Q(171), 
                           ZN => n76);
   U82 : AOI22_X1 port map( A1 => n269, A2 => Q(203), B1 => n268, B2 => Q(43), 
                           ZN => n77);
   U83 : NAND4_X1 port map( A1 => n74, A2 => n75, A3 => n76, A4 => n77, ZN => 
                           n78);
   U84 : AOI22_X1 port map( A1 => n240, A2 => Q(1003), B1 => n239, B2 => Q(939)
                           , ZN => n79);
   U85 : AOI22_X1 port map( A1 => n242, A2 => Q(971), B1 => n241, B2 => Q(907),
                           ZN => n80);
   U86 : AOI222_X1 port map( A1 => n244, A2 => Q(811), B1 => n245, B2 => Q(107)
                           , C1 => n243, C2 => Q(747), ZN => n81);
   U87 : NAND3_X1 port map( A1 => n79, A2 => n80, A3 => n81, ZN => n82);
   U88 : AOI22_X1 port map( A1 => n247, A2 => Q(843), B1 => n246, B2 => Q(715),
                           ZN => n83);
   U89 : AOI22_X1 port map( A1 => n249, A2 => Q(779), B1 => n248, B2 => Q(875),
                           ZN => n84);
   U90 : NAND4_X1 port map( A1 => n309, A2 => n310, A3 => n83, A4 => n84, ZN =>
                           n85);
   U91 : OR4_X1 port map( A1 => n73, A2 => n78, A3 => n82, A4 => n85, ZN => 
                           Y(11));
   U92 : AOI22_X1 port map( A1 => n255, A2 => Q(487), B1 => n254, B2 => Q(551),
                           ZN => n86);
   U93 : AOI22_X1 port map( A1 => n257, A2 => Q(647), B1 => n256, B2 => Q(455),
                           ZN => n87);
   U94 : AOI22_X1 port map( A1 => n259, A2 => Q(359), B1 => n258, B2 => Q(295),
                           ZN => n88);
   U95 : AOI22_X1 port map( A1 => n261, A2 => Q(391), B1 => n260, B2 => Q(263),
                           ZN => n89);
   U96 : NAND4_X1 port map( A1 => n86, A2 => n87, A3 => n88, A4 => n89, ZN => 
                           n90);
   U97 : AOI22_X1 port map( A1 => n263, A2 => Q(327), B1 => n262, B2 => Q(423),
                           ZN => n91);
   U98 : AOI22_X1 port map( A1 => n265, A2 => Q(231), B1 => n264, B2 => Q(135),
                           ZN => n92);
   U99 : AOI22_X1 port map( A1 => n267, A2 => Q(71), B1 => n266, B2 => Q(167), 
                           ZN => n93);
   U100 : AOI22_X1 port map( A1 => n269, A2 => Q(199), B1 => n268, B2 => Q(39),
                           ZN => n94);
   U101 : NAND4_X1 port map( A1 => n91, A2 => n92, A3 => n93, A4 => n94, ZN => 
                           n95);
   U102 : AOI22_X1 port map( A1 => n240, A2 => Q(999), B1 => n239, B2 => Q(935)
                           , ZN => n96);
   U103 : AOI22_X1 port map( A1 => n242, A2 => Q(967), B1 => n241, B2 => Q(903)
                           , ZN => n97);
   U104 : AOI222_X1 port map( A1 => n244, A2 => Q(807), B1 => n245, B2 => 
                           Q(103), C1 => n243, C2 => Q(743), ZN => n98);
   U105 : NAND3_X1 port map( A1 => n96, A2 => n97, A3 => n98, ZN => n99);
   U106 : AOI22_X1 port map( A1 => n247, A2 => Q(839), B1 => n246, B2 => Q(711)
                           , ZN => n100);
   U107 : AOI22_X1 port map( A1 => n249, A2 => Q(775), B1 => n248, B2 => Q(871)
                           , ZN => n101);
   U108 : NAND4_X1 port map( A1 => n669, A2 => n670, A3 => n100, A4 => n101, ZN
                           => n102);
   U109 : OR4_X1 port map( A1 => n90, A2 => n95, A3 => n99, A4 => n102, ZN => 
                           Y(7));
   U110 : AOI22_X1 port map( A1 => n255, A2 => Q(488), B1 => n254, B2 => Q(552)
                           , ZN => n103);
   U111 : AOI22_X1 port map( A1 => n257, A2 => Q(648), B1 => n256, B2 => Q(456)
                           , ZN => n104);
   U112 : AOI22_X1 port map( A1 => n259, A2 => Q(360), B1 => n258, B2 => Q(296)
                           , ZN => n105);
   U113 : AOI22_X1 port map( A1 => n261, A2 => Q(392), B1 => n260, B2 => Q(264)
                           , ZN => n106);
   U114 : NAND4_X1 port map( A1 => n103, A2 => n104, A3 => n105, A4 => n106, ZN
                           => n107);
   U115 : AOI22_X1 port map( A1 => n263, A2 => Q(328), B1 => n262, B2 => Q(424)
                           , ZN => n108);
   U116 : AOI22_X1 port map( A1 => n265, A2 => Q(232), B1 => n264, B2 => Q(136)
                           , ZN => n109);
   U117 : AOI22_X1 port map( A1 => n267, A2 => Q(72), B1 => n266, B2 => Q(168),
                           ZN => n110);
   U118 : AOI22_X1 port map( A1 => n269, A2 => Q(200), B1 => n268, B2 => Q(40),
                           ZN => n111);
   U119 : NAND4_X1 port map( A1 => n108, A2 => n109, A3 => n110, A4 => n111, ZN
                           => n112);
   U120 : AOI22_X1 port map( A1 => n240, A2 => Q(1000), B1 => n239, B2 => 
                           Q(936), ZN => n113);
   U121 : AOI22_X1 port map( A1 => n242, A2 => Q(968), B1 => n241, B2 => Q(904)
                           , ZN => n114);
   U122 : AOI222_X1 port map( A1 => n244, A2 => Q(808), B1 => n245, B2 => 
                           Q(104), C1 => n243, C2 => Q(744), ZN => n115);
   U123 : NAND3_X1 port map( A1 => n113, A2 => n114, A3 => n115, ZN => n116);
   U124 : AOI22_X1 port map( A1 => n247, A2 => Q(840), B1 => n246, B2 => Q(712)
                           , ZN => n117);
   U125 : AOI22_X1 port map( A1 => n249, A2 => Q(776), B1 => n248, B2 => Q(872)
                           , ZN => n118);
   U126 : NAND4_X1 port map( A1 => n671, A2 => n672, A3 => n117, A4 => n118, ZN
                           => n119);
   U127 : OR4_X1 port map( A1 => n107, A2 => n112, A3 => n116, A4 => n119, ZN 
                           => Y(8));
   U128 : AOI22_X1 port map( A1 => n255, A2 => Q(485), B1 => n254, B2 => Q(549)
                           , ZN => n120);
   U129 : AOI22_X1 port map( A1 => n257, A2 => Q(645), B1 => n256, B2 => Q(453)
                           , ZN => n121);
   U130 : AOI22_X1 port map( A1 => n259, A2 => Q(357), B1 => n258, B2 => Q(293)
                           , ZN => n122);
   U131 : AOI22_X1 port map( A1 => n261, A2 => Q(389), B1 => n260, B2 => Q(261)
                           , ZN => n123);
   U132 : NAND4_X1 port map( A1 => n120, A2 => n121, A3 => n122, A4 => n123, ZN
                           => n124);
   U133 : AOI22_X1 port map( A1 => n263, A2 => Q(325), B1 => n262, B2 => Q(421)
                           , ZN => n125);
   U134 : AOI22_X1 port map( A1 => n265, A2 => Q(229), B1 => n264, B2 => Q(133)
                           , ZN => n126);
   U135 : AOI22_X1 port map( A1 => n267, A2 => Q(69), B1 => n266, B2 => Q(165),
                           ZN => n127);
   U136 : AOI22_X1 port map( A1 => n269, A2 => Q(197), B1 => n268, B2 => Q(37),
                           ZN => n128);
   U137 : NAND4_X1 port map( A1 => n125, A2 => n126, A3 => n127, A4 => n128, ZN
                           => n129);
   U138 : AOI22_X1 port map( A1 => n240, A2 => Q(997), B1 => n239, B2 => Q(933)
                           , ZN => n130);
   U139 : AOI22_X1 port map( A1 => n242, A2 => Q(965), B1 => n241, B2 => Q(901)
                           , ZN => n131);
   U140 : AOI222_X1 port map( A1 => n244, A2 => Q(805), B1 => n245, B2 => 
                           Q(101), C1 => n243, C2 => Q(741), ZN => n132);
   U141 : NAND3_X1 port map( A1 => n130, A2 => n131, A3 => n132, ZN => n133);
   U142 : AOI22_X1 port map( A1 => n247, A2 => Q(837), B1 => n246, B2 => Q(709)
                           , ZN => n134);
   U143 : AOI22_X1 port map( A1 => n249, A2 => Q(773), B1 => n248, B2 => Q(869)
                           , ZN => n135);
   U144 : NAND4_X1 port map( A1 => n665, A2 => n666, A3 => n134, A4 => n135, ZN
                           => n136);
   U145 : OR4_X1 port map( A1 => n124, A2 => n129, A3 => n133, A4 => n136, ZN 
                           => Y(5));
   U146 : AOI22_X1 port map( A1 => n255, A2 => Q(486), B1 => n254, B2 => Q(550)
                           , ZN => n137);
   U147 : AOI22_X1 port map( A1 => n257, A2 => Q(646), B1 => n256, B2 => Q(454)
                           , ZN => n138);
   U148 : AOI22_X1 port map( A1 => n259, A2 => Q(358), B1 => n258, B2 => Q(294)
                           , ZN => n139);
   U149 : AOI22_X1 port map( A1 => n261, A2 => Q(390), B1 => n260, B2 => Q(262)
                           , ZN => n140);
   U150 : NAND4_X1 port map( A1 => n137, A2 => n138, A3 => n139, A4 => n140, ZN
                           => n141);
   U151 : AOI22_X1 port map( A1 => n263, A2 => Q(326), B1 => n262, B2 => Q(422)
                           , ZN => n142);
   U152 : AOI22_X1 port map( A1 => n265, A2 => Q(230), B1 => n264, B2 => Q(134)
                           , ZN => n143);
   U153 : AOI22_X1 port map( A1 => n267, A2 => Q(70), B1 => n266, B2 => Q(166),
                           ZN => n144);
   U154 : AOI22_X1 port map( A1 => n269, A2 => Q(198), B1 => n268, B2 => Q(38),
                           ZN => n145);
   U155 : NAND4_X1 port map( A1 => n142, A2 => n143, A3 => n144, A4 => n145, ZN
                           => n146);
   U156 : AOI22_X1 port map( A1 => n240, A2 => Q(998), B1 => n239, B2 => Q(934)
                           , ZN => n147);
   U157 : AOI22_X1 port map( A1 => n242, A2 => Q(966), B1 => n241, B2 => Q(902)
                           , ZN => n148);
   U158 : AOI222_X1 port map( A1 => n244, A2 => Q(806), B1 => n245, B2 => 
                           Q(102), C1 => n243, C2 => Q(742), ZN => n149);
   U159 : NAND3_X1 port map( A1 => n147, A2 => n148, A3 => n149, ZN => n150);
   U160 : AOI22_X1 port map( A1 => n247, A2 => Q(838), B1 => n246, B2 => Q(710)
                           , ZN => n151);
   U161 : AOI22_X1 port map( A1 => n249, A2 => Q(774), B1 => n248, B2 => Q(870)
                           , ZN => n152);
   U162 : NAND4_X1 port map( A1 => n667, A2 => n668, A3 => n151, A4 => n152, ZN
                           => n153);
   U163 : OR4_X1 port map( A1 => n141, A2 => n146, A3 => n150, A4 => n153, ZN 
                           => Y(6));
   U164 : AOI22_X1 port map( A1 => n255, A2 => Q(483), B1 => n254, B2 => Q(547)
                           , ZN => n154);
   U165 : AOI22_X1 port map( A1 => n257, A2 => Q(643), B1 => n256, B2 => Q(451)
                           , ZN => n155);
   U166 : AOI22_X1 port map( A1 => n259, A2 => Q(355), B1 => n258, B2 => Q(291)
                           , ZN => n156);
   U167 : AOI22_X1 port map( A1 => n261, A2 => Q(387), B1 => n260, B2 => Q(259)
                           , ZN => n157);
   U168 : NAND4_X1 port map( A1 => n154, A2 => n155, A3 => n156, A4 => n157, ZN
                           => n158);
   U169 : AOI22_X1 port map( A1 => n263, A2 => Q(323), B1 => n262, B2 => Q(419)
                           , ZN => n159);
   U170 : AOI22_X1 port map( A1 => n265, A2 => Q(227), B1 => n264, B2 => Q(131)
                           , ZN => n160);
   U171 : AOI22_X1 port map( A1 => n267, A2 => Q(67), B1 => n266, B2 => Q(163),
                           ZN => n161);
   U172 : AOI22_X1 port map( A1 => n269, A2 => Q(195), B1 => n268, B2 => Q(35),
                           ZN => n162);
   U173 : NAND4_X1 port map( A1 => n159, A2 => n160, A3 => n161, A4 => n162, ZN
                           => n163);
   U174 : AOI22_X1 port map( A1 => n240, A2 => Q(995), B1 => n239, B2 => Q(931)
                           , ZN => n164);
   U175 : AOI22_X1 port map( A1 => n242, A2 => Q(963), B1 => n241, B2 => Q(899)
                           , ZN => n165);
   U176 : AOI222_X1 port map( A1 => n244, A2 => Q(803), B1 => n245, B2 => Q(99)
                           , C1 => n243, C2 => Q(739), ZN => n166);
   U177 : NAND3_X1 port map( A1 => n164, A2 => n165, A3 => n166, ZN => n167);
   U178 : AOI22_X1 port map( A1 => n247, A2 => Q(835), B1 => n246, B2 => Q(707)
                           , ZN => n168);
   U179 : AOI22_X1 port map( A1 => n249, A2 => Q(771), B1 => n248, B2 => Q(867)
                           , ZN => n169);
   U180 : NAND4_X1 port map( A1 => n661, A2 => n662, A3 => n168, A4 => n169, ZN
                           => n170);
   U181 : OR4_X1 port map( A1 => n158, A2 => n163, A3 => n167, A4 => n170, ZN 
                           => Y(3));
   U182 : AOI22_X1 port map( A1 => n255, A2 => Q(484), B1 => n254, B2 => Q(548)
                           , ZN => n171);
   U183 : AOI22_X1 port map( A1 => n257, A2 => Q(644), B1 => n256, B2 => Q(452)
                           , ZN => n172);
   U184 : AOI22_X1 port map( A1 => n259, A2 => Q(356), B1 => n258, B2 => Q(292)
                           , ZN => n173);
   U185 : AOI22_X1 port map( A1 => n261, A2 => Q(388), B1 => n260, B2 => Q(260)
                           , ZN => n174);
   U186 : NAND4_X1 port map( A1 => n171, A2 => n172, A3 => n173, A4 => n174, ZN
                           => n175);
   U187 : AOI22_X1 port map( A1 => n263, A2 => Q(324), B1 => n262, B2 => Q(420)
                           , ZN => n176);
   U188 : AOI22_X1 port map( A1 => n265, A2 => Q(228), B1 => n264, B2 => Q(132)
                           , ZN => n177);
   U189 : AOI22_X1 port map( A1 => n267, A2 => Q(68), B1 => n266, B2 => Q(164),
                           ZN => n178);
   U190 : AOI22_X1 port map( A1 => n269, A2 => Q(196), B1 => n268, B2 => Q(36),
                           ZN => n179);
   U191 : NAND4_X1 port map( A1 => n176, A2 => n177, A3 => n178, A4 => n179, ZN
                           => n180);
   U192 : AOI22_X1 port map( A1 => n240, A2 => Q(996), B1 => n239, B2 => Q(932)
                           , ZN => n181);
   U193 : AOI22_X1 port map( A1 => n242, A2 => Q(964), B1 => n241, B2 => Q(900)
                           , ZN => n182);
   U194 : AOI222_X1 port map( A1 => n244, A2 => Q(804), B1 => n245, B2 => 
                           Q(100), C1 => n243, C2 => Q(740), ZN => n183);
   U195 : NAND3_X1 port map( A1 => n181, A2 => n182, A3 => n183, ZN => n184);
   U196 : AOI22_X1 port map( A1 => n247, A2 => Q(836), B1 => n246, B2 => Q(708)
                           , ZN => n185);
   U197 : AOI22_X1 port map( A1 => n249, A2 => Q(772), B1 => n248, B2 => Q(868)
                           , ZN => n186);
   U198 : NAND4_X1 port map( A1 => n663, A2 => n664, A3 => n185, A4 => n186, ZN
                           => n187);
   U199 : OR4_X1 port map( A1 => n175, A2 => n180, A3 => n184, A4 => n187, ZN 
                           => Y(4));
   U200 : AOI22_X1 port map( A1 => n690, A2 => Q(546), B1 => n691, B2 => Q(482)
                           , ZN => n188);
   U201 : AOI22_X1 port map( A1 => n692, A2 => Q(450), B1 => n693, B2 => Q(642)
                           , ZN => n189);
   U202 : AOI22_X1 port map( A1 => n694, A2 => Q(290), B1 => n695, B2 => Q(354)
                           , ZN => n190);
   U203 : AOI22_X1 port map( A1 => n696, A2 => Q(258), B1 => n697, B2 => Q(386)
                           , ZN => n191);
   U204 : NAND4_X1 port map( A1 => n188, A2 => n189, A3 => n190, A4 => n191, ZN
                           => n192);
   U205 : AOI22_X1 port map( A1 => n698, A2 => Q(418), B1 => n699, B2 => Q(322)
                           , ZN => n193);
   U206 : AOI22_X1 port map( A1 => n700, A2 => Q(130), B1 => n701, B2 => Q(226)
                           , ZN => n194);
   U207 : AOI22_X1 port map( A1 => n702, A2 => Q(162), B1 => n703, B2 => Q(66),
                           ZN => n195);
   U208 : AOI22_X1 port map( A1 => n704, A2 => Q(34), B1 => n705, B2 => Q(194),
                           ZN => n196);
   U209 : NAND4_X1 port map( A1 => n193, A2 => n194, A3 => n195, A4 => n196, ZN
                           => n197);
   U210 : AOI22_X1 port map( A1 => n673, A2 => Q(930), B1 => n674, B2 => Q(994)
                           , ZN => n198);
   U211 : AOI22_X1 port map( A1 => n675, A2 => Q(898), B1 => n676, B2 => Q(962)
                           , ZN => n199);
   U212 : AOI222_X1 port map( A1 => n677, A2 => Q(738), B1 => n678, B2 => 
                           Q(802), C1 => n679, C2 => Q(98), ZN => n200);
   U213 : NAND3_X1 port map( A1 => n198, A2 => n199, A3 => n200, ZN => n201);
   U214 : AOI22_X1 port map( A1 => n680, A2 => Q(706), B1 => n681, B2 => Q(834)
                           , ZN => n202);
   U215 : AOI22_X1 port map( A1 => n682, A2 => Q(866), B1 => n683, B2 => Q(770)
                           , ZN => n203);
   U216 : NAND4_X1 port map( A1 => n637, A2 => n638, A3 => n202, A4 => n203, ZN
                           => n204);
   U217 : OR4_X1 port map( A1 => n192, A2 => n197, A3 => n201, A4 => n204, ZN 
                           => Y(2));
   U218 : AOI22_X1 port map( A1 => n255, A2 => Q(511), B1 => n254, B2 => Q(575)
                           , ZN => n205);
   U219 : AOI22_X1 port map( A1 => n257, A2 => Q(671), B1 => n256, B2 => Q(479)
                           , ZN => n206);
   U220 : AOI22_X1 port map( A1 => n259, A2 => Q(383), B1 => n258, B2 => Q(319)
                           , ZN => n207);
   U221 : AOI22_X1 port map( A1 => n261, A2 => Q(415), B1 => n260, B2 => Q(287)
                           , ZN => n208);
   U222 : NAND4_X1 port map( A1 => n205, A2 => n206, A3 => n207, A4 => n208, ZN
                           => n209);
   U223 : AOI22_X1 port map( A1 => n263, A2 => Q(351), B1 => n262, B2 => Q(447)
                           , ZN => n210);
   U224 : AOI22_X1 port map( A1 => n265, A2 => Q(255), B1 => n264, B2 => Q(159)
                           , ZN => n211);
   U225 : AOI22_X1 port map( A1 => n267, A2 => Q(95), B1 => n266, B2 => Q(191),
                           ZN => n212);
   U226 : AOI22_X1 port map( A1 => n269, A2 => Q(223), B1 => n268, B2 => Q(63),
                           ZN => n213);
   U227 : NAND4_X1 port map( A1 => n210, A2 => n211, A3 => n212, A4 => n213, ZN
                           => n214);
   U228 : AOI22_X1 port map( A1 => n240, A2 => Q(1023), B1 => n239, B2 => 
                           Q(959), ZN => n215);
   U229 : AOI22_X1 port map( A1 => n242, A2 => Q(991), B1 => n241, B2 => Q(927)
                           , ZN => n216);
   U230 : AOI222_X1 port map( A1 => n244, A2 => Q(831), B1 => n245, B2 => 
                           Q(127), C1 => n243, C2 => Q(767), ZN => n217);
   U231 : NAND3_X1 port map( A1 => n215, A2 => n216, A3 => n217, ZN => n218);
   U232 : AOI22_X1 port map( A1 => n247, A2 => Q(863), B1 => n246, B2 => Q(735)
                           , ZN => n219);
   U233 : AOI22_X1 port map( A1 => n249, A2 => Q(799), B1 => n248, B2 => Q(895)
                           , ZN => n220);
   U234 : NAND4_X1 port map( A1 => n659, A2 => n660, A3 => n219, A4 => n220, ZN
                           => n221);
   U235 : OR4_X1 port map( A1 => n209, A2 => n214, A3 => n218, A4 => n221, ZN 
                           => Y(31));
   U236 : AOI22_X1 port map( A1 => n255, A2 => Q(480), B1 => n254, B2 => Q(544)
                           , ZN => n222);
   U237 : AOI22_X1 port map( A1 => n257, A2 => Q(640), B1 => n256, B2 => Q(448)
                           , ZN => n223);
   U238 : AOI22_X1 port map( A1 => n259, A2 => Q(352), B1 => n258, B2 => Q(288)
                           , ZN => n224);
   U239 : AOI22_X1 port map( A1 => n261, A2 => Q(384), B1 => n260, B2 => Q(256)
                           , ZN => n225);
   U240 : NAND4_X1 port map( A1 => n222, A2 => n223, A3 => n224, A4 => n225, ZN
                           => n226);
   U241 : AOI22_X1 port map( A1 => n263, A2 => Q(320), B1 => n262, B2 => Q(416)
                           , ZN => n227);
   U242 : AOI22_X1 port map( A1 => n265, A2 => Q(224), B1 => n264, B2 => Q(128)
                           , ZN => n228);
   U243 : AOI22_X1 port map( A1 => n267, A2 => Q(64), B1 => n266, B2 => Q(160),
                           ZN => n229);
   U244 : AOI22_X1 port map( A1 => n269, A2 => Q(192), B1 => n268, B2 => Q(32),
                           ZN => n230);
   U245 : NAND4_X1 port map( A1 => n227, A2 => n228, A3 => n229, A4 => n230, ZN
                           => n231);
   U246 : AOI22_X1 port map( A1 => n240, A2 => Q(992), B1 => n239, B2 => Q(928)
                           , ZN => n232);
   U247 : AOI22_X1 port map( A1 => n242, A2 => Q(960), B1 => n241, B2 => Q(896)
                           , ZN => n233);
   U248 : AOI222_X1 port map( A1 => n244, A2 => Q(800), B1 => n245, B2 => Q(96)
                           , C1 => n243, C2 => Q(736), ZN => n234);
   U249 : NAND3_X1 port map( A1 => n232, A2 => n233, A3 => n234, ZN => n235);
   U250 : AOI22_X1 port map( A1 => n247, A2 => Q(832), B1 => n246, B2 => Q(704)
                           , ZN => n236);
   U251 : AOI22_X1 port map( A1 => n249, A2 => Q(768), B1 => n248, B2 => Q(864)
                           , ZN => n237);
   U252 : NAND4_X1 port map( A1 => n274, A2 => n275, A3 => n236, A4 => n237, ZN
                           => n238);
   U253 : OR4_X1 port map( A1 => n226, A2 => n231, A3 => n235, A4 => n238, ZN 
                           => Y(0));
   U254 : OR4_X1 port map( A1 => n472, A2 => n471, A3 => n470, A4 => n469, ZN 
                           => Y(1));
   U255 : OR4_X1 port map( A1 => n308, A2 => n307, A3 => n306, A4 => n305, ZN 
                           => Y(10));
   U256 : OR4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN 
                           => Y(12));
   U257 : OR4_X1 port map( A1 => n352, A2 => n351, A3 => n350, A4 => n349, ZN 
                           => Y(14));
   U258 : OR4_X1 port map( A1 => n372, A2 => n371, A3 => n370, A4 => n369, ZN 
                           => Y(15));
   U259 : OR4_X1 port map( A1 => n392, A2 => n391, A3 => n390, A4 => n389, ZN 
                           => Y(16));
   U260 : OR4_X1 port map( A1 => n412, A2 => n411, A3 => n410, A4 => n409, ZN 
                           => Y(17));
   U261 : OR4_X1 port map( A1 => n432, A2 => n431, A3 => n430, A4 => n429, ZN 
                           => Y(18));
   U262 : OR4_X1 port map( A1 => n452, A2 => n451, A3 => n450, A4 => n449, ZN 
                           => Y(19));
   U263 : OR4_X1 port map( A1 => n494, A2 => n493, A3 => n492, A4 => n491, ZN 
                           => Y(21));
   U264 : OR4_X1 port map( A1 => n516, A2 => n515, A3 => n514, A4 => n513, ZN 
                           => Y(23));
   U265 : OR4_X1 port map( A1 => n536, A2 => n535, A3 => n534, A4 => n533, ZN 
                           => Y(24));
   U266 : OR4_X1 port map( A1 => n556, A2 => n555, A3 => n554, A4 => n553, ZN 
                           => Y(25));
   U267 : OR4_X1 port map( A1 => n576, A2 => n575, A3 => n574, A4 => n573, ZN 
                           => Y(26));
   U268 : OR4_X1 port map( A1 => n596, A2 => n595, A3 => n594, A4 => n593, ZN 
                           => Y(27));
   U269 : OR4_X1 port map( A1 => n616, A2 => n615, A3 => n614, A4 => n613, ZN 
                           => Y(28));
   U270 : OR4_X1 port map( A1 => n636, A2 => n635, A3 => n634, A4 => n633, ZN 
                           => Y(29));
   U271 : BUF_X1 port map( A => n704, Z => n268);
   U272 : BUF_X1 port map( A => n705, Z => n269);
   U273 : BUF_X1 port map( A => n702, Z => n266);
   U274 : BUF_X1 port map( A => n703, Z => n267);
   U275 : BUF_X1 port map( A => n700, Z => n264);
   U276 : BUF_X1 port map( A => n701, Z => n265);
   U277 : BUF_X1 port map( A => n698, Z => n262);
   U278 : BUF_X1 port map( A => n699, Z => n263);
   U279 : BUF_X1 port map( A => n696, Z => n260);
   U280 : BUF_X1 port map( A => n697, Z => n261);
   U281 : BUF_X1 port map( A => n694, Z => n258);
   U282 : BUF_X1 port map( A => n695, Z => n259);
   U283 : BUF_X1 port map( A => n692, Z => n256);
   U284 : BUF_X1 port map( A => n693, Z => n257);
   U285 : BUF_X1 port map( A => n690, Z => n254);
   U286 : BUF_X1 port map( A => n691, Z => n255);
   U287 : BUF_X1 port map( A => n686, Z => n252);
   U288 : BUF_X1 port map( A => n687, Z => n253);
   U289 : BUF_X1 port map( A => n684, Z => n250);
   U290 : BUF_X1 port map( A => n685, Z => n251);
   U291 : BUF_X1 port map( A => n682, Z => n248);
   U292 : BUF_X1 port map( A => n683, Z => n249);
   U293 : BUF_X1 port map( A => n680, Z => n246);
   U294 : BUF_X1 port map( A => n681, Z => n247);
   U295 : BUF_X1 port map( A => n679, Z => n245);
   U296 : BUF_X1 port map( A => n677, Z => n243);
   U297 : BUF_X1 port map( A => n678, Z => n244);
   U298 : BUF_X1 port map( A => n675, Z => n241);
   U299 : BUF_X1 port map( A => n676, Z => n242);
   U300 : BUF_X1 port map( A => n673, Z => n239);
   U301 : BUF_X1 port map( A => n674, Z => n240);
   U302 : OR4_X1 port map( A1 => n658, A2 => n657, A3 => n656, A4 => n655, ZN 
                           => Y(30));
   U303 : OR2_X1 port map( A1 => S(1), A2 => S(2), ZN => n287);
   U304 : OR2_X1 port map( A1 => n270, A2 => S(1), ZN => n284);
   U305 : NAND2_X1 port map( A1 => S(1), A2 => S(2), ZN => n286);
   U306 : NAND3_X1 port map( A1 => S(3), A2 => S(4), A3 => S(0), ZN => n273);
   U307 : NOR2_X1 port map( A1 => n286, A2 => n273, ZN => n674);
   U308 : INV_X1 port map( A => S(2), ZN => n270);
   U309 : NOR2_X1 port map( A1 => n273, A2 => n284, ZN => n673);
   U310 : INV_X1 port map( A => S(0), ZN => n271);
   U311 : NAND3_X1 port map( A1 => S(4), A2 => S(3), A3 => n271, ZN => n272);
   U312 : NOR2_X1 port map( A1 => n286, A2 => n272, ZN => n676);
   U313 : NOR2_X1 port map( A1 => n284, A2 => n272, ZN => n675);
   U314 : NOR2_X1 port map( A1 => n273, A2 => n287, ZN => n678);
   U315 : INV_X1 port map( A => S(3), ZN => n281);
   U316 : NAND3_X1 port map( A1 => S(4), A2 => S(0), A3 => n281, ZN => n277);
   U317 : NOR2_X1 port map( A1 => n286, A2 => n277, ZN => n677);
   U318 : NAND2_X1 port map( A1 => S(1), A2 => n270, ZN => n283);
   U319 : INV_X1 port map( A => S(4), ZN => n276);
   U320 : NAND3_X1 port map( A1 => S(0), A2 => n281, A3 => n276, ZN => n288);
   U321 : NOR2_X1 port map( A1 => n283, A2 => n288, ZN => n679);
   U322 : NOR2_X1 port map( A1 => n283, A2 => n272, ZN => n681);
   U323 : NAND3_X1 port map( A1 => S(4), A2 => n281, A3 => n271, ZN => n278);
   U324 : NOR2_X1 port map( A1 => n286, A2 => n278, ZN => n680);
   U325 : NOR2_X1 port map( A1 => n272, A2 => n287, ZN => n683);
   U326 : NOR2_X1 port map( A1 => n283, A2 => n273, ZN => n682);
   U327 : NOR2_X1 port map( A1 => n284, A2 => n277, ZN => n685);
   U328 : NOR2_X1 port map( A1 => n283, A2 => n278, ZN => n684);
   U329 : AOI22_X1 port map( A1 => n251, A2 => Q(672), B1 => n250, B2 => Q(576)
                           , ZN => n275);
   U330 : NOR2_X1 port map( A1 => n287, A2 => n278, ZN => n687);
   U331 : NOR2_X1 port map( A1 => n283, A2 => n277, ZN => n686);
   U332 : AOI22_X1 port map( A1 => n253, A2 => Q(512), B1 => n252, B2 => Q(608)
                           , ZN => n274);
   U333 : NAND3_X1 port map( A1 => S(3), A2 => S(0), A3 => n276, ZN => n280);
   U334 : NOR2_X1 port map( A1 => n286, A2 => n280, ZN => n691);
   U335 : NOR2_X1 port map( A1 => n287, A2 => n277, ZN => n690);
   U336 : NOR2_X1 port map( A1 => n284, A2 => n278, ZN => n693);
   U337 : NOR2_X1 port map( A1 => S(4), A2 => S(0), ZN => n282);
   U338 : NAND2_X1 port map( A1 => S(3), A2 => n282, ZN => n279);
   U339 : NOR2_X1 port map( A1 => n286, A2 => n279, ZN => n692);
   U340 : NOR2_X1 port map( A1 => n283, A2 => n280, ZN => n695);
   U341 : NOR2_X1 port map( A1 => n287, A2 => n280, ZN => n694);
   U342 : NOR2_X1 port map( A1 => n284, A2 => n279, ZN => n697);
   U343 : NOR2_X1 port map( A1 => n287, A2 => n279, ZN => n696);
   U344 : NOR2_X1 port map( A1 => n283, A2 => n279, ZN => n699);
   U345 : NOR2_X1 port map( A1 => n284, A2 => n280, ZN => n698);
   U346 : NOR2_X1 port map( A1 => n288, A2 => n286, ZN => n701);
   U347 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => n285);
   U348 : NOR2_X1 port map( A1 => n284, A2 => n285, ZN => n700);
   U349 : NOR2_X1 port map( A1 => n283, A2 => n285, ZN => n703);
   U350 : NOR2_X1 port map( A1 => n288, A2 => n284, ZN => n702);
   U351 : NOR2_X1 port map( A1 => n286, A2 => n285, ZN => n705);
   U352 : NOR2_X1 port map( A1 => n288, A2 => n287, ZN => n704);
   U353 : AOI22_X1 port map( A1 => n674, A2 => Q(1002), B1 => n673, B2 => 
                           Q(938), ZN => n292);
   U354 : AOI22_X1 port map( A1 => n676, A2 => Q(970), B1 => n675, B2 => Q(906)
                           , ZN => n291);
   U355 : AOI22_X1 port map( A1 => n678, A2 => Q(810), B1 => n677, B2 => Q(746)
                           , ZN => n290);
   U356 : NAND2_X1 port map( A1 => n679, A2 => Q(106), ZN => n289);
   U357 : NAND4_X1 port map( A1 => n292, A2 => n291, A3 => n290, A4 => n289, ZN
                           => n308);
   U358 : AOI22_X1 port map( A1 => n681, A2 => Q(842), B1 => n680, B2 => Q(714)
                           , ZN => n296);
   U359 : AOI22_X1 port map( A1 => n683, A2 => Q(778), B1 => n682, B2 => Q(874)
                           , ZN => n295);
   U360 : AOI22_X1 port map( A1 => n685, A2 => Q(682), B1 => n684, B2 => Q(586)
                           , ZN => n294);
   U361 : AOI22_X1 port map( A1 => n687, A2 => Q(522), B1 => n686, B2 => Q(618)
                           , ZN => n293);
   U362 : NAND4_X1 port map( A1 => n296, A2 => n295, A3 => n294, A4 => n293, ZN
                           => n307);
   U363 : AOI22_X1 port map( A1 => n691, A2 => Q(490), B1 => n690, B2 => Q(554)
                           , ZN => n300);
   U364 : AOI22_X1 port map( A1 => n693, A2 => Q(650), B1 => n692, B2 => Q(458)
                           , ZN => n299);
   U365 : AOI22_X1 port map( A1 => n695, A2 => Q(362), B1 => n694, B2 => Q(298)
                           , ZN => n298);
   U366 : AOI22_X1 port map( A1 => n697, A2 => Q(394), B1 => n696, B2 => Q(266)
                           , ZN => n297);
   U367 : NAND4_X1 port map( A1 => n300, A2 => n299, A3 => n298, A4 => n297, ZN
                           => n306);
   U368 : AOI22_X1 port map( A1 => n699, A2 => Q(330), B1 => n698, B2 => Q(426)
                           , ZN => n304);
   U369 : AOI22_X1 port map( A1 => n701, A2 => Q(234), B1 => n700, B2 => Q(138)
                           , ZN => n303);
   U370 : AOI22_X1 port map( A1 => n703, A2 => Q(74), B1 => n702, B2 => Q(170),
                           ZN => n302);
   U371 : AOI22_X1 port map( A1 => n705, A2 => Q(202), B1 => n704, B2 => Q(42),
                           ZN => n301);
   U372 : NAND4_X1 port map( A1 => n304, A2 => n303, A3 => n302, A4 => n301, ZN
                           => n305);
   U373 : AOI22_X1 port map( A1 => n251, A2 => Q(683), B1 => n250, B2 => Q(587)
                           , ZN => n310);
   U374 : AOI22_X1 port map( A1 => n253, A2 => Q(523), B1 => n252, B2 => Q(619)
                           , ZN => n309);
   U375 : AOI22_X1 port map( A1 => n674, A2 => Q(1004), B1 => n673, B2 => 
                           Q(940), ZN => n314);
   U376 : AOI22_X1 port map( A1 => n676, A2 => Q(972), B1 => n675, B2 => Q(908)
                           , ZN => n313);
   U377 : AOI22_X1 port map( A1 => n678, A2 => Q(812), B1 => n677, B2 => Q(748)
                           , ZN => n312);
   U378 : NAND2_X1 port map( A1 => n679, A2 => Q(108), ZN => n311);
   U379 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => n330);
   U380 : AOI22_X1 port map( A1 => n681, A2 => Q(844), B1 => n680, B2 => Q(716)
                           , ZN => n318);
   U381 : AOI22_X1 port map( A1 => n683, A2 => Q(780), B1 => n682, B2 => Q(876)
                           , ZN => n317);
   U382 : AOI22_X1 port map( A1 => n685, A2 => Q(684), B1 => n684, B2 => Q(588)
                           , ZN => n316);
   U383 : AOI22_X1 port map( A1 => n687, A2 => Q(524), B1 => n686, B2 => Q(620)
                           , ZN => n315);
   U384 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => n329);
   U385 : AOI22_X1 port map( A1 => n691, A2 => Q(492), B1 => n690, B2 => Q(556)
                           , ZN => n322);
   U386 : AOI22_X1 port map( A1 => n693, A2 => Q(652), B1 => n692, B2 => Q(460)
                           , ZN => n321);
   U387 : AOI22_X1 port map( A1 => n695, A2 => Q(364), B1 => n694, B2 => Q(300)
                           , ZN => n320);
   U388 : AOI22_X1 port map( A1 => n697, A2 => Q(396), B1 => n696, B2 => Q(268)
                           , ZN => n319);
   U389 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => n328);
   U390 : AOI22_X1 port map( A1 => n699, A2 => Q(332), B1 => n698, B2 => Q(428)
                           , ZN => n326);
   U391 : AOI22_X1 port map( A1 => n701, A2 => Q(236), B1 => n700, B2 => Q(140)
                           , ZN => n325);
   U392 : AOI22_X1 port map( A1 => n703, A2 => Q(76), B1 => n702, B2 => Q(172),
                           ZN => n324);
   U393 : AOI22_X1 port map( A1 => n705, A2 => Q(204), B1 => n704, B2 => Q(44),
                           ZN => n323);
   U394 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => n327);
   U395 : AOI22_X1 port map( A1 => n251, A2 => Q(685), B1 => n250, B2 => Q(589)
                           , ZN => n332);
   U396 : AOI22_X1 port map( A1 => n253, A2 => Q(525), B1 => n252, B2 => Q(621)
                           , ZN => n331);
   U397 : AOI22_X1 port map( A1 => n674, A2 => Q(1006), B1 => n673, B2 => 
                           Q(942), ZN => n336);
   U398 : AOI22_X1 port map( A1 => n676, A2 => Q(974), B1 => n675, B2 => Q(910)
                           , ZN => n335);
   U399 : AOI22_X1 port map( A1 => n678, A2 => Q(814), B1 => n677, B2 => Q(750)
                           , ZN => n334);
   U400 : NAND2_X1 port map( A1 => n679, A2 => Q(110), ZN => n333);
   U401 : NAND4_X1 port map( A1 => n336, A2 => n335, A3 => n334, A4 => n333, ZN
                           => n352);
   U402 : AOI22_X1 port map( A1 => n681, A2 => Q(846), B1 => n680, B2 => Q(718)
                           , ZN => n340);
   U403 : AOI22_X1 port map( A1 => n683, A2 => Q(782), B1 => n682, B2 => Q(878)
                           , ZN => n339);
   U404 : AOI22_X1 port map( A1 => n685, A2 => Q(686), B1 => n684, B2 => Q(590)
                           , ZN => n338);
   U405 : AOI22_X1 port map( A1 => n687, A2 => Q(526), B1 => n686, B2 => Q(622)
                           , ZN => n337);
   U406 : NAND4_X1 port map( A1 => n340, A2 => n339, A3 => n338, A4 => n337, ZN
                           => n351);
   U407 : AOI22_X1 port map( A1 => n691, A2 => Q(494), B1 => n690, B2 => Q(558)
                           , ZN => n344);
   U408 : AOI22_X1 port map( A1 => n693, A2 => Q(654), B1 => n692, B2 => Q(462)
                           , ZN => n343);
   U409 : AOI22_X1 port map( A1 => n695, A2 => Q(366), B1 => n694, B2 => Q(302)
                           , ZN => n342);
   U410 : AOI22_X1 port map( A1 => n697, A2 => Q(398), B1 => n696, B2 => Q(270)
                           , ZN => n341);
   U411 : NAND4_X1 port map( A1 => n344, A2 => n343, A3 => n342, A4 => n341, ZN
                           => n350);
   U412 : AOI22_X1 port map( A1 => n699, A2 => Q(334), B1 => n698, B2 => Q(430)
                           , ZN => n348);
   U413 : AOI22_X1 port map( A1 => n701, A2 => Q(238), B1 => n700, B2 => Q(142)
                           , ZN => n347);
   U414 : AOI22_X1 port map( A1 => n703, A2 => Q(78), B1 => n702, B2 => Q(174),
                           ZN => n346);
   U415 : AOI22_X1 port map( A1 => n705, A2 => Q(206), B1 => n704, B2 => Q(46),
                           ZN => n345);
   U416 : NAND4_X1 port map( A1 => n348, A2 => n347, A3 => n346, A4 => n345, ZN
                           => n349);
   U417 : AOI22_X1 port map( A1 => n674, A2 => Q(1007), B1 => n673, B2 => 
                           Q(943), ZN => n356);
   U418 : AOI22_X1 port map( A1 => n676, A2 => Q(975), B1 => n675, B2 => Q(911)
                           , ZN => n355);
   U419 : AOI22_X1 port map( A1 => n678, A2 => Q(815), B1 => n677, B2 => Q(751)
                           , ZN => n354);
   U420 : NAND2_X1 port map( A1 => n679, A2 => Q(111), ZN => n353);
   U421 : NAND4_X1 port map( A1 => n356, A2 => n355, A3 => n354, A4 => n353, ZN
                           => n372);
   U422 : AOI22_X1 port map( A1 => n681, A2 => Q(847), B1 => n680, B2 => Q(719)
                           , ZN => n360);
   U423 : AOI22_X1 port map( A1 => n683, A2 => Q(783), B1 => n682, B2 => Q(879)
                           , ZN => n359);
   U424 : AOI22_X1 port map( A1 => n685, A2 => Q(687), B1 => n684, B2 => Q(591)
                           , ZN => n358);
   U425 : AOI22_X1 port map( A1 => n687, A2 => Q(527), B1 => n686, B2 => Q(623)
                           , ZN => n357);
   U426 : NAND4_X1 port map( A1 => n360, A2 => n359, A3 => n358, A4 => n357, ZN
                           => n371);
   U427 : AOI22_X1 port map( A1 => n691, A2 => Q(495), B1 => n690, B2 => Q(559)
                           , ZN => n364);
   U428 : AOI22_X1 port map( A1 => n693, A2 => Q(655), B1 => n692, B2 => Q(463)
                           , ZN => n363);
   U429 : AOI22_X1 port map( A1 => n695, A2 => Q(367), B1 => n694, B2 => Q(303)
                           , ZN => n362);
   U430 : AOI22_X1 port map( A1 => n697, A2 => Q(399), B1 => n696, B2 => Q(271)
                           , ZN => n361);
   U431 : NAND4_X1 port map( A1 => n364, A2 => n363, A3 => n362, A4 => n361, ZN
                           => n370);
   U432 : AOI22_X1 port map( A1 => n699, A2 => Q(335), B1 => n698, B2 => Q(431)
                           , ZN => n368);
   U433 : AOI22_X1 port map( A1 => n701, A2 => Q(239), B1 => n700, B2 => Q(143)
                           , ZN => n367);
   U434 : AOI22_X1 port map( A1 => n703, A2 => Q(79), B1 => n702, B2 => Q(175),
                           ZN => n366);
   U435 : AOI22_X1 port map( A1 => n705, A2 => Q(207), B1 => n704, B2 => Q(47),
                           ZN => n365);
   U436 : NAND4_X1 port map( A1 => n368, A2 => n367, A3 => n366, A4 => n365, ZN
                           => n369);
   U437 : AOI22_X1 port map( A1 => n674, A2 => Q(1008), B1 => n673, B2 => 
                           Q(944), ZN => n376);
   U438 : AOI22_X1 port map( A1 => n676, A2 => Q(976), B1 => n675, B2 => Q(912)
                           , ZN => n375);
   U439 : AOI22_X1 port map( A1 => n678, A2 => Q(816), B1 => n677, B2 => Q(752)
                           , ZN => n374);
   U440 : NAND2_X1 port map( A1 => n679, A2 => Q(112), ZN => n373);
   U441 : NAND4_X1 port map( A1 => n376, A2 => n375, A3 => n374, A4 => n373, ZN
                           => n392);
   U442 : AOI22_X1 port map( A1 => n681, A2 => Q(848), B1 => n680, B2 => Q(720)
                           , ZN => n380);
   U443 : AOI22_X1 port map( A1 => n683, A2 => Q(784), B1 => n682, B2 => Q(880)
                           , ZN => n379);
   U444 : AOI22_X1 port map( A1 => n685, A2 => Q(688), B1 => n684, B2 => Q(592)
                           , ZN => n378);
   U445 : AOI22_X1 port map( A1 => n687, A2 => Q(528), B1 => n686, B2 => Q(624)
                           , ZN => n377);
   U446 : NAND4_X1 port map( A1 => n380, A2 => n379, A3 => n378, A4 => n377, ZN
                           => n391);
   U447 : AOI22_X1 port map( A1 => n691, A2 => Q(496), B1 => n690, B2 => Q(560)
                           , ZN => n384);
   U448 : AOI22_X1 port map( A1 => n693, A2 => Q(656), B1 => n692, B2 => Q(464)
                           , ZN => n383);
   U449 : AOI22_X1 port map( A1 => n695, A2 => Q(368), B1 => n694, B2 => Q(304)
                           , ZN => n382);
   U450 : AOI22_X1 port map( A1 => n697, A2 => Q(400), B1 => n696, B2 => Q(272)
                           , ZN => n381);
   U451 : NAND4_X1 port map( A1 => n384, A2 => n383, A3 => n382, A4 => n381, ZN
                           => n390);
   U452 : AOI22_X1 port map( A1 => n699, A2 => Q(336), B1 => n698, B2 => Q(432)
                           , ZN => n388);
   U453 : AOI22_X1 port map( A1 => n701, A2 => Q(240), B1 => n700, B2 => Q(144)
                           , ZN => n387);
   U454 : AOI22_X1 port map( A1 => n703, A2 => Q(80), B1 => n702, B2 => Q(176),
                           ZN => n386);
   U455 : AOI22_X1 port map( A1 => n705, A2 => Q(208), B1 => n704, B2 => Q(48),
                           ZN => n385);
   U456 : NAND4_X1 port map( A1 => n388, A2 => n387, A3 => n386, A4 => n385, ZN
                           => n389);
   U457 : AOI22_X1 port map( A1 => n674, A2 => Q(1009), B1 => n673, B2 => 
                           Q(945), ZN => n396);
   U458 : AOI22_X1 port map( A1 => n676, A2 => Q(977), B1 => n675, B2 => Q(913)
                           , ZN => n395);
   U459 : AOI22_X1 port map( A1 => n678, A2 => Q(817), B1 => n677, B2 => Q(753)
                           , ZN => n394);
   U460 : NAND2_X1 port map( A1 => n679, A2 => Q(113), ZN => n393);
   U461 : NAND4_X1 port map( A1 => n396, A2 => n395, A3 => n394, A4 => n393, ZN
                           => n412);
   U462 : AOI22_X1 port map( A1 => n681, A2 => Q(849), B1 => n680, B2 => Q(721)
                           , ZN => n400);
   U463 : AOI22_X1 port map( A1 => n683, A2 => Q(785), B1 => n682, B2 => Q(881)
                           , ZN => n399);
   U464 : AOI22_X1 port map( A1 => n685, A2 => Q(689), B1 => n684, B2 => Q(593)
                           , ZN => n398);
   U465 : AOI22_X1 port map( A1 => n687, A2 => Q(529), B1 => n686, B2 => Q(625)
                           , ZN => n397);
   U466 : NAND4_X1 port map( A1 => n400, A2 => n399, A3 => n398, A4 => n397, ZN
                           => n411);
   U467 : AOI22_X1 port map( A1 => n691, A2 => Q(497), B1 => n690, B2 => Q(561)
                           , ZN => n404);
   U468 : AOI22_X1 port map( A1 => n693, A2 => Q(657), B1 => n692, B2 => Q(465)
                           , ZN => n403);
   U469 : AOI22_X1 port map( A1 => n695, A2 => Q(369), B1 => n694, B2 => Q(305)
                           , ZN => n402);
   U470 : AOI22_X1 port map( A1 => n697, A2 => Q(401), B1 => n696, B2 => Q(273)
                           , ZN => n401);
   U471 : NAND4_X1 port map( A1 => n404, A2 => n403, A3 => n402, A4 => n401, ZN
                           => n410);
   U472 : AOI22_X1 port map( A1 => n699, A2 => Q(337), B1 => n698, B2 => Q(433)
                           , ZN => n408);
   U473 : AOI22_X1 port map( A1 => n701, A2 => Q(241), B1 => n700, B2 => Q(145)
                           , ZN => n407);
   U474 : AOI22_X1 port map( A1 => n703, A2 => Q(81), B1 => n702, B2 => Q(177),
                           ZN => n406);
   U475 : AOI22_X1 port map( A1 => n705, A2 => Q(209), B1 => n704, B2 => Q(49),
                           ZN => n405);
   U476 : NAND4_X1 port map( A1 => n408, A2 => n407, A3 => n406, A4 => n405, ZN
                           => n409);
   U477 : AOI22_X1 port map( A1 => n674, A2 => Q(1010), B1 => n673, B2 => 
                           Q(946), ZN => n416);
   U478 : AOI22_X1 port map( A1 => n676, A2 => Q(978), B1 => n675, B2 => Q(914)
                           , ZN => n415);
   U479 : AOI22_X1 port map( A1 => n678, A2 => Q(818), B1 => n677, B2 => Q(754)
                           , ZN => n414);
   U480 : NAND2_X1 port map( A1 => n679, A2 => Q(114), ZN => n413);
   U481 : NAND4_X1 port map( A1 => n416, A2 => n415, A3 => n414, A4 => n413, ZN
                           => n432);
   U482 : AOI22_X1 port map( A1 => n681, A2 => Q(850), B1 => n680, B2 => Q(722)
                           , ZN => n420);
   U483 : AOI22_X1 port map( A1 => n683, A2 => Q(786), B1 => n682, B2 => Q(882)
                           , ZN => n419);
   U484 : AOI22_X1 port map( A1 => n685, A2 => Q(690), B1 => n684, B2 => Q(594)
                           , ZN => n418);
   U485 : AOI22_X1 port map( A1 => n687, A2 => Q(530), B1 => n686, B2 => Q(626)
                           , ZN => n417);
   U486 : NAND4_X1 port map( A1 => n420, A2 => n419, A3 => n418, A4 => n417, ZN
                           => n431);
   U487 : AOI22_X1 port map( A1 => n691, A2 => Q(498), B1 => n690, B2 => Q(562)
                           , ZN => n424);
   U488 : AOI22_X1 port map( A1 => n693, A2 => Q(658), B1 => n692, B2 => Q(466)
                           , ZN => n423);
   U489 : AOI22_X1 port map( A1 => n695, A2 => Q(370), B1 => n694, B2 => Q(306)
                           , ZN => n422);
   U490 : AOI22_X1 port map( A1 => n697, A2 => Q(402), B1 => n696, B2 => Q(274)
                           , ZN => n421);
   U491 : NAND4_X1 port map( A1 => n424, A2 => n423, A3 => n422, A4 => n421, ZN
                           => n430);
   U492 : AOI22_X1 port map( A1 => n699, A2 => Q(338), B1 => n698, B2 => Q(434)
                           , ZN => n428);
   U493 : AOI22_X1 port map( A1 => n701, A2 => Q(242), B1 => n700, B2 => Q(146)
                           , ZN => n427);
   U494 : AOI22_X1 port map( A1 => n703, A2 => Q(82), B1 => n702, B2 => Q(178),
                           ZN => n426);
   U495 : AOI22_X1 port map( A1 => n705, A2 => Q(210), B1 => n704, B2 => Q(50),
                           ZN => n425);
   U496 : NAND4_X1 port map( A1 => n428, A2 => n427, A3 => n426, A4 => n425, ZN
                           => n429);
   U497 : AOI22_X1 port map( A1 => n674, A2 => Q(1011), B1 => n673, B2 => 
                           Q(947), ZN => n436);
   U498 : AOI22_X1 port map( A1 => n676, A2 => Q(979), B1 => n675, B2 => Q(915)
                           , ZN => n435);
   U499 : AOI22_X1 port map( A1 => n678, A2 => Q(819), B1 => n677, B2 => Q(755)
                           , ZN => n434);
   U500 : NAND2_X1 port map( A1 => n679, A2 => Q(115), ZN => n433);
   U501 : NAND4_X1 port map( A1 => n436, A2 => n435, A3 => n434, A4 => n433, ZN
                           => n452);
   U502 : AOI22_X1 port map( A1 => n681, A2 => Q(851), B1 => n680, B2 => Q(723)
                           , ZN => n440);
   U503 : AOI22_X1 port map( A1 => n683, A2 => Q(787), B1 => n682, B2 => Q(883)
                           , ZN => n439);
   U504 : AOI22_X1 port map( A1 => n685, A2 => Q(691), B1 => n684, B2 => Q(595)
                           , ZN => n438);
   U505 : AOI22_X1 port map( A1 => n687, A2 => Q(531), B1 => n686, B2 => Q(627)
                           , ZN => n437);
   U506 : NAND4_X1 port map( A1 => n440, A2 => n439, A3 => n438, A4 => n437, ZN
                           => n451);
   U507 : AOI22_X1 port map( A1 => n691, A2 => Q(499), B1 => n690, B2 => Q(563)
                           , ZN => n444);
   U508 : AOI22_X1 port map( A1 => n693, A2 => Q(659), B1 => n692, B2 => Q(467)
                           , ZN => n443);
   U509 : AOI22_X1 port map( A1 => n695, A2 => Q(371), B1 => n694, B2 => Q(307)
                           , ZN => n442);
   U510 : AOI22_X1 port map( A1 => n697, A2 => Q(403), B1 => n696, B2 => Q(275)
                           , ZN => n441);
   U511 : NAND4_X1 port map( A1 => n444, A2 => n443, A3 => n442, A4 => n441, ZN
                           => n450);
   U512 : AOI22_X1 port map( A1 => n699, A2 => Q(339), B1 => n698, B2 => Q(435)
                           , ZN => n448);
   U513 : AOI22_X1 port map( A1 => n701, A2 => Q(243), B1 => n700, B2 => Q(147)
                           , ZN => n447);
   U514 : AOI22_X1 port map( A1 => n703, A2 => Q(83), B1 => n702, B2 => Q(179),
                           ZN => n446);
   U515 : AOI22_X1 port map( A1 => n705, A2 => Q(211), B1 => n704, B2 => Q(51),
                           ZN => n445);
   U516 : NAND4_X1 port map( A1 => n448, A2 => n447, A3 => n446, A4 => n445, ZN
                           => n449);
   U517 : AOI22_X1 port map( A1 => n674, A2 => Q(993), B1 => n673, B2 => Q(929)
                           , ZN => n456);
   U518 : AOI22_X1 port map( A1 => n676, A2 => Q(961), B1 => n675, B2 => Q(897)
                           , ZN => n455);
   U519 : AOI22_X1 port map( A1 => n678, A2 => Q(801), B1 => n677, B2 => Q(737)
                           , ZN => n454);
   U520 : NAND2_X1 port map( A1 => n679, A2 => Q(97), ZN => n453);
   U521 : NAND4_X1 port map( A1 => n456, A2 => n455, A3 => n454, A4 => n453, ZN
                           => n472);
   U522 : AOI22_X1 port map( A1 => n681, A2 => Q(833), B1 => n680, B2 => Q(705)
                           , ZN => n460);
   U523 : AOI22_X1 port map( A1 => n683, A2 => Q(769), B1 => n682, B2 => Q(865)
                           , ZN => n459);
   U524 : AOI22_X1 port map( A1 => n685, A2 => Q(673), B1 => n684, B2 => Q(577)
                           , ZN => n458);
   U525 : AOI22_X1 port map( A1 => n687, A2 => Q(513), B1 => n686, B2 => Q(609)
                           , ZN => n457);
   U526 : NAND4_X1 port map( A1 => n460, A2 => n459, A3 => n458, A4 => n457, ZN
                           => n471);
   U527 : AOI22_X1 port map( A1 => n691, A2 => Q(481), B1 => n690, B2 => Q(545)
                           , ZN => n464);
   U528 : AOI22_X1 port map( A1 => n693, A2 => Q(641), B1 => n692, B2 => Q(449)
                           , ZN => n463);
   U529 : AOI22_X1 port map( A1 => n695, A2 => Q(353), B1 => n694, B2 => Q(289)
                           , ZN => n462);
   U530 : AOI22_X1 port map( A1 => n697, A2 => Q(385), B1 => n696, B2 => Q(257)
                           , ZN => n461);
   U531 : NAND4_X1 port map( A1 => n464, A2 => n463, A3 => n462, A4 => n461, ZN
                           => n470);
   U532 : AOI22_X1 port map( A1 => n699, A2 => Q(321), B1 => n698, B2 => Q(417)
                           , ZN => n468);
   U533 : AOI22_X1 port map( A1 => n701, A2 => Q(225), B1 => n700, B2 => Q(129)
                           , ZN => n467);
   U534 : AOI22_X1 port map( A1 => n703, A2 => Q(65), B1 => n702, B2 => Q(161),
                           ZN => n466);
   U535 : AOI22_X1 port map( A1 => n705, A2 => Q(193), B1 => n704, B2 => Q(33),
                           ZN => n465);
   U536 : NAND4_X1 port map( A1 => n468, A2 => n467, A3 => n466, A4 => n465, ZN
                           => n469);
   U537 : AOI22_X1 port map( A1 => n251, A2 => Q(692), B1 => n250, B2 => Q(596)
                           , ZN => n474);
   U538 : AOI22_X1 port map( A1 => n253, A2 => Q(532), B1 => n252, B2 => Q(628)
                           , ZN => n473);
   U539 : AOI22_X1 port map( A1 => n240, A2 => Q(1013), B1 => n239, B2 => 
                           Q(949), ZN => n478);
   U540 : AOI22_X1 port map( A1 => n242, A2 => Q(981), B1 => n241, B2 => Q(917)
                           , ZN => n477);
   U541 : AOI22_X1 port map( A1 => n244, A2 => Q(821), B1 => n243, B2 => Q(757)
                           , ZN => n476);
   U542 : NAND2_X1 port map( A1 => n245, A2 => Q(117), ZN => n475);
   U543 : NAND4_X1 port map( A1 => n478, A2 => n477, A3 => n476, A4 => n475, ZN
                           => n494);
   U544 : AOI22_X1 port map( A1 => n247, A2 => Q(853), B1 => n246, B2 => Q(725)
                           , ZN => n482);
   U545 : AOI22_X1 port map( A1 => n249, A2 => Q(789), B1 => n248, B2 => Q(885)
                           , ZN => n481);
   U546 : AOI22_X1 port map( A1 => n251, A2 => Q(693), B1 => n250, B2 => Q(597)
                           , ZN => n480);
   U547 : AOI22_X1 port map( A1 => n253, A2 => Q(533), B1 => n252, B2 => Q(629)
                           , ZN => n479);
   U548 : NAND4_X1 port map( A1 => n482, A2 => n481, A3 => n480, A4 => n479, ZN
                           => n493);
   U549 : AOI22_X1 port map( A1 => n255, A2 => Q(501), B1 => n254, B2 => Q(565)
                           , ZN => n486);
   U550 : AOI22_X1 port map( A1 => n257, A2 => Q(661), B1 => n256, B2 => Q(469)
                           , ZN => n485);
   U551 : AOI22_X1 port map( A1 => n259, A2 => Q(373), B1 => n258, B2 => Q(309)
                           , ZN => n484);
   U552 : AOI22_X1 port map( A1 => n261, A2 => Q(405), B1 => n260, B2 => Q(277)
                           , ZN => n483);
   U553 : NAND4_X1 port map( A1 => n486, A2 => n485, A3 => n484, A4 => n483, ZN
                           => n492);
   U554 : AOI22_X1 port map( A1 => n263, A2 => Q(341), B1 => n262, B2 => Q(437)
                           , ZN => n490);
   U555 : AOI22_X1 port map( A1 => n265, A2 => Q(245), B1 => n264, B2 => Q(149)
                           , ZN => n489);
   U556 : AOI22_X1 port map( A1 => n267, A2 => Q(85), B1 => n266, B2 => Q(181),
                           ZN => n488);
   U557 : AOI22_X1 port map( A1 => n269, A2 => Q(213), B1 => n268, B2 => Q(53),
                           ZN => n487);
   U558 : NAND4_X1 port map( A1 => n490, A2 => n489, A3 => n488, A4 => n487, ZN
                           => n491);
   U559 : AOI22_X1 port map( A1 => n251, A2 => Q(694), B1 => n250, B2 => Q(598)
                           , ZN => n496);
   U560 : AOI22_X1 port map( A1 => n253, A2 => Q(534), B1 => n252, B2 => Q(630)
                           , ZN => n495);
   U561 : AOI22_X1 port map( A1 => n240, A2 => Q(1015), B1 => n239, B2 => 
                           Q(951), ZN => n500);
   U562 : AOI22_X1 port map( A1 => n242, A2 => Q(983), B1 => n241, B2 => Q(919)
                           , ZN => n499);
   U563 : AOI22_X1 port map( A1 => n244, A2 => Q(823), B1 => n243, B2 => Q(759)
                           , ZN => n498);
   U564 : NAND2_X1 port map( A1 => n245, A2 => Q(119), ZN => n497);
   U565 : NAND4_X1 port map( A1 => n500, A2 => n499, A3 => n498, A4 => n497, ZN
                           => n516);
   U566 : AOI22_X1 port map( A1 => n247, A2 => Q(855), B1 => n246, B2 => Q(727)
                           , ZN => n504);
   U567 : AOI22_X1 port map( A1 => n249, A2 => Q(791), B1 => n248, B2 => Q(887)
                           , ZN => n503);
   U568 : AOI22_X1 port map( A1 => n251, A2 => Q(695), B1 => n250, B2 => Q(599)
                           , ZN => n502);
   U569 : AOI22_X1 port map( A1 => n253, A2 => Q(535), B1 => n252, B2 => Q(631)
                           , ZN => n501);
   U570 : NAND4_X1 port map( A1 => n504, A2 => n503, A3 => n502, A4 => n501, ZN
                           => n515);
   U571 : AOI22_X1 port map( A1 => n255, A2 => Q(503), B1 => n254, B2 => Q(567)
                           , ZN => n508);
   U572 : AOI22_X1 port map( A1 => n257, A2 => Q(663), B1 => n256, B2 => Q(471)
                           , ZN => n507);
   U573 : AOI22_X1 port map( A1 => n259, A2 => Q(375), B1 => n258, B2 => Q(311)
                           , ZN => n506);
   U574 : AOI22_X1 port map( A1 => n261, A2 => Q(407), B1 => n260, B2 => Q(279)
                           , ZN => n505);
   U575 : NAND4_X1 port map( A1 => n508, A2 => n507, A3 => n506, A4 => n505, ZN
                           => n514);
   U576 : AOI22_X1 port map( A1 => n263, A2 => Q(343), B1 => n262, B2 => Q(439)
                           , ZN => n512);
   U577 : AOI22_X1 port map( A1 => n265, A2 => Q(247), B1 => n264, B2 => Q(151)
                           , ZN => n511);
   U578 : AOI22_X1 port map( A1 => n267, A2 => Q(87), B1 => n266, B2 => Q(183),
                           ZN => n510);
   U579 : AOI22_X1 port map( A1 => n269, A2 => Q(215), B1 => n268, B2 => Q(55),
                           ZN => n509);
   U580 : NAND4_X1 port map( A1 => n512, A2 => n511, A3 => n510, A4 => n509, ZN
                           => n513);
   U581 : AOI22_X1 port map( A1 => n240, A2 => Q(1016), B1 => n239, B2 => 
                           Q(952), ZN => n520);
   U582 : AOI22_X1 port map( A1 => n242, A2 => Q(984), B1 => n241, B2 => Q(920)
                           , ZN => n519);
   U583 : AOI22_X1 port map( A1 => n244, A2 => Q(824), B1 => n243, B2 => Q(760)
                           , ZN => n518);
   U584 : NAND2_X1 port map( A1 => n245, A2 => Q(120), ZN => n517);
   U585 : NAND4_X1 port map( A1 => n520, A2 => n519, A3 => n518, A4 => n517, ZN
                           => n536);
   U586 : AOI22_X1 port map( A1 => n247, A2 => Q(856), B1 => n246, B2 => Q(728)
                           , ZN => n524);
   U587 : AOI22_X1 port map( A1 => n249, A2 => Q(792), B1 => n248, B2 => Q(888)
                           , ZN => n523);
   U588 : AOI22_X1 port map( A1 => n251, A2 => Q(696), B1 => n250, B2 => Q(600)
                           , ZN => n522);
   U589 : AOI22_X1 port map( A1 => n253, A2 => Q(536), B1 => n252, B2 => Q(632)
                           , ZN => n521);
   U590 : NAND4_X1 port map( A1 => n524, A2 => n523, A3 => n522, A4 => n521, ZN
                           => n535);
   U591 : AOI22_X1 port map( A1 => n255, A2 => Q(504), B1 => n254, B2 => Q(568)
                           , ZN => n528);
   U592 : AOI22_X1 port map( A1 => n257, A2 => Q(664), B1 => n256, B2 => Q(472)
                           , ZN => n527);
   U593 : AOI22_X1 port map( A1 => n259, A2 => Q(376), B1 => n258, B2 => Q(312)
                           , ZN => n526);
   U594 : AOI22_X1 port map( A1 => n261, A2 => Q(408), B1 => n260, B2 => Q(280)
                           , ZN => n525);
   U595 : NAND4_X1 port map( A1 => n528, A2 => n527, A3 => n526, A4 => n525, ZN
                           => n534);
   U596 : AOI22_X1 port map( A1 => n263, A2 => Q(344), B1 => n262, B2 => Q(440)
                           , ZN => n532);
   U597 : AOI22_X1 port map( A1 => n265, A2 => Q(248), B1 => n264, B2 => Q(152)
                           , ZN => n531);
   U598 : AOI22_X1 port map( A1 => n267, A2 => Q(88), B1 => n266, B2 => Q(184),
                           ZN => n530);
   U599 : AOI22_X1 port map( A1 => n269, A2 => Q(216), B1 => n268, B2 => Q(56),
                           ZN => n529);
   U600 : NAND4_X1 port map( A1 => n532, A2 => n531, A3 => n530, A4 => n529, ZN
                           => n533);
   U601 : AOI22_X1 port map( A1 => n240, A2 => Q(1017), B1 => n239, B2 => 
                           Q(953), ZN => n540);
   U602 : AOI22_X1 port map( A1 => n242, A2 => Q(985), B1 => n241, B2 => Q(921)
                           , ZN => n539);
   U603 : AOI22_X1 port map( A1 => n244, A2 => Q(825), B1 => n243, B2 => Q(761)
                           , ZN => n538);
   U604 : NAND2_X1 port map( A1 => n245, A2 => Q(121), ZN => n537);
   U605 : NAND4_X1 port map( A1 => n540, A2 => n539, A3 => n538, A4 => n537, ZN
                           => n556);
   U606 : AOI22_X1 port map( A1 => n247, A2 => Q(857), B1 => n246, B2 => Q(729)
                           , ZN => n544);
   U607 : AOI22_X1 port map( A1 => n249, A2 => Q(793), B1 => n248, B2 => Q(889)
                           , ZN => n543);
   U608 : AOI22_X1 port map( A1 => n251, A2 => Q(697), B1 => n250, B2 => Q(601)
                           , ZN => n542);
   U609 : AOI22_X1 port map( A1 => n253, A2 => Q(537), B1 => n252, B2 => Q(633)
                           , ZN => n541);
   U610 : NAND4_X1 port map( A1 => n544, A2 => n543, A3 => n542, A4 => n541, ZN
                           => n555);
   U611 : AOI22_X1 port map( A1 => n255, A2 => Q(505), B1 => n254, B2 => Q(569)
                           , ZN => n548);
   U612 : AOI22_X1 port map( A1 => n257, A2 => Q(665), B1 => n256, B2 => Q(473)
                           , ZN => n547);
   U613 : AOI22_X1 port map( A1 => n259, A2 => Q(377), B1 => n258, B2 => Q(313)
                           , ZN => n546);
   U614 : AOI22_X1 port map( A1 => n261, A2 => Q(409), B1 => n260, B2 => Q(281)
                           , ZN => n545);
   U615 : NAND4_X1 port map( A1 => n548, A2 => n547, A3 => n546, A4 => n545, ZN
                           => n554);
   U616 : AOI22_X1 port map( A1 => n263, A2 => Q(345), B1 => n262, B2 => Q(441)
                           , ZN => n552);
   U617 : AOI22_X1 port map( A1 => n265, A2 => Q(249), B1 => n264, B2 => Q(153)
                           , ZN => n551);
   U618 : AOI22_X1 port map( A1 => n267, A2 => Q(89), B1 => n266, B2 => Q(185),
                           ZN => n550);
   U619 : AOI22_X1 port map( A1 => n269, A2 => Q(217), B1 => n268, B2 => Q(57),
                           ZN => n549);
   U620 : NAND4_X1 port map( A1 => n552, A2 => n551, A3 => n550, A4 => n549, ZN
                           => n553);
   U621 : AOI22_X1 port map( A1 => n240, A2 => Q(1018), B1 => n239, B2 => 
                           Q(954), ZN => n560);
   U622 : AOI22_X1 port map( A1 => n242, A2 => Q(986), B1 => n241, B2 => Q(922)
                           , ZN => n559);
   U623 : AOI22_X1 port map( A1 => n244, A2 => Q(826), B1 => n243, B2 => Q(762)
                           , ZN => n558);
   U624 : NAND2_X1 port map( A1 => n245, A2 => Q(122), ZN => n557);
   U625 : NAND4_X1 port map( A1 => n560, A2 => n559, A3 => n558, A4 => n557, ZN
                           => n576);
   U626 : AOI22_X1 port map( A1 => n247, A2 => Q(858), B1 => n246, B2 => Q(730)
                           , ZN => n564);
   U627 : AOI22_X1 port map( A1 => n249, A2 => Q(794), B1 => n248, B2 => Q(890)
                           , ZN => n563);
   U628 : AOI22_X1 port map( A1 => n251, A2 => Q(698), B1 => n250, B2 => Q(602)
                           , ZN => n562);
   U629 : AOI22_X1 port map( A1 => n253, A2 => Q(538), B1 => n252, B2 => Q(634)
                           , ZN => n561);
   U630 : NAND4_X1 port map( A1 => n564, A2 => n563, A3 => n562, A4 => n561, ZN
                           => n575);
   U631 : AOI22_X1 port map( A1 => n255, A2 => Q(506), B1 => n254, B2 => Q(570)
                           , ZN => n568);
   U632 : AOI22_X1 port map( A1 => n257, A2 => Q(666), B1 => n256, B2 => Q(474)
                           , ZN => n567);
   U633 : AOI22_X1 port map( A1 => n259, A2 => Q(378), B1 => n258, B2 => Q(314)
                           , ZN => n566);
   U634 : AOI22_X1 port map( A1 => n261, A2 => Q(410), B1 => n260, B2 => Q(282)
                           , ZN => n565);
   U635 : NAND4_X1 port map( A1 => n568, A2 => n567, A3 => n566, A4 => n565, ZN
                           => n574);
   U636 : AOI22_X1 port map( A1 => n263, A2 => Q(346), B1 => n262, B2 => Q(442)
                           , ZN => n572);
   U637 : AOI22_X1 port map( A1 => n265, A2 => Q(250), B1 => n264, B2 => Q(154)
                           , ZN => n571);
   U638 : AOI22_X1 port map( A1 => n267, A2 => Q(90), B1 => n266, B2 => Q(186),
                           ZN => n570);
   U639 : AOI22_X1 port map( A1 => n269, A2 => Q(218), B1 => n268, B2 => Q(58),
                           ZN => n569);
   U640 : NAND4_X1 port map( A1 => n572, A2 => n571, A3 => n570, A4 => n569, ZN
                           => n573);
   U641 : AOI22_X1 port map( A1 => n240, A2 => Q(1019), B1 => n239, B2 => 
                           Q(955), ZN => n580);
   U642 : AOI22_X1 port map( A1 => n242, A2 => Q(987), B1 => n241, B2 => Q(923)
                           , ZN => n579);
   U643 : AOI22_X1 port map( A1 => n244, A2 => Q(827), B1 => n243, B2 => Q(763)
                           , ZN => n578);
   U644 : NAND2_X1 port map( A1 => n245, A2 => Q(123), ZN => n577);
   U645 : NAND4_X1 port map( A1 => n580, A2 => n579, A3 => n578, A4 => n577, ZN
                           => n596);
   U646 : AOI22_X1 port map( A1 => n247, A2 => Q(859), B1 => n246, B2 => Q(731)
                           , ZN => n584);
   U647 : AOI22_X1 port map( A1 => n249, A2 => Q(795), B1 => n248, B2 => Q(891)
                           , ZN => n583);
   U648 : AOI22_X1 port map( A1 => n251, A2 => Q(699), B1 => n250, B2 => Q(603)
                           , ZN => n582);
   U649 : AOI22_X1 port map( A1 => n253, A2 => Q(539), B1 => n252, B2 => Q(635)
                           , ZN => n581);
   U650 : NAND4_X1 port map( A1 => n584, A2 => n583, A3 => n582, A4 => n581, ZN
                           => n595);
   U651 : AOI22_X1 port map( A1 => n255, A2 => Q(507), B1 => n254, B2 => Q(571)
                           , ZN => n588);
   U652 : AOI22_X1 port map( A1 => n257, A2 => Q(667), B1 => n256, B2 => Q(475)
                           , ZN => n587);
   U653 : AOI22_X1 port map( A1 => n259, A2 => Q(379), B1 => n258, B2 => Q(315)
                           , ZN => n586);
   U654 : AOI22_X1 port map( A1 => n261, A2 => Q(411), B1 => n260, B2 => Q(283)
                           , ZN => n585);
   U655 : NAND4_X1 port map( A1 => n588, A2 => n587, A3 => n586, A4 => n585, ZN
                           => n594);
   U656 : AOI22_X1 port map( A1 => n263, A2 => Q(347), B1 => n262, B2 => Q(443)
                           , ZN => n592);
   U657 : AOI22_X1 port map( A1 => n265, A2 => Q(251), B1 => n264, B2 => Q(155)
                           , ZN => n591);
   U658 : AOI22_X1 port map( A1 => n267, A2 => Q(91), B1 => n266, B2 => Q(187),
                           ZN => n590);
   U659 : AOI22_X1 port map( A1 => n269, A2 => Q(219), B1 => n268, B2 => Q(59),
                           ZN => n589);
   U660 : NAND4_X1 port map( A1 => n592, A2 => n591, A3 => n590, A4 => n589, ZN
                           => n593);
   U661 : AOI22_X1 port map( A1 => n240, A2 => Q(1020), B1 => n673, B2 => 
                           Q(956), ZN => n600);
   U662 : AOI22_X1 port map( A1 => n242, A2 => Q(988), B1 => n675, B2 => Q(924)
                           , ZN => n599);
   U663 : AOI22_X1 port map( A1 => n244, A2 => Q(828), B1 => n677, B2 => Q(764)
                           , ZN => n598);
   U664 : NAND2_X1 port map( A1 => n245, A2 => Q(124), ZN => n597);
   U665 : NAND4_X1 port map( A1 => n600, A2 => n599, A3 => n598, A4 => n597, ZN
                           => n616);
   U666 : AOI22_X1 port map( A1 => n247, A2 => Q(860), B1 => n680, B2 => Q(732)
                           , ZN => n604);
   U667 : AOI22_X1 port map( A1 => n249, A2 => Q(796), B1 => n682, B2 => Q(892)
                           , ZN => n603);
   U668 : AOI22_X1 port map( A1 => n251, A2 => Q(700), B1 => n684, B2 => Q(604)
                           , ZN => n602);
   U669 : AOI22_X1 port map( A1 => n253, A2 => Q(540), B1 => n686, B2 => Q(636)
                           , ZN => n601);
   U670 : NAND4_X1 port map( A1 => n604, A2 => n603, A3 => n602, A4 => n601, ZN
                           => n615);
   U671 : AOI22_X1 port map( A1 => n255, A2 => Q(508), B1 => n690, B2 => Q(572)
                           , ZN => n608);
   U672 : AOI22_X1 port map( A1 => n257, A2 => Q(668), B1 => n692, B2 => Q(476)
                           , ZN => n607);
   U673 : AOI22_X1 port map( A1 => n259, A2 => Q(380), B1 => n694, B2 => Q(316)
                           , ZN => n606);
   U674 : AOI22_X1 port map( A1 => n261, A2 => Q(412), B1 => n696, B2 => Q(284)
                           , ZN => n605);
   U675 : NAND4_X1 port map( A1 => n608, A2 => n607, A3 => n606, A4 => n605, ZN
                           => n614);
   U676 : AOI22_X1 port map( A1 => n263, A2 => Q(348), B1 => n698, B2 => Q(444)
                           , ZN => n612);
   U677 : AOI22_X1 port map( A1 => n265, A2 => Q(252), B1 => n700, B2 => Q(156)
                           , ZN => n611);
   U678 : AOI22_X1 port map( A1 => n267, A2 => Q(92), B1 => n702, B2 => Q(188),
                           ZN => n610);
   U679 : AOI22_X1 port map( A1 => n269, A2 => Q(220), B1 => n704, B2 => Q(60),
                           ZN => n609);
   U680 : NAND4_X1 port map( A1 => n612, A2 => n611, A3 => n610, A4 => n609, ZN
                           => n613);
   U681 : AOI22_X1 port map( A1 => n240, A2 => Q(1021), B1 => n239, B2 => 
                           Q(957), ZN => n620);
   U682 : AOI22_X1 port map( A1 => n242, A2 => Q(989), B1 => n241, B2 => Q(925)
                           , ZN => n619);
   U683 : AOI22_X1 port map( A1 => n244, A2 => Q(829), B1 => n243, B2 => Q(765)
                           , ZN => n618);
   U684 : NAND2_X1 port map( A1 => n245, A2 => Q(125), ZN => n617);
   U685 : NAND4_X1 port map( A1 => n620, A2 => n619, A3 => n618, A4 => n617, ZN
                           => n636);
   U686 : AOI22_X1 port map( A1 => n247, A2 => Q(861), B1 => n246, B2 => Q(733)
                           , ZN => n624);
   U687 : AOI22_X1 port map( A1 => n249, A2 => Q(797), B1 => n248, B2 => Q(893)
                           , ZN => n623);
   U688 : AOI22_X1 port map( A1 => n251, A2 => Q(701), B1 => n250, B2 => Q(605)
                           , ZN => n622);
   U689 : AOI22_X1 port map( A1 => n253, A2 => Q(541), B1 => n252, B2 => Q(637)
                           , ZN => n621);
   U690 : NAND4_X1 port map( A1 => n624, A2 => n623, A3 => n622, A4 => n621, ZN
                           => n635);
   U691 : AOI22_X1 port map( A1 => n255, A2 => Q(509), B1 => n254, B2 => Q(573)
                           , ZN => n628);
   U692 : AOI22_X1 port map( A1 => n257, A2 => Q(669), B1 => n256, B2 => Q(477)
                           , ZN => n627);
   U693 : AOI22_X1 port map( A1 => n259, A2 => Q(381), B1 => n258, B2 => Q(317)
                           , ZN => n626);
   U694 : AOI22_X1 port map( A1 => n261, A2 => Q(413), B1 => n260, B2 => Q(285)
                           , ZN => n625);
   U695 : NAND4_X1 port map( A1 => n628, A2 => n627, A3 => n626, A4 => n625, ZN
                           => n634);
   U696 : AOI22_X1 port map( A1 => n263, A2 => Q(349), B1 => n262, B2 => Q(445)
                           , ZN => n632);
   U697 : AOI22_X1 port map( A1 => n265, A2 => Q(253), B1 => n264, B2 => Q(157)
                           , ZN => n631);
   U698 : AOI22_X1 port map( A1 => n267, A2 => Q(93), B1 => n266, B2 => Q(189),
                           ZN => n630);
   U699 : AOI22_X1 port map( A1 => n269, A2 => Q(221), B1 => n268, B2 => Q(61),
                           ZN => n629);
   U700 : NAND4_X1 port map( A1 => n632, A2 => n631, A3 => n630, A4 => n629, ZN
                           => n633);
   U701 : AOI22_X1 port map( A1 => n685, A2 => Q(674), B1 => n684, B2 => Q(578)
                           , ZN => n638);
   U702 : AOI22_X1 port map( A1 => n687, A2 => Q(514), B1 => n686, B2 => Q(610)
                           , ZN => n637);
   U703 : AOI22_X1 port map( A1 => n674, A2 => Q(1022), B1 => n673, B2 => 
                           Q(958), ZN => n642);
   U704 : AOI22_X1 port map( A1 => n676, A2 => Q(990), B1 => n675, B2 => Q(926)
                           , ZN => n641);
   U705 : AOI22_X1 port map( A1 => n678, A2 => Q(830), B1 => n677, B2 => Q(766)
                           , ZN => n640);
   U706 : NAND2_X1 port map( A1 => n679, A2 => Q(126), ZN => n639);
   U707 : NAND4_X1 port map( A1 => n642, A2 => n641, A3 => n640, A4 => n639, ZN
                           => n658);
   U708 : AOI22_X1 port map( A1 => n681, A2 => Q(862), B1 => n680, B2 => Q(734)
                           , ZN => n646);
   U709 : AOI22_X1 port map( A1 => n683, A2 => Q(798), B1 => n682, B2 => Q(894)
                           , ZN => n645);
   U710 : AOI22_X1 port map( A1 => n685, A2 => Q(702), B1 => n684, B2 => Q(606)
                           , ZN => n644);
   U711 : AOI22_X1 port map( A1 => n687, A2 => Q(542), B1 => n686, B2 => Q(638)
                           , ZN => n643);
   U712 : NAND4_X1 port map( A1 => n646, A2 => n645, A3 => n644, A4 => n643, ZN
                           => n657);
   U713 : AOI22_X1 port map( A1 => n691, A2 => Q(510), B1 => n690, B2 => Q(574)
                           , ZN => n650);
   U714 : AOI22_X1 port map( A1 => n693, A2 => Q(670), B1 => n692, B2 => Q(478)
                           , ZN => n649);
   U715 : AOI22_X1 port map( A1 => n695, A2 => Q(382), B1 => n694, B2 => Q(318)
                           , ZN => n648);
   U716 : AOI22_X1 port map( A1 => n697, A2 => Q(414), B1 => n696, B2 => Q(286)
                           , ZN => n647);
   U717 : NAND4_X1 port map( A1 => n650, A2 => n649, A3 => n648, A4 => n647, ZN
                           => n656);
   U718 : AOI22_X1 port map( A1 => n699, A2 => Q(350), B1 => n698, B2 => Q(446)
                           , ZN => n654);
   U719 : AOI22_X1 port map( A1 => n701, A2 => Q(254), B1 => n700, B2 => Q(158)
                           , ZN => n653);
   U720 : AOI22_X1 port map( A1 => n703, A2 => Q(94), B1 => n702, B2 => Q(190),
                           ZN => n652);
   U721 : AOI22_X1 port map( A1 => n705, A2 => Q(222), B1 => n704, B2 => Q(62),
                           ZN => n651);
   U722 : NAND4_X1 port map( A1 => n654, A2 => n653, A3 => n652, A4 => n651, ZN
                           => n655);
   U723 : AOI22_X1 port map( A1 => n251, A2 => Q(703), B1 => n250, B2 => Q(607)
                           , ZN => n660);
   U724 : AOI22_X1 port map( A1 => n253, A2 => Q(543), B1 => n252, B2 => Q(639)
                           , ZN => n659);
   U725 : AOI22_X1 port map( A1 => n251, A2 => Q(675), B1 => n250, B2 => Q(579)
                           , ZN => n662);
   U726 : AOI22_X1 port map( A1 => n253, A2 => Q(515), B1 => n252, B2 => Q(611)
                           , ZN => n661);
   U727 : AOI22_X1 port map( A1 => n251, A2 => Q(676), B1 => n250, B2 => Q(580)
                           , ZN => n664);
   U728 : AOI22_X1 port map( A1 => n253, A2 => Q(516), B1 => n252, B2 => Q(612)
                           , ZN => n663);
   U729 : AOI22_X1 port map( A1 => n251, A2 => Q(677), B1 => n250, B2 => Q(581)
                           , ZN => n666);
   U730 : AOI22_X1 port map( A1 => n253, A2 => Q(517), B1 => n252, B2 => Q(613)
                           , ZN => n665);
   U731 : AOI22_X1 port map( A1 => n251, A2 => Q(678), B1 => n250, B2 => Q(582)
                           , ZN => n668);
   U732 : AOI22_X1 port map( A1 => n253, A2 => Q(518), B1 => n252, B2 => Q(614)
                           , ZN => n667);
   U733 : AOI22_X1 port map( A1 => n251, A2 => Q(679), B1 => n250, B2 => Q(583)
                           , ZN => n670);
   U734 : AOI22_X1 port map( A1 => n253, A2 => Q(519), B1 => n252, B2 => Q(615)
                           , ZN => n669);
   U735 : AOI22_X1 port map( A1 => n251, A2 => Q(680), B1 => n250, B2 => Q(584)
                           , ZN => n672);
   U736 : AOI22_X1 port map( A1 => n253, A2 => Q(520), B1 => n252, B2 => Q(616)
                           , ZN => n671);
   U737 : AOI22_X1 port map( A1 => n251, A2 => Q(681), B1 => n250, B2 => Q(585)
                           , ZN => n689);
   U738 : AOI22_X1 port map( A1 => n253, A2 => Q(521), B1 => n252, B2 => Q(617)
                           , ZN => n688);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32.all;

entity select_block_NBIT_DATA32_N8_F5 is

   port( regs : in std_logic_vector (2559 downto 0);  win : in std_logic_vector
         (4 downto 0);  curr_proc_regs : out std_logic_vector (767 downto 0));

end select_block_NBIT_DATA32_N8_F5;

architecture SYN_behav of select_block_NBIT_DATA32_N8_F5 is

   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
      n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, 
      n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, 
      n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
      n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
      n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, 
      n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
      n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
      n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
      n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
      n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, 
      n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, 
      n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
      n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
      n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
      n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
      n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
      n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
      n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
      n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
      n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
      n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
      n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
      n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
      n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
      n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
      n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
      n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
      n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
      n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, 
      n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, 
      n2213, n2214, n2215 : std_logic;

begin
   
   U2 : CLKBUF_X3 port map( A => n2211, Z => n5);
   U3 : BUF_X1 port map( A => n2128, Z => n16);
   U4 : INV_X1 port map( A => n16, ZN => n2);
   U5 : BUF_X1 port map( A => n2215, Z => n6);
   U6 : INV_X2 port map( A => n58, ZN => n1);
   U7 : BUF_X1 port map( A => n2128, Z => n12);
   U8 : INV_X2 port map( A => n57, ZN => n3);
   U9 : BUF_X4 port map( A => n74, Z => n73);
   U10 : INV_X2 port map( A => n15, ZN => n4);
   U11 : BUF_X1 port map( A => n78, Z => n11);
   U12 : CLKBUF_X3 port map( A => n2211, Z => n74);
   U13 : BUF_X2 port map( A => n2211, Z => n69);
   U14 : BUF_X1 port map( A => n2215, Z => n13);
   U15 : INV_X2 port map( A => n132, ZN => n7);
   U16 : INV_X2 port map( A => n9, ZN => n8);
   U17 : BUF_X2 port map( A => n58, Z => n9);
   U18 : BUF_X2 port map( A => n5, Z => n71);
   U19 : BUF_X2 port map( A => n5, Z => n66);
   U20 : BUF_X2 port map( A => n57, Z => n10);
   U21 : BUF_X2 port map( A => n2201, Z => n40);
   U22 : BUF_X2 port map( A => n2128, Z => n15);
   U23 : BUF_X2 port map( A => n2215, Z => n77);
   U24 : NAND2_X2 port map( A1 => n135, A2 => win(1), ZN => n2201);
   U25 : INV_X2 port map( A => win(4), ZN => n132);
   U26 : BUF_X1 port map( A => n78, Z => n103);
   U27 : INV_X1 port map( A => n77, ZN => n92);
   U28 : INV_X1 port map( A => n77, ZN => n91);
   U29 : BUF_X1 port map( A => n10, Z => n58);
   U30 : BUF_X1 port map( A => n2215, Z => n78);
   U31 : BUF_X1 port map( A => n2201, Z => n57);
   U32 : INV_X1 port map( A => n132, ZN => n104);
   U33 : INV_X1 port map( A => n132, ZN => n131);
   U34 : BUF_X2 port map( A => n2211, Z => n68);
   U35 : BUF_X2 port map( A => n66, Z => n72);
   U36 : BUF_X2 port map( A => n2211, Z => n63);
   U37 : BUF_X1 port map( A => n68, Z => n67);
   U38 : BUF_X1 port map( A => n73, Z => n64);
   U39 : BUF_X1 port map( A => n71, Z => n60);
   U40 : BUF_X1 port map( A => n73, Z => n65);
   U41 : BUF_X1 port map( A => n72, Z => n70);
   U42 : BUF_X1 port map( A => n2211, Z => n62);
   U43 : BUF_X1 port map( A => n2211, Z => n61);
   U44 : BUF_X1 port map( A => n73, Z => n76);
   U45 : BUF_X1 port map( A => n66, Z => n75);
   U46 : BUF_X1 port map( A => n2201, Z => n59);
   U47 : INV_X1 port map( A => n132, ZN => n105);
   U48 : BUF_X1 port map( A => n2128, Z => n14);
   U49 : INV_X1 port map( A => n16, ZN => n17);
   U50 : INV_X1 port map( A => n16, ZN => n18);
   U51 : INV_X1 port map( A => n16, ZN => n19);
   U52 : INV_X1 port map( A => n16, ZN => n20);
   U53 : INV_X1 port map( A => n16, ZN => n21);
   U54 : INV_X1 port map( A => n16, ZN => n22);
   U55 : INV_X1 port map( A => n16, ZN => n23);
   U56 : INV_X1 port map( A => n16, ZN => n24);
   U57 : INV_X1 port map( A => n16, ZN => n25);
   U58 : INV_X1 port map( A => n16, ZN => n26);
   U59 : INV_X1 port map( A => n16, ZN => n27);
   U60 : INV_X1 port map( A => n15, ZN => n28);
   U61 : INV_X1 port map( A => n15, ZN => n29);
   U62 : INV_X1 port map( A => n15, ZN => n30);
   U63 : INV_X1 port map( A => n15, ZN => n31);
   U64 : INV_X1 port map( A => n15, ZN => n32);
   U65 : INV_X1 port map( A => n15, ZN => n33);
   U66 : INV_X1 port map( A => n15, ZN => n34);
   U67 : INV_X1 port map( A => n15, ZN => n35);
   U68 : INV_X1 port map( A => n15, ZN => n36);
   U69 : INV_X1 port map( A => n15, ZN => n37);
   U70 : INV_X1 port map( A => n15, ZN => n38);
   U71 : INV_X1 port map( A => n15, ZN => n39);
   U72 : INV_X1 port map( A => n2201, ZN => n41);
   U73 : INV_X1 port map( A => n2201, ZN => n42);
   U74 : INV_X1 port map( A => n57, ZN => n43);
   U75 : INV_X1 port map( A => n57, ZN => n44);
   U76 : INV_X1 port map( A => n57, ZN => n45);
   U77 : INV_X1 port map( A => n10, ZN => n46);
   U78 : INV_X1 port map( A => n10, ZN => n47);
   U79 : INV_X1 port map( A => n10, ZN => n48);
   U80 : INV_X1 port map( A => n10, ZN => n49);
   U81 : INV_X1 port map( A => n10, ZN => n50);
   U82 : INV_X1 port map( A => n10, ZN => n51);
   U83 : INV_X1 port map( A => n10, ZN => n52);
   U84 : INV_X1 port map( A => n57, ZN => n53);
   U85 : INV_X1 port map( A => n57, ZN => n54);
   U86 : INV_X1 port map( A => n10, ZN => n55);
   U87 : INV_X1 port map( A => n57, ZN => n56);
   U88 : INV_X1 port map( A => n77, ZN => n79);
   U89 : INV_X1 port map( A => n77, ZN => n80);
   U90 : INV_X1 port map( A => n77, ZN => n81);
   U91 : INV_X1 port map( A => n77, ZN => n82);
   U92 : INV_X1 port map( A => n77, ZN => n83);
   U93 : INV_X1 port map( A => n77, ZN => n84);
   U94 : INV_X1 port map( A => n77, ZN => n85);
   U95 : INV_X1 port map( A => n77, ZN => n86);
   U96 : INV_X1 port map( A => n77, ZN => n87);
   U97 : INV_X1 port map( A => n77, ZN => n88);
   U98 : INV_X1 port map( A => n77, ZN => n89);
   U99 : INV_X1 port map( A => n77, ZN => n90);
   U100 : INV_X1 port map( A => n77, ZN => n93);
   U101 : INV_X1 port map( A => n77, ZN => n94);
   U102 : INV_X1 port map( A => n77, ZN => n95);
   U103 : INV_X1 port map( A => n77, ZN => n96);
   U104 : INV_X1 port map( A => n77, ZN => n97);
   U105 : INV_X1 port map( A => n77, ZN => n98);
   U106 : INV_X1 port map( A => n77, ZN => n99);
   U107 : INV_X1 port map( A => n77, ZN => n100);
   U108 : INV_X1 port map( A => n77, ZN => n101);
   U109 : INV_X1 port map( A => n77, ZN => n102);
   U110 : INV_X1 port map( A => n132, ZN => n106);
   U111 : INV_X1 port map( A => n132, ZN => n107);
   U112 : INV_X1 port map( A => n132, ZN => n108);
   U113 : INV_X1 port map( A => n132, ZN => n109);
   U114 : INV_X1 port map( A => n132, ZN => n110);
   U115 : INV_X1 port map( A => n132, ZN => n111);
   U116 : INV_X1 port map( A => n132, ZN => n112);
   U117 : INV_X1 port map( A => n132, ZN => n113);
   U118 : INV_X1 port map( A => n132, ZN => n114);
   U119 : INV_X1 port map( A => n132, ZN => n115);
   U120 : INV_X1 port map( A => n132, ZN => n116);
   U121 : INV_X1 port map( A => n132, ZN => n117);
   U122 : INV_X1 port map( A => n132, ZN => n118);
   U123 : INV_X1 port map( A => n132, ZN => n119);
   U124 : INV_X1 port map( A => n132, ZN => n120);
   U125 : INV_X1 port map( A => n132, ZN => n121);
   U126 : INV_X1 port map( A => n132, ZN => n122);
   U127 : INV_X1 port map( A => n132, ZN => n123);
   U128 : INV_X1 port map( A => n132, ZN => n124);
   U129 : INV_X1 port map( A => n132, ZN => n125);
   U130 : INV_X1 port map( A => n132, ZN => n126);
   U131 : INV_X1 port map( A => n132, ZN => n127);
   U132 : INV_X1 port map( A => n132, ZN => n128);
   U133 : INV_X1 port map( A => n132, ZN => n129);
   U134 : INV_X1 port map( A => n132, ZN => n130);
   U135 : NOR3_X1 port map( A1 => win(3), A2 => n131, A3 => win(2), ZN => n135)
                           ;
   U136 : INV_X1 port map( A => regs(512), ZN => n1310);
   U137 : INV_X1 port map( A => win(3), ZN => n133);
   U138 : NOR2_X1 port map( A1 => n104, A2 => n133, ZN => n2211);
   U139 : AOI22_X1 port map( A1 => n125, A2 => regs(2048), B1 => n60, B2 => 
                           regs(1536), ZN => n137);
   U140 : NAND3_X1 port map( A1 => n133, A2 => n132, A3 => win(2), ZN => n2215)
                           ;
   U141 : INV_X1 port map( A => win(1), ZN => n134);
   U142 : NAND3_X1 port map( A1 => n135, A2 => win(0), A3 => n134, ZN => n2128)
                           ;
   U143 : AOI22_X1 port map( A1 => n79, A2 => regs(1024), B1 => n21, B2 => 
                           regs(0), ZN => n136);
   U144 : OAI211_X1 port map( C1 => n57, C2 => n1310, A => n137, B => n136, ZN 
                           => curr_proc_regs(0));
   U145 : INV_X1 port map( A => regs(1124), ZN => n1617);
   U146 : AOI22_X1 port map( A1 => n125, A2 => regs(2148), B1 => n60, B2 => 
                           regs(1636), ZN => n139);
   U147 : AOI22_X1 port map( A1 => n42, A2 => regs(612), B1 => n21, B2 => 
                           regs(100), ZN => n138);
   U148 : OAI211_X1 port map( C1 => n2215, C2 => n1617, A => n139, B => n138, 
                           ZN => curr_proc_regs(100));
   U149 : INV_X1 port map( A => regs(613), ZN => n1620);
   U150 : AOI22_X1 port map( A1 => n124, A2 => regs(2149), B1 => n60, B2 => 
                           regs(1637), ZN => n141);
   U151 : AOI22_X1 port map( A1 => n96, A2 => regs(1125), B1 => n21, B2 => 
                           regs(101), ZN => n140);
   U152 : OAI211_X1 port map( C1 => n10, C2 => n1620, A => n141, B => n140, ZN 
                           => curr_proc_regs(101));
   U153 : INV_X1 port map( A => regs(614), ZN => n1623);
   U154 : AOI22_X1 port map( A1 => n113, A2 => regs(2150), B1 => n60, B2 => 
                           regs(1638), ZN => n143);
   U155 : AOI22_X1 port map( A1 => n89, A2 => regs(1126), B1 => n21, B2 => 
                           regs(102), ZN => n142);
   U156 : OAI211_X1 port map( C1 => n9, C2 => n1623, A => n143, B => n142, ZN 
                           => curr_proc_regs(102));
   U157 : INV_X1 port map( A => regs(615), ZN => n1626);
   U158 : AOI22_X1 port map( A1 => n114, A2 => regs(2151), B1 => n60, B2 => 
                           regs(1639), ZN => n145);
   U159 : AOI22_X1 port map( A1 => n88, A2 => regs(1127), B1 => n35, B2 => 
                           regs(103), ZN => n144);
   U160 : OAI211_X1 port map( C1 => n2201, C2 => n1626, A => n145, B => n144, 
                           ZN => curr_proc_regs(103));
   U161 : INV_X1 port map( A => regs(616), ZN => n1629);
   U162 : AOI22_X1 port map( A1 => n125, A2 => regs(2152), B1 => n60, B2 => 
                           regs(1640), ZN => n147);
   U163 : AOI22_X1 port map( A1 => n89, A2 => regs(1128), B1 => n39, B2 => 
                           regs(104), ZN => n146);
   U164 : OAI211_X1 port map( C1 => n10, C2 => n1629, A => n147, B => n146, ZN 
                           => curr_proc_regs(104));
   U165 : INV_X1 port map( A => regs(617), ZN => n1632);
   U166 : AOI22_X1 port map( A1 => n124, A2 => regs(2153), B1 => n60, B2 => 
                           regs(1641), ZN => n149);
   U167 : AOI22_X1 port map( A1 => n89, A2 => regs(1129), B1 => n38, B2 => 
                           regs(105), ZN => n148);
   U168 : OAI211_X1 port map( C1 => n10, C2 => n1632, A => n149, B => n148, ZN 
                           => curr_proc_regs(105));
   U169 : INV_X1 port map( A => regs(618), ZN => n1635);
   U170 : AOI22_X1 port map( A1 => n112, A2 => regs(2154), B1 => n60, B2 => 
                           regs(1642), ZN => n151);
   U171 : AOI22_X1 port map( A1 => n88, A2 => regs(1130), B1 => n37, B2 => 
                           regs(106), ZN => n150);
   U172 : OAI211_X1 port map( C1 => n10, C2 => n1635, A => n151, B => n150, ZN 
                           => curr_proc_regs(106));
   U173 : INV_X1 port map( A => regs(1131), ZN => n1638);
   U174 : AOI22_X1 port map( A1 => n117, A2 => regs(2155), B1 => n60, B2 => 
                           regs(1643), ZN => n153);
   U175 : AOI22_X1 port map( A1 => n49, A2 => regs(619), B1 => n36, B2 => 
                           regs(107), ZN => n152);
   U176 : OAI211_X1 port map( C1 => n77, C2 => n1638, A => n153, B => n152, ZN 
                           => curr_proc_regs(107));
   U177 : INV_X1 port map( A => regs(620), ZN => n1644);
   U178 : AOI22_X1 port map( A1 => n125, A2 => regs(2156), B1 => n60, B2 => 
                           regs(1644), ZN => n155);
   U179 : AOI22_X1 port map( A1 => n89, A2 => regs(1132), B1 => n34, B2 => 
                           regs(108), ZN => n154);
   U180 : OAI211_X1 port map( C1 => n9, C2 => n1644, A => n155, B => n154, ZN 
                           => curr_proc_regs(108));
   U181 : INV_X1 port map( A => regs(1133), ZN => n1647);
   U182 : AOI22_X1 port map( A1 => n124, A2 => regs(2157), B1 => n60, B2 => 
                           regs(1645), ZN => n157);
   U183 : AOI22_X1 port map( A1 => n42, A2 => regs(621), B1 => n33, B2 => 
                           regs(109), ZN => n156);
   U184 : OAI211_X1 port map( C1 => n77, C2 => n1647, A => n157, B => n156, ZN 
                           => curr_proc_regs(109));
   U185 : INV_X1 port map( A => regs(522), ZN => n1339);
   U186 : AOI22_X1 port map( A1 => n109, A2 => regs(2058), B1 => n60, B2 => 
                           regs(1546), ZN => n159);
   U187 : AOI22_X1 port map( A1 => n89, A2 => regs(1034), B1 => n31, B2 => 
                           regs(10), ZN => n158);
   U188 : OAI211_X1 port map( C1 => n10, C2 => n1339, A => n159, B => n158, ZN 
                           => curr_proc_regs(10));
   U189 : INV_X1 port map( A => regs(622), ZN => n1650);
   U190 : AOI22_X1 port map( A1 => n120, A2 => regs(2158), B1 => n68, B2 => 
                           regs(1646), ZN => n161);
   U191 : AOI22_X1 port map( A1 => n88, A2 => regs(1134), B1 => n22, B2 => 
                           regs(110), ZN => n160);
   U192 : OAI211_X1 port map( C1 => n10, C2 => n1650, A => n161, B => n160, ZN 
                           => curr_proc_regs(110));
   U193 : INV_X1 port map( A => regs(623), ZN => n1653);
   U194 : AOI22_X1 port map( A1 => n124, A2 => regs(2159), B1 => n68, B2 => 
                           regs(1647), ZN => n163);
   U195 : AOI22_X1 port map( A1 => n88, A2 => regs(1135), B1 => n22, B2 => 
                           regs(111), ZN => n162);
   U196 : OAI211_X1 port map( C1 => n9, C2 => n1653, A => n163, B => n162, ZN 
                           => curr_proc_regs(111));
   U197 : INV_X1 port map( A => regs(624), ZN => n1656);
   U198 : AOI22_X1 port map( A1 => n115, A2 => regs(2160), B1 => n68, B2 => 
                           regs(1648), ZN => n165);
   U199 : AOI22_X1 port map( A1 => n95, A2 => regs(1136), B1 => n22, B2 => 
                           regs(112), ZN => n164);
   U200 : OAI211_X1 port map( C1 => n10, C2 => n1656, A => n165, B => n164, ZN 
                           => curr_proc_regs(112));
   U201 : INV_X1 port map( A => regs(625), ZN => n1659);
   U202 : AOI22_X1 port map( A1 => n104, A2 => regs(2161), B1 => n72, B2 => 
                           regs(1649), ZN => n167);
   U203 : AOI22_X1 port map( A1 => n88, A2 => regs(1137), B1 => n22, B2 => 
                           regs(113), ZN => n166);
   U204 : OAI211_X1 port map( C1 => n9, C2 => n1659, A => n167, B => n166, ZN 
                           => curr_proc_regs(113));
   U205 : INV_X1 port map( A => regs(626), ZN => n1662);
   U206 : AOI22_X1 port map( A1 => n125, A2 => regs(2162), B1 => n70, B2 => 
                           regs(1650), ZN => n169);
   U207 : AOI22_X1 port map( A1 => n88, A2 => regs(1138), B1 => n21, B2 => 
                           regs(114), ZN => n168);
   U208 : OAI211_X1 port map( C1 => n9, C2 => n1662, A => n169, B => n168, ZN 
                           => curr_proc_regs(114));
   U209 : INV_X1 port map( A => regs(627), ZN => n1665);
   U210 : AOI22_X1 port map( A1 => n128, A2 => regs(2163), B1 => n74, B2 => 
                           regs(1651), ZN => n171);
   U211 : AOI22_X1 port map( A1 => n88, A2 => regs(1139), B1 => n21, B2 => 
                           regs(115), ZN => n170);
   U212 : OAI211_X1 port map( C1 => n9, C2 => n1665, A => n171, B => n170, ZN 
                           => curr_proc_regs(115));
   U213 : INV_X1 port map( A => regs(628), ZN => n1668);
   U214 : AOI22_X1 port map( A1 => n113, A2 => regs(2164), B1 => n65, B2 => 
                           regs(1652), ZN => n173);
   U215 : AOI22_X1 port map( A1 => n88, A2 => regs(1140), B1 => n21, B2 => 
                           regs(116), ZN => n172);
   U216 : OAI211_X1 port map( C1 => n9, C2 => n1668, A => n173, B => n172, ZN 
                           => curr_proc_regs(116));
   U217 : INV_X1 port map( A => regs(629), ZN => n1671);
   U218 : AOI22_X1 port map( A1 => n112, A2 => regs(2165), B1 => n69, B2 => 
                           regs(1653), ZN => n175);
   U219 : AOI22_X1 port map( A1 => n88, A2 => regs(1141), B1 => n21, B2 => 
                           regs(117), ZN => n174);
   U220 : OAI211_X1 port map( C1 => n9, C2 => n1671, A => n175, B => n174, ZN 
                           => curr_proc_regs(117));
   U221 : INV_X1 port map( A => regs(630), ZN => n1677);
   U222 : AOI22_X1 port map( A1 => n109, A2 => regs(2166), B1 => n67, B2 => 
                           regs(1654), ZN => n177);
   U223 : AOI22_X1 port map( A1 => n92, A2 => regs(1142), B1 => n21, B2 => 
                           regs(118), ZN => n176);
   U224 : OAI211_X1 port map( C1 => n9, C2 => n1677, A => n177, B => n176, ZN 
                           => curr_proc_regs(118));
   U225 : INV_X1 port map( A => regs(1143), ZN => n1680);
   U226 : AOI22_X1 port map( A1 => n115, A2 => regs(2167), B1 => n72, B2 => 
                           regs(1655), ZN => n179);
   U227 : AOI22_X1 port map( A1 => n42, A2 => regs(631), B1 => n21, B2 => 
                           regs(119), ZN => n178);
   U228 : OAI211_X1 port map( C1 => n2215, C2 => n1680, A => n179, B => n178, 
                           ZN => curr_proc_regs(119));
   U229 : INV_X1 port map( A => regs(523), ZN => n1342);
   U230 : AOI22_X1 port map( A1 => n114, A2 => regs(2059), B1 => n66, B2 => 
                           regs(1547), ZN => n181);
   U231 : AOI22_X1 port map( A1 => n98, A2 => regs(1035), B1 => n21, B2 => 
                           regs(11), ZN => n180);
   U232 : OAI211_X1 port map( C1 => n9, C2 => n1342, A => n181, B => n180, ZN 
                           => curr_proc_regs(11));
   U233 : INV_X1 port map( A => regs(1144), ZN => n1683);
   U234 : AOI22_X1 port map( A1 => n117, A2 => regs(2168), B1 => n66, B2 => 
                           regs(1656), ZN => n183);
   U235 : AOI22_X1 port map( A1 => n42, A2 => regs(632), B1 => n21, B2 => 
                           regs(120), ZN => n182);
   U236 : OAI211_X1 port map( C1 => n77, C2 => n1683, A => n183, B => n182, ZN 
                           => curr_proc_regs(120));
   U237 : INV_X1 port map( A => regs(633), ZN => n1686);
   U238 : AOI22_X1 port map( A1 => n120, A2 => regs(2169), B1 => n63, B2 => 
                           regs(1657), ZN => n185);
   U239 : AOI22_X1 port map( A1 => n94, A2 => regs(1145), B1 => n23, B2 => 
                           regs(121), ZN => n184);
   U240 : OAI211_X1 port map( C1 => n2201, C2 => n1686, A => n185, B => n184, 
                           ZN => curr_proc_regs(121));
   U241 : INV_X1 port map( A => regs(1146), ZN => n1689);
   U242 : AOI22_X1 port map( A1 => n114, A2 => regs(2170), B1 => n63, B2 => 
                           regs(1658), ZN => n187);
   U243 : AOI22_X1 port map( A1 => n42, A2 => regs(634), B1 => n23, B2 => 
                           regs(122), ZN => n186);
   U244 : OAI211_X1 port map( C1 => n77, C2 => n1689, A => n187, B => n186, ZN 
                           => curr_proc_regs(122));
   U245 : INV_X1 port map( A => regs(635), ZN => n1692);
   U246 : AOI22_X1 port map( A1 => n117, A2 => regs(2171), B1 => n63, B2 => 
                           regs(1659), ZN => n189);
   U247 : AOI22_X1 port map( A1 => n94, A2 => regs(1147), B1 => n23, B2 => 
                           regs(123), ZN => n188);
   U248 : OAI211_X1 port map( C1 => n2201, C2 => n1692, A => n189, B => n188, 
                           ZN => curr_proc_regs(123));
   U249 : INV_X1 port map( A => regs(1148), ZN => n1695);
   U250 : AOI22_X1 port map( A1 => n120, A2 => regs(2172), B1 => n63, B2 => 
                           regs(1660), ZN => n191);
   U251 : AOI22_X1 port map( A1 => n42, A2 => regs(636), B1 => n23, B2 => 
                           regs(124), ZN => n190);
   U252 : OAI211_X1 port map( C1 => n77, C2 => n1695, A => n191, B => n190, ZN 
                           => curr_proc_regs(124));
   U253 : INV_X1 port map( A => regs(1149), ZN => n1698);
   U254 : AOI22_X1 port map( A1 => n105, A2 => regs(2173), B1 => n63, B2 => 
                           regs(1661), ZN => n193);
   U255 : AOI22_X1 port map( A1 => n42, A2 => regs(637), B1 => n22, B2 => 
                           regs(125), ZN => n192);
   U256 : OAI211_X1 port map( C1 => n2215, C2 => n1698, A => n193, B => n192, 
                           ZN => curr_proc_regs(125));
   U257 : INV_X1 port map( A => regs(1150), ZN => n1701);
   U258 : AOI22_X1 port map( A1 => n122, A2 => regs(2174), B1 => n63, B2 => 
                           regs(1662), ZN => n195);
   U259 : AOI22_X1 port map( A1 => n42, A2 => regs(638), B1 => n22, B2 => 
                           regs(126), ZN => n194);
   U260 : OAI211_X1 port map( C1 => n77, C2 => n1701, A => n195, B => n194, ZN 
                           => curr_proc_regs(126));
   U261 : INV_X1 port map( A => regs(1151), ZN => n1704);
   U262 : AOI22_X1 port map( A1 => n124, A2 => regs(2175), B1 => n63, B2 => 
                           regs(1663), ZN => n197);
   U263 : AOI22_X1 port map( A1 => n42, A2 => regs(639), B1 => n22, B2 => 
                           regs(127), ZN => n196);
   U264 : OAI211_X1 port map( C1 => n77, C2 => n1704, A => n197, B => n196, ZN 
                           => curr_proc_regs(127));
   U265 : INV_X1 port map( A => regs(1152), ZN => n1710);
   U266 : AOI22_X1 port map( A1 => n104, A2 => regs(2176), B1 => n5, B2 => 
                           regs(1664), ZN => n199);
   U267 : AOI22_X1 port map( A1 => n42, A2 => regs(640), B1 => n22, B2 => 
                           regs(128), ZN => n198);
   U268 : OAI211_X1 port map( C1 => n77, C2 => n1710, A => n199, B => n198, ZN 
                           => curr_proc_regs(128));
   U269 : INV_X1 port map( A => regs(641), ZN => n1713);
   U270 : AOI22_X1 port map( A1 => n125, A2 => regs(2177), B1 => n63, B2 => 
                           regs(1665), ZN => n201);
   U271 : AOI22_X1 port map( A1 => n91, A2 => regs(1153), B1 => n22, B2 => 
                           regs(129), ZN => n200);
   U272 : OAI211_X1 port map( C1 => n2201, C2 => n1713, A => n201, B => n200, 
                           ZN => curr_proc_regs(129));
   U273 : INV_X1 port map( A => regs(524), ZN => n1345);
   U274 : AOI22_X1 port map( A1 => n128, A2 => regs(2060), B1 => n60, B2 => 
                           regs(1548), ZN => n203);
   U275 : AOI22_X1 port map( A1 => n88, A2 => regs(1036), B1 => n22, B2 => 
                           regs(12), ZN => n202);
   U276 : OAI211_X1 port map( C1 => n2201, C2 => n1345, A => n203, B => n202, 
                           ZN => curr_proc_regs(12));
   U277 : INV_X1 port map( A => regs(1154), ZN => n1716);
   U278 : AOI22_X1 port map( A1 => n113, A2 => regs(2178), B1 => n64, B2 => 
                           regs(1666), ZN => n205);
   U279 : AOI22_X1 port map( A1 => n42, A2 => regs(642), B1 => n22, B2 => 
                           regs(130), ZN => n204);
   U280 : OAI211_X1 port map( C1 => n77, C2 => n1716, A => n205, B => n204, ZN 
                           => curr_proc_regs(130));
   U281 : INV_X1 port map( A => regs(1155), ZN => n1719);
   U282 : AOI22_X1 port map( A1 => n112, A2 => regs(2179), B1 => n62, B2 => 
                           regs(1667), ZN => n207);
   U283 : AOI22_X1 port map( A1 => n44, A2 => regs(643), B1 => n22, B2 => 
                           regs(131), ZN => n206);
   U284 : OAI211_X1 port map( C1 => n77, C2 => n1719, A => n207, B => n206, ZN 
                           => curr_proc_regs(131));
   U285 : INV_X1 port map( A => regs(1156), ZN => n1722);
   U286 : AOI22_X1 port map( A1 => n109, A2 => regs(2180), B1 => n73, B2 => 
                           regs(1668), ZN => n209);
   U287 : AOI22_X1 port map( A1 => n44, A2 => regs(644), B1 => n24, B2 => 
                           regs(132), ZN => n208);
   U288 : OAI211_X1 port map( C1 => n77, C2 => n1722, A => n209, B => n208, ZN 
                           => curr_proc_regs(132));
   U289 : INV_X1 port map( A => regs(1157), ZN => n1725);
   U290 : AOI22_X1 port map( A1 => n124, A2 => regs(2181), B1 => n74, B2 => 
                           regs(1669), ZN => n211);
   U291 : AOI22_X1 port map( A1 => n49, A2 => regs(645), B1 => n24, B2 => 
                           regs(133), ZN => n210);
   U292 : OAI211_X1 port map( C1 => n77, C2 => n1725, A => n211, B => n210, ZN 
                           => curr_proc_regs(133));
   U293 : INV_X1 port map( A => regs(1158), ZN => n1728);
   U294 : AOI22_X1 port map( A1 => n124, A2 => regs(2182), B1 => n68, B2 => 
                           regs(1670), ZN => n213);
   U295 : AOI22_X1 port map( A1 => n41, A2 => regs(646), B1 => n24, B2 => 
                           regs(134), ZN => n212);
   U296 : OAI211_X1 port map( C1 => n77, C2 => n1728, A => n213, B => n212, ZN 
                           => curr_proc_regs(134));
   U297 : INV_X1 port map( A => regs(647), ZN => n1731);
   U298 : AOI22_X1 port map( A1 => n124, A2 => regs(2183), B1 => n72, B2 => 
                           regs(1671), ZN => n215);
   U299 : AOI22_X1 port map( A1 => n88, A2 => regs(1159), B1 => n24, B2 => 
                           regs(135), ZN => n214);
   U300 : OAI211_X1 port map( C1 => n9, C2 => n1731, A => n215, B => n214, ZN 
                           => curr_proc_regs(135));
   U301 : INV_X1 port map( A => regs(648), ZN => n1734);
   U302 : AOI22_X1 port map( A1 => n124, A2 => regs(2184), B1 => n72, B2 => 
                           regs(1672), ZN => n217);
   U303 : AOI22_X1 port map( A1 => n100, A2 => regs(1160), B1 => n23, B2 => 
                           regs(136), ZN => n216);
   U304 : OAI211_X1 port map( C1 => n58, C2 => n1734, A => n217, B => n216, ZN 
                           => curr_proc_regs(136));
   U305 : INV_X1 port map( A => regs(1161), ZN => n1737);
   U306 : AOI22_X1 port map( A1 => n124, A2 => regs(2185), B1 => n68, B2 => 
                           regs(1673), ZN => n219);
   U307 : AOI22_X1 port map( A1 => n41, A2 => regs(649), B1 => n23, B2 => 
                           regs(137), ZN => n218);
   U308 : OAI211_X1 port map( C1 => n77, C2 => n1737, A => n219, B => n218, ZN 
                           => curr_proc_regs(137));
   U309 : INV_X1 port map( A => regs(650), ZN => n1743);
   U310 : AOI22_X1 port map( A1 => n124, A2 => regs(2186), B1 => n70, B2 => 
                           regs(1674), ZN => n221);
   U311 : AOI22_X1 port map( A1 => n88, A2 => regs(1162), B1 => n23, B2 => 
                           regs(138), ZN => n220);
   U312 : OAI211_X1 port map( C1 => n2201, C2 => n1743, A => n221, B => n220, 
                           ZN => curr_proc_regs(138));
   U313 : INV_X1 port map( A => regs(1163), ZN => n1746);
   U314 : AOI22_X1 port map( A1 => n124, A2 => regs(2187), B1 => n74, B2 => 
                           regs(1675), ZN => n223);
   U315 : AOI22_X1 port map( A1 => n41, A2 => regs(651), B1 => n23, B2 => 
                           regs(139), ZN => n222);
   U316 : OAI211_X1 port map( C1 => n77, C2 => n1746, A => n223, B => n222, ZN 
                           => curr_proc_regs(139));
   U317 : INV_X1 port map( A => regs(525), ZN => n1348);
   U318 : AOI22_X1 port map( A1 => n124, A2 => regs(2061), B1 => n65, B2 => 
                           regs(1549), ZN => n225);
   U319 : AOI22_X1 port map( A1 => n100, A2 => regs(1037), B1 => n23, B2 => 
                           regs(13), ZN => n224);
   U320 : OAI211_X1 port map( C1 => n9, C2 => n1348, A => n225, B => n224, ZN 
                           => curr_proc_regs(13));
   U321 : INV_X1 port map( A => regs(652), ZN => n1749);
   U322 : AOI22_X1 port map( A1 => n124, A2 => regs(2188), B1 => n69, B2 => 
                           regs(1676), ZN => n227);
   U323 : AOI22_X1 port map( A1 => n98, A2 => regs(1164), B1 => n23, B2 => 
                           regs(140), ZN => n226);
   U324 : OAI211_X1 port map( C1 => n57, C2 => n1749, A => n227, B => n226, ZN 
                           => curr_proc_regs(140));
   U325 : INV_X1 port map( A => regs(1165), ZN => n1752);
   U326 : AOI22_X1 port map( A1 => n124, A2 => regs(2189), B1 => n5, B2 => 
                           regs(1677), ZN => n229);
   U327 : AOI22_X1 port map( A1 => n41, A2 => regs(653), B1 => n23, B2 => 
                           regs(141), ZN => n228);
   U328 : OAI211_X1 port map( C1 => n77, C2 => n1752, A => n229, B => n228, ZN 
                           => curr_proc_regs(141));
   U329 : INV_X1 port map( A => regs(654), ZN => n1755);
   U330 : AOI22_X1 port map( A1 => n124, A2 => regs(2190), B1 => n67, B2 => 
                           regs(1678), ZN => n231);
   U331 : AOI22_X1 port map( A1 => n96, A2 => regs(1166), B1 => n23, B2 => 
                           regs(142), ZN => n230);
   U332 : OAI211_X1 port map( C1 => n10, C2 => n1755, A => n231, B => n230, ZN 
                           => curr_proc_regs(142));
   U333 : INV_X1 port map( A => regs(1167), ZN => n1758);
   U334 : AOI22_X1 port map( A1 => n124, A2 => regs(2191), B1 => n61, B2 => 
                           regs(1679), ZN => n233);
   U335 : AOI22_X1 port map( A1 => n41, A2 => regs(655), B1 => n4, B2 => 
                           regs(143), ZN => n232);
   U336 : OAI211_X1 port map( C1 => n13, C2 => n1758, A => n233, B => n232, ZN 
                           => curr_proc_regs(143));
   U337 : INV_X1 port map( A => regs(1168), ZN => n1761);
   U338 : AOI22_X1 port map( A1 => n105, A2 => regs(2192), B1 => n61, B2 => 
                           regs(1680), ZN => n235);
   U339 : AOI22_X1 port map( A1 => n41, A2 => regs(656), B1 => n4, B2 => 
                           regs(144), ZN => n234);
   U340 : OAI211_X1 port map( C1 => n13, C2 => n1761, A => n235, B => n234, ZN 
                           => curr_proc_regs(144));
   U341 : INV_X1 port map( A => regs(657), ZN => n1764);
   U342 : AOI22_X1 port map( A1 => n7, A2 => regs(2193), B1 => n61, B2 => 
                           regs(1681), ZN => n237);
   U343 : AOI22_X1 port map( A1 => n92, A2 => regs(1169), B1 => n4, B2 => 
                           regs(145), ZN => n236);
   U344 : OAI211_X1 port map( C1 => n9, C2 => n1764, A => n237, B => n236, ZN 
                           => curr_proc_regs(145));
   U345 : INV_X1 port map( A => regs(1170), ZN => n1767);
   U346 : AOI22_X1 port map( A1 => n122, A2 => regs(2194), B1 => n61, B2 => 
                           regs(1682), ZN => n239);
   U347 : AOI22_X1 port map( A1 => n41, A2 => regs(658), B1 => n4, B2 => 
                           regs(146), ZN => n238);
   U348 : OAI211_X1 port map( C1 => n13, C2 => n1767, A => n239, B => n238, ZN 
                           => curr_proc_regs(146));
   U349 : INV_X1 port map( A => regs(1171), ZN => n1770);
   U350 : AOI22_X1 port map( A1 => n123, A2 => regs(2195), B1 => n61, B2 => 
                           regs(1683), ZN => n241);
   U351 : AOI22_X1 port map( A1 => n41, A2 => regs(659), B1 => n24, B2 => 
                           regs(147), ZN => n240);
   U352 : OAI211_X1 port map( C1 => n13, C2 => n1770, A => n241, B => n240, ZN 
                           => curr_proc_regs(147));
   U353 : INV_X1 port map( A => regs(660), ZN => n1776);
   U354 : AOI22_X1 port map( A1 => n105, A2 => regs(2196), B1 => n61, B2 => 
                           regs(1684), ZN => n243);
   U355 : AOI22_X1 port map( A1 => n94, A2 => regs(1172), B1 => n24, B2 => 
                           regs(148), ZN => n242);
   U356 : OAI211_X1 port map( C1 => n57, C2 => n1776, A => n243, B => n242, ZN 
                           => curr_proc_regs(148));
   U357 : INV_X1 port map( A => regs(1173), ZN => n1779);
   U358 : AOI22_X1 port map( A1 => n123, A2 => regs(2197), B1 => n61, B2 => 
                           regs(1685), ZN => n245);
   U359 : AOI22_X1 port map( A1 => n41, A2 => regs(661), B1 => n24, B2 => 
                           regs(149), ZN => n244);
   U360 : OAI211_X1 port map( C1 => n13, C2 => n1779, A => n245, B => n244, ZN 
                           => curr_proc_regs(149));
   U361 : INV_X1 port map( A => regs(1038), ZN => n1351);
   U362 : AOI22_X1 port map( A1 => n7, A2 => regs(2062), B1 => n61, B2 => 
                           regs(1550), ZN => n247);
   U363 : AOI22_X1 port map( A1 => n53, A2 => regs(526), B1 => n24, B2 => 
                           regs(14), ZN => n246);
   U364 : OAI211_X1 port map( C1 => n13, C2 => n1351, A => n247, B => n246, ZN 
                           => curr_proc_regs(14));
   U365 : INV_X1 port map( A => regs(1174), ZN => n1782);
   U366 : AOI22_X1 port map( A1 => n104, A2 => regs(2198), B1 => n61, B2 => 
                           regs(1686), ZN => n249);
   U367 : AOI22_X1 port map( A1 => n53, A2 => regs(662), B1 => n24, B2 => 
                           regs(150), ZN => n248);
   U368 : OAI211_X1 port map( C1 => n13, C2 => n1782, A => n249, B => n248, ZN 
                           => curr_proc_regs(150));
   U369 : INV_X1 port map( A => regs(1175), ZN => n1785);
   U370 : AOI22_X1 port map( A1 => n105, A2 => regs(2199), B1 => n61, B2 => 
                           regs(1687), ZN => n251);
   U371 : AOI22_X1 port map( A1 => n53, A2 => regs(663), B1 => n24, B2 => 
                           regs(151), ZN => n250);
   U372 : OAI211_X1 port map( C1 => n13, C2 => n1785, A => n251, B => n250, ZN 
                           => curr_proc_regs(151));
   U373 : INV_X1 port map( A => regs(664), ZN => n1788);
   U374 : AOI22_X1 port map( A1 => n7, A2 => regs(2200), B1 => n61, B2 => 
                           regs(1688), ZN => n253);
   U375 : AOI22_X1 port map( A1 => n94, A2 => regs(1176), B1 => n24, B2 => 
                           regs(152), ZN => n252);
   U376 : OAI211_X1 port map( C1 => n10, C2 => n1788, A => n253, B => n252, ZN 
                           => curr_proc_regs(152));
   U377 : INV_X1 port map( A => regs(665), ZN => n1791);
   U378 : AOI22_X1 port map( A1 => n122, A2 => regs(2201), B1 => n61, B2 => 
                           regs(1689), ZN => n255);
   U379 : AOI22_X1 port map( A1 => n89, A2 => regs(1177), B1 => n24, B2 => 
                           regs(153), ZN => n254);
   U380 : OAI211_X1 port map( C1 => n10, C2 => n1791, A => n255, B => n254, ZN 
                           => curr_proc_regs(153));
   U381 : INV_X1 port map( A => regs(666), ZN => n1794);
   U382 : AOI22_X1 port map( A1 => n123, A2 => regs(2202), B1 => n62, B2 => 
                           regs(1690), ZN => n257);
   U383 : AOI22_X1 port map( A1 => n95, A2 => regs(1178), B1 => n25, B2 => 
                           regs(154), ZN => n256);
   U384 : OAI211_X1 port map( C1 => n58, C2 => n1794, A => n257, B => n256, ZN 
                           => curr_proc_regs(154));
   U385 : INV_X1 port map( A => regs(667), ZN => n1797);
   U386 : AOI22_X1 port map( A1 => n122, A2 => regs(2203), B1 => n62, B2 => 
                           regs(1691), ZN => n259);
   U387 : AOI22_X1 port map( A1 => n98, A2 => regs(1179), B1 => n25, B2 => 
                           regs(155), ZN => n258);
   U388 : OAI211_X1 port map( C1 => n57, C2 => n1797, A => n259, B => n258, ZN 
                           => curr_proc_regs(155));
   U389 : INV_X1 port map( A => regs(668), ZN => n1800);
   U390 : AOI22_X1 port map( A1 => n104, A2 => regs(2204), B1 => n62, B2 => 
                           regs(1692), ZN => n261);
   U391 : AOI22_X1 port map( A1 => n89, A2 => regs(1180), B1 => n25, B2 => 
                           regs(156), ZN => n260);
   U392 : OAI211_X1 port map( C1 => n59, C2 => n1800, A => n261, B => n260, ZN 
                           => curr_proc_regs(156));
   U393 : INV_X1 port map( A => regs(669), ZN => n1803);
   U394 : AOI22_X1 port map( A1 => n105, A2 => regs(2205), B1 => n62, B2 => 
                           regs(1693), ZN => n263);
   U395 : AOI22_X1 port map( A1 => n100, A2 => regs(1181), B1 => n25, B2 => 
                           regs(157), ZN => n262);
   U396 : OAI211_X1 port map( C1 => n59, C2 => n1803, A => n263, B => n262, ZN 
                           => curr_proc_regs(157));
   U397 : INV_X1 port map( A => regs(1182), ZN => n1809);
   U398 : AOI22_X1 port map( A1 => n7, A2 => regs(2206), B1 => n62, B2 => 
                           regs(1694), ZN => n265);
   U399 : AOI22_X1 port map( A1 => n53, A2 => regs(670), B1 => n4, B2 => 
                           regs(158), ZN => n264);
   U400 : OAI211_X1 port map( C1 => n13, C2 => n1809, A => n265, B => n264, ZN 
                           => curr_proc_regs(158));
   U401 : INV_X1 port map( A => regs(1183), ZN => n1812);
   U402 : AOI22_X1 port map( A1 => n122, A2 => regs(2207), B1 => n62, B2 => 
                           regs(1695), ZN => n267);
   U403 : AOI22_X1 port map( A1 => n53, A2 => regs(671), B1 => n4, B2 => 
                           regs(159), ZN => n266);
   U404 : OAI211_X1 port map( C1 => n13, C2 => n1812, A => n267, B => n266, ZN 
                           => curr_proc_regs(159));
   U405 : INV_X1 port map( A => regs(1039), ZN => n1354);
   U406 : AOI22_X1 port map( A1 => n123, A2 => regs(2063), B1 => n62, B2 => 
                           regs(1551), ZN => n269);
   U407 : AOI22_X1 port map( A1 => n41, A2 => regs(527), B1 => n4, B2 => 
                           regs(15), ZN => n268);
   U408 : OAI211_X1 port map( C1 => n13, C2 => n1354, A => n269, B => n268, ZN 
                           => curr_proc_regs(15));
   U409 : INV_X1 port map( A => regs(1184), ZN => n1815);
   U410 : AOI22_X1 port map( A1 => n123, A2 => regs(2208), B1 => n62, B2 => 
                           regs(1696), ZN => n271);
   U411 : AOI22_X1 port map( A1 => n42, A2 => regs(672), B1 => n4, B2 => 
                           regs(160), ZN => n270);
   U412 : OAI211_X1 port map( C1 => n13, C2 => n1815, A => n271, B => n270, ZN 
                           => curr_proc_regs(160));
   U413 : INV_X1 port map( A => regs(673), ZN => n1818);
   U414 : AOI22_X1 port map( A1 => n104, A2 => regs(2209), B1 => n62, B2 => 
                           regs(1697), ZN => n273);
   U415 : AOI22_X1 port map( A1 => n98, A2 => regs(1185), B1 => n4, B2 => 
                           regs(161), ZN => n272);
   U416 : OAI211_X1 port map( C1 => n58, C2 => n1818, A => n273, B => n272, ZN 
                           => curr_proc_regs(161));
   U417 : INV_X1 port map( A => regs(1186), ZN => n1821);
   U418 : AOI22_X1 port map( A1 => n104, A2 => regs(2210), B1 => n62, B2 => 
                           regs(1698), ZN => n275);
   U419 : AOI22_X1 port map( A1 => n53, A2 => regs(674), B1 => n4, B2 => 
                           regs(162), ZN => n274);
   U420 : OAI211_X1 port map( C1 => n13, C2 => n1821, A => n275, B => n274, ZN 
                           => curr_proc_regs(162));
   U421 : INV_X1 port map( A => regs(1187), ZN => n1824);
   U422 : AOI22_X1 port map( A1 => n105, A2 => regs(2211), B1 => n62, B2 => 
                           regs(1699), ZN => n277);
   U423 : AOI22_X1 port map( A1 => n54, A2 => regs(675), B1 => n4, B2 => 
                           regs(163), ZN => n276);
   U424 : OAI211_X1 port map( C1 => n13, C2 => n1824, A => n277, B => n276, ZN 
                           => curr_proc_regs(163));
   U425 : INV_X1 port map( A => regs(676), ZN => n1827);
   U426 : AOI22_X1 port map( A1 => n7, A2 => regs(2212), B1 => n62, B2 => 
                           regs(1700), ZN => n279);
   U427 : AOI22_X1 port map( A1 => n92, A2 => regs(1188), B1 => n4, B2 => 
                           regs(164), ZN => n278);
   U428 : OAI211_X1 port map( C1 => n57, C2 => n1827, A => n279, B => n278, ZN 
                           => curr_proc_regs(164));
   U429 : INV_X1 port map( A => regs(1189), ZN => n1830);
   U430 : AOI22_X1 port map( A1 => n122, A2 => regs(2213), B1 => n62, B2 => 
                           regs(1701), ZN => n281);
   U431 : AOI22_X1 port map( A1 => n43, A2 => regs(677), B1 => n26, B2 => 
                           regs(165), ZN => n280);
   U432 : OAI211_X1 port map( C1 => n2215, C2 => n1830, A => n281, B => n280, 
                           ZN => curr_proc_regs(165));
   U433 : INV_X1 port map( A => regs(678), ZN => n1833);
   U434 : AOI22_X1 port map( A1 => n105, A2 => regs(2214), B1 => n73, B2 => 
                           regs(1702), ZN => n283);
   U435 : AOI22_X1 port map( A1 => n95, A2 => regs(1190), B1 => n26, B2 => 
                           regs(166), ZN => n282);
   U436 : OAI211_X1 port map( C1 => n57, C2 => n1833, A => n283, B => n282, ZN 
                           => curr_proc_regs(166));
   U437 : INV_X1 port map( A => regs(679), ZN => n1836);
   U438 : AOI22_X1 port map( A1 => n7, A2 => regs(2215), B1 => n61, B2 => 
                           regs(1703), ZN => n285);
   U439 : AOI22_X1 port map( A1 => n95, A2 => regs(1191), B1 => n26, B2 => 
                           regs(167), ZN => n284);
   U440 : OAI211_X1 port map( C1 => n10, C2 => n1836, A => n285, B => n284, ZN 
                           => curr_proc_regs(167));
   U441 : INV_X1 port map( A => regs(680), ZN => n1842);
   U442 : AOI22_X1 port map( A1 => n122, A2 => regs(2216), B1 => n62, B2 => 
                           regs(1704), ZN => n287);
   U443 : AOI22_X1 port map( A1 => n96, A2 => regs(1192), B1 => n26, B2 => 
                           regs(168), ZN => n286);
   U444 : OAI211_X1 port map( C1 => n9, C2 => n1842, A => n287, B => n286, ZN 
                           => curr_proc_regs(168));
   U445 : INV_X1 port map( A => regs(1193), ZN => n1845);
   U446 : AOI22_X1 port map( A1 => n123, A2 => regs(2217), B1 => n69, B2 => 
                           regs(1705), ZN => n289);
   U447 : AOI22_X1 port map( A1 => n43, A2 => regs(681), B1 => n25, B2 => 
                           regs(169), ZN => n288);
   U448 : OAI211_X1 port map( C1 => n13, C2 => n1845, A => n289, B => n288, ZN 
                           => curr_proc_regs(169));
   U449 : INV_X1 port map( A => regs(1040), ZN => n1357);
   U450 : AOI22_X1 port map( A1 => n104, A2 => regs(2064), B1 => n61, B2 => 
                           regs(1552), ZN => n291);
   U451 : AOI22_X1 port map( A1 => n41, A2 => regs(528), B1 => n25, B2 => 
                           regs(16), ZN => n290);
   U452 : OAI211_X1 port map( C1 => n2215, C2 => n1357, A => n291, B => n290, 
                           ZN => curr_proc_regs(16));
   U453 : INV_X1 port map( A => regs(1194), ZN => n1848);
   U454 : AOI22_X1 port map( A1 => n104, A2 => regs(2218), B1 => n62, B2 => 
                           regs(1706), ZN => n293);
   U455 : AOI22_X1 port map( A1 => n3, A2 => regs(682), B1 => n25, B2 => 
                           regs(170), ZN => n292);
   U456 : OAI211_X1 port map( C1 => n13, C2 => n1848, A => n293, B => n292, ZN 
                           => curr_proc_regs(170));
   U457 : INV_X1 port map( A => regs(1195), ZN => n1851);
   U458 : AOI22_X1 port map( A1 => n105, A2 => regs(2219), B1 => n72, B2 => 
                           regs(1707), ZN => n295);
   U459 : AOI22_X1 port map( A1 => n1, A2 => regs(683), B1 => n25, B2 => 
                           regs(171), ZN => n294);
   U460 : OAI211_X1 port map( C1 => n2215, C2 => n1851, A => n295, B => n294, 
                           ZN => curr_proc_regs(171));
   U461 : INV_X1 port map( A => regs(1196), ZN => n1854);
   U462 : AOI22_X1 port map( A1 => n7, A2 => regs(2220), B1 => n61, B2 => 
                           regs(1708), ZN => n297);
   U463 : AOI22_X1 port map( A1 => n8, A2 => regs(684), B1 => n25, B2 => 
                           regs(172), ZN => n296);
   U464 : OAI211_X1 port map( C1 => n13, C2 => n1854, A => n297, B => n296, ZN 
                           => curr_proc_regs(172));
   U465 : INV_X1 port map( A => regs(1197), ZN => n1857);
   U466 : AOI22_X1 port map( A1 => n122, A2 => regs(2221), B1 => n62, B2 => 
                           regs(1709), ZN => n299);
   U467 : AOI22_X1 port map( A1 => n3, A2 => regs(685), B1 => n25, B2 => 
                           regs(173), ZN => n298);
   U468 : OAI211_X1 port map( C1 => n2215, C2 => n1857, A => n299, B => n298, 
                           ZN => curr_proc_regs(173));
   U469 : INV_X1 port map( A => regs(686), ZN => n1860);
   U470 : AOI22_X1 port map( A1 => n123, A2 => regs(2222), B1 => n68, B2 => 
                           regs(1710), ZN => n301);
   U471 : AOI22_X1 port map( A1 => n91, A2 => regs(1198), B1 => n25, B2 => 
                           regs(174), ZN => n300);
   U472 : OAI211_X1 port map( C1 => n59, C2 => n1860, A => n301, B => n300, ZN 
                           => curr_proc_regs(174));
   U473 : INV_X1 port map( A => regs(687), ZN => n1863);
   U474 : AOI22_X1 port map( A1 => n105, A2 => regs(2223), B1 => n61, B2 => 
                           regs(1711), ZN => n303);
   U475 : AOI22_X1 port map( A1 => n100, A2 => regs(1199), B1 => n25, B2 => 
                           regs(175), ZN => n302);
   U476 : OAI211_X1 port map( C1 => n10, C2 => n1863, A => n303, B => n302, ZN 
                           => curr_proc_regs(175));
   U477 : INV_X1 port map( A => regs(1200), ZN => n1866);
   U478 : AOI22_X1 port map( A1 => n104, A2 => regs(2224), B1 => n61, B2 => 
                           regs(1712), ZN => n305);
   U479 : AOI22_X1 port map( A1 => n1, A2 => regs(688), B1 => n26, B2 => 
                           regs(176), ZN => n304);
   U480 : OAI211_X1 port map( C1 => n11, C2 => n1866, A => n305, B => n304, ZN 
                           => curr_proc_regs(176));
   U481 : INV_X1 port map( A => regs(689), ZN => n1869);
   U482 : AOI22_X1 port map( A1 => n7, A2 => regs(2225), B1 => n62, B2 => 
                           regs(1713), ZN => n307);
   U483 : AOI22_X1 port map( A1 => n91, A2 => regs(1201), B1 => n25, B2 => 
                           regs(177), ZN => n306);
   U484 : OAI211_X1 port map( C1 => n58, C2 => n1869, A => n307, B => n306, ZN 
                           => curr_proc_regs(177));
   U485 : INV_X1 port map( A => regs(1202), ZN => n1875);
   U486 : AOI22_X1 port map( A1 => n122, A2 => regs(2226), B1 => n74, B2 => 
                           regs(1714), ZN => n309);
   U487 : AOI22_X1 port map( A1 => n53, A2 => regs(690), B1 => n39, B2 => 
                           regs(178), ZN => n308);
   U488 : OAI211_X1 port map( C1 => n11, C2 => n1875, A => n309, B => n308, ZN 
                           => curr_proc_regs(178));
   U489 : INV_X1 port map( A => regs(691), ZN => n1878);
   U490 : AOI22_X1 port map( A1 => n123, A2 => regs(2227), B1 => n62, B2 => 
                           regs(1715), ZN => n311);
   U491 : AOI22_X1 port map( A1 => n89, A2 => regs(1203), B1 => n4, B2 => 
                           regs(179), ZN => n310);
   U492 : OAI211_X1 port map( C1 => n10, C2 => n1878, A => n311, B => n310, ZN 
                           => curr_proc_regs(179));
   U493 : INV_X1 port map( A => regs(1041), ZN => n1360);
   U494 : AOI22_X1 port map( A1 => n104, A2 => regs(2065), B1 => n61, B2 => 
                           regs(1553), ZN => n313);
   U495 : AOI22_X1 port map( A1 => n53, A2 => regs(529), B1 => n26, B2 => 
                           regs(17), ZN => n312);
   U496 : OAI211_X1 port map( C1 => n6, C2 => n1360, A => n313, B => n312, ZN 
                           => curr_proc_regs(17));
   U497 : INV_X1 port map( A => regs(692), ZN => n1881);
   U498 : AOI22_X1 port map( A1 => n105, A2 => regs(2228), B1 => n62, B2 => 
                           regs(1716), ZN => n315);
   U499 : AOI22_X1 port map( A1 => n98, A2 => regs(1204), B1 => n26, B2 => 
                           regs(180), ZN => n314);
   U500 : OAI211_X1 port map( C1 => n9, C2 => n1881, A => n315, B => n314, ZN 
                           => curr_proc_regs(180));
   U501 : INV_X1 port map( A => regs(693), ZN => n1884);
   U502 : AOI22_X1 port map( A1 => n7, A2 => regs(2229), B1 => n71, B2 => 
                           regs(1717), ZN => n317);
   U503 : AOI22_X1 port map( A1 => n96, A2 => regs(1205), B1 => n26, B2 => 
                           regs(181), ZN => n316);
   U504 : OAI211_X1 port map( C1 => n2201, C2 => n1884, A => n317, B => n316, 
                           ZN => curr_proc_regs(181));
   U505 : INV_X1 port map( A => regs(694), ZN => n1887);
   U506 : AOI22_X1 port map( A1 => n122, A2 => regs(2230), B1 => n71, B2 => 
                           regs(1718), ZN => n319);
   U507 : AOI22_X1 port map( A1 => n88, A2 => regs(1206), B1 => n26, B2 => 
                           regs(182), ZN => n318);
   U508 : OAI211_X1 port map( C1 => n9, C2 => n1887, A => n319, B => n318, ZN 
                           => curr_proc_regs(182));
   U509 : INV_X1 port map( A => regs(695), ZN => n1890);
   U510 : AOI22_X1 port map( A1 => n123, A2 => regs(2231), B1 => n61, B2 => 
                           regs(1719), ZN => n321);
   U511 : AOI22_X1 port map( A1 => n94, A2 => regs(1207), B1 => n26, B2 => 
                           regs(183), ZN => n320);
   U512 : OAI211_X1 port map( C1 => n9, C2 => n1890, A => n321, B => n320, ZN 
                           => curr_proc_regs(183));
   U513 : INV_X1 port map( A => regs(696), ZN => n1893);
   U514 : AOI22_X1 port map( A1 => n104, A2 => regs(2232), B1 => n62, B2 => 
                           regs(1720), ZN => n323);
   U515 : AOI22_X1 port map( A1 => n95, A2 => regs(1208), B1 => n26, B2 => 
                           regs(184), ZN => n322);
   U516 : OAI211_X1 port map( C1 => n2201, C2 => n1893, A => n323, B => n322, 
                           ZN => curr_proc_regs(184));
   U517 : INV_X1 port map( A => regs(697), ZN => n1896);
   U518 : AOI22_X1 port map( A1 => n105, A2 => regs(2233), B1 => n5, B2 => 
                           regs(1721), ZN => n325);
   U519 : AOI22_X1 port map( A1 => n89, A2 => regs(1209), B1 => n26, B2 => 
                           regs(185), ZN => n324);
   U520 : OAI211_X1 port map( C1 => n9, C2 => n1896, A => n325, B => n324, ZN 
                           => curr_proc_regs(185));
   U521 : INV_X1 port map( A => regs(1210), ZN => n1899);
   U522 : AOI22_X1 port map( A1 => n125, A2 => regs(2234), B1 => n61, B2 => 
                           regs(1722), ZN => n327);
   U523 : AOI22_X1 port map( A1 => n53, A2 => regs(698), B1 => n26, B2 => 
                           regs(186), ZN => n326);
   U524 : OAI211_X1 port map( C1 => n2215, C2 => n1899, A => n327, B => n326, 
                           ZN => curr_proc_regs(186));
   U525 : INV_X1 port map( A => regs(1211), ZN => n1902);
   U526 : AOI22_X1 port map( A1 => n122, A2 => regs(2235), B1 => n73, B2 => 
                           regs(1723), ZN => n329);
   U527 : AOI22_X1 port map( A1 => n53, A2 => regs(699), B1 => n35, B2 => 
                           regs(187), ZN => n328);
   U528 : OAI211_X1 port map( C1 => n11, C2 => n1902, A => n329, B => n328, ZN 
                           => curr_proc_regs(187));
   U529 : INV_X1 port map( A => regs(700), ZN => n1911);
   U530 : AOI22_X1 port map( A1 => n123, A2 => regs(2236), B1 => n61, B2 => 
                           regs(1724), ZN => n331);
   U531 : AOI22_X1 port map( A1 => n88, A2 => regs(1212), B1 => n39, B2 => 
                           regs(188), ZN => n330);
   U532 : OAI211_X1 port map( C1 => n58, C2 => n1911, A => n331, B => n330, ZN 
                           => curr_proc_regs(188));
   U533 : INV_X1 port map( A => regs(701), ZN => n1914);
   U534 : AOI22_X1 port map( A1 => n123, A2 => regs(2237), B1 => n62, B2 => 
                           regs(1725), ZN => n333);
   U535 : AOI22_X1 port map( A1 => n100, A2 => regs(1213), B1 => n4, B2 => 
                           regs(189), ZN => n332);
   U536 : OAI211_X1 port map( C1 => n9, C2 => n1914, A => n333, B => n332, ZN 
                           => curr_proc_regs(189));
   U537 : INV_X1 port map( A => regs(1042), ZN => n1365);
   U538 : AOI22_X1 port map( A1 => n123, A2 => regs(2066), B1 => n61, B2 => 
                           regs(1554), ZN => n335);
   U539 : AOI22_X1 port map( A1 => n53, A2 => regs(530), B1 => n28, B2 => 
                           regs(18), ZN => n334);
   U540 : OAI211_X1 port map( C1 => n2215, C2 => n1365, A => n335, B => n334, 
                           ZN => curr_proc_regs(18));
   U541 : INV_X1 port map( A => regs(702), ZN => n1917);
   U542 : AOI22_X1 port map( A1 => n123, A2 => regs(2238), B1 => n62, B2 => 
                           regs(1726), ZN => n337);
   U543 : AOI22_X1 port map( A1 => n92, A2 => regs(1214), B1 => n21, B2 => 
                           regs(190), ZN => n336);
   U544 : OAI211_X1 port map( C1 => n9, C2 => n1917, A => n337, B => n336, ZN 
                           => curr_proc_regs(190));
   U545 : INV_X1 port map( A => regs(703), ZN => n1920);
   U546 : AOI22_X1 port map( A1 => n123, A2 => regs(2239), B1 => n5, B2 => 
                           regs(1727), ZN => n339);
   U547 : AOI22_X1 port map( A1 => n94, A2 => regs(1215), B1 => n22, B2 => 
                           regs(191), ZN => n338);
   U548 : OAI211_X1 port map( C1 => n9, C2 => n1920, A => n339, B => n338, ZN 
                           => curr_proc_regs(191));
   U549 : INV_X1 port map( A => regs(1216), ZN => n1923);
   U550 : AOI22_X1 port map( A1 => n123, A2 => regs(2240), B1 => n62, B2 => 
                           regs(1728), ZN => n341);
   U551 : AOI22_X1 port map( A1 => n53, A2 => regs(704), B1 => n23, B2 => 
                           regs(192), ZN => n340);
   U552 : OAI211_X1 port map( C1 => n78, C2 => n1923, A => n341, B => n340, ZN 
                           => curr_proc_regs(192));
   U553 : INV_X1 port map( A => regs(1217), ZN => n1926);
   U554 : AOI22_X1 port map( A1 => n123, A2 => regs(2241), B1 => n66, B2 => 
                           regs(1729), ZN => n343);
   U555 : AOI22_X1 port map( A1 => n53, A2 => regs(705), B1 => n24, B2 => 
                           regs(193), ZN => n342);
   U556 : OAI211_X1 port map( C1 => n103, C2 => n1926, A => n343, B => n342, ZN
                           => curr_proc_regs(193));
   U557 : INV_X1 port map( A => regs(1218), ZN => n1929);
   U558 : AOI22_X1 port map( A1 => n123, A2 => regs(2242), B1 => n61, B2 => 
                           regs(1730), ZN => n345);
   U559 : AOI22_X1 port map( A1 => n46, A2 => regs(706), B1 => n17, B2 => 
                           regs(194), ZN => n344);
   U560 : OAI211_X1 port map( C1 => n103, C2 => n1929, A => n345, B => n344, ZN
                           => curr_proc_regs(194));
   U561 : INV_X1 port map( A => regs(1219), ZN => n1932);
   U562 : AOI22_X1 port map( A1 => n123, A2 => regs(2243), B1 => n62, B2 => 
                           regs(1731), ZN => n347);
   U563 : AOI22_X1 port map( A1 => n43, A2 => regs(707), B1 => n18, B2 => 
                           regs(195), ZN => n346);
   U564 : OAI211_X1 port map( C1 => n78, C2 => n1932, A => n347, B => n346, ZN 
                           => curr_proc_regs(195));
   U565 : INV_X1 port map( A => regs(708), ZN => n1935);
   U566 : AOI22_X1 port map( A1 => n123, A2 => regs(2244), B1 => n66, B2 => 
                           regs(1732), ZN => n349);
   U567 : AOI22_X1 port map( A1 => n95, A2 => regs(1220), B1 => n19, B2 => 
                           regs(196), ZN => n348);
   U568 : OAI211_X1 port map( C1 => n9, C2 => n1935, A => n349, B => n348, ZN 
                           => curr_proc_regs(196));
   U569 : INV_X1 port map( A => regs(1221), ZN => n1938);
   U570 : AOI22_X1 port map( A1 => n123, A2 => regs(2245), B1 => n5, B2 => 
                           regs(1733), ZN => n351);
   U571 : AOI22_X1 port map( A1 => n43, A2 => regs(709), B1 => n27, B2 => 
                           regs(197), ZN => n350);
   U572 : OAI211_X1 port map( C1 => n103, C2 => n1938, A => n351, B => n350, ZN
                           => curr_proc_regs(197));
   U573 : INV_X1 port map( A => regs(1222), ZN => n1944);
   U574 : AOI22_X1 port map( A1 => n123, A2 => regs(2246), B1 => n63, B2 => 
                           regs(1734), ZN => n353);
   U575 : AOI22_X1 port map( A1 => n43, A2 => regs(710), B1 => n27, B2 => 
                           regs(198), ZN => n352);
   U576 : OAI211_X1 port map( C1 => n78, C2 => n1944, A => n353, B => n352, ZN 
                           => curr_proc_regs(198));
   U577 : INV_X1 port map( A => regs(711), ZN => n1947);
   U578 : AOI22_X1 port map( A1 => n122, A2 => regs(2247), B1 => n74, B2 => 
                           regs(1735), ZN => n355);
   U579 : AOI22_X1 port map( A1 => n89, A2 => regs(1223), B1 => n27, B2 => 
                           regs(199), ZN => n354);
   U580 : OAI211_X1 port map( C1 => n9, C2 => n1947, A => n355, B => n354, ZN 
                           => curr_proc_regs(199));
   U581 : INV_X1 port map( A => regs(531), ZN => n1368);
   U582 : AOI22_X1 port map( A1 => n122, A2 => regs(2067), B1 => n70, B2 => 
                           regs(1555), ZN => n357);
   U583 : AOI22_X1 port map( A1 => n88, A2 => regs(1043), B1 => n27, B2 => 
                           regs(19), ZN => n356);
   U584 : OAI211_X1 port map( C1 => n9, C2 => n1368, A => n357, B => n356, ZN 
                           => curr_proc_regs(19));
   U585 : INV_X1 port map( A => regs(513), ZN => n1313);
   U586 : AOI22_X1 port map( A1 => n122, A2 => regs(2049), B1 => n74, B2 => 
                           regs(1537), ZN => n359);
   U587 : AOI22_X1 port map( A1 => n98, A2 => regs(1025), B1 => n27, B2 => 
                           regs(1), ZN => n358);
   U588 : OAI211_X1 port map( C1 => n9, C2 => n1313, A => n359, B => n358, ZN 
                           => curr_proc_regs(1));
   U589 : INV_X1 port map( A => regs(1224), ZN => n1950);
   U590 : AOI22_X1 port map( A1 => n122, A2 => regs(2248), B1 => n61, B2 => 
                           regs(1736), ZN => n361);
   U591 : AOI22_X1 port map( A1 => n43, A2 => regs(712), B1 => n23, B2 => 
                           regs(200), ZN => n360);
   U592 : OAI211_X1 port map( C1 => n103, C2 => n1950, A => n361, B => n360, ZN
                           => curr_proc_regs(200));
   U593 : INV_X1 port map( A => regs(1225), ZN => n1953);
   U594 : AOI22_X1 port map( A1 => n122, A2 => regs(2249), B1 => n62, B2 => 
                           regs(1737), ZN => n363);
   U595 : AOI22_X1 port map( A1 => n43, A2 => regs(713), B1 => n24, B2 => 
                           regs(201), ZN => n362);
   U596 : OAI211_X1 port map( C1 => n78, C2 => n1953, A => n363, B => n362, ZN 
                           => curr_proc_regs(201));
   U597 : INV_X1 port map( A => regs(714), ZN => n1956);
   U598 : AOI22_X1 port map( A1 => n122, A2 => regs(2250), B1 => n65, B2 => 
                           regs(1738), ZN => n365);
   U599 : AOI22_X1 port map( A1 => n100, A2 => regs(1226), B1 => n17, B2 => 
                           regs(202), ZN => n364);
   U600 : OAI211_X1 port map( C1 => n9, C2 => n1956, A => n365, B => n364, ZN 
                           => curr_proc_regs(202));
   U601 : INV_X1 port map( A => regs(715), ZN => n1959);
   U602 : AOI22_X1 port map( A1 => n122, A2 => regs(2251), B1 => n69, B2 => 
                           regs(1739), ZN => n367);
   U603 : AOI22_X1 port map( A1 => n96, A2 => regs(1227), B1 => n18, B2 => 
                           regs(203), ZN => n366);
   U604 : OAI211_X1 port map( C1 => n58, C2 => n1959, A => n367, B => n366, ZN 
                           => curr_proc_regs(203));
   U605 : INV_X1 port map( A => regs(1228), ZN => n1962);
   U606 : AOI22_X1 port map( A1 => n122, A2 => regs(2252), B1 => n67, B2 => 
                           regs(1740), ZN => n369);
   U607 : AOI22_X1 port map( A1 => n43, A2 => regs(716), B1 => n19, B2 => 
                           regs(204), ZN => n368);
   U608 : OAI211_X1 port map( C1 => n6, C2 => n1962, A => n369, B => n368, ZN 
                           => curr_proc_regs(204));
   U609 : INV_X1 port map( A => regs(1229), ZN => n1965);
   U610 : AOI22_X1 port map( A1 => n122, A2 => regs(2253), B1 => n61, B2 => 
                           regs(1741), ZN => n371);
   U611 : AOI22_X1 port map( A1 => n43, A2 => regs(717), B1 => n27, B2 => 
                           regs(205), ZN => n370);
   U612 : OAI211_X1 port map( C1 => n6, C2 => n1965, A => n371, B => n370, ZN 
                           => curr_proc_regs(205));
   U613 : INV_X1 port map( A => regs(718), ZN => n1968);
   U614 : AOI22_X1 port map( A1 => n122, A2 => regs(2254), B1 => n76, B2 => 
                           regs(1742), ZN => n373);
   U615 : AOI22_X1 port map( A1 => n91, A2 => regs(1230), B1 => n26, B2 => 
                           regs(206), ZN => n372);
   U616 : OAI211_X1 port map( C1 => n58, C2 => n1968, A => n373, B => n372, ZN 
                           => curr_proc_regs(206));
   U617 : INV_X1 port map( A => regs(719), ZN => n1971);
   U618 : AOI22_X1 port map( A1 => n122, A2 => regs(2255), B1 => n75, B2 => 
                           regs(1743), ZN => n375);
   U619 : AOI22_X1 port map( A1 => n92, A2 => regs(1231), B1 => n25, B2 => 
                           regs(207), ZN => n374);
   U620 : OAI211_X1 port map( C1 => n10, C2 => n1971, A => n375, B => n374, ZN 
                           => curr_proc_regs(207));
   U621 : INV_X1 port map( A => regs(1232), ZN => n1977);
   U622 : AOI22_X1 port map( A1 => n122, A2 => regs(2256), B1 => n63, B2 => 
                           regs(1744), ZN => n377);
   U623 : AOI22_X1 port map( A1 => n43, A2 => regs(720), B1 => n28, B2 => 
                           regs(208), ZN => n376);
   U624 : OAI211_X1 port map( C1 => n6, C2 => n1977, A => n377, B => n376, ZN 
                           => curr_proc_regs(208));
   U625 : INV_X1 port map( A => regs(1233), ZN => n1980);
   U626 : AOI22_X1 port map( A1 => n7, A2 => regs(2257), B1 => n63, B2 => 
                           regs(1745), ZN => n379);
   U627 : AOI22_X1 port map( A1 => n43, A2 => regs(721), B1 => n29, B2 => 
                           regs(209), ZN => n378);
   U628 : OAI211_X1 port map( C1 => n6, C2 => n1980, A => n379, B => n378, ZN 
                           => curr_proc_regs(209));
   U629 : INV_X1 port map( A => regs(1044), ZN => n1371);
   U630 : AOI22_X1 port map( A1 => n7, A2 => regs(2068), B1 => n63, B2 => 
                           regs(1556), ZN => n381);
   U631 : AOI22_X1 port map( A1 => n43, A2 => regs(532), B1 => n30, B2 => 
                           regs(20), ZN => n380);
   U632 : OAI211_X1 port map( C1 => n6, C2 => n1371, A => n381, B => n380, ZN 
                           => curr_proc_regs(20));
   U633 : INV_X1 port map( A => regs(1234), ZN => n1983);
   U634 : AOI22_X1 port map( A1 => n7, A2 => regs(2258), B1 => n63, B2 => 
                           regs(1746), ZN => n383);
   U635 : AOI22_X1 port map( A1 => n43, A2 => regs(722), B1 => n32, B2 => 
                           regs(210), ZN => n382);
   U636 : OAI211_X1 port map( C1 => n6, C2 => n1983, A => n383, B => n382, ZN 
                           => curr_proc_regs(210));
   U637 : INV_X1 port map( A => regs(1235), ZN => n1986);
   U638 : AOI22_X1 port map( A1 => n7, A2 => regs(2259), B1 => n63, B2 => 
                           regs(1747), ZN => n385);
   U639 : AOI22_X1 port map( A1 => n47, A2 => regs(723), B1 => n27, B2 => 
                           regs(211), ZN => n384);
   U640 : OAI211_X1 port map( C1 => n6, C2 => n1986, A => n385, B => n384, ZN 
                           => curr_proc_regs(211));
   U641 : INV_X1 port map( A => regs(724), ZN => n1989);
   U642 : AOI22_X1 port map( A1 => n7, A2 => regs(2260), B1 => n63, B2 => 
                           regs(1748), ZN => n387);
   U643 : AOI22_X1 port map( A1 => n96, A2 => regs(1236), B1 => n27, B2 => 
                           regs(212), ZN => n386);
   U644 : OAI211_X1 port map( C1 => n9, C2 => n1989, A => n387, B => n386, ZN 
                           => curr_proc_regs(212));
   U645 : INV_X1 port map( A => regs(1237), ZN => n1992);
   U646 : AOI22_X1 port map( A1 => n7, A2 => regs(2261), B1 => n63, B2 => 
                           regs(1749), ZN => n389);
   U647 : AOI22_X1 port map( A1 => n46, A2 => regs(725), B1 => n27, B2 => 
                           regs(213), ZN => n388);
   U648 : OAI211_X1 port map( C1 => n6, C2 => n1992, A => n389, B => n388, ZN 
                           => curr_proc_regs(213));
   U649 : INV_X1 port map( A => regs(1238), ZN => n1995);
   U650 : AOI22_X1 port map( A1 => n7, A2 => regs(2262), B1 => n63, B2 => 
                           regs(1750), ZN => n391);
   U651 : AOI22_X1 port map( A1 => n46, A2 => regs(726), B1 => n27, B2 => 
                           regs(214), ZN => n390);
   U652 : OAI211_X1 port map( C1 => n78, C2 => n1995, A => n391, B => n390, ZN 
                           => curr_proc_regs(214));
   U653 : INV_X1 port map( A => regs(1239), ZN => n1998);
   U654 : AOI22_X1 port map( A1 => n7, A2 => regs(2263), B1 => n63, B2 => 
                           regs(1751), ZN => n393);
   U655 : AOI22_X1 port map( A1 => n47, A2 => regs(727), B1 => n27, B2 => 
                           regs(215), ZN => n392);
   U656 : OAI211_X1 port map( C1 => n11, C2 => n1998, A => n393, B => n392, ZN 
                           => curr_proc_regs(215));
   U657 : INV_X1 port map( A => regs(1240), ZN => n2001);
   U658 : AOI22_X1 port map( A1 => n7, A2 => regs(2264), B1 => n63, B2 => 
                           regs(1752), ZN => n395);
   U659 : AOI22_X1 port map( A1 => n46, A2 => regs(728), B1 => n27, B2 => 
                           regs(216), ZN => n394);
   U660 : OAI211_X1 port map( C1 => n2215, C2 => n2001, A => n395, B => n394, 
                           ZN => curr_proc_regs(216));
   U661 : INV_X1 port map( A => regs(1241), ZN => n2004);
   U662 : AOI22_X1 port map( A1 => n7, A2 => regs(2265), B1 => n63, B2 => 
                           regs(1753), ZN => n397);
   U663 : AOI22_X1 port map( A1 => n52, A2 => regs(729), B1 => n27, B2 => 
                           regs(217), ZN => n396);
   U664 : OAI211_X1 port map( C1 => n78, C2 => n2004, A => n397, B => n396, ZN 
                           => curr_proc_regs(217));
   U665 : INV_X1 port map( A => regs(1242), ZN => n2010);
   U666 : AOI22_X1 port map( A1 => n7, A2 => regs(2266), B1 => n63, B2 => 
                           regs(1754), ZN => n399);
   U667 : AOI22_X1 port map( A1 => n51, A2 => regs(730), B1 => n27, B2 => 
                           regs(218), ZN => n398);
   U668 : OAI211_X1 port map( C1 => n6, C2 => n2010, A => n399, B => n398, ZN 
                           => curr_proc_regs(218));
   U669 : INV_X1 port map( A => regs(731), ZN => n2013);
   U670 : AOI22_X1 port map( A1 => n7, A2 => regs(2267), B1 => n64, B2 => 
                           regs(1755), ZN => n401);
   U671 : AOI22_X1 port map( A1 => n94, A2 => regs(1243), B1 => n28, B2 => 
                           regs(219), ZN => n400);
   U672 : OAI211_X1 port map( C1 => n9, C2 => n2013, A => n401, B => n400, ZN 
                           => curr_proc_regs(219));
   U673 : INV_X1 port map( A => regs(533), ZN => n1374);
   U674 : AOI22_X1 port map( A1 => win(4), A2 => regs(2069), B1 => n72, B2 => 
                           regs(1557), ZN => n403);
   U675 : AOI22_X1 port map( A1 => n95, A2 => regs(1045), B1 => n28, B2 => 
                           regs(21), ZN => n402);
   U676 : OAI211_X1 port map( C1 => n9, C2 => n1374, A => n403, B => n402, ZN 
                           => curr_proc_regs(21));
   U677 : INV_X1 port map( A => regs(732), ZN => n2016);
   U678 : AOI22_X1 port map( A1 => n119, A2 => regs(2268), B1 => n63, B2 => 
                           regs(1756), ZN => n405);
   U679 : AOI22_X1 port map( A1 => n88, A2 => regs(1244), B1 => n28, B2 => 
                           regs(220), ZN => n404);
   U680 : OAI211_X1 port map( C1 => n2201, C2 => n2016, A => n405, B => n404, 
                           ZN => curr_proc_regs(220));
   U681 : INV_X1 port map( A => regs(1245), ZN => n2019);
   U682 : AOI22_X1 port map( A1 => n120, A2 => regs(2269), B1 => n63, B2 => 
                           regs(1757), ZN => n407);
   U683 : AOI22_X1 port map( A1 => n50, A2 => regs(733), B1 => n28, B2 => 
                           regs(221), ZN => n406);
   U684 : OAI211_X1 port map( C1 => n6, C2 => n2019, A => n407, B => n406, ZN 
                           => curr_proc_regs(221));
   U685 : INV_X1 port map( A => regs(734), ZN => n2022);
   U686 : AOI22_X1 port map( A1 => n121, A2 => regs(2270), B1 => n60, B2 => 
                           regs(1758), ZN => n409);
   U687 : AOI22_X1 port map( A1 => n100, A2 => regs(1246), B1 => n18, B2 => 
                           regs(222), ZN => n408);
   U688 : OAI211_X1 port map( C1 => n9, C2 => n2022, A => n409, B => n408, ZN 
                           => curr_proc_regs(222));
   U689 : INV_X1 port map( A => regs(735), ZN => n2025);
   U690 : AOI22_X1 port map( A1 => win(4), A2 => regs(2271), B1 => n64, B2 => 
                           regs(1759), ZN => n411);
   U691 : AOI22_X1 port map( A1 => n98, A2 => regs(1247), B1 => n19, B2 => 
                           regs(223), ZN => n410);
   U692 : OAI211_X1 port map( C1 => n9, C2 => n2025, A => n411, B => n410, ZN 
                           => curr_proc_regs(223));
   U693 : INV_X1 port map( A => regs(1248), ZN => n2028);
   U694 : AOI22_X1 port map( A1 => win(4), A2 => regs(2272), B1 => n2211, B2 =>
                           regs(1760), ZN => n413);
   U695 : AOI22_X1 port map( A1 => n49, A2 => regs(736), B1 => n27, B2 => 
                           regs(224), ZN => n412);
   U696 : OAI211_X1 port map( C1 => n11, C2 => n2028, A => n413, B => n412, ZN 
                           => curr_proc_regs(224));
   U697 : INV_X1 port map( A => regs(1249), ZN => n2031);
   U698 : AOI22_X1 port map( A1 => win(4), A2 => regs(2273), B1 => n63, B2 => 
                           regs(1761), ZN => n415);
   U699 : AOI22_X1 port map( A1 => n48, A2 => regs(737), B1 => n26, B2 => 
                           regs(225), ZN => n414);
   U700 : OAI211_X1 port map( C1 => n11, C2 => n2031, A => n415, B => n414, ZN 
                           => curr_proc_regs(225));
   U701 : INV_X1 port map( A => regs(738), ZN => n2034);
   U702 : AOI22_X1 port map( A1 => n119, A2 => regs(2274), B1 => n60, B2 => 
                           regs(1762), ZN => n417);
   U703 : AOI22_X1 port map( A1 => n100, A2 => regs(1250), B1 => n25, B2 => 
                           regs(226), ZN => n416);
   U704 : OAI211_X1 port map( C1 => n9, C2 => n2034, A => n417, B => n416, ZN 
                           => curr_proc_regs(226));
   U705 : INV_X1 port map( A => regs(1251), ZN => n2037);
   U706 : AOI22_X1 port map( A1 => n120, A2 => regs(2275), B1 => n60, B2 => 
                           regs(1763), ZN => n419);
   U707 : AOI22_X1 port map( A1 => n47, A2 => regs(739), B1 => n32, B2 => 
                           regs(227), ZN => n418);
   U708 : OAI211_X1 port map( C1 => n11, C2 => n2037, A => n419, B => n418, ZN 
                           => curr_proc_regs(227));
   U709 : INV_X1 port map( A => regs(1252), ZN => n2043);
   U710 : AOI22_X1 port map( A1 => n121, A2 => regs(2276), B1 => n64, B2 => 
                           regs(1764), ZN => n421);
   U711 : AOI22_X1 port map( A1 => n49, A2 => regs(740), B1 => n35, B2 => 
                           regs(228), ZN => n420);
   U712 : OAI211_X1 port map( C1 => n11, C2 => n2043, A => n421, B => n420, ZN 
                           => curr_proc_regs(228));
   U713 : INV_X1 port map( A => regs(1253), ZN => n2046);
   U714 : AOI22_X1 port map( A1 => n119, A2 => regs(2277), B1 => n72, B2 => 
                           regs(1765), ZN => n423);
   U715 : AOI22_X1 port map( A1 => n48, A2 => regs(741), B1 => n37, B2 => 
                           regs(229), ZN => n422);
   U716 : OAI211_X1 port map( C1 => n11, C2 => n2046, A => n423, B => n422, ZN 
                           => curr_proc_regs(229));
   U717 : INV_X1 port map( A => regs(534), ZN => n1377);
   U718 : AOI22_X1 port map( A1 => n119, A2 => regs(2070), B1 => n69, B2 => 
                           regs(1558), ZN => n425);
   U719 : AOI22_X1 port map( A1 => n83, A2 => regs(1046), B1 => n29, B2 => 
                           regs(22), ZN => n424);
   U720 : OAI211_X1 port map( C1 => n9, C2 => n1377, A => n425, B => n424, ZN 
                           => curr_proc_regs(22));
   U721 : INV_X1 port map( A => regs(1254), ZN => n2049);
   U722 : AOI22_X1 port map( A1 => n120, A2 => regs(2278), B1 => n5, B2 => 
                           regs(1766), ZN => n427);
   U723 : AOI22_X1 port map( A1 => n47, A2 => regs(742), B1 => n29, B2 => 
                           regs(230), ZN => n426);
   U724 : OAI211_X1 port map( C1 => n11, C2 => n2049, A => n427, B => n426, ZN 
                           => curr_proc_regs(230));
   U725 : INV_X1 port map( A => regs(1255), ZN => n2052);
   U726 : AOI22_X1 port map( A1 => n121, A2 => regs(2279), B1 => n74, B2 => 
                           regs(1767), ZN => n429);
   U727 : AOI22_X1 port map( A1 => n50, A2 => regs(743), B1 => n29, B2 => 
                           regs(231), ZN => n428);
   U728 : OAI211_X1 port map( C1 => n11, C2 => n2052, A => n429, B => n428, ZN 
                           => curr_proc_regs(231));
   U729 : INV_X1 port map( A => regs(1256), ZN => n2055);
   U730 : AOI22_X1 port map( A1 => n120, A2 => regs(2280), B1 => n71, B2 => 
                           regs(1768), ZN => n431);
   U731 : AOI22_X1 port map( A1 => n46, A2 => regs(744), B1 => n29, B2 => 
                           regs(232), ZN => n430);
   U732 : OAI211_X1 port map( C1 => n78, C2 => n2055, A => n431, B => n430, ZN 
                           => curr_proc_regs(232));
   U733 : INV_X1 port map( A => regs(1257), ZN => n2058);
   U734 : AOI22_X1 port map( A1 => win(4), A2 => regs(2281), B1 => n68, B2 => 
                           regs(1769), ZN => n433);
   U735 : AOI22_X1 port map( A1 => n46, A2 => regs(745), B1 => n28, B2 => 
                           regs(233), ZN => n432);
   U736 : OAI211_X1 port map( C1 => n78, C2 => n2058, A => n433, B => n432, ZN 
                           => curr_proc_regs(233));
   U737 : INV_X1 port map( A => regs(1258), ZN => n2061);
   U738 : AOI22_X1 port map( A1 => n119, A2 => regs(2282), B1 => n66, B2 => 
                           regs(1770), ZN => n435);
   U739 : AOI22_X1 port map( A1 => n48, A2 => regs(746), B1 => n28, B2 => 
                           regs(234), ZN => n434);
   U740 : OAI211_X1 port map( C1 => n103, C2 => n2061, A => n435, B => n434, ZN
                           => curr_proc_regs(234));
   U741 : INV_X1 port map( A => regs(747), ZN => n2064);
   U742 : AOI22_X1 port map( A1 => n120, A2 => regs(2283), B1 => n72, B2 => 
                           regs(1771), ZN => n437);
   U743 : AOI22_X1 port map( A1 => n97, A2 => regs(1259), B1 => n28, B2 => 
                           regs(235), ZN => n436);
   U744 : OAI211_X1 port map( C1 => n9, C2 => n2064, A => n437, B => n436, ZN 
                           => curr_proc_regs(235));
   U745 : INV_X1 port map( A => regs(748), ZN => n2067);
   U746 : AOI22_X1 port map( A1 => n121, A2 => regs(2284), B1 => n63, B2 => 
                           regs(1772), ZN => n439);
   U747 : AOI22_X1 port map( A1 => n93, A2 => regs(1260), B1 => n28, B2 => 
                           regs(236), ZN => n438);
   U748 : OAI211_X1 port map( C1 => n9, C2 => n2067, A => n439, B => n438, ZN 
                           => curr_proc_regs(236));
   U749 : INV_X1 port map( A => regs(1261), ZN => n2070);
   U750 : AOI22_X1 port map( A1 => n121, A2 => regs(2285), B1 => n70, B2 => 
                           regs(1773), ZN => n441);
   U751 : AOI22_X1 port map( A1 => n52, A2 => regs(749), B1 => n28, B2 => 
                           regs(237), ZN => n440);
   U752 : OAI211_X1 port map( C1 => n78, C2 => n2070, A => n441, B => n440, ZN 
                           => curr_proc_regs(237));
   U753 : INV_X1 port map( A => regs(750), ZN => n2076);
   U754 : AOI22_X1 port map( A1 => win(4), A2 => regs(2286), B1 => n74, B2 => 
                           regs(1774), ZN => n443);
   U755 : AOI22_X1 port map( A1 => n83, A2 => regs(1262), B1 => n28, B2 => 
                           regs(238), ZN => n442);
   U756 : OAI211_X1 port map( C1 => n9, C2 => n2076, A => n443, B => n442, ZN 
                           => curr_proc_regs(238));
   U757 : INV_X1 port map( A => regs(751), ZN => n2079);
   U758 : AOI22_X1 port map( A1 => n119, A2 => regs(2287), B1 => n65, B2 => 
                           regs(1775), ZN => n445);
   U759 : AOI22_X1 port map( A1 => n98, A2 => regs(1263), B1 => n28, B2 => 
                           regs(239), ZN => n444);
   U760 : OAI211_X1 port map( C1 => n10, C2 => n2079, A => n445, B => n444, ZN 
                           => curr_proc_regs(239));
   U761 : INV_X1 port map( A => regs(1047), ZN => n1380);
   U762 : AOI22_X1 port map( A1 => n120, A2 => regs(2071), B1 => n69, B2 => 
                           regs(1559), ZN => n447);
   U763 : AOI22_X1 port map( A1 => n51, A2 => regs(535), B1 => n28, B2 => 
                           regs(23), ZN => n446);
   U764 : OAI211_X1 port map( C1 => n103, C2 => n1380, A => n447, B => n446, ZN
                           => curr_proc_regs(23));
   U765 : INV_X1 port map( A => regs(1264), ZN => n2082);
   U766 : AOI22_X1 port map( A1 => n121, A2 => regs(2288), B1 => n63, B2 => 
                           regs(1776), ZN => n449);
   U767 : AOI22_X1 port map( A1 => n50, A2 => regs(752), B1 => n30, B2 => 
                           regs(240), ZN => n448);
   U768 : OAI211_X1 port map( C1 => n78, C2 => n2082, A => n449, B => n448, ZN 
                           => curr_proc_regs(240));
   U769 : INV_X1 port map( A => regs(753), ZN => n2085);
   U770 : AOI22_X1 port map( A1 => win(4), A2 => regs(2289), B1 => n63, B2 => 
                           regs(1777), ZN => n451);
   U771 : AOI22_X1 port map( A1 => n97, A2 => regs(1265), B1 => n30, B2 => 
                           regs(241), ZN => n450);
   U772 : OAI211_X1 port map( C1 => n10, C2 => n2085, A => n451, B => n450, ZN 
                           => curr_proc_regs(241));
   U773 : INV_X1 port map( A => regs(1266), ZN => n2088);
   U774 : AOI22_X1 port map( A1 => n119, A2 => regs(2290), B1 => n64, B2 => 
                           regs(1778), ZN => n453);
   U775 : AOI22_X1 port map( A1 => n49, A2 => regs(754), B1 => n30, B2 => 
                           regs(242), ZN => n452);
   U776 : OAI211_X1 port map( C1 => n103, C2 => n2088, A => n453, B => n452, ZN
                           => curr_proc_regs(242));
   U777 : INV_X1 port map( A => regs(755), ZN => n2091);
   U778 : AOI22_X1 port map( A1 => n120, A2 => regs(2291), B1 => n60, B2 => 
                           regs(1779), ZN => n455);
   U779 : AOI22_X1 port map( A1 => n99, A2 => regs(1267), B1 => n30, B2 => 
                           regs(243), ZN => n454);
   U780 : OAI211_X1 port map( C1 => n10, C2 => n2091, A => n455, B => n454, ZN 
                           => curr_proc_regs(243));
   U781 : INV_X1 port map( A => regs(756), ZN => n2094);
   U782 : AOI22_X1 port map( A1 => n121, A2 => regs(2292), B1 => n64, B2 => 
                           regs(1780), ZN => n457);
   U783 : AOI22_X1 port map( A1 => n81, A2 => regs(1268), B1 => n29, B2 => 
                           regs(244), ZN => n456);
   U784 : OAI211_X1 port map( C1 => n10, C2 => n2094, A => n457, B => n456, ZN 
                           => curr_proc_regs(244));
   U785 : INV_X1 port map( A => regs(1269), ZN => n2097);
   U786 : AOI22_X1 port map( A1 => win(4), A2 => regs(2293), B1 => n73, B2 => 
                           regs(1781), ZN => n459);
   U787 : AOI22_X1 port map( A1 => n48, A2 => regs(757), B1 => n29, B2 => 
                           regs(245), ZN => n458);
   U788 : OAI211_X1 port map( C1 => n2215, C2 => n2097, A => n459, B => n458, 
                           ZN => curr_proc_regs(245));
   U789 : INV_X1 port map( A => regs(1270), ZN => n2100);
   U790 : AOI22_X1 port map( A1 => n119, A2 => regs(2294), B1 => n71, B2 => 
                           regs(1782), ZN => n461);
   U791 : AOI22_X1 port map( A1 => n50, A2 => regs(758), B1 => n29, B2 => 
                           regs(246), ZN => n460);
   U792 : OAI211_X1 port map( C1 => n103, C2 => n2100, A => n461, B => n460, ZN
                           => curr_proc_regs(246));
   U793 : INV_X1 port map( A => regs(759), ZN => n2103);
   U794 : AOI22_X1 port map( A1 => n120, A2 => regs(2295), B1 => n63, B2 => 
                           regs(1783), ZN => n463);
   U795 : AOI22_X1 port map( A1 => n86, A2 => regs(1271), B1 => n29, B2 => 
                           regs(247), ZN => n462);
   U796 : OAI211_X1 port map( C1 => n10, C2 => n2103, A => n463, B => n462, ZN 
                           => curr_proc_regs(247));
   U797 : INV_X1 port map( A => regs(760), ZN => n2109);
   U798 : AOI22_X1 port map( A1 => n121, A2 => regs(2296), B1 => n63, B2 => 
                           regs(1784), ZN => n465);
   U799 : AOI22_X1 port map( A1 => n87, A2 => regs(1272), B1 => n29, B2 => 
                           regs(248), ZN => n464);
   U800 : OAI211_X1 port map( C1 => n10, C2 => n2109, A => n465, B => n464, ZN 
                           => curr_proc_regs(248));
   U801 : INV_X1 port map( A => regs(761), ZN => n2112);
   U802 : AOI22_X1 port map( A1 => win(4), A2 => regs(2297), B1 => n60, B2 => 
                           regs(1785), ZN => n467);
   U803 : AOI22_X1 port map( A1 => n82, A2 => regs(1273), B1 => n29, B2 => 
                           regs(249), ZN => n466);
   U804 : OAI211_X1 port map( C1 => n10, C2 => n2112, A => n467, B => n466, ZN 
                           => curr_proc_regs(249));
   U805 : INV_X1 port map( A => regs(536), ZN => n1383);
   U806 : AOI22_X1 port map( A1 => n119, A2 => regs(2072), B1 => n64, B2 => 
                           regs(1560), ZN => n469);
   U807 : AOI22_X1 port map( A1 => n84, A2 => regs(1048), B1 => n29, B2 => 
                           regs(24), ZN => n468);
   U808 : OAI211_X1 port map( C1 => n10, C2 => n1383, A => n469, B => n468, ZN 
                           => curr_proc_regs(24));
   U809 : INV_X1 port map( A => regs(762), ZN => n2115);
   U810 : AOI22_X1 port map( A1 => n120, A2 => regs(2298), B1 => n68, B2 => 
                           regs(1786), ZN => n471);
   U811 : AOI22_X1 port map( A1 => n81, A2 => regs(1274), B1 => n29, B2 => 
                           regs(250), ZN => n470);
   U812 : OAI211_X1 port map( C1 => n10, C2 => n2115, A => n471, B => n470, ZN 
                           => curr_proc_regs(250));
   U813 : INV_X1 port map( A => regs(1275), ZN => n2118);
   U814 : AOI22_X1 port map( A1 => n121, A2 => regs(2299), B1 => n66, B2 => 
                           regs(1787), ZN => n473);
   U815 : AOI22_X1 port map( A1 => n52, A2 => regs(763), B1 => n31, B2 => 
                           regs(251), ZN => n472);
   U816 : OAI211_X1 port map( C1 => n11, C2 => n2118, A => n473, B => n472, ZN 
                           => curr_proc_regs(251));
   U817 : INV_X1 port map( A => regs(1276), ZN => n2121);
   U818 : AOI22_X1 port map( A1 => n121, A2 => regs(2300), B1 => n5, B2 => 
                           regs(1788), ZN => n475);
   U819 : AOI22_X1 port map( A1 => n48, A2 => regs(764), B1 => n31, B2 => 
                           regs(252), ZN => n474);
   U820 : OAI211_X1 port map( C1 => n2215, C2 => n2121, A => n475, B => n474, 
                           ZN => curr_proc_regs(252));
   U821 : INV_X1 port map( A => regs(765), ZN => n2124);
   U822 : AOI22_X1 port map( A1 => n121, A2 => regs(2301), B1 => n74, B2 => 
                           regs(1789), ZN => n477);
   U823 : AOI22_X1 port map( A1 => n80, A2 => regs(1277), B1 => n31, B2 => 
                           regs(253), ZN => n476);
   U824 : OAI211_X1 port map( C1 => n10, C2 => n2124, A => n477, B => n476, ZN 
                           => curr_proc_regs(253));
   U825 : INV_X1 port map( A => regs(766), ZN => n2127);
   U826 : AOI22_X1 port map( A1 => n121, A2 => regs(2302), B1 => n71, B2 => 
                           regs(1790), ZN => n479);
   U827 : AOI22_X1 port map( A1 => n85, A2 => regs(1278), B1 => n31, B2 => 
                           regs(254), ZN => n478);
   U828 : OAI211_X1 port map( C1 => n10, C2 => n2127, A => n479, B => n478, ZN 
                           => curr_proc_regs(254));
   U829 : INV_X1 port map( A => regs(1279), ZN => n2131);
   U830 : AOI22_X1 port map( A1 => n121, A2 => regs(2303), B1 => n5, B2 => 
                           regs(1791), ZN => n481);
   U831 : AOI22_X1 port map( A1 => n47, A2 => regs(767), B1 => n30, B2 => 
                           regs(255), ZN => n480);
   U832 : OAI211_X1 port map( C1 => n13, C2 => n2131, A => n481, B => n480, ZN 
                           => curr_proc_regs(255));
   U833 : NAND2_X1 port map( A1 => regs(768), A2 => n1, ZN => n484);
   U834 : AOI22_X1 port map( A1 => n86, A2 => regs(1280), B1 => n30, B2 => 
                           regs(256), ZN => n483);
   U835 : AOI22_X1 port map( A1 => n121, A2 => regs(2304), B1 => n72, B2 => 
                           regs(1792), ZN => n482);
   U836 : NAND3_X1 port map( A1 => n484, A2 => n483, A3 => n482, ZN => 
                           curr_proc_regs(256));
   U837 : NAND2_X1 port map( A1 => regs(1281), A2 => n90, ZN => n487);
   U838 : AOI22_X1 port map( A1 => n46, A2 => regs(769), B1 => n30, B2 => 
                           regs(257), ZN => n486);
   U839 : AOI22_X1 port map( A1 => n121, A2 => regs(2305), B1 => n69, B2 => 
                           regs(1793), ZN => n485);
   U840 : NAND3_X1 port map( A1 => n487, A2 => n486, A3 => n485, ZN => 
                           curr_proc_regs(257));
   U841 : NAND2_X1 port map( A1 => regs(1282), A2 => n89, ZN => n490);
   U842 : AOI22_X1 port map( A1 => n51, A2 => regs(770), B1 => n30, B2 => 
                           regs(258), ZN => n489);
   U843 : AOI22_X1 port map( A1 => n121, A2 => regs(2306), B1 => n74, B2 => 
                           regs(1794), ZN => n488);
   U844 : NAND3_X1 port map( A1 => n490, A2 => n489, A3 => n488, ZN => 
                           curr_proc_regs(258));
   U845 : NAND2_X1 port map( A1 => regs(1283), A2 => n89, ZN => n493);
   U846 : AOI22_X1 port map( A1 => n47, A2 => regs(771), B1 => n30, B2 => 
                           regs(259), ZN => n492);
   U847 : AOI22_X1 port map( A1 => n121, A2 => regs(2307), B1 => n71, B2 => 
                           regs(1795), ZN => n491);
   U848 : NAND3_X1 port map( A1 => n493, A2 => n492, A3 => n491, ZN => 
                           curr_proc_regs(259));
   U849 : INV_X1 port map( A => regs(1049), ZN => n1386);
   U850 : AOI22_X1 port map( A1 => n121, A2 => regs(2073), B1 => n5, B2 => 
                           regs(1561), ZN => n495);
   U851 : AOI22_X1 port map( A1 => n47, A2 => regs(537), B1 => n30, B2 => 
                           regs(25), ZN => n494);
   U852 : OAI211_X1 port map( C1 => n6, C2 => n1386, A => n495, B => n494, ZN 
                           => curr_proc_regs(25));
   U853 : NAND2_X1 port map( A1 => regs(1284), A2 => n89, ZN => n498);
   U854 : AOI22_X1 port map( A1 => n49, A2 => regs(772), B1 => n30, B2 => 
                           regs(260), ZN => n497);
   U855 : AOI22_X1 port map( A1 => n121, A2 => regs(2308), B1 => n63, B2 => 
                           regs(1796), ZN => n496);
   U856 : NAND3_X1 port map( A1 => n498, A2 => n497, A3 => n496, ZN => 
                           curr_proc_regs(260));
   U857 : NAND2_X1 port map( A1 => regs(1285), A2 => n90, ZN => n501);
   U858 : AOI22_X1 port map( A1 => n52, A2 => regs(773), B1 => n30, B2 => 
                           regs(261), ZN => n500);
   U859 : AOI22_X1 port map( A1 => n121, A2 => regs(2309), B1 => n63, B2 => 
                           regs(1797), ZN => n499);
   U860 : NAND3_X1 port map( A1 => n501, A2 => n500, A3 => n499, ZN => 
                           curr_proc_regs(261));
   U861 : NAND2_X1 port map( A1 => regs(1286), A2 => n89, ZN => n504);
   U862 : AOI22_X1 port map( A1 => n51, A2 => regs(774), B1 => n32, B2 => 
                           regs(262), ZN => n503);
   U863 : AOI22_X1 port map( A1 => n121, A2 => regs(2310), B1 => n72, B2 => 
                           regs(1798), ZN => n502);
   U864 : NAND3_X1 port map( A1 => n504, A2 => n503, A3 => n502, ZN => 
                           curr_proc_regs(262));
   U865 : NAND2_X1 port map( A1 => regs(775), A2 => n1, ZN => n507);
   U866 : AOI22_X1 port map( A1 => n87, A2 => regs(1287), B1 => n32, B2 => 
                           regs(263), ZN => n506);
   U867 : AOI22_X1 port map( A1 => win(4), A2 => regs(2311), B1 => n71, B2 => 
                           regs(1799), ZN => n505);
   U868 : NAND3_X1 port map( A1 => n507, A2 => n506, A3 => n505, ZN => 
                           curr_proc_regs(263));
   U869 : NAND2_X1 port map( A1 => regs(1288), A2 => n90, ZN => n510);
   U870 : AOI22_X1 port map( A1 => n50, A2 => regs(776), B1 => n32, B2 => 
                           regs(264), ZN => n509);
   U871 : AOI22_X1 port map( A1 => win(4), A2 => regs(2312), B1 => n68, B2 => 
                           regs(1800), ZN => n508);
   U872 : NAND3_X1 port map( A1 => n510, A2 => n509, A3 => n508, ZN => 
                           curr_proc_regs(264));
   U873 : NAND2_X1 port map( A1 => regs(1289), A2 => n90, ZN => n513);
   U874 : AOI22_X1 port map( A1 => n50, A2 => regs(777), B1 => n32, B2 => 
                           regs(265), ZN => n512);
   U875 : AOI22_X1 port map( A1 => win(4), A2 => regs(2313), B1 => n74, B2 => 
                           regs(1801), ZN => n511);
   U876 : NAND3_X1 port map( A1 => n513, A2 => n512, A3 => n511, ZN => 
                           curr_proc_regs(265));
   U877 : NAND2_X1 port map( A1 => regs(778), A2 => n8, ZN => n516);
   U878 : AOI22_X1 port map( A1 => n87, A2 => regs(1290), B1 => n31, B2 => 
                           regs(266), ZN => n515);
   U879 : AOI22_X1 port map( A1 => win(4), A2 => regs(2314), B1 => n65, B2 => 
                           regs(1802), ZN => n514);
   U880 : NAND3_X1 port map( A1 => n516, A2 => n515, A3 => n514, ZN => 
                           curr_proc_regs(266));
   U881 : NAND2_X1 port map( A1 => regs(779), A2 => n45, ZN => n519);
   U882 : AOI22_X1 port map( A1 => n87, A2 => regs(1291), B1 => n31, B2 => 
                           regs(267), ZN => n518);
   U883 : AOI22_X1 port map( A1 => win(4), A2 => regs(2315), B1 => n69, B2 => 
                           regs(1803), ZN => n517);
   U884 : NAND3_X1 port map( A1 => n519, A2 => n518, A3 => n517, ZN => 
                           curr_proc_regs(267));
   U885 : NAND2_X1 port map( A1 => regs(780), A2 => n1, ZN => n522);
   U886 : AOI22_X1 port map( A1 => n87, A2 => regs(1292), B1 => n31, B2 => 
                           regs(268), ZN => n521);
   U887 : AOI22_X1 port map( A1 => win(4), A2 => regs(2316), B1 => n71, B2 => 
                           regs(1804), ZN => n520);
   U888 : NAND3_X1 port map( A1 => n522, A2 => n521, A3 => n520, ZN => 
                           curr_proc_regs(268));
   U889 : NAND2_X1 port map( A1 => regs(781), A2 => n1, ZN => n525);
   U890 : AOI22_X1 port map( A1 => n87, A2 => regs(1293), B1 => n31, B2 => 
                           regs(269), ZN => n524);
   U891 : AOI22_X1 port map( A1 => win(4), A2 => regs(2317), B1 => n5, B2 => 
                           regs(1805), ZN => n523);
   U892 : NAND3_X1 port map( A1 => n525, A2 => n524, A3 => n523, ZN => 
                           curr_proc_regs(269));
   U893 : INV_X1 port map( A => regs(1050), ZN => n1389);
   U894 : AOI22_X1 port map( A1 => win(4), A2 => regs(2074), B1 => n74, B2 => 
                           regs(1562), ZN => n527);
   U895 : AOI22_X1 port map( A1 => n49, A2 => regs(538), B1 => n31, B2 => 
                           regs(26), ZN => n526);
   U896 : OAI211_X1 port map( C1 => n2215, C2 => n1389, A => n527, B => n526, 
                           ZN => curr_proc_regs(26));
   U897 : NAND2_X1 port map( A1 => regs(1294), A2 => n90, ZN => n530);
   U898 : AOI22_X1 port map( A1 => n51, A2 => regs(782), B1 => n31, B2 => 
                           regs(270), ZN => n529);
   U899 : AOI22_X1 port map( A1 => win(4), A2 => regs(2318), B1 => n66, B2 => 
                           regs(1806), ZN => n528);
   U900 : NAND3_X1 port map( A1 => n530, A2 => n529, A3 => n528, ZN => 
                           curr_proc_regs(270));
   U901 : NAND2_X1 port map( A1 => regs(1295), A2 => n90, ZN => n533);
   U902 : AOI22_X1 port map( A1 => n52, A2 => regs(783), B1 => n31, B2 => 
                           regs(271), ZN => n532);
   U903 : AOI22_X1 port map( A1 => win(4), A2 => regs(2319), B1 => n71, B2 => 
                           regs(1807), ZN => n531);
   U904 : NAND3_X1 port map( A1 => n533, A2 => n532, A3 => n531, ZN => 
                           curr_proc_regs(271));
   U905 : NAND2_X1 port map( A1 => regs(784), A2 => n1, ZN => n536);
   U906 : AOI22_X1 port map( A1 => n87, A2 => regs(1296), B1 => n31, B2 => 
                           regs(272), ZN => n535);
   U907 : AOI22_X1 port map( A1 => n7, A2 => regs(2320), B1 => n5, B2 => 
                           regs(1808), ZN => n534);
   U908 : NAND3_X1 port map( A1 => n536, A2 => n535, A3 => n534, ZN => 
                           curr_proc_regs(272));
   U909 : NAND2_X1 port map( A1 => regs(785), A2 => n1, ZN => n539);
   U910 : AOI22_X1 port map( A1 => n96, A2 => regs(1297), B1 => n4, B2 => 
                           regs(273), ZN => n538);
   U911 : AOI22_X1 port map( A1 => n7, A2 => regs(2321), B1 => n73, B2 => 
                           regs(1809), ZN => n537);
   U912 : NAND3_X1 port map( A1 => n539, A2 => n538, A3 => n537, ZN => 
                           curr_proc_regs(273));
   U913 : NAND2_X1 port map( A1 => regs(1298), A2 => n90, ZN => n542);
   U914 : AOI22_X1 port map( A1 => n51, A2 => regs(786), B1 => n4, B2 => 
                           regs(274), ZN => n541);
   U915 : AOI22_X1 port map( A1 => n131, A2 => regs(2322), B1 => n73, B2 => 
                           regs(1810), ZN => n540);
   U916 : NAND3_X1 port map( A1 => n542, A2 => n541, A3 => n540, ZN => 
                           curr_proc_regs(274));
   U917 : NAND2_X1 port map( A1 => regs(787), A2 => n1, ZN => n545);
   U918 : AOI22_X1 port map( A1 => n99, A2 => regs(1299), B1 => n4, B2 => 
                           regs(275), ZN => n544);
   U919 : AOI22_X1 port map( A1 => n131, A2 => regs(2323), B1 => n73, B2 => 
                           regs(1811), ZN => n543);
   U920 : NAND3_X1 port map( A1 => n545, A2 => n544, A3 => n543, ZN => 
                           curr_proc_regs(275));
   U921 : NAND2_X1 port map( A1 => regs(1300), A2 => n90, ZN => n548);
   U922 : AOI22_X1 port map( A1 => n50, A2 => regs(788), B1 => n4, B2 => 
                           regs(276), ZN => n547);
   U923 : AOI22_X1 port map( A1 => n131, A2 => regs(2324), B1 => n73, B2 => 
                           regs(1812), ZN => n546);
   U924 : NAND3_X1 port map( A1 => n548, A2 => n547, A3 => n546, ZN => 
                           curr_proc_regs(276));
   U925 : NAND2_X1 port map( A1 => regs(789), A2 => n1, ZN => n551);
   U926 : AOI22_X1 port map( A1 => n89, A2 => regs(1301), B1 => n32, B2 => 
                           regs(277), ZN => n550);
   U927 : AOI22_X1 port map( A1 => n131, A2 => regs(2325), B1 => n73, B2 => 
                           regs(1813), ZN => n549);
   U928 : NAND3_X1 port map( A1 => n551, A2 => n550, A3 => n549, ZN => 
                           curr_proc_regs(277));
   U929 : NAND2_X1 port map( A1 => regs(1302), A2 => n90, ZN => n554);
   U930 : AOI22_X1 port map( A1 => n41, A2 => regs(790), B1 => n32, B2 => 
                           regs(278), ZN => n553);
   U931 : AOI22_X1 port map( A1 => n131, A2 => regs(2326), B1 => n73, B2 => 
                           regs(1814), ZN => n552);
   U932 : NAND3_X1 port map( A1 => n554, A2 => n553, A3 => n552, ZN => 
                           curr_proc_regs(278));
   U933 : NAND2_X1 port map( A1 => regs(791), A2 => n1, ZN => n557);
   U934 : AOI22_X1 port map( A1 => n93, A2 => regs(1303), B1 => n32, B2 => 
                           regs(279), ZN => n556);
   U935 : AOI22_X1 port map( A1 => n131, A2 => regs(2327), B1 => n73, B2 => 
                           regs(1815), ZN => n555);
   U936 : NAND3_X1 port map( A1 => n557, A2 => n556, A3 => n555, ZN => 
                           curr_proc_regs(279));
   U937 : INV_X1 port map( A => regs(1051), ZN => n1392);
   U938 : AOI22_X1 port map( A1 => n131, A2 => regs(2075), B1 => n73, B2 => 
                           regs(1563), ZN => n559);
   U939 : AOI22_X1 port map( A1 => n48, A2 => regs(539), B1 => n32, B2 => 
                           regs(27), ZN => n558);
   U940 : OAI211_X1 port map( C1 => n103, C2 => n1392, A => n559, B => n558, ZN
                           => curr_proc_regs(27));
   U941 : NAND2_X1 port map( A1 => regs(792), A2 => n51, ZN => n562);
   U942 : AOI22_X1 port map( A1 => n99, A2 => regs(1304), B1 => n32, B2 => 
                           regs(280), ZN => n561);
   U943 : AOI22_X1 port map( A1 => n131, A2 => regs(2328), B1 => n73, B2 => 
                           regs(1816), ZN => n560);
   U944 : NAND3_X1 port map( A1 => n562, A2 => n561, A3 => n560, ZN => 
                           curr_proc_regs(280));
   U945 : NAND2_X1 port map( A1 => regs(793), A2 => n50, ZN => n565);
   U946 : AOI22_X1 port map( A1 => n86, A2 => regs(1305), B1 => n32, B2 => 
                           regs(281), ZN => n564);
   U947 : AOI22_X1 port map( A1 => n131, A2 => regs(2329), B1 => n73, B2 => 
                           regs(1817), ZN => n563);
   U948 : NAND3_X1 port map( A1 => n565, A2 => n564, A3 => n563, ZN => 
                           curr_proc_regs(281));
   U949 : NAND2_X1 port map( A1 => regs(1306), A2 => n90, ZN => n568);
   U950 : AOI22_X1 port map( A1 => n47, A2 => regs(794), B1 => n32, B2 => 
                           regs(282), ZN => n567);
   U951 : AOI22_X1 port map( A1 => n131, A2 => regs(2330), B1 => n73, B2 => 
                           regs(1818), ZN => n566);
   U952 : NAND3_X1 port map( A1 => n568, A2 => n567, A3 => n566, ZN => 
                           curr_proc_regs(282));
   U953 : NAND2_X1 port map( A1 => regs(1307), A2 => n90, ZN => n571);
   U954 : AOI22_X1 port map( A1 => n46, A2 => regs(795), B1 => n32, B2 => 
                           regs(283), ZN => n570);
   U955 : AOI22_X1 port map( A1 => n131, A2 => regs(2331), B1 => n73, B2 => 
                           regs(1819), ZN => n569);
   U956 : NAND3_X1 port map( A1 => n571, A2 => n570, A3 => n569, ZN => 
                           curr_proc_regs(283));
   U957 : NAND2_X1 port map( A1 => regs(1308), A2 => n90, ZN => n574);
   U958 : AOI22_X1 port map( A1 => n48, A2 => regs(796), B1 => n4, B2 => 
                           regs(284), ZN => n573);
   U959 : AOI22_X1 port map( A1 => n131, A2 => regs(2332), B1 => n73, B2 => 
                           regs(1820), ZN => n572);
   U960 : NAND3_X1 port map( A1 => n574, A2 => n573, A3 => n572, ZN => 
                           curr_proc_regs(284));
   U961 : NAND2_X1 port map( A1 => regs(797), A2 => n53, ZN => n577);
   U962 : AOI22_X1 port map( A1 => n86, A2 => regs(1309), B1 => n4, B2 => 
                           regs(285), ZN => n576);
   U963 : AOI22_X1 port map( A1 => n130, A2 => regs(2333), B1 => n73, B2 => 
                           regs(1821), ZN => n575);
   U964 : NAND3_X1 port map( A1 => n577, A2 => n576, A3 => n575, ZN => 
                           curr_proc_regs(285));
   U965 : NAND2_X1 port map( A1 => regs(798), A2 => n42, ZN => n580);
   U966 : AOI22_X1 port map( A1 => n86, A2 => regs(1310), B1 => n4, B2 => 
                           regs(286), ZN => n579);
   U967 : AOI22_X1 port map( A1 => n7, A2 => regs(2334), B1 => n73, B2 => 
                           regs(1822), ZN => n578);
   U968 : NAND3_X1 port map( A1 => n580, A2 => n579, A3 => n578, ZN => 
                           curr_proc_regs(286));
   U969 : NAND2_X1 port map( A1 => regs(1311), A2 => n91, ZN => n583);
   U970 : AOI22_X1 port map( A1 => n48, A2 => regs(799), B1 => n4, B2 => 
                           regs(287), ZN => n582);
   U971 : AOI22_X1 port map( A1 => n7, A2 => regs(2335), B1 => n73, B2 => 
                           regs(1823), ZN => n581);
   U972 : NAND3_X1 port map( A1 => n583, A2 => n582, A3 => n581, ZN => 
                           curr_proc_regs(287));
   U973 : NAND2_X1 port map( A1 => regs(800), A2 => n8, ZN => n586);
   U974 : AOI22_X1 port map( A1 => n86, A2 => regs(1312), B1 => n4, B2 => 
                           regs(288), ZN => n585);
   U975 : AOI22_X1 port map( A1 => n131, A2 => regs(2336), B1 => n73, B2 => 
                           regs(1824), ZN => n584);
   U976 : NAND3_X1 port map( A1 => n586, A2 => n585, A3 => n584, ZN => 
                           curr_proc_regs(288));
   U977 : NAND2_X1 port map( A1 => regs(801), A2 => n55, ZN => n589);
   U978 : AOI22_X1 port map( A1 => n100, A2 => regs(1313), B1 => n4, B2 => 
                           regs(289), ZN => n588);
   U979 : AOI22_X1 port map( A1 => n131, A2 => regs(2337), B1 => n73, B2 => 
                           regs(1825), ZN => n587);
   U980 : NAND3_X1 port map( A1 => n589, A2 => n588, A3 => n587, ZN => 
                           curr_proc_regs(289));
   U981 : INV_X1 port map( A => regs(540), ZN => n1397);
   U982 : AOI22_X1 port map( A1 => n130, A2 => regs(2076), B1 => n73, B2 => 
                           regs(1564), ZN => n591);
   U983 : AOI22_X1 port map( A1 => n86, A2 => regs(1052), B1 => n4, B2 => 
                           regs(28), ZN => n590);
   U984 : OAI211_X1 port map( C1 => n10, C2 => n1397, A => n591, B => n590, ZN 
                           => curr_proc_regs(28));
   U985 : NAND2_X1 port map( A1 => regs(802), A2 => n44, ZN => n594);
   U986 : AOI22_X1 port map( A1 => n86, A2 => regs(1314), B1 => n4, B2 => 
                           regs(290), ZN => n593);
   U987 : AOI22_X1 port map( A1 => n7, A2 => regs(2338), B1 => n73, B2 => 
                           regs(1826), ZN => n592);
   U988 : NAND3_X1 port map( A1 => n594, A2 => n593, A3 => n592, ZN => 
                           curr_proc_regs(290));
   U989 : NAND2_X1 port map( A1 => regs(803), A2 => n53, ZN => n597);
   U990 : AOI22_X1 port map( A1 => n86, A2 => regs(1315), B1 => n4, B2 => 
                           regs(291), ZN => n596);
   U991 : AOI22_X1 port map( A1 => n131, A2 => regs(2339), B1 => n73, B2 => 
                           regs(1827), ZN => n595);
   U992 : NAND3_X1 port map( A1 => n597, A2 => n596, A3 => n595, ZN => 
                           curr_proc_regs(291));
   U993 : NAND2_X1 port map( A1 => regs(804), A2 => n1, ZN => n600);
   U994 : AOI22_X1 port map( A1 => n86, A2 => regs(1316), B1 => n4, B2 => 
                           regs(292), ZN => n599);
   U995 : AOI22_X1 port map( A1 => n130, A2 => regs(2340), B1 => n73, B2 => 
                           regs(1828), ZN => n598);
   U996 : NAND3_X1 port map( A1 => n600, A2 => n599, A3 => n598, ZN => 
                           curr_proc_regs(292));
   U997 : NAND2_X1 port map( A1 => regs(1317), A2 => n97, ZN => n603);
   U998 : AOI22_X1 port map( A1 => n51, A2 => regs(805), B1 => n4, B2 => 
                           regs(293), ZN => n602);
   U999 : AOI22_X1 port map( A1 => n131, A2 => regs(2341), B1 => n73, B2 => 
                           regs(1829), ZN => n601);
   U1000 : NAND3_X1 port map( A1 => n603, A2 => n602, A3 => n601, ZN => 
                           curr_proc_regs(293));
   U1001 : NAND2_X1 port map( A1 => regs(806), A2 => n1, ZN => n606);
   U1002 : AOI22_X1 port map( A1 => n86, A2 => regs(1318), B1 => n4, B2 => 
                           regs(294), ZN => n605);
   U1003 : AOI22_X1 port map( A1 => n130, A2 => regs(2342), B1 => n73, B2 => 
                           regs(1830), ZN => n604);
   U1004 : NAND3_X1 port map( A1 => n606, A2 => n605, A3 => n604, ZN => 
                           curr_proc_regs(294));
   U1005 : NAND2_X1 port map( A1 => regs(1319), A2 => n97, ZN => n609);
   U1006 : AOI22_X1 port map( A1 => n50, A2 => regs(807), B1 => n33, B2 => 
                           regs(295), ZN => n608);
   U1007 : AOI22_X1 port map( A1 => n7, A2 => regs(2343), B1 => n73, B2 => 
                           regs(1831), ZN => n607);
   U1008 : NAND3_X1 port map( A1 => n609, A2 => n608, A3 => n607, ZN => 
                           curr_proc_regs(295));
   U1009 : NAND2_X1 port map( A1 => regs(808), A2 => n1, ZN => n612);
   U1010 : AOI22_X1 port map( A1 => n86, A2 => regs(1320), B1 => n33, B2 => 
                           regs(296), ZN => n611);
   U1011 : AOI22_X1 port map( A1 => n130, A2 => regs(2344), B1 => n2211, B2 => 
                           regs(1832), ZN => n610);
   U1012 : NAND3_X1 port map( A1 => n612, A2 => n611, A3 => n610, ZN => 
                           curr_proc_regs(296));
   U1013 : NAND2_X1 port map( A1 => regs(809), A2 => n1, ZN => n615);
   U1014 : AOI22_X1 port map( A1 => n97, A2 => regs(1321), B1 => n33, B2 => 
                           regs(297), ZN => n614);
   U1015 : AOI22_X1 port map( A1 => n7, A2 => regs(2345), B1 => n73, B2 => 
                           regs(1833), ZN => n613);
   U1016 : NAND3_X1 port map( A1 => n615, A2 => n614, A3 => n613, ZN => 
                           curr_proc_regs(297));
   U1017 : NAND2_X1 port map( A1 => regs(1322), A2 => n97, ZN => n618);
   U1018 : AOI22_X1 port map( A1 => n51, A2 => regs(810), B1 => n33, B2 => 
                           regs(298), ZN => n617);
   U1019 : AOI22_X1 port map( A1 => n7, A2 => regs(2346), B1 => n73, B2 => 
                           regs(1834), ZN => n616);
   U1020 : NAND3_X1 port map( A1 => n618, A2 => n617, A3 => n616, ZN => 
                           curr_proc_regs(298));
   U1021 : NAND2_X1 port map( A1 => regs(811), A2 => n1, ZN => n621);
   U1022 : AOI22_X1 port map( A1 => n90, A2 => regs(1323), B1 => n4, B2 => 
                           regs(299), ZN => n620);
   U1023 : AOI22_X1 port map( A1 => n131, A2 => regs(2347), B1 => n71, B2 => 
                           regs(1835), ZN => n619);
   U1024 : NAND3_X1 port map( A1 => n621, A2 => n620, A3 => n619, ZN => 
                           curr_proc_regs(299));
   U1025 : INV_X1 port map( A => regs(1053), ZN => n1400);
   U1026 : AOI22_X1 port map( A1 => n130, A2 => regs(2077), B1 => n73, B2 => 
                           regs(1565), ZN => n623);
   U1027 : AOI22_X1 port map( A1 => n50, A2 => regs(541), B1 => n4, B2 => 
                           regs(29), ZN => n622);
   U1028 : OAI211_X1 port map( C1 => n2215, C2 => n1400, A => n623, B => n622, 
                           ZN => curr_proc_regs(29));
   U1029 : INV_X1 port map( A => regs(514), ZN => n1316);
   U1030 : AOI22_X1 port map( A1 => n7, A2 => regs(2050), B1 => n73, B2 => 
                           regs(1538), ZN => n625);
   U1031 : AOI22_X1 port map( A1 => n83, A2 => regs(1026), B1 => n4, B2 => 
                           regs(2), ZN => n624);
   U1032 : OAI211_X1 port map( C1 => n10, C2 => n1316, A => n625, B => n624, ZN
                           => curr_proc_regs(2));
   U1033 : NAND2_X1 port map( A1 => regs(812), A2 => n1, ZN => n628);
   U1034 : AOI22_X1 port map( A1 => n90, A2 => regs(1324), B1 => n4, B2 => 
                           regs(300), ZN => n627);
   U1035 : AOI22_X1 port map( A1 => n131, A2 => regs(2348), B1 => n69, B2 => 
                           regs(1836), ZN => n626);
   U1036 : NAND3_X1 port map( A1 => n628, A2 => n627, A3 => n626, ZN => 
                           curr_proc_regs(300));
   U1037 : NAND2_X1 port map( A1 => regs(813), A2 => n1, ZN => n631);
   U1038 : AOI22_X1 port map( A1 => n93, A2 => regs(1325), B1 => n4, B2 => 
                           regs(301), ZN => n630);
   U1039 : AOI22_X1 port map( A1 => n131, A2 => regs(2349), B1 => n73, B2 => 
                           regs(1837), ZN => n629);
   U1040 : NAND3_X1 port map( A1 => n631, A2 => n630, A3 => n629, ZN => 
                           curr_proc_regs(301));
   U1041 : NAND2_X1 port map( A1 => regs(814), A2 => n1, ZN => n634);
   U1042 : AOI22_X1 port map( A1 => n97, A2 => regs(1326), B1 => n4, B2 => 
                           regs(302), ZN => n633);
   U1043 : AOI22_X1 port map( A1 => n130, A2 => regs(2350), B1 => n73, B2 => 
                           regs(1838), ZN => n632);
   U1044 : NAND3_X1 port map( A1 => n634, A2 => n633, A3 => n632, ZN => 
                           curr_proc_regs(302));
   U1045 : NAND2_X1 port map( A1 => regs(815), A2 => n1, ZN => n637);
   U1046 : AOI22_X1 port map( A1 => n99, A2 => regs(1327), B1 => n4, B2 => 
                           regs(303), ZN => n636);
   U1047 : AOI22_X1 port map( A1 => n7, A2 => regs(2351), B1 => n72, B2 => 
                           regs(1839), ZN => n635);
   U1048 : NAND3_X1 port map( A1 => n637, A2 => n636, A3 => n635, ZN => 
                           curr_proc_regs(303));
   U1049 : NAND2_X1 port map( A1 => regs(1328), A2 => n97, ZN => n640);
   U1050 : AOI22_X1 port map( A1 => n49, A2 => regs(816), B1 => n4, B2 => 
                           regs(304), ZN => n639);
   U1051 : AOI22_X1 port map( A1 => n130, A2 => regs(2352), B1 => n73, B2 => 
                           regs(1840), ZN => n638);
   U1052 : NAND3_X1 port map( A1 => n640, A2 => n639, A3 => n638, ZN => 
                           curr_proc_regs(304));
   U1053 : NAND2_X1 port map( A1 => regs(817), A2 => n1, ZN => n643);
   U1054 : AOI22_X1 port map( A1 => n87, A2 => regs(1329), B1 => n34, B2 => 
                           regs(305), ZN => n642);
   U1055 : AOI22_X1 port map( A1 => n131, A2 => regs(2353), B1 => n73, B2 => 
                           regs(1841), ZN => n641);
   U1056 : NAND3_X1 port map( A1 => n643, A2 => n642, A3 => n641, ZN => 
                           curr_proc_regs(305));
   U1057 : NAND2_X1 port map( A1 => regs(1330), A2 => n97, ZN => n646);
   U1058 : AOI22_X1 port map( A1 => n48, A2 => regs(818), B1 => n34, B2 => 
                           regs(306), ZN => n645);
   U1059 : AOI22_X1 port map( A1 => n130, A2 => regs(2354), B1 => n73, B2 => 
                           regs(1842), ZN => n644);
   U1060 : NAND3_X1 port map( A1 => n646, A2 => n645, A3 => n644, ZN => 
                           curr_proc_regs(306));
   U1061 : NAND2_X1 port map( A1 => regs(1331), A2 => n97, ZN => n649);
   U1062 : AOI22_X1 port map( A1 => n47, A2 => regs(819), B1 => n34, B2 => 
                           regs(307), ZN => n648);
   U1063 : AOI22_X1 port map( A1 => n7, A2 => regs(2355), B1 => n74, B2 => 
                           regs(1843), ZN => n647);
   U1064 : NAND3_X1 port map( A1 => n649, A2 => n648, A3 => n647, ZN => 
                           curr_proc_regs(307));
   U1065 : NAND2_X1 port map( A1 => regs(820), A2 => n45, ZN => n652);
   U1066 : AOI22_X1 port map( A1 => n87, A2 => regs(1332), B1 => n34, B2 => 
                           regs(308), ZN => n651);
   U1067 : AOI22_X1 port map( A1 => n131, A2 => regs(2356), B1 => n73, B2 => 
                           regs(1844), ZN => n650);
   U1068 : NAND3_X1 port map( A1 => n652, A2 => n651, A3 => n650, ZN => 
                           curr_proc_regs(308));
   U1069 : NAND2_X1 port map( A1 => regs(821), A2 => n41, ZN => n655);
   U1070 : AOI22_X1 port map( A1 => n87, A2 => regs(1333), B1 => n33, B2 => 
                           regs(309), ZN => n654);
   U1071 : AOI22_X1 port map( A1 => n130, A2 => regs(2357), B1 => n73, B2 => 
                           regs(1845), ZN => n653);
   U1072 : NAND3_X1 port map( A1 => n655, A2 => n654, A3 => n653, ZN => 
                           curr_proc_regs(309));
   U1073 : INV_X1 port map( A => regs(1054), ZN => n1403);
   U1074 : AOI22_X1 port map( A1 => n7, A2 => regs(2078), B1 => n73, B2 => 
                           regs(1566), ZN => n657);
   U1075 : AOI22_X1 port map( A1 => n46, A2 => regs(542), B1 => n33, B2 => 
                           regs(30), ZN => n656);
   U1076 : OAI211_X1 port map( C1 => n11, C2 => n1403, A => n657, B => n656, ZN
                           => curr_proc_regs(30));
   U1077 : NAND2_X1 port map( A1 => regs(822), A2 => n56, ZN => n660);
   U1078 : AOI22_X1 port map( A1 => n87, A2 => regs(1334), B1 => n33, B2 => 
                           regs(310), ZN => n659);
   U1079 : AOI22_X1 port map( A1 => n131, A2 => regs(2358), B1 => n71, B2 => 
                           regs(1846), ZN => n658);
   U1080 : NAND3_X1 port map( A1 => n660, A2 => n659, A3 => n658, ZN => 
                           curr_proc_regs(310));
   U1081 : NAND2_X1 port map( A1 => regs(823), A2 => n3, ZN => n663);
   U1082 : AOI22_X1 port map( A1 => n87, A2 => regs(1335), B1 => n33, B2 => 
                           regs(311), ZN => n662);
   U1083 : AOI22_X1 port map( A1 => n130, A2 => regs(2359), B1 => n5, B2 => 
                           regs(1847), ZN => n661);
   U1084 : NAND3_X1 port map( A1 => n663, A2 => n662, A3 => n661, ZN => 
                           curr_proc_regs(311));
   U1085 : NAND2_X1 port map( A1 => regs(824), A2 => n8, ZN => n666);
   U1086 : AOI22_X1 port map( A1 => n87, A2 => regs(1336), B1 => n33, B2 => 
                           regs(312), ZN => n665);
   U1087 : AOI22_X1 port map( A1 => n7, A2 => regs(2360), B1 => n73, B2 => 
                           regs(1848), ZN => n664);
   U1088 : NAND3_X1 port map( A1 => n666, A2 => n665, A3 => n664, ZN => 
                           curr_proc_regs(312));
   U1089 : NAND2_X1 port map( A1 => regs(1337), A2 => n96, ZN => n669);
   U1090 : AOI22_X1 port map( A1 => n49, A2 => regs(825), B1 => n33, B2 => 
                           regs(313), ZN => n668);
   U1091 : AOI22_X1 port map( A1 => n131, A2 => regs(2361), B1 => n73, B2 => 
                           regs(1849), ZN => n667);
   U1092 : NAND3_X1 port map( A1 => n669, A2 => n668, A3 => n667, ZN => 
                           curr_proc_regs(313));
   U1093 : NAND2_X1 port map( A1 => regs(826), A2 => n41, ZN => n672);
   U1094 : AOI22_X1 port map( A1 => n87, A2 => regs(1338), B1 => n33, B2 => 
                           regs(314), ZN => n671);
   U1095 : AOI22_X1 port map( A1 => n130, A2 => regs(2362), B1 => n68, B2 => 
                           regs(1850), ZN => n670);
   U1096 : NAND3_X1 port map( A1 => n672, A2 => n671, A3 => n670, ZN => 
                           curr_proc_regs(314));
   U1097 : NAND2_X1 port map( A1 => regs(1339), A2 => n95, ZN => n675);
   U1098 : AOI22_X1 port map( A1 => n52, A2 => regs(827), B1 => n33, B2 => 
                           regs(315), ZN => n674);
   U1099 : AOI22_X1 port map( A1 => n7, A2 => regs(2363), B1 => n73, B2 => 
                           regs(1851), ZN => n673);
   U1100 : NAND3_X1 port map( A1 => n675, A2 => n674, A3 => n673, ZN => 
                           curr_proc_regs(315));
   U1101 : NAND2_X1 port map( A1 => regs(1340), A2 => n94, ZN => n678);
   U1102 : AOI22_X1 port map( A1 => n52, A2 => regs(828), B1 => n35, B2 => 
                           regs(316), ZN => n677);
   U1103 : AOI22_X1 port map( A1 => n131, A2 => regs(2364), B1 => n61, B2 => 
                           regs(1852), ZN => n676);
   U1104 : NAND3_X1 port map( A1 => n678, A2 => n677, A3 => n676, ZN => 
                           curr_proc_regs(316));
   U1105 : NAND2_X1 port map( A1 => regs(1341), A2 => n94, ZN => n681);
   U1106 : AOI22_X1 port map( A1 => n51, A2 => regs(829), B1 => n35, B2 => 
                           regs(317), ZN => n680);
   U1107 : AOI22_X1 port map( A1 => n130, A2 => regs(2365), B1 => n73, B2 => 
                           regs(1853), ZN => n679);
   U1108 : NAND3_X1 port map( A1 => n681, A2 => n680, A3 => n679, ZN => 
                           curr_proc_regs(317));
   U1109 : NAND2_X1 port map( A1 => regs(1342), A2 => n94, ZN => n684);
   U1110 : AOI22_X1 port map( A1 => n3, A2 => regs(830), B1 => n35, B2 => 
                           regs(318), ZN => n683);
   U1111 : AOI22_X1 port map( A1 => n7, A2 => regs(2366), B1 => n73, B2 => 
                           regs(1854), ZN => n682);
   U1112 : NAND3_X1 port map( A1 => n684, A2 => n683, A3 => n682, ZN => 
                           curr_proc_regs(318));
   U1113 : NAND2_X1 port map( A1 => regs(831), A2 => n54, ZN => n687);
   U1114 : AOI22_X1 port map( A1 => n85, A2 => regs(1343), B1 => n35, B2 => 
                           regs(319), ZN => n686);
   U1115 : AOI22_X1 port map( A1 => n7, A2 => regs(2367), B1 => n73, B2 => 
                           regs(1855), ZN => n685);
   U1116 : NAND3_X1 port map( A1 => n687, A2 => n686, A3 => n685, ZN => 
                           curr_proc_regs(319));
   U1117 : INV_X1 port map( A => regs(543), ZN => n1406);
   U1118 : AOI22_X1 port map( A1 => n7, A2 => regs(2079), B1 => n73, B2 => 
                           regs(1567), ZN => n689);
   U1119 : AOI22_X1 port map( A1 => n80, A2 => regs(1055), B1 => n34, B2 => 
                           regs(31), ZN => n688);
   U1120 : OAI211_X1 port map( C1 => n10, C2 => n1406, A => n689, B => n688, ZN
                           => curr_proc_regs(31));
   U1121 : NAND2_X1 port map( A1 => regs(1344), A2 => n94, ZN => n692);
   U1122 : AOI22_X1 port map( A1 => n44, A2 => regs(832), B1 => n34, B2 => 
                           regs(320), ZN => n691);
   U1123 : AOI22_X1 port map( A1 => n7, A2 => regs(2368), B1 => n74, B2 => 
                           regs(1856), ZN => n690);
   U1124 : NAND3_X1 port map( A1 => n692, A2 => n691, A3 => n690, ZN => 
                           curr_proc_regs(320));
   U1125 : NAND2_X1 port map( A1 => regs(1345), A2 => n94, ZN => n695);
   U1126 : AOI22_X1 port map( A1 => n43, A2 => regs(833), B1 => n34, B2 => 
                           regs(321), ZN => n694);
   U1127 : AOI22_X1 port map( A1 => n7, A2 => regs(2369), B1 => n73, B2 => 
                           regs(1857), ZN => n693);
   U1128 : NAND3_X1 port map( A1 => n695, A2 => n694, A3 => n693, ZN => 
                           curr_proc_regs(321));
   U1129 : NAND2_X1 port map( A1 => regs(834), A2 => n54, ZN => n698);
   U1130 : AOI22_X1 port map( A1 => n83, A2 => regs(1346), B1 => n34, B2 => 
                           regs(322), ZN => n697);
   U1131 : AOI22_X1 port map( A1 => n7, A2 => regs(2370), B1 => n66, B2 => 
                           regs(1858), ZN => n696);
   U1132 : NAND3_X1 port map( A1 => n698, A2 => n697, A3 => n696, ZN => 
                           curr_proc_regs(322));
   U1133 : NAND2_X1 port map( A1 => regs(835), A2 => n53, ZN => n701);
   U1134 : AOI22_X1 port map( A1 => n93, A2 => regs(1347), B1 => n34, B2 => 
                           regs(323), ZN => n700);
   U1135 : AOI22_X1 port map( A1 => n7, A2 => regs(2371), B1 => n73, B2 => 
                           regs(1859), ZN => n699);
   U1136 : NAND3_X1 port map( A1 => n701, A2 => n700, A3 => n699, ZN => 
                           curr_proc_regs(323));
   U1137 : NAND2_X1 port map( A1 => regs(1348), A2 => n93, ZN => n704);
   U1138 : AOI22_X1 port map( A1 => n54, A2 => regs(836), B1 => n34, B2 => 
                           regs(324), ZN => n703);
   U1139 : AOI22_X1 port map( A1 => n127, A2 => regs(2372), B1 => n73, B2 => 
                           regs(1860), ZN => n702);
   U1140 : NAND3_X1 port map( A1 => n704, A2 => n703, A3 => n702, ZN => 
                           curr_proc_regs(324));
   U1141 : NAND2_X1 port map( A1 => regs(837), A2 => n45, ZN => n707);
   U1142 : AOI22_X1 port map( A1 => n90, A2 => regs(1349), B1 => n34, B2 => 
                           regs(325), ZN => n706);
   U1143 : AOI22_X1 port map( A1 => n7, A2 => regs(2373), B1 => n66, B2 => 
                           regs(1861), ZN => n705);
   U1144 : NAND3_X1 port map( A1 => n707, A2 => n706, A3 => n705, ZN => 
                           curr_proc_regs(325));
   U1145 : NAND2_X1 port map( A1 => regs(838), A2 => n56, ZN => n710);
   U1146 : AOI22_X1 port map( A1 => n99, A2 => regs(1350), B1 => n34, B2 => 
                           regs(326), ZN => n709);
   U1147 : AOI22_X1 port map( A1 => n7, A2 => regs(2374), B1 => n5, B2 => 
                           regs(1862), ZN => n708);
   U1148 : NAND3_X1 port map( A1 => n710, A2 => n709, A3 => n708, ZN => 
                           curr_proc_regs(326));
   U1149 : NAND2_X1 port map( A1 => regs(1351), A2 => n93, ZN => n713);
   U1150 : AOI22_X1 port map( A1 => n53, A2 => regs(839), B1 => n36, B2 => 
                           regs(327), ZN => n712);
   U1151 : AOI22_X1 port map( A1 => n7, A2 => regs(2375), B1 => n63, B2 => 
                           regs(1863), ZN => n711);
   U1152 : NAND3_X1 port map( A1 => n713, A2 => n712, A3 => n711, ZN => 
                           curr_proc_regs(327));
   U1153 : NAND2_X1 port map( A1 => regs(1352), A2 => n93, ZN => n716);
   U1154 : AOI22_X1 port map( A1 => n55, A2 => regs(840), B1 => n36, B2 => 
                           regs(328), ZN => n715);
   U1155 : AOI22_X1 port map( A1 => n7, A2 => regs(2376), B1 => n68, B2 => 
                           regs(1864), ZN => n714);
   U1156 : NAND3_X1 port map( A1 => n716, A2 => n715, A3 => n714, ZN => 
                           curr_proc_regs(328));
   U1157 : NAND2_X1 port map( A1 => regs(841), A2 => n41, ZN => n719);
   U1158 : AOI22_X1 port map( A1 => n91, A2 => regs(1353), B1 => n36, B2 => 
                           regs(329), ZN => n718);
   U1159 : AOI22_X1 port map( A1 => n130, A2 => regs(2377), B1 => n68, B2 => 
                           regs(1865), ZN => n717);
   U1160 : NAND3_X1 port map( A1 => n719, A2 => n718, A3 => n717, ZN => 
                           curr_proc_regs(329));
   U1161 : INV_X1 port map( A => regs(544), ZN => n1409);
   U1162 : AOI22_X1 port map( A1 => n130, A2 => regs(2080), B1 => n70, B2 => 
                           regs(1568), ZN => n721);
   U1163 : AOI22_X1 port map( A1 => n96, A2 => regs(1056), B1 => n36, B2 => 
                           regs(32), ZN => n720);
   U1164 : OAI211_X1 port map( C1 => n58, C2 => n1409, A => n721, B => n720, ZN
                           => curr_proc_regs(32));
   U1165 : NAND2_X1 port map( A1 => regs(1354), A2 => n94, ZN => n724);
   U1166 : AOI22_X1 port map( A1 => n52, A2 => regs(842), B1 => n35, B2 => 
                           regs(330), ZN => n723);
   U1167 : AOI22_X1 port map( A1 => n130, A2 => regs(2378), B1 => n73, B2 => 
                           regs(1866), ZN => n722);
   U1168 : NAND3_X1 port map( A1 => n724, A2 => n723, A3 => n722, ZN => 
                           curr_proc_regs(330));
   U1169 : NAND2_X1 port map( A1 => regs(843), A2 => n56, ZN => n727);
   U1170 : AOI22_X1 port map( A1 => n89, A2 => regs(1355), B1 => n35, B2 => 
                           regs(331), ZN => n726);
   U1171 : AOI22_X1 port map( A1 => n130, A2 => regs(2379), B1 => n73, B2 => 
                           regs(1867), ZN => n725);
   U1172 : NAND3_X1 port map( A1 => n727, A2 => n726, A3 => n725, ZN => 
                           curr_proc_regs(331));
   U1173 : NAND2_X1 port map( A1 => regs(1356), A2 => n91, ZN => n730);
   U1174 : AOI22_X1 port map( A1 => n50, A2 => regs(844), B1 => n35, B2 => 
                           regs(332), ZN => n729);
   U1175 : AOI22_X1 port map( A1 => n130, A2 => regs(2380), B1 => n74, B2 => 
                           regs(1868), ZN => n728);
   U1176 : NAND3_X1 port map( A1 => n730, A2 => n729, A3 => n728, ZN => 
                           curr_proc_regs(332));
   U1177 : NAND2_X1 port map( A1 => regs(845), A2 => n42, ZN => n733);
   U1178 : AOI22_X1 port map( A1 => n92, A2 => regs(1357), B1 => n35, B2 => 
                           regs(333), ZN => n732);
   U1179 : AOI22_X1 port map( A1 => n130, A2 => regs(2381), B1 => n65, B2 => 
                           regs(1869), ZN => n731);
   U1180 : NAND3_X1 port map( A1 => n733, A2 => n732, A3 => n731, ZN => 
                           curr_proc_regs(333));
   U1181 : NAND2_X1 port map( A1 => regs(846), A2 => n3, ZN => n736);
   U1182 : AOI22_X1 port map( A1 => n91, A2 => regs(1358), B1 => n35, B2 => 
                           regs(334), ZN => n735);
   U1183 : AOI22_X1 port map( A1 => n130, A2 => regs(2382), B1 => n69, B2 => 
                           regs(1870), ZN => n734);
   U1184 : NAND3_X1 port map( A1 => n736, A2 => n735, A3 => n734, ZN => 
                           curr_proc_regs(334));
   U1185 : NAND2_X1 port map( A1 => regs(847), A2 => n44, ZN => n739);
   U1186 : AOI22_X1 port map( A1 => n98, A2 => regs(1359), B1 => n35, B2 => 
                           regs(335), ZN => n738);
   U1187 : AOI22_X1 port map( A1 => n130, A2 => regs(2383), B1 => n67, B2 => 
                           regs(1871), ZN => n737);
   U1188 : NAND3_X1 port map( A1 => n739, A2 => n738, A3 => n737, ZN => 
                           curr_proc_regs(335));
   U1189 : NAND2_X1 port map( A1 => regs(1360), A2 => n94, ZN => n742);
   U1190 : AOI22_X1 port map( A1 => n50, A2 => regs(848), B1 => n35, B2 => 
                           regs(336), ZN => n741);
   U1191 : AOI22_X1 port map( A1 => n130, A2 => regs(2384), B1 => n72, B2 => 
                           regs(1872), ZN => n740);
   U1192 : NAND3_X1 port map( A1 => n742, A2 => n741, A3 => n740, ZN => 
                           curr_proc_regs(336));
   U1193 : NAND2_X1 port map( A1 => regs(849), A2 => n42, ZN => n745);
   U1194 : AOI22_X1 port map( A1 => n98, A2 => regs(1361), B1 => n35, B2 => 
                           regs(337), ZN => n744);
   U1195 : AOI22_X1 port map( A1 => n130, A2 => regs(2385), B1 => n75, B2 => 
                           regs(1873), ZN => n743);
   U1196 : NAND3_X1 port map( A1 => n745, A2 => n744, A3 => n743, ZN => 
                           curr_proc_regs(337));
   U1197 : NAND2_X1 port map( A1 => regs(1362), A2 => n92, ZN => n748);
   U1198 : AOI22_X1 port map( A1 => n47, A2 => regs(850), B1 => n37, B2 => 
                           regs(338), ZN => n747);
   U1199 : AOI22_X1 port map( A1 => n130, A2 => regs(2386), B1 => n60, B2 => 
                           regs(1874), ZN => n746);
   U1200 : NAND3_X1 port map( A1 => n748, A2 => n747, A3 => n746, ZN => 
                           curr_proc_regs(338));
   U1201 : NAND2_X1 port map( A1 => regs(1363), A2 => n92, ZN => n751);
   U1202 : AOI22_X1 port map( A1 => n49, A2 => regs(851), B1 => n37, B2 => 
                           regs(339), ZN => n750);
   U1203 : AOI22_X1 port map( A1 => n130, A2 => regs(2387), B1 => n64, B2 => 
                           regs(1875), ZN => n749);
   U1204 : NAND3_X1 port map( A1 => n751, A2 => n750, A3 => n749, ZN => 
                           curr_proc_regs(339));
   U1205 : INV_X1 port map( A => regs(1057), ZN => n1412);
   U1206 : AOI22_X1 port map( A1 => n129, A2 => regs(2081), B1 => n73, B2 => 
                           regs(1569), ZN => n753);
   U1207 : AOI22_X1 port map( A1 => n46, A2 => regs(545), B1 => n37, B2 => 
                           regs(33), ZN => n752);
   U1208 : OAI211_X1 port map( C1 => n13, C2 => n1412, A => n753, B => n752, ZN
                           => curr_proc_regs(33));
   U1209 : NAND2_X1 port map( A1 => regs(1364), A2 => n92, ZN => n756);
   U1210 : AOI22_X1 port map( A1 => n49, A2 => regs(852), B1 => n37, B2 => 
                           regs(340), ZN => n755);
   U1211 : AOI22_X1 port map( A1 => n126, A2 => regs(2388), B1 => n60, B2 => 
                           regs(1876), ZN => n754);
   U1212 : NAND3_X1 port map( A1 => n756, A2 => n755, A3 => n754, ZN => 
                           curr_proc_regs(340));
   U1213 : NAND2_X1 port map( A1 => regs(1365), A2 => n92, ZN => n759);
   U1214 : AOI22_X1 port map( A1 => n50, A2 => regs(853), B1 => n36, B2 => 
                           regs(341), ZN => n758);
   U1215 : AOI22_X1 port map( A1 => n129, A2 => regs(2389), B1 => n64, B2 => 
                           regs(1877), ZN => n757);
   U1216 : NAND3_X1 port map( A1 => n759, A2 => n758, A3 => n757, ZN => 
                           curr_proc_regs(341));
   U1217 : NAND2_X1 port map( A1 => regs(1366), A2 => n91, ZN => n762);
   U1218 : AOI22_X1 port map( A1 => n51, A2 => regs(854), B1 => n36, B2 => 
                           regs(342), ZN => n761);
   U1219 : AOI22_X1 port map( A1 => n128, A2 => regs(2390), B1 => n63, B2 => 
                           regs(1878), ZN => n760);
   U1220 : NAND3_X1 port map( A1 => n762, A2 => n761, A3 => n760, ZN => 
                           curr_proc_regs(342));
   U1221 : NAND2_X1 port map( A1 => regs(855), A2 => n43, ZN => n765);
   U1222 : AOI22_X1 port map( A1 => n92, A2 => regs(1367), B1 => n36, B2 => 
                           regs(343), ZN => n764);
   U1223 : AOI22_X1 port map( A1 => n129, A2 => regs(2391), B1 => n60, B2 => 
                           regs(1879), ZN => n763);
   U1224 : NAND3_X1 port map( A1 => n765, A2 => n764, A3 => n763, ZN => 
                           curr_proc_regs(343));
   U1225 : NAND2_X1 port map( A1 => regs(856), A2 => n49, ZN => n768);
   U1226 : AOI22_X1 port map( A1 => n91, A2 => regs(1368), B1 => n36, B2 => 
                           regs(344), ZN => n767);
   U1227 : AOI22_X1 port map( A1 => n129, A2 => regs(2392), B1 => n60, B2 => 
                           regs(1880), ZN => n766);
   U1228 : NAND3_X1 port map( A1 => n768, A2 => n767, A3 => n766, ZN => 
                           curr_proc_regs(344));
   U1229 : NAND2_X1 port map( A1 => regs(1369), A2 => n95, ZN => n771);
   U1230 : AOI22_X1 port map( A1 => n49, A2 => regs(857), B1 => n36, B2 => 
                           regs(345), ZN => n770);
   U1231 : AOI22_X1 port map( A1 => n129, A2 => regs(2393), B1 => n64, B2 => 
                           regs(1881), ZN => n769);
   U1232 : NAND3_X1 port map( A1 => n771, A2 => n770, A3 => n769, ZN => 
                           curr_proc_regs(345));
   U1233 : NAND2_X1 port map( A1 => regs(1370), A2 => n91, ZN => n774);
   U1234 : AOI22_X1 port map( A1 => n46, A2 => regs(858), B1 => n36, B2 => 
                           regs(346), ZN => n773);
   U1235 : AOI22_X1 port map( A1 => n126, A2 => regs(2394), B1 => n74, B2 => 
                           regs(1882), ZN => n772);
   U1236 : NAND3_X1 port map( A1 => n774, A2 => n773, A3 => n772, ZN => 
                           curr_proc_regs(346));
   U1237 : NAND2_X1 port map( A1 => regs(859), A2 => n1, ZN => n777);
   U1238 : AOI22_X1 port map( A1 => n100, A2 => regs(1371), B1 => n36, B2 => 
                           regs(347), ZN => n776);
   U1239 : AOI22_X1 port map( A1 => n127, A2 => regs(2395), B1 => n63, B2 => 
                           regs(1883), ZN => n775);
   U1240 : NAND3_X1 port map( A1 => n777, A2 => n776, A3 => n775, ZN => 
                           curr_proc_regs(347));
   U1241 : NAND2_X1 port map( A1 => regs(860), A2 => n1, ZN => n780);
   U1242 : AOI22_X1 port map( A1 => n95, A2 => regs(1372), B1 => n36, B2 => 
                           regs(348), ZN => n779);
   U1243 : AOI22_X1 port map( A1 => n128, A2 => regs(2396), B1 => n71, B2 => 
                           regs(1884), ZN => n778);
   U1244 : NAND3_X1 port map( A1 => n780, A2 => n779, A3 => n778, ZN => 
                           curr_proc_regs(348));
   U1245 : NAND2_X1 port map( A1 => regs(861), A2 => n1, ZN => n783);
   U1246 : AOI22_X1 port map( A1 => n94, A2 => regs(1373), B1 => n38, B2 => 
                           regs(349), ZN => n782);
   U1247 : AOI22_X1 port map( A1 => n126, A2 => regs(2397), B1 => n64, B2 => 
                           regs(1885), ZN => n781);
   U1248 : NAND3_X1 port map( A1 => n783, A2 => n782, A3 => n781, ZN => 
                           curr_proc_regs(349));
   U1249 : INV_X1 port map( A => regs(546), ZN => n1415);
   U1250 : AOI22_X1 port map( A1 => n126, A2 => regs(2082), B1 => n64, B2 => 
                           regs(1570), ZN => n785);
   U1251 : AOI22_X1 port map( A1 => n89, A2 => regs(1058), B1 => n38, B2 => 
                           regs(34), ZN => n784);
   U1252 : OAI211_X1 port map( C1 => n58, C2 => n1415, A => n785, B => n784, ZN
                           => curr_proc_regs(34));
   U1253 : NAND2_X1 port map( A1 => regs(862), A2 => n8, ZN => n788);
   U1254 : AOI22_X1 port map( A1 => n92, A2 => regs(1374), B1 => n38, B2 => 
                           regs(350), ZN => n787);
   U1255 : AOI22_X1 port map( A1 => n129, A2 => regs(2398), B1 => n64, B2 => 
                           regs(1886), ZN => n786);
   U1256 : NAND3_X1 port map( A1 => n788, A2 => n787, A3 => n786, ZN => 
                           curr_proc_regs(350));
   U1257 : NAND2_X1 port map( A1 => regs(863), A2 => n3, ZN => n791);
   U1258 : AOI22_X1 port map( A1 => n96, A2 => regs(1375), B1 => n38, B2 => 
                           regs(351), ZN => n790);
   U1259 : AOI22_X1 port map( A1 => n129, A2 => regs(2399), B1 => n64, B2 => 
                           regs(1887), ZN => n789);
   U1260 : NAND3_X1 port map( A1 => n791, A2 => n790, A3 => n789, ZN => 
                           curr_proc_regs(351));
   U1261 : NAND2_X1 port map( A1 => regs(864), A2 => n42, ZN => n794);
   U1262 : AOI22_X1 port map( A1 => n98, A2 => regs(1376), B1 => n37, B2 => 
                           regs(352), ZN => n793);
   U1263 : AOI22_X1 port map( A1 => n129, A2 => regs(2400), B1 => n64, B2 => 
                           regs(1888), ZN => n792);
   U1264 : NAND3_X1 port map( A1 => n794, A2 => n793, A3 => n792, ZN => 
                           curr_proc_regs(352));
   U1265 : NAND2_X1 port map( A1 => regs(1377), A2 => n92, ZN => n797);
   U1266 : AOI22_X1 port map( A1 => n54, A2 => regs(865), B1 => n37, B2 => 
                           regs(353), ZN => n796);
   U1267 : AOI22_X1 port map( A1 => n129, A2 => regs(2401), B1 => n64, B2 => 
                           regs(1889), ZN => n795);
   U1268 : NAND3_X1 port map( A1 => n797, A2 => n796, A3 => n795, ZN => 
                           curr_proc_regs(353));
   U1269 : NAND2_X1 port map( A1 => regs(866), A2 => n43, ZN => n800);
   U1270 : AOI22_X1 port map( A1 => n88, A2 => regs(1378), B1 => n37, B2 => 
                           regs(354), ZN => n799);
   U1271 : AOI22_X1 port map( A1 => n129, A2 => regs(2402), B1 => n64, B2 => 
                           regs(1890), ZN => n798);
   U1272 : NAND3_X1 port map( A1 => n800, A2 => n799, A3 => n798, ZN => 
                           curr_proc_regs(354));
   U1273 : NAND2_X1 port map( A1 => regs(867), A2 => n44, ZN => n803);
   U1274 : AOI22_X1 port map( A1 => n94, A2 => regs(1379), B1 => n37, B2 => 
                           regs(355), ZN => n802);
   U1275 : AOI22_X1 port map( A1 => n129, A2 => regs(2403), B1 => n64, B2 => 
                           regs(1891), ZN => n801);
   U1276 : NAND3_X1 port map( A1 => n803, A2 => n802, A3 => n801, ZN => 
                           curr_proc_regs(355));
   U1277 : NAND2_X1 port map( A1 => regs(868), A2 => n55, ZN => n806);
   U1278 : AOI22_X1 port map( A1 => n91, A2 => regs(1380), B1 => n37, B2 => 
                           regs(356), ZN => n805);
   U1279 : AOI22_X1 port map( A1 => n129, A2 => regs(2404), B1 => n64, B2 => 
                           regs(1892), ZN => n804);
   U1280 : NAND3_X1 port map( A1 => n806, A2 => n805, A3 => n804, ZN => 
                           curr_proc_regs(356));
   U1281 : NAND2_X1 port map( A1 => regs(869), A2 => n43, ZN => n809);
   U1282 : AOI22_X1 port map( A1 => n96, A2 => regs(1381), B1 => n37, B2 => 
                           regs(357), ZN => n808);
   U1283 : AOI22_X1 port map( A1 => n129, A2 => regs(2405), B1 => n64, B2 => 
                           regs(1893), ZN => n807);
   U1284 : NAND3_X1 port map( A1 => n809, A2 => n808, A3 => n807, ZN => 
                           curr_proc_regs(357));
   U1285 : NAND2_X1 port map( A1 => regs(870), A2 => n56, ZN => n812);
   U1286 : AOI22_X1 port map( A1 => n88, A2 => regs(1382), B1 => n37, B2 => 
                           regs(358), ZN => n811);
   U1287 : AOI22_X1 port map( A1 => n129, A2 => regs(2406), B1 => n64, B2 => 
                           regs(1894), ZN => n810);
   U1288 : NAND3_X1 port map( A1 => n812, A2 => n811, A3 => n810, ZN => 
                           curr_proc_regs(358));
   U1289 : NAND2_X1 port map( A1 => regs(871), A2 => n1, ZN => n815);
   U1290 : AOI22_X1 port map( A1 => n95, A2 => regs(1383), B1 => n37, B2 => 
                           regs(359), ZN => n814);
   U1291 : AOI22_X1 port map( A1 => n129, A2 => regs(2407), B1 => n64, B2 => 
                           regs(1895), ZN => n813);
   U1292 : NAND3_X1 port map( A1 => n815, A2 => n814, A3 => n813, ZN => 
                           curr_proc_regs(359));
   U1293 : INV_X1 port map( A => regs(1059), ZN => n1418);
   U1294 : AOI22_X1 port map( A1 => n127, A2 => regs(2083), B1 => n74, B2 => 
                           regs(1571), ZN => n817);
   U1295 : AOI22_X1 port map( A1 => n47, A2 => regs(547), B1 => n39, B2 => 
                           regs(35), ZN => n816);
   U1296 : OAI211_X1 port map( C1 => n6, C2 => n1418, A => n817, B => n816, ZN 
                           => curr_proc_regs(35));
   U1297 : NAND2_X1 port map( A1 => regs(872), A2 => n54, ZN => n820);
   U1298 : AOI22_X1 port map( A1 => n91, A2 => regs(1384), B1 => n39, B2 => 
                           regs(360), ZN => n819);
   U1299 : AOI22_X1 port map( A1 => n128, A2 => regs(2408), B1 => n69, B2 => 
                           regs(1896), ZN => n818);
   U1300 : NAND3_X1 port map( A1 => n820, A2 => n819, A3 => n818, ZN => 
                           curr_proc_regs(360));
   U1301 : NAND2_X1 port map( A1 => regs(1385), A2 => n95, ZN => n823);
   U1302 : AOI22_X1 port map( A1 => n52, A2 => regs(873), B1 => n39, B2 => 
                           regs(361), ZN => n822);
   U1303 : AOI22_X1 port map( A1 => n127, A2 => regs(2409), B1 => n73, B2 => 
                           regs(1897), ZN => n821);
   U1304 : NAND3_X1 port map( A1 => n823, A2 => n822, A3 => n821, ZN => 
                           curr_proc_regs(361));
   U1305 : NAND2_X1 port map( A1 => regs(1386), A2 => n95, ZN => n826);
   U1306 : AOI22_X1 port map( A1 => n46, A2 => regs(874), B1 => n39, B2 => 
                           regs(362), ZN => n825);
   U1307 : AOI22_X1 port map( A1 => n129, A2 => regs(2410), B1 => n71, B2 => 
                           regs(1898), ZN => n824);
   U1308 : NAND3_X1 port map( A1 => n826, A2 => n825, A3 => n824, ZN => 
                           curr_proc_regs(362));
   U1309 : NAND2_X1 port map( A1 => regs(875), A2 => n3, ZN => n829);
   U1310 : AOI22_X1 port map( A1 => n89, A2 => regs(1387), B1 => n38, B2 => 
                           regs(363), ZN => n828);
   U1311 : AOI22_X1 port map( A1 => n126, A2 => regs(2411), B1 => n5, B2 => 
                           regs(1899), ZN => n827);
   U1312 : NAND3_X1 port map( A1 => n829, A2 => n828, A3 => n827, ZN => 
                           curr_proc_regs(363));
   U1313 : NAND2_X1 port map( A1 => regs(876), A2 => n44, ZN => n832);
   U1314 : AOI22_X1 port map( A1 => n92, A2 => regs(1388), B1 => n38, B2 => 
                           regs(364), ZN => n831);
   U1315 : AOI22_X1 port map( A1 => n127, A2 => regs(2412), B1 => n68, B2 => 
                           regs(1900), ZN => n830);
   U1316 : NAND3_X1 port map( A1 => n832, A2 => n831, A3 => n830, ZN => 
                           curr_proc_regs(364));
   U1317 : NAND2_X1 port map( A1 => regs(877), A2 => n8, ZN => n835);
   U1318 : AOI22_X1 port map( A1 => n96, A2 => regs(1389), B1 => n38, B2 => 
                           regs(365), ZN => n834);
   U1319 : AOI22_X1 port map( A1 => n128, A2 => regs(2413), B1 => n72, B2 => 
                           regs(1901), ZN => n833);
   U1320 : NAND3_X1 port map( A1 => n835, A2 => n834, A3 => n833, ZN => 
                           curr_proc_regs(365));
   U1321 : NAND2_X1 port map( A1 => regs(1390), A2 => n96, ZN => n838);
   U1322 : AOI22_X1 port map( A1 => n46, A2 => regs(878), B1 => n38, B2 => 
                           regs(366), ZN => n837);
   U1323 : AOI22_X1 port map( A1 => n128, A2 => regs(2414), B1 => n70, B2 => 
                           regs(1902), ZN => n836);
   U1324 : NAND3_X1 port map( A1 => n838, A2 => n837, A3 => n836, ZN => 
                           curr_proc_regs(366));
   U1325 : NAND2_X1 port map( A1 => regs(1391), A2 => n95, ZN => n841);
   U1326 : AOI22_X1 port map( A1 => n41, A2 => regs(879), B1 => n38, B2 => 
                           regs(367), ZN => n840);
   U1327 : AOI22_X1 port map( A1 => n129, A2 => regs(2415), B1 => n74, B2 => 
                           regs(1903), ZN => n839);
   U1328 : NAND3_X1 port map( A1 => n841, A2 => n840, A3 => n839, ZN => 
                           curr_proc_regs(367));
   U1329 : NAND2_X1 port map( A1 => regs(1392), A2 => n97, ZN => n844);
   U1330 : AOI22_X1 port map( A1 => n48, A2 => regs(880), B1 => n38, B2 => 
                           regs(368), ZN => n843);
   U1331 : AOI22_X1 port map( A1 => n126, A2 => regs(2416), B1 => n65, B2 => 
                           regs(1904), ZN => n842);
   U1332 : NAND3_X1 port map( A1 => n844, A2 => n843, A3 => n842, ZN => 
                           curr_proc_regs(368));
   U1333 : NAND2_X1 port map( A1 => regs(1393), A2 => n96, ZN => n847);
   U1334 : AOI22_X1 port map( A1 => n41, A2 => regs(881), B1 => n38, B2 => 
                           regs(369), ZN => n846);
   U1335 : AOI22_X1 port map( A1 => n127, A2 => regs(2417), B1 => n69, B2 => 
                           regs(1905), ZN => n845);
   U1336 : NAND3_X1 port map( A1 => n847, A2 => n846, A3 => n845, ZN => 
                           curr_proc_regs(369));
   U1337 : INV_X1 port map( A => regs(1060), ZN => n1421);
   U1338 : AOI22_X1 port map( A1 => n128, A2 => regs(2084), B1 => n66, B2 => 
                           regs(1572), ZN => n849);
   U1339 : AOI22_X1 port map( A1 => n46, A2 => regs(548), B1 => n38, B2 => 
                           regs(36), ZN => n848);
   U1340 : OAI211_X1 port map( C1 => n78, C2 => n1421, A => n849, B => n848, ZN
                           => curr_proc_regs(36));
   U1341 : NAND2_X1 port map( A1 => regs(1394), A2 => n97, ZN => n852);
   U1342 : AOI22_X1 port map( A1 => n47, A2 => regs(882), B1 => n28, B2 => 
                           regs(370), ZN => n851);
   U1343 : AOI22_X1 port map( A1 => n129, A2 => regs(2418), B1 => n63, B2 => 
                           regs(1906), ZN => n850);
   U1344 : NAND3_X1 port map( A1 => n852, A2 => n851, A3 => n850, ZN => 
                           curr_proc_regs(370));
   U1345 : NAND2_X1 port map( A1 => regs(883), A2 => n8, ZN => n855);
   U1346 : AOI22_X1 port map( A1 => n88, A2 => regs(1395), B1 => n29, B2 => 
                           regs(371), ZN => n854);
   U1347 : AOI22_X1 port map( A1 => n126, A2 => regs(2419), B1 => n64, B2 => 
                           regs(1907), ZN => n853);
   U1348 : NAND3_X1 port map( A1 => n855, A2 => n854, A3 => n853, ZN => 
                           curr_proc_regs(371));
   U1349 : NAND2_X1 port map( A1 => regs(1396), A2 => n98, ZN => n858);
   U1350 : AOI22_X1 port map( A1 => n52, A2 => regs(884), B1 => n30, B2 => 
                           regs(372), ZN => n857);
   U1351 : AOI22_X1 port map( A1 => n127, A2 => regs(2420), B1 => n60, B2 => 
                           regs(1908), ZN => n856);
   U1352 : NAND3_X1 port map( A1 => n858, A2 => n857, A3 => n856, ZN => 
                           curr_proc_regs(372));
   U1353 : NAND2_X1 port map( A1 => regs(885), A2 => n8, ZN => n861);
   U1354 : AOI22_X1 port map( A1 => n89, A2 => regs(1397), B1 => n32, B2 => 
                           regs(373), ZN => n860);
   U1355 : AOI22_X1 port map( A1 => n128, A2 => regs(2421), B1 => n64, B2 => 
                           regs(1909), ZN => n859);
   U1356 : NAND3_X1 port map( A1 => n861, A2 => n860, A3 => n859, ZN => 
                           curr_proc_regs(373));
   U1357 : NAND2_X1 port map( A1 => regs(886), A2 => n8, ZN => n864);
   U1358 : AOI22_X1 port map( A1 => n88, A2 => regs(1398), B1 => n39, B2 => 
                           regs(374), ZN => n863);
   U1359 : AOI22_X1 port map( A1 => n129, A2 => regs(2422), B1 => n5, B2 => 
                           regs(1910), ZN => n862);
   U1360 : NAND3_X1 port map( A1 => n864, A2 => n863, A3 => n862, ZN => 
                           curr_proc_regs(374));
   U1361 : NAND2_X1 port map( A1 => regs(887), A2 => n56, ZN => n867);
   U1362 : AOI22_X1 port map( A1 => n100, A2 => regs(1399), B1 => n39, B2 => 
                           regs(375), ZN => n866);
   U1363 : AOI22_X1 port map( A1 => n126, A2 => regs(2423), B1 => n71, B2 => 
                           regs(1911), ZN => n865);
   U1364 : NAND3_X1 port map( A1 => n867, A2 => n866, A3 => n865, ZN => 
                           curr_proc_regs(375));
   U1365 : NAND2_X1 port map( A1 => regs(1400), A2 => n97, ZN => n870);
   U1366 : AOI22_X1 port map( A1 => n52, A2 => regs(888), B1 => n39, B2 => 
                           regs(376), ZN => n869);
   U1367 : AOI22_X1 port map( A1 => n127, A2 => regs(2424), B1 => n74, B2 => 
                           regs(1912), ZN => n868);
   U1368 : NAND3_X1 port map( A1 => n870, A2 => n869, A3 => n868, ZN => 
                           curr_proc_regs(376));
   U1369 : NAND2_X1 port map( A1 => regs(889), A2 => n56, ZN => n873);
   U1370 : AOI22_X1 port map( A1 => n89, A2 => regs(1401), B1 => n39, B2 => 
                           regs(377), ZN => n872);
   U1371 : AOI22_X1 port map( A1 => n128, A2 => regs(2425), B1 => n74, B2 => 
                           regs(1913), ZN => n871);
   U1372 : NAND3_X1 port map( A1 => n873, A2 => n872, A3 => n871, ZN => 
                           curr_proc_regs(377));
   U1373 : NAND2_X1 port map( A1 => regs(890), A2 => n8, ZN => n876);
   U1374 : AOI22_X1 port map( A1 => n88, A2 => regs(1402), B1 => n39, B2 => 
                           regs(378), ZN => n875);
   U1375 : AOI22_X1 port map( A1 => n129, A2 => regs(2426), B1 => n63, B2 => 
                           regs(1914), ZN => n874);
   U1376 : NAND3_X1 port map( A1 => n876, A2 => n875, A3 => n874, ZN => 
                           curr_proc_regs(378));
   U1377 : NAND2_X1 port map( A1 => regs(1403), A2 => n97, ZN => n879);
   U1378 : AOI22_X1 port map( A1 => n42, A2 => regs(891), B1 => n39, B2 => 
                           regs(379), ZN => n878);
   U1379 : AOI22_X1 port map( A1 => n126, A2 => regs(2427), B1 => n63, B2 => 
                           regs(1915), ZN => n877);
   U1380 : NAND3_X1 port map( A1 => n879, A2 => n878, A3 => n877, ZN => 
                           curr_proc_regs(379));
   U1381 : INV_X1 port map( A => regs(549), ZN => n1424);
   U1382 : AOI22_X1 port map( A1 => n127, A2 => regs(2085), B1 => n2211, B2 => 
                           regs(1573), ZN => n881);
   U1383 : AOI22_X1 port map( A1 => n89, A2 => regs(1061), B1 => n39, B2 => 
                           regs(37), ZN => n880);
   U1384 : OAI211_X1 port map( C1 => n58, C2 => n1424, A => n881, B => n880, ZN
                           => curr_proc_regs(37));
   U1385 : NAND2_X1 port map( A1 => regs(1404), A2 => n98, ZN => n884);
   U1386 : AOI22_X1 port map( A1 => n48, A2 => regs(892), B1 => n39, B2 => 
                           regs(380), ZN => n883);
   U1387 : AOI22_X1 port map( A1 => n128, A2 => regs(2428), B1 => n5, B2 => 
                           regs(1916), ZN => n882);
   U1388 : NAND3_X1 port map( A1 => n884, A2 => n883, A3 => n882, ZN => 
                           curr_proc_regs(380));
   U1389 : NAND2_X1 port map( A1 => regs(893), A2 => n56, ZN => n887);
   U1390 : AOI22_X1 port map( A1 => n89, A2 => regs(1405), B1 => n24, B2 => 
                           regs(381), ZN => n886);
   U1391 : AOI22_X1 port map( A1 => n128, A2 => regs(2429), B1 => n74, B2 => 
                           regs(1917), ZN => n885);
   U1392 : NAND3_X1 port map( A1 => n887, A2 => n886, A3 => n885, ZN => 
                           curr_proc_regs(381));
   U1393 : NAND2_X1 port map( A1 => regs(1406), A2 => n91, ZN => n890);
   U1394 : AOI22_X1 port map( A1 => n52, A2 => regs(894), B1 => n17, B2 => 
                           regs(382), ZN => n889);
   U1395 : AOI22_X1 port map( A1 => n128, A2 => regs(2430), B1 => n5, B2 => 
                           regs(1918), ZN => n888);
   U1396 : NAND3_X1 port map( A1 => n890, A2 => n889, A3 => n888, ZN => 
                           curr_proc_regs(382));
   U1397 : NAND2_X1 port map( A1 => regs(895), A2 => n8, ZN => n893);
   U1398 : AOI22_X1 port map( A1 => n80, A2 => regs(1407), B1 => n18, B2 => 
                           regs(383), ZN => n892);
   U1399 : AOI22_X1 port map( A1 => n128, A2 => regs(2431), B1 => n68, B2 => 
                           regs(1919), ZN => n891);
   U1400 : NAND3_X1 port map( A1 => n893, A2 => n892, A3 => n891, ZN => 
                           curr_proc_regs(383));
   U1401 : NAND2_X1 port map( A1 => regs(1408), A2 => n95, ZN => n896);
   U1402 : AOI22_X1 port map( A1 => n42, A2 => regs(896), B1 => n19, B2 => 
                           regs(384), ZN => n895);
   U1403 : AOI22_X1 port map( A1 => n128, A2 => regs(2432), B1 => n72, B2 => 
                           regs(1920), ZN => n894);
   U1404 : NAND3_X1 port map( A1 => n896, A2 => n895, A3 => n894, ZN => 
                           curr_proc_regs(384));
   U1405 : NAND2_X1 port map( A1 => regs(897), A2 => n56, ZN => n899);
   U1406 : AOI22_X1 port map( A1 => n82, A2 => regs(1409), B1 => n27, B2 => 
                           regs(385), ZN => n898);
   U1407 : AOI22_X1 port map( A1 => n128, A2 => regs(2433), B1 => n72, B2 => 
                           regs(1921), ZN => n897);
   U1408 : NAND3_X1 port map( A1 => n899, A2 => n898, A3 => n897, ZN => 
                           curr_proc_regs(385));
   U1409 : NAND2_X1 port map( A1 => regs(898), A2 => n3, ZN => n902);
   U1410 : AOI22_X1 port map( A1 => n84, A2 => regs(1410), B1 => n26, B2 => 
                           regs(386), ZN => n901);
   U1411 : AOI22_X1 port map( A1 => n128, A2 => regs(2434), B1 => n72, B2 => 
                           regs(1922), ZN => n900);
   U1412 : NAND3_X1 port map( A1 => n902, A2 => n901, A3 => n900, ZN => 
                           curr_proc_regs(386));
   U1413 : NAND2_X1 port map( A1 => regs(899), A2 => n8, ZN => n905);
   U1414 : AOI22_X1 port map( A1 => n81, A2 => regs(1411), B1 => n25, B2 => 
                           regs(387), ZN => n904);
   U1415 : AOI22_X1 port map( A1 => n128, A2 => regs(2435), B1 => n2211, B2 => 
                           regs(1923), ZN => n903);
   U1416 : NAND3_X1 port map( A1 => n905, A2 => n904, A3 => n903, ZN => 
                           curr_proc_regs(387));
   U1417 : NAND2_X1 port map( A1 => regs(1412), A2 => n98, ZN => n908);
   U1418 : AOI22_X1 port map( A1 => n51, A2 => regs(900), B1 => n28, B2 => 
                           regs(388), ZN => n907);
   U1419 : AOI22_X1 port map( A1 => n128, A2 => regs(2436), B1 => n74, B2 => 
                           regs(1924), ZN => n906);
   U1420 : NAND3_X1 port map( A1 => n908, A2 => n907, A3 => n906, ZN => 
                           curr_proc_regs(388));
   U1421 : NAND2_X1 port map( A1 => regs(1413), A2 => n97, ZN => n911);
   U1422 : AOI22_X1 port map( A1 => n48, A2 => regs(901), B1 => n29, B2 => 
                           regs(389), ZN => n910);
   U1423 : AOI22_X1 port map( A1 => n128, A2 => regs(2437), B1 => n5, B2 => 
                           regs(1925), ZN => n909);
   U1424 : NAND3_X1 port map( A1 => n911, A2 => n910, A3 => n909, ZN => 
                           curr_proc_regs(389));
   U1425 : INV_X1 port map( A => regs(550), ZN => n1429);
   U1426 : AOI22_X1 port map( A1 => n128, A2 => regs(2086), B1 => n74, B2 => 
                           regs(1574), ZN => n913);
   U1427 : AOI22_X1 port map( A1 => n80, A2 => regs(1062), B1 => n35, B2 => 
                           regs(38), ZN => n912);
   U1428 : OAI211_X1 port map( C1 => n58, C2 => n1429, A => n913, B => n912, ZN
                           => curr_proc_regs(38));
   U1429 : NAND2_X1 port map( A1 => regs(1414), A2 => n98, ZN => n916);
   U1430 : AOI22_X1 port map( A1 => n51, A2 => regs(902), B1 => n37, B2 => 
                           regs(390), ZN => n915);
   U1431 : AOI22_X1 port map( A1 => n128, A2 => regs(2438), B1 => n5, B2 => 
                           regs(1926), ZN => n914);
   U1432 : NAND3_X1 port map( A1 => n916, A2 => n915, A3 => n914, ZN => 
                           curr_proc_regs(390));
   U1433 : NAND2_X1 port map( A1 => regs(903), A2 => n8, ZN => n919);
   U1434 : AOI22_X1 port map( A1 => n85, A2 => regs(1415), B1 => n21, B2 => 
                           regs(391), ZN => n918);
   U1435 : AOI22_X1 port map( A1 => n128, A2 => regs(2439), B1 => n68, B2 => 
                           regs(1927), ZN => n917);
   U1436 : NAND3_X1 port map( A1 => n919, A2 => n918, A3 => n917, ZN => 
                           curr_proc_regs(391));
   U1437 : NAND2_X1 port map( A1 => regs(904), A2 => n56, ZN => n922);
   U1438 : AOI22_X1 port map( A1 => n86, A2 => regs(1416), B1 => n17, B2 => 
                           regs(392), ZN => n921);
   U1439 : AOI22_X1 port map( A1 => n127, A2 => regs(2440), B1 => n60, B2 => 
                           regs(1928), ZN => n920);
   U1440 : NAND3_X1 port map( A1 => n922, A2 => n921, A3 => n920, ZN => 
                           curr_proc_regs(392));
   U1441 : NAND2_X1 port map( A1 => regs(905), A2 => n8, ZN => n925);
   U1442 : AOI22_X1 port map( A1 => n87, A2 => regs(1417), B1 => n17, B2 => 
                           regs(393), ZN => n924);
   U1443 : AOI22_X1 port map( A1 => n127, A2 => regs(2441), B1 => n64, B2 => 
                           regs(1929), ZN => n923);
   U1444 : NAND3_X1 port map( A1 => n925, A2 => n924, A3 => n923, ZN => 
                           curr_proc_regs(393));
   U1445 : NAND2_X1 port map( A1 => regs(1418), A2 => n98, ZN => n928);
   U1446 : AOI22_X1 port map( A1 => n47, A2 => regs(906), B1 => n17, B2 => 
                           regs(394), ZN => n927);
   U1447 : AOI22_X1 port map( A1 => n127, A2 => regs(2442), B1 => n69, B2 => 
                           regs(1930), ZN => n926);
   U1448 : NAND3_X1 port map( A1 => n928, A2 => n927, A3 => n926, ZN => 
                           curr_proc_regs(394));
   U1449 : NAND2_X1 port map( A1 => regs(907), A2 => n53, ZN => n931);
   U1450 : AOI22_X1 port map( A1 => n82, A2 => regs(1419), B1 => n17, B2 => 
                           regs(395), ZN => n930);
   U1451 : AOI22_X1 port map( A1 => n127, A2 => regs(2443), B1 => n72, B2 => 
                           regs(1931), ZN => n929);
   U1452 : NAND3_X1 port map( A1 => n931, A2 => n930, A3 => n929, ZN => 
                           curr_proc_regs(395));
   U1453 : NAND2_X1 port map( A1 => regs(908), A2 => n8, ZN => n934);
   U1454 : AOI22_X1 port map( A1 => n87, A2 => regs(1420), B1 => n17, B2 => 
                           regs(396), ZN => n933);
   U1455 : AOI22_X1 port map( A1 => n127, A2 => regs(2444), B1 => n5, B2 => 
                           regs(1932), ZN => n932);
   U1456 : NAND3_X1 port map( A1 => n934, A2 => n933, A3 => n932, ZN => 
                           curr_proc_regs(396));
   U1457 : NAND2_X1 port map( A1 => regs(909), A2 => n8, ZN => n937);
   U1458 : AOI22_X1 port map( A1 => n84, A2 => regs(1421), B1 => n17, B2 => 
                           regs(397), ZN => n936);
   U1459 : AOI22_X1 port map( A1 => n127, A2 => regs(2445), B1 => n66, B2 => 
                           regs(1933), ZN => n935);
   U1460 : NAND3_X1 port map( A1 => n937, A2 => n936, A3 => n935, ZN => 
                           curr_proc_regs(397));
   U1461 : NAND2_X1 port map( A1 => regs(910), A2 => n56, ZN => n940);
   U1462 : AOI22_X1 port map( A1 => n80, A2 => regs(1422), B1 => n17, B2 => 
                           regs(398), ZN => n939);
   U1463 : AOI22_X1 port map( A1 => n127, A2 => regs(2446), B1 => n66, B2 => 
                           regs(1934), ZN => n938);
   U1464 : NAND3_X1 port map( A1 => n940, A2 => n939, A3 => n938, ZN => 
                           curr_proc_regs(398));
   U1465 : NAND2_X1 port map( A1 => regs(1423), A2 => n98, ZN => n943);
   U1466 : AOI22_X1 port map( A1 => n47, A2 => regs(911), B1 => n17, B2 => 
                           regs(399), ZN => n942);
   U1467 : AOI22_X1 port map( A1 => n127, A2 => regs(2447), B1 => n63, B2 => 
                           regs(1935), ZN => n941);
   U1468 : NAND3_X1 port map( A1 => n943, A2 => n942, A3 => n941, ZN => 
                           curr_proc_regs(399));
   U1469 : INV_X1 port map( A => regs(551), ZN => n1432);
   U1470 : AOI22_X1 port map( A1 => n127, A2 => regs(2087), B1 => n60, B2 => 
                           regs(1575), ZN => n945);
   U1471 : AOI22_X1 port map( A1 => n82, A2 => regs(1063), B1 => n17, B2 => 
                           regs(39), ZN => n944);
   U1472 : OAI211_X1 port map( C1 => n58, C2 => n1432, A => n945, B => n944, ZN
                           => curr_proc_regs(39));
   U1473 : INV_X1 port map( A => regs(515), ZN => n1319);
   U1474 : AOI22_X1 port map( A1 => n127, A2 => regs(2051), B1 => n60, B2 => 
                           regs(1539), ZN => n947);
   U1475 : AOI22_X1 port map( A1 => n93, A2 => regs(1027), B1 => n17, B2 => 
                           regs(3), ZN => n946);
   U1476 : OAI211_X1 port map( C1 => n58, C2 => n1319, A => n947, B => n946, ZN
                           => curr_proc_regs(3));
   U1477 : NAND2_X1 port map( A1 => regs(912), A2 => n8, ZN => n950);
   U1478 : AOI22_X1 port map( A1 => n90, A2 => regs(1424), B1 => n17, B2 => 
                           regs(400), ZN => n949);
   U1479 : AOI22_X1 port map( A1 => n127, A2 => regs(2448), B1 => n64, B2 => 
                           regs(1936), ZN => n948);
   U1480 : NAND3_X1 port map( A1 => n950, A2 => n949, A3 => n948, ZN => 
                           curr_proc_regs(400));
   U1481 : NAND2_X1 port map( A1 => regs(913), A2 => n56, ZN => n953);
   U1482 : AOI22_X1 port map( A1 => n83, A2 => regs(1425), B1 => n17, B2 => 
                           regs(401), ZN => n952);
   U1483 : AOI22_X1 port map( A1 => n127, A2 => regs(2449), B1 => n74, B2 => 
                           regs(1937), ZN => n951);
   U1484 : NAND3_X1 port map( A1 => n953, A2 => n952, A3 => n951, ZN => 
                           curr_proc_regs(401));
   U1485 : NAND2_X1 port map( A1 => regs(1426), A2 => n97, ZN => n956);
   U1486 : AOI22_X1 port map( A1 => n47, A2 => regs(914), B1 => n2, B2 => 
                           regs(402), ZN => n955);
   U1487 : AOI22_X1 port map( A1 => n126, A2 => regs(2450), B1 => n68, B2 => 
                           regs(1938), ZN => n954);
   U1488 : NAND3_X1 port map( A1 => n956, A2 => n955, A3 => n954, ZN => 
                           curr_proc_regs(402));
   U1489 : NAND2_X1 port map( A1 => regs(1427), A2 => n96, ZN => n959);
   U1490 : AOI22_X1 port map( A1 => n47, A2 => regs(915), B1 => n2, B2 => 
                           regs(403), ZN => n958);
   U1491 : AOI22_X1 port map( A1 => n126, A2 => regs(2451), B1 => n74, B2 => 
                           regs(1939), ZN => n957);
   U1492 : NAND3_X1 port map( A1 => n959, A2 => n958, A3 => n957, ZN => 
                           curr_proc_regs(403));
   U1493 : NAND2_X1 port map( A1 => regs(1428), A2 => n96, ZN => n962);
   U1494 : AOI22_X1 port map( A1 => n47, A2 => regs(916), B1 => n2, B2 => 
                           regs(404), ZN => n961);
   U1495 : AOI22_X1 port map( A1 => n126, A2 => regs(2452), B1 => n74, B2 => 
                           regs(1940), ZN => n960);
   U1496 : NAND3_X1 port map( A1 => n962, A2 => n961, A3 => n960, ZN => 
                           curr_proc_regs(404));
   U1497 : NAND2_X1 port map( A1 => regs(917), A2 => n8, ZN => n965);
   U1498 : AOI22_X1 port map( A1 => n99, A2 => regs(1429), B1 => n2, B2 => 
                           regs(405), ZN => n964);
   U1499 : AOI22_X1 port map( A1 => n126, A2 => regs(2453), B1 => n69, B2 => 
                           regs(1941), ZN => n963);
   U1500 : NAND3_X1 port map( A1 => n965, A2 => n964, A3 => n963, ZN => 
                           curr_proc_regs(405));
   U1501 : NAND2_X1 port map( A1 => regs(1430), A2 => n96, ZN => n968);
   U1502 : AOI22_X1 port map( A1 => n47, A2 => regs(918), B1 => n2, B2 => 
                           regs(406), ZN => n967);
   U1503 : AOI22_X1 port map( A1 => n126, A2 => regs(2454), B1 => n72, B2 => 
                           regs(1942), ZN => n966);
   U1504 : NAND3_X1 port map( A1 => n968, A2 => n967, A3 => n966, ZN => 
                           curr_proc_regs(406));
   U1505 : NAND2_X1 port map( A1 => regs(919), A2 => n56, ZN => n971);
   U1506 : AOI22_X1 port map( A1 => n97, A2 => regs(1431), B1 => n2, B2 => 
                           regs(407), ZN => n970);
   U1507 : AOI22_X1 port map( A1 => n126, A2 => regs(2455), B1 => n70, B2 => 
                           regs(1943), ZN => n969);
   U1508 : NAND3_X1 port map( A1 => n971, A2 => n970, A3 => n969, ZN => 
                           curr_proc_regs(407));
   U1509 : NAND2_X1 port map( A1 => regs(1432), A2 => n96, ZN => n974);
   U1510 : AOI22_X1 port map( A1 => n47, A2 => regs(920), B1 => n2, B2 => 
                           regs(408), ZN => n973);
   U1511 : AOI22_X1 port map( A1 => n126, A2 => regs(2456), B1 => n65, B2 => 
                           regs(1944), ZN => n972);
   U1512 : NAND3_X1 port map( A1 => n974, A2 => n973, A3 => n972, ZN => 
                           curr_proc_regs(408));
   U1513 : NAND2_X1 port map( A1 => regs(921), A2 => n8, ZN => n977);
   U1514 : AOI22_X1 port map( A1 => n83, A2 => regs(1433), B1 => n2, B2 => 
                           regs(409), ZN => n976);
   U1515 : AOI22_X1 port map( A1 => n126, A2 => regs(2457), B1 => n72, B2 => 
                           regs(1945), ZN => n975);
   U1516 : NAND3_X1 port map( A1 => n977, A2 => n976, A3 => n975, ZN => 
                           curr_proc_regs(409));
   U1517 : INV_X1 port map( A => regs(552), ZN => n1435);
   U1518 : AOI22_X1 port map( A1 => n126, A2 => regs(2088), B1 => n5, B2 => 
                           regs(1576), ZN => n979);
   U1519 : AOI22_X1 port map( A1 => n90, A2 => regs(1064), B1 => n2, B2 => 
                           regs(40), ZN => n978);
   U1520 : OAI211_X1 port map( C1 => n58, C2 => n1435, A => n979, B => n978, ZN
                           => curr_proc_regs(40));
   U1521 : NAND2_X1 port map( A1 => regs(1434), A2 => n95, ZN => n982);
   U1522 : AOI22_X1 port map( A1 => n47, A2 => regs(922), B1 => n2, B2 => 
                           regs(410), ZN => n981);
   U1523 : AOI22_X1 port map( A1 => n126, A2 => regs(2458), B1 => n69, B2 => 
                           regs(1946), ZN => n980);
   U1524 : NAND3_X1 port map( A1 => n982, A2 => n981, A3 => n980, ZN => 
                           curr_proc_regs(410));
   U1525 : NAND2_X1 port map( A1 => regs(1435), A2 => n95, ZN => n985);
   U1526 : AOI22_X1 port map( A1 => n48, A2 => regs(923), B1 => n2, B2 => 
                           regs(411), ZN => n984);
   U1527 : AOI22_X1 port map( A1 => n126, A2 => regs(2459), B1 => n66, B2 => 
                           regs(1947), ZN => n983);
   U1528 : NAND3_X1 port map( A1 => n985, A2 => n984, A3 => n983, ZN => 
                           curr_proc_regs(411));
   U1529 : NAND2_X1 port map( A1 => regs(924), A2 => n8, ZN => n988);
   U1530 : AOI22_X1 port map( A1 => n90, A2 => regs(1436), B1 => n2, B2 => 
                           regs(412), ZN => n987);
   U1531 : AOI22_X1 port map( A1 => n126, A2 => regs(2460), B1 => n72, B2 => 
                           regs(1948), ZN => n986);
   U1532 : NAND3_X1 port map( A1 => n988, A2 => n987, A3 => n986, ZN => 
                           curr_proc_regs(412));
   U1533 : NAND2_X1 port map( A1 => regs(1437), A2 => n95, ZN => n991);
   U1534 : AOI22_X1 port map( A1 => n54, A2 => regs(925), B1 => n18, B2 => 
                           regs(413), ZN => n990);
   U1535 : AOI22_X1 port map( A1 => n125, A2 => regs(2461), B1 => n65, B2 => 
                           regs(1949), ZN => n989);
   U1536 : NAND3_X1 port map( A1 => n991, A2 => n990, A3 => n989, ZN => 
                           curr_proc_regs(413));
   U1537 : NAND2_X1 port map( A1 => regs(1438), A2 => n95, ZN => n994);
   U1538 : AOI22_X1 port map( A1 => n46, A2 => regs(926), B1 => n18, B2 => 
                           regs(414), ZN => n993);
   U1539 : AOI22_X1 port map( A1 => n124, A2 => regs(2462), B1 => n65, B2 => 
                           regs(1950), ZN => n992);
   U1540 : NAND3_X1 port map( A1 => n994, A2 => n993, A3 => n992, ZN => 
                           curr_proc_regs(414));
   U1541 : NAND2_X1 port map( A1 => regs(927), A2 => n56, ZN => n997);
   U1542 : AOI22_X1 port map( A1 => n99, A2 => regs(1439), B1 => n18, B2 => 
                           regs(415), ZN => n996);
   U1543 : AOI22_X1 port map( A1 => n105, A2 => regs(2463), B1 => n65, B2 => 
                           regs(1951), ZN => n995);
   U1544 : NAND3_X1 port map( A1 => n997, A2 => n996, A3 => n995, ZN => 
                           curr_proc_regs(415));
   U1545 : NAND2_X1 port map( A1 => regs(1440), A2 => n94, ZN => n1000);
   U1546 : AOI22_X1 port map( A1 => n46, A2 => regs(928), B1 => n18, B2 => 
                           regs(416), ZN => n999);
   U1547 : AOI22_X1 port map( A1 => n125, A2 => regs(2464), B1 => n65, B2 => 
                           regs(1952), ZN => n998);
   U1548 : NAND3_X1 port map( A1 => n1000, A2 => n999, A3 => n998, ZN => 
                           curr_proc_regs(416));
   U1549 : NAND2_X1 port map( A1 => regs(929), A2 => n56, ZN => n1003);
   U1550 : AOI22_X1 port map( A1 => n97, A2 => regs(1441), B1 => n18, B2 => 
                           regs(417), ZN => n1002);
   U1551 : AOI22_X1 port map( A1 => n125, A2 => regs(2465), B1 => n65, B2 => 
                           regs(1953), ZN => n1001);
   U1552 : NAND3_X1 port map( A1 => n1003, A2 => n1002, A3 => n1001, ZN => 
                           curr_proc_regs(417));
   U1553 : NAND2_X1 port map( A1 => regs(1442), A2 => n94, ZN => n1006);
   U1554 : AOI22_X1 port map( A1 => n46, A2 => regs(930), B1 => n18, B2 => 
                           regs(418), ZN => n1005);
   U1555 : AOI22_X1 port map( A1 => n125, A2 => regs(2466), B1 => n65, B2 => 
                           regs(1954), ZN => n1004);
   U1556 : NAND3_X1 port map( A1 => n1006, A2 => n1005, A3 => n1004, ZN => 
                           curr_proc_regs(418));
   U1557 : NAND2_X1 port map( A1 => regs(1443), A2 => n93, ZN => n1009);
   U1558 : AOI22_X1 port map( A1 => n46, A2 => regs(931), B1 => n18, B2 => 
                           regs(419), ZN => n1008);
   U1559 : AOI22_X1 port map( A1 => n125, A2 => regs(2467), B1 => n65, B2 => 
                           regs(1955), ZN => n1007);
   U1560 : NAND3_X1 port map( A1 => n1009, A2 => n1008, A3 => n1007, ZN => 
                           curr_proc_regs(419));
   U1561 : INV_X1 port map( A => regs(1065), ZN => n1438);
   U1562 : AOI22_X1 port map( A1 => n124, A2 => regs(2089), B1 => n65, B2 => 
                           regs(1577), ZN => n1011);
   U1563 : AOI22_X1 port map( A1 => n46, A2 => regs(553), B1 => n18, B2 => 
                           regs(41), ZN => n1010);
   U1564 : OAI211_X1 port map( C1 => n2215, C2 => n1438, A => n1011, B => n1010
                           , ZN => curr_proc_regs(41));
   U1565 : NAND2_X1 port map( A1 => regs(1444), A2 => n93, ZN => n1014);
   U1566 : AOI22_X1 port map( A1 => n46, A2 => regs(932), B1 => n18, B2 => 
                           regs(420), ZN => n1013);
   U1567 : AOI22_X1 port map( A1 => n122, A2 => regs(2468), B1 => n65, B2 => 
                           regs(1956), ZN => n1012);
   U1568 : NAND3_X1 port map( A1 => n1014, A2 => n1013, A3 => n1012, ZN => 
                           curr_proc_regs(420));
   U1569 : NAND2_X1 port map( A1 => regs(933), A2 => n8, ZN => n1017);
   U1570 : AOI22_X1 port map( A1 => n93, A2 => regs(1445), B1 => n18, B2 => 
                           regs(421), ZN => n1016);
   U1571 : AOI22_X1 port map( A1 => n128, A2 => regs(2469), B1 => n65, B2 => 
                           regs(1957), ZN => n1015);
   U1572 : NAND3_X1 port map( A1 => n1017, A2 => n1016, A3 => n1015, ZN => 
                           curr_proc_regs(421));
   U1573 : NAND2_X1 port map( A1 => regs(1446), A2 => n93, ZN => n1020);
   U1574 : AOI22_X1 port map( A1 => n46, A2 => regs(934), B1 => n18, B2 => 
                           regs(422), ZN => n1019);
   U1575 : AOI22_X1 port map( A1 => n124, A2 => regs(2470), B1 => n65, B2 => 
                           regs(1958), ZN => n1018);
   U1576 : NAND3_X1 port map( A1 => n1020, A2 => n1019, A3 => n1018, ZN => 
                           curr_proc_regs(422));
   U1577 : NAND2_X1 port map( A1 => regs(1447), A2 => n93, ZN => n1023);
   U1578 : AOI22_X1 port map( A1 => n46, A2 => regs(935), B1 => n18, B2 => 
                           regs(423), ZN => n1022);
   U1579 : AOI22_X1 port map( A1 => n124, A2 => regs(2471), B1 => n65, B2 => 
                           regs(1959), ZN => n1021);
   U1580 : NAND3_X1 port map( A1 => n1023, A2 => n1022, A3 => n1021, ZN => 
                           curr_proc_regs(423));
   U1581 : NAND2_X1 port map( A1 => regs(1448), A2 => n93, ZN => n1026);
   U1582 : AOI22_X1 port map( A1 => n46, A2 => regs(936), B1 => n2, B2 => 
                           regs(424), ZN => n1025);
   U1583 : AOI22_X1 port map( A1 => n124, A2 => regs(2472), B1 => n5, B2 => 
                           regs(1960), ZN => n1024);
   U1584 : NAND3_X1 port map( A1 => n1026, A2 => n1025, A3 => n1024, ZN => 
                           curr_proc_regs(424));
   U1585 : NAND2_X1 port map( A1 => regs(1449), A2 => n92, ZN => n1029);
   U1586 : AOI22_X1 port map( A1 => n46, A2 => regs(937), B1 => n2, B2 => 
                           regs(425), ZN => n1028);
   U1587 : AOI22_X1 port map( A1 => n113, A2 => regs(2473), B1 => n5, B2 => 
                           regs(1961), ZN => n1027);
   U1588 : NAND3_X1 port map( A1 => n1029, A2 => n1028, A3 => n1027, ZN => 
                           curr_proc_regs(425));
   U1589 : NAND2_X1 port map( A1 => regs(938), A2 => n56, ZN => n1032);
   U1590 : AOI22_X1 port map( A1 => n90, A2 => regs(1450), B1 => n2, B2 => 
                           regs(426), ZN => n1031);
   U1591 : AOI22_X1 port map( A1 => n104, A2 => regs(2474), B1 => n5, B2 => 
                           regs(1962), ZN => n1030);
   U1592 : NAND3_X1 port map( A1 => n1032, A2 => n1031, A3 => n1030, ZN => 
                           curr_proc_regs(426));
   U1593 : NAND2_X1 port map( A1 => regs(1451), A2 => n88, ZN => n1035);
   U1594 : AOI22_X1 port map( A1 => n47, A2 => regs(939), B1 => n2, B2 => 
                           regs(427), ZN => n1034);
   U1595 : AOI22_X1 port map( A1 => n125, A2 => regs(2475), B1 => n5, B2 => 
                           regs(1963), ZN => n1033);
   U1596 : NAND3_X1 port map( A1 => n1035, A2 => n1034, A3 => n1033, ZN => 
                           curr_proc_regs(427));
   U1597 : NAND2_X1 port map( A1 => regs(1452), A2 => n100, ZN => n1038);
   U1598 : AOI22_X1 port map( A1 => n55, A2 => regs(940), B1 => n2, B2 => 
                           regs(428), ZN => n1037);
   U1599 : AOI22_X1 port map( A1 => n124, A2 => regs(2476), B1 => n5, B2 => 
                           regs(1964), ZN => n1036);
   U1600 : NAND3_X1 port map( A1 => n1038, A2 => n1037, A3 => n1036, ZN => 
                           curr_proc_regs(428));
   U1601 : NAND2_X1 port map( A1 => regs(941), A2 => n8, ZN => n1041);
   U1602 : AOI22_X1 port map( A1 => n82, A2 => regs(1453), B1 => n2, B2 => 
                           regs(429), ZN => n1040);
   U1603 : AOI22_X1 port map( A1 => n125, A2 => regs(2477), B1 => n5, B2 => 
                           regs(1965), ZN => n1039);
   U1604 : NAND3_X1 port map( A1 => n1041, A2 => n1040, A3 => n1039, ZN => 
                           curr_proc_regs(429));
   U1605 : INV_X1 port map( A => regs(1066), ZN => n1441);
   U1606 : AOI22_X1 port map( A1 => n112, A2 => regs(2090), B1 => n5, B2 => 
                           regs(1578), ZN => n1043);
   U1607 : AOI22_X1 port map( A1 => n55, A2 => regs(554), B1 => n2, B2 => 
                           regs(42), ZN => n1042);
   U1608 : OAI211_X1 port map( C1 => n2215, C2 => n1441, A => n1043, B => n1042
                           , ZN => curr_proc_regs(42));
   U1609 : NAND2_X1 port map( A1 => regs(942), A2 => n8, ZN => n1046);
   U1610 : AOI22_X1 port map( A1 => n84, A2 => regs(1454), B1 => n2, B2 => 
                           regs(430), ZN => n1045);
   U1611 : AOI22_X1 port map( A1 => n109, A2 => regs(2478), B1 => n5, B2 => 
                           regs(1966), ZN => n1044);
   U1612 : NAND3_X1 port map( A1 => n1046, A2 => n1045, A3 => n1044, ZN => 
                           curr_proc_regs(430));
   U1613 : NAND2_X1 port map( A1 => regs(1455), A2 => n98, ZN => n1049);
   U1614 : AOI22_X1 port map( A1 => n55, A2 => regs(943), B1 => n2, B2 => 
                           regs(431), ZN => n1048);
   U1615 : AOI22_X1 port map( A1 => n125, A2 => regs(2479), B1 => n5, B2 => 
                           regs(1967), ZN => n1047);
   U1616 : NAND3_X1 port map( A1 => n1049, A2 => n1048, A3 => n1047, ZN => 
                           curr_proc_regs(431));
   U1617 : NAND2_X1 port map( A1 => regs(1456), A2 => n92, ZN => n1052);
   U1618 : AOI22_X1 port map( A1 => n55, A2 => regs(944), B1 => n2, B2 => 
                           regs(432), ZN => n1051);
   U1619 : AOI22_X1 port map( A1 => n124, A2 => regs(2480), B1 => n5, B2 => 
                           regs(1968), ZN => n1050);
   U1620 : NAND3_X1 port map( A1 => n1052, A2 => n1051, A3 => n1050, ZN => 
                           curr_proc_regs(432));
   U1621 : NAND2_X1 port map( A1 => regs(945), A2 => n1, ZN => n1055);
   U1622 : AOI22_X1 port map( A1 => n81, A2 => regs(1457), B1 => n2, B2 => 
                           regs(433), ZN => n1054);
   U1623 : AOI22_X1 port map( A1 => n128, A2 => regs(2481), B1 => n5, B2 => 
                           regs(1969), ZN => n1053);
   U1624 : NAND3_X1 port map( A1 => n1055, A2 => n1054, A3 => n1053, ZN => 
                           curr_proc_regs(433));
   U1625 : NAND2_X1 port map( A1 => regs(1458), A2 => n92, ZN => n1058);
   U1626 : AOI22_X1 port map( A1 => n55, A2 => regs(946), B1 => n2, B2 => 
                           regs(434), ZN => n1057);
   U1627 : AOI22_X1 port map( A1 => n115, A2 => regs(2482), B1 => n5, B2 => 
                           regs(1970), ZN => n1056);
   U1628 : NAND3_X1 port map( A1 => n1058, A2 => n1057, A3 => n1056, ZN => 
                           curr_proc_regs(434));
   U1629 : NAND2_X1 port map( A1 => regs(947), A2 => n8, ZN => n1061);
   U1630 : AOI22_X1 port map( A1 => n80, A2 => regs(1459), B1 => n37, B2 => 
                           regs(435), ZN => n1060);
   U1631 : AOI22_X1 port map( A1 => n125, A2 => regs(2483), B1 => n5, B2 => 
                           regs(1971), ZN => n1059);
   U1632 : NAND3_X1 port map( A1 => n1061, A2 => n1060, A3 => n1059, ZN => 
                           curr_proc_regs(435));
   U1633 : NAND2_X1 port map( A1 => regs(948), A2 => n8, ZN => n1064);
   U1634 : AOI22_X1 port map( A1 => n85, A2 => regs(1460), B1 => n36, B2 => 
                           regs(436), ZN => n1063);
   U1635 : AOI22_X1 port map( A1 => n125, A2 => regs(2484), B1 => n74, B2 => 
                           regs(1972), ZN => n1062);
   U1636 : NAND3_X1 port map( A1 => n1064, A2 => n1063, A3 => n1062, ZN => 
                           curr_proc_regs(436));
   U1637 : NAND2_X1 port map( A1 => regs(1461), A2 => n92, ZN => n1067);
   U1638 : AOI22_X1 port map( A1 => n55, A2 => regs(949), B1 => n34, B2 => 
                           regs(437), ZN => n1066);
   U1639 : AOI22_X1 port map( A1 => n125, A2 => regs(2485), B1 => n69, B2 => 
                           regs(1973), ZN => n1065);
   U1640 : NAND3_X1 port map( A1 => n1067, A2 => n1066, A3 => n1065, ZN => 
                           curr_proc_regs(437));
   U1641 : NAND2_X1 port map( A1 => regs(1462), A2 => n91, ZN => n1070);
   U1642 : AOI22_X1 port map( A1 => n54, A2 => regs(950), B1 => n33, B2 => 
                           regs(438), ZN => n1069);
   U1643 : AOI22_X1 port map( A1 => n125, A2 => regs(2486), B1 => n71, B2 => 
                           regs(1974), ZN => n1068);
   U1644 : NAND3_X1 port map( A1 => n1070, A2 => n1069, A3 => n1068, ZN => 
                           curr_proc_regs(438));
   U1645 : NAND2_X1 port map( A1 => regs(951), A2 => n44, ZN => n1073);
   U1646 : AOI22_X1 port map( A1 => n86, A2 => regs(1463), B1 => n31, B2 => 
                           regs(439), ZN => n1072);
   U1647 : AOI22_X1 port map( A1 => n125, A2 => regs(2487), B1 => n68, B2 => 
                           regs(1975), ZN => n1071);
   U1648 : NAND3_X1 port map( A1 => n1073, A2 => n1072, A3 => n1071, ZN => 
                           curr_proc_regs(439));
   U1649 : INV_X1 port map( A => regs(1067), ZN => n1444);
   U1650 : AOI22_X1 port map( A1 => n125, A2 => regs(2091), B1 => n5, B2 => 
                           regs(1579), ZN => n1075);
   U1651 : AOI22_X1 port map( A1 => n54, A2 => regs(555), B1 => n20, B2 => 
                           regs(43), ZN => n1074);
   U1652 : OAI211_X1 port map( C1 => n11, C2 => n1444, A => n1075, B => n1074, 
                           ZN => curr_proc_regs(43));
   U1653 : NAND2_X1 port map( A1 => regs(952), A2 => n45, ZN => n1078);
   U1654 : AOI22_X1 port map( A1 => n87, A2 => regs(1464), B1 => n21, B2 => 
                           regs(440), ZN => n1077);
   U1655 : AOI22_X1 port map( A1 => n125, A2 => regs(2488), B1 => n71, B2 => 
                           regs(1976), ZN => n1076);
   U1656 : NAND3_X1 port map( A1 => n1078, A2 => n1077, A3 => n1076, ZN => 
                           curr_proc_regs(440));
   U1657 : NAND2_X1 port map( A1 => regs(1465), A2 => n91, ZN => n1081);
   U1658 : AOI22_X1 port map( A1 => n54, A2 => regs(953), B1 => n22, B2 => 
                           regs(441), ZN => n1080);
   U1659 : AOI22_X1 port map( A1 => n125, A2 => regs(2489), B1 => n68, B2 => 
                           regs(1977), ZN => n1079);
   U1660 : NAND3_X1 port map( A1 => n1081, A2 => n1080, A3 => n1079, ZN => 
                           curr_proc_regs(441));
   U1661 : NAND2_X1 port map( A1 => regs(954), A2 => n45, ZN => n1084);
   U1662 : AOI22_X1 port map( A1 => n81, A2 => regs(1466), B1 => n23, B2 => 
                           regs(442), ZN => n1083);
   U1663 : AOI22_X1 port map( A1 => n125, A2 => regs(2490), B1 => n5, B2 => 
                           regs(1978), ZN => n1082);
   U1664 : NAND3_X1 port map( A1 => n1084, A2 => n1083, A3 => n1082, ZN => 
                           curr_proc_regs(442));
   U1665 : NAND2_X1 port map( A1 => regs(955), A2 => n53, ZN => n1087);
   U1666 : AOI22_X1 port map( A1 => n82, A2 => regs(1467), B1 => n24, B2 => 
                           regs(443), ZN => n1086);
   U1667 : AOI22_X1 port map( A1 => n125, A2 => regs(2491), B1 => n74, B2 => 
                           regs(1979), ZN => n1085);
   U1668 : NAND3_X1 port map( A1 => n1087, A2 => n1086, A3 => n1085, ZN => 
                           curr_proc_regs(443));
   U1669 : NAND2_X1 port map( A1 => regs(956), A2 => n55, ZN => n1090);
   U1670 : AOI22_X1 port map( A1 => n82, A2 => regs(1468), B1 => n17, B2 => 
                           regs(444), ZN => n1089);
   U1671 : AOI22_X1 port map( A1 => n129, A2 => regs(2492), B1 => n69, B2 => 
                           regs(1980), ZN => n1088);
   U1672 : NAND3_X1 port map( A1 => n1090, A2 => n1089, A3 => n1088, ZN => 
                           curr_proc_regs(444));
   U1673 : NAND2_X1 port map( A1 => regs(957), A2 => n56, ZN => n1093);
   U1674 : AOI22_X1 port map( A1 => n85, A2 => regs(1469), B1 => n18, B2 => 
                           regs(445), ZN => n1092);
   U1675 : AOI22_X1 port map( A1 => n121, A2 => regs(2493), B1 => n71, B2 => 
                           regs(1981), ZN => n1091);
   U1676 : NAND3_X1 port map( A1 => n1093, A2 => n1092, A3 => n1091, ZN => 
                           curr_proc_regs(445));
   U1677 : NAND2_X1 port map( A1 => regs(1470), A2 => n91, ZN => n1096);
   U1678 : AOI22_X1 port map( A1 => n54, A2 => regs(958), B1 => n28, B2 => 
                           regs(446), ZN => n1095);
   U1679 : AOI22_X1 port map( A1 => n123, A2 => regs(2494), B1 => n66, B2 => 
                           regs(1982), ZN => n1094);
   U1680 : NAND3_X1 port map( A1 => n1096, A2 => n1095, A3 => n1094, ZN => 
                           curr_proc_regs(446));
   U1681 : NAND2_X1 port map( A1 => regs(959), A2 => n42, ZN => n1099);
   U1682 : AOI22_X1 port map( A1 => n84, A2 => regs(1471), B1 => n29, B2 => 
                           regs(447), ZN => n1098);
   U1683 : AOI22_X1 port map( A1 => n110, A2 => regs(2495), B1 => n66, B2 => 
                           regs(1983), ZN => n1097);
   U1684 : NAND3_X1 port map( A1 => n1099, A2 => n1098, A3 => n1097, ZN => 
                           curr_proc_regs(447));
   U1685 : NAND2_X1 port map( A1 => regs(960), A2 => n3, ZN => n1102);
   U1686 : AOI22_X1 port map( A1 => n81, A2 => regs(1472), B1 => n30, B2 => 
                           regs(448), ZN => n1101);
   U1687 : AOI22_X1 port map( A1 => n111, A2 => regs(2496), B1 => n66, B2 => 
                           regs(1984), ZN => n1100);
   U1688 : NAND3_X1 port map( A1 => n1102, A2 => n1101, A3 => n1100, ZN => 
                           curr_proc_regs(448));
   U1689 : NAND2_X1 port map( A1 => regs(961), A2 => n45, ZN => n1105);
   U1690 : AOI22_X1 port map( A1 => n80, A2 => regs(1473), B1 => n32, B2 => 
                           regs(449), ZN => n1104);
   U1691 : AOI22_X1 port map( A1 => n112, A2 => regs(2497), B1 => n66, B2 => 
                           regs(1985), ZN => n1103);
   U1692 : NAND3_X1 port map( A1 => n1105, A2 => n1104, A3 => n1103, ZN => 
                           curr_proc_regs(449));
   U1693 : INV_X1 port map( A => regs(556), ZN => n1447);
   U1694 : AOI22_X1 port map( A1 => n113, A2 => regs(2092), B1 => n66, B2 => 
                           regs(1580), ZN => n1107);
   U1695 : AOI22_X1 port map( A1 => n85, A2 => regs(1068), B1 => n35, B2 => 
                           regs(44), ZN => n1106);
   U1696 : OAI211_X1 port map( C1 => n9, C2 => n1447, A => n1107, B => n1106, 
                           ZN => curr_proc_regs(44));
   U1697 : NAND2_X1 port map( A1 => regs(962), A2 => n56, ZN => n1110);
   U1698 : AOI22_X1 port map( A1 => n86, A2 => regs(1474), B1 => n39, B2 => 
                           regs(450), ZN => n1109);
   U1699 : AOI22_X1 port map( A1 => n110, A2 => regs(2498), B1 => n66, B2 => 
                           regs(1986), ZN => n1108);
   U1700 : NAND3_X1 port map( A1 => n1110, A2 => n1109, A3 => n1108, ZN => 
                           curr_proc_regs(450));
   U1701 : NAND2_X1 port map( A1 => regs(1475), A2 => n91, ZN => n1113);
   U1702 : AOI22_X1 port map( A1 => n54, A2 => regs(963), B1 => n38, B2 => 
                           regs(451), ZN => n1112);
   U1703 : AOI22_X1 port map( A1 => n110, A2 => regs(2499), B1 => n66, B2 => 
                           regs(1987), ZN => n1111);
   U1704 : NAND3_X1 port map( A1 => n1113, A2 => n1112, A3 => n1111, ZN => 
                           curr_proc_regs(451));
   U1705 : NAND2_X1 port map( A1 => regs(1476), A2 => n91, ZN => n1116);
   U1706 : AOI22_X1 port map( A1 => n54, A2 => regs(964), B1 => n37, B2 => 
                           regs(452), ZN => n1115);
   U1707 : AOI22_X1 port map( A1 => n110, A2 => regs(2500), B1 => n66, B2 => 
                           regs(1988), ZN => n1114);
   U1708 : NAND3_X1 port map( A1 => n1116, A2 => n1115, A3 => n1114, ZN => 
                           curr_proc_regs(452));
   U1709 : NAND2_X1 port map( A1 => regs(1477), A2 => n91, ZN => n1119);
   U1710 : AOI22_X1 port map( A1 => n3, A2 => regs(965), B1 => n36, B2 => 
                           regs(453), ZN => n1118);
   U1711 : AOI22_X1 port map( A1 => n111, A2 => regs(2501), B1 => n66, B2 => 
                           regs(1989), ZN => n1117);
   U1712 : NAND3_X1 port map( A1 => n1119, A2 => n1118, A3 => n1117, ZN => 
                           curr_proc_regs(453));
   U1713 : NAND2_X1 port map( A1 => regs(1478), A2 => n91, ZN => n1122);
   U1714 : AOI22_X1 port map( A1 => n56, A2 => regs(966), B1 => n34, B2 => 
                           regs(454), ZN => n1121);
   U1715 : AOI22_X1 port map( A1 => n112, A2 => regs(2502), B1 => n66, B2 => 
                           regs(1990), ZN => n1120);
   U1716 : NAND3_X1 port map( A1 => n1122, A2 => n1121, A3 => n1120, ZN => 
                           curr_proc_regs(454));
   U1717 : NAND2_X1 port map( A1 => regs(967), A2 => n45, ZN => n1125);
   U1718 : AOI22_X1 port map( A1 => n87, A2 => regs(1479), B1 => n33, B2 => 
                           regs(455), ZN => n1124);
   U1719 : AOI22_X1 port map( A1 => n113, A2 => regs(2503), B1 => n66, B2 => 
                           regs(1991), ZN => n1123);
   U1720 : NAND3_X1 port map( A1 => n1125, A2 => n1124, A3 => n1123, ZN => 
                           curr_proc_regs(455));
   U1721 : NAND2_X1 port map( A1 => regs(968), A2 => n8, ZN => n1128);
   U1722 : AOI22_X1 port map( A1 => n80, A2 => regs(1480), B1 => n31, B2 => 
                           regs(456), ZN => n1127);
   U1723 : AOI22_X1 port map( A1 => n111, A2 => regs(2504), B1 => n66, B2 => 
                           regs(1992), ZN => n1126);
   U1724 : NAND3_X1 port map( A1 => n1128, A2 => n1127, A3 => n1126, ZN => 
                           curr_proc_regs(456));
   U1725 : NAND2_X1 port map( A1 => regs(1481), A2 => n92, ZN => n1131);
   U1726 : AOI22_X1 port map( A1 => n1, A2 => regs(969), B1 => n25, B2 => 
                           regs(457), ZN => n1130);
   U1727 : AOI22_X1 port map( A1 => n111, A2 => regs(2505), B1 => n67, B2 => 
                           regs(1993), ZN => n1129);
   U1728 : NAND3_X1 port map( A1 => n1131, A2 => n1130, A3 => n1129, ZN => 
                           curr_proc_regs(457));
   U1729 : NAND2_X1 port map( A1 => regs(1482), A2 => n92, ZN => n1134);
   U1730 : AOI22_X1 port map( A1 => n1, A2 => regs(970), B1 => n30, B2 => 
                           regs(458), ZN => n1133);
   U1731 : AOI22_X1 port map( A1 => n112, A2 => regs(2506), B1 => n67, B2 => 
                           regs(1994), ZN => n1132);
   U1732 : NAND3_X1 port map( A1 => n1134, A2 => n1133, A3 => n1132, ZN => 
                           curr_proc_regs(458));
   U1733 : NAND2_X1 port map( A1 => regs(1483), A2 => n92, ZN => n1137);
   U1734 : AOI22_X1 port map( A1 => n8, A2 => regs(971), B1 => n32, B2 => 
                           regs(459), ZN => n1136);
   U1735 : AOI22_X1 port map( A1 => n113, A2 => regs(2507), B1 => n67, B2 => 
                           regs(1995), ZN => n1135);
   U1736 : NAND3_X1 port map( A1 => n1137, A2 => n1136, A3 => n1135, ZN => 
                           curr_proc_regs(459));
   U1737 : INV_X1 port map( A => regs(557), ZN => n1450);
   U1738 : AOI22_X1 port map( A1 => n112, A2 => regs(2093), B1 => n67, B2 => 
                           regs(1581), ZN => n1139);
   U1739 : AOI22_X1 port map( A1 => n84, A2 => regs(1069), B1 => n38, B2 => 
                           regs(45), ZN => n1138);
   U1740 : OAI211_X1 port map( C1 => n2201, C2 => n1450, A => n1139, B => n1138
                           , ZN => curr_proc_regs(45));
   U1741 : NAND2_X1 port map( A1 => regs(1484), A2 => n92, ZN => n1142);
   U1742 : AOI22_X1 port map( A1 => n43, A2 => regs(972), B1 => n34, B2 => 
                           regs(460), ZN => n1141);
   U1743 : AOI22_X1 port map( A1 => n110, A2 => regs(2508), B1 => n67, B2 => 
                           regs(1996), ZN => n1140);
   U1744 : NAND3_X1 port map( A1 => n1142, A2 => n1141, A3 => n1140, ZN => 
                           curr_proc_regs(460));
   U1745 : NAND2_X1 port map( A1 => regs(973), A2 => n1, ZN => n1145);
   U1746 : AOI22_X1 port map( A1 => n84, A2 => regs(1485), B1 => n28, B2 => 
                           regs(461), ZN => n1144);
   U1747 : AOI22_X1 port map( A1 => n111, A2 => regs(2509), B1 => n67, B2 => 
                           regs(1997), ZN => n1143);
   U1748 : NAND3_X1 port map( A1 => n1145, A2 => n1144, A3 => n1143, ZN => 
                           curr_proc_regs(461));
   U1749 : NAND2_X1 port map( A1 => regs(974), A2 => n1, ZN => n1148);
   U1750 : AOI22_X1 port map( A1 => n86, A2 => regs(1486), B1 => n29, B2 => 
                           regs(462), ZN => n1147);
   U1751 : AOI22_X1 port map( A1 => n112, A2 => regs(2510), B1 => n67, B2 => 
                           regs(1998), ZN => n1146);
   U1752 : NAND3_X1 port map( A1 => n1148, A2 => n1147, A3 => n1146, ZN => 
                           curr_proc_regs(462));
   U1753 : NAND2_X1 port map( A1 => regs(975), A2 => n56, ZN => n1151);
   U1754 : AOI22_X1 port map( A1 => n82, A2 => regs(1487), B1 => n30, B2 => 
                           regs(463), ZN => n1150);
   U1755 : AOI22_X1 port map( A1 => n113, A2 => regs(2511), B1 => n67, B2 => 
                           regs(1999), ZN => n1149);
   U1756 : NAND3_X1 port map( A1 => n1151, A2 => n1150, A3 => n1149, ZN => 
                           curr_proc_regs(463));
   U1757 : NAND2_X1 port map( A1 => regs(1488), A2 => n95, ZN => n1154);
   U1758 : AOI22_X1 port map( A1 => n55, A2 => regs(976), B1 => n32, B2 => 
                           regs(464), ZN => n1153);
   U1759 : AOI22_X1 port map( A1 => n113, A2 => regs(2512), B1 => n67, B2 => 
                           regs(2000), ZN => n1152);
   U1760 : NAND3_X1 port map( A1 => n1154, A2 => n1153, A3 => n1152, ZN => 
                           curr_proc_regs(464));
   U1761 : NAND2_X1 port map( A1 => regs(977), A2 => n44, ZN => n1157);
   U1762 : AOI22_X1 port map( A1 => n84, A2 => regs(1489), B1 => n35, B2 => 
                           regs(465), ZN => n1156);
   U1763 : AOI22_X1 port map( A1 => n110, A2 => regs(2513), B1 => n67, B2 => 
                           regs(2001), ZN => n1155);
   U1764 : NAND3_X1 port map( A1 => n1157, A2 => n1156, A3 => n1155, ZN => 
                           curr_proc_regs(465));
   U1765 : NAND2_X1 port map( A1 => regs(1490), A2 => n92, ZN => n1160);
   U1766 : AOI22_X1 port map( A1 => n55, A2 => regs(978), B1 => n39, B2 => 
                           regs(466), ZN => n1159);
   U1767 : AOI22_X1 port map( A1 => n111, A2 => regs(2514), B1 => n67, B2 => 
                           regs(2002), ZN => n1158);
   U1768 : NAND3_X1 port map( A1 => n1160, A2 => n1159, A3 => n1158, ZN => 
                           curr_proc_regs(466));
   U1769 : NAND2_X1 port map( A1 => regs(979), A2 => n45, ZN => n1163);
   U1770 : AOI22_X1 port map( A1 => n81, A2 => regs(1491), B1 => n38, B2 => 
                           regs(467), ZN => n1162);
   U1771 : AOI22_X1 port map( A1 => n112, A2 => regs(2515), B1 => n67, B2 => 
                           regs(2003), ZN => n1161);
   U1772 : NAND3_X1 port map( A1 => n1163, A2 => n1162, A3 => n1161, ZN => 
                           curr_proc_regs(467));
   U1773 : NAND2_X1 port map( A1 => regs(1492), A2 => n91, ZN => n1166);
   U1774 : AOI22_X1 port map( A1 => n55, A2 => regs(980), B1 => n19, B2 => 
                           regs(468), ZN => n1165);
   U1775 : AOI22_X1 port map( A1 => n113, A2 => regs(2516), B1 => n73, B2 => 
                           regs(2004), ZN => n1164);
   U1776 : NAND3_X1 port map( A1 => n1166, A2 => n1165, A3 => n1164, ZN => 
                           curr_proc_regs(468));
   U1777 : NAND2_X1 port map( A1 => regs(981), A2 => n1, ZN => n1169);
   U1778 : AOI22_X1 port map( A1 => n87, A2 => regs(1493), B1 => n19, B2 => 
                           regs(469), ZN => n1168);
   U1779 : AOI22_X1 port map( A1 => n110, A2 => regs(2517), B1 => n71, B2 => 
                           regs(2005), ZN => n1167);
   U1780 : NAND3_X1 port map( A1 => n1169, A2 => n1168, A3 => n1167, ZN => 
                           curr_proc_regs(469));
   U1781 : INV_X1 port map( A => regs(558), ZN => n1453);
   U1782 : AOI22_X1 port map( A1 => n111, A2 => regs(2094), B1 => n72, B2 => 
                           regs(1582), ZN => n1171);
   U1783 : AOI22_X1 port map( A1 => n85, A2 => regs(1070), B1 => n19, B2 => 
                           regs(46), ZN => n1170);
   U1784 : OAI211_X1 port map( C1 => n2201, C2 => n1453, A => n1171, B => n1170
                           , ZN => curr_proc_regs(46));
   U1785 : NAND2_X1 port map( A1 => regs(982), A2 => n54, ZN => n1174);
   U1786 : AOI22_X1 port map( A1 => n81, A2 => regs(1494), B1 => n19, B2 => 
                           regs(470), ZN => n1173);
   U1787 : AOI22_X1 port map( A1 => n112, A2 => regs(2518), B1 => n69, B2 => 
                           regs(2006), ZN => n1172);
   U1788 : NAND3_X1 port map( A1 => n1174, A2 => n1173, A3 => n1172, ZN => 
                           curr_proc_regs(470));
   U1789 : NAND2_X1 port map( A1 => regs(1495), A2 => n89, ZN => n1177);
   U1790 : AOI22_X1 port map( A1 => n55, A2 => regs(983), B1 => n19, B2 => 
                           regs(471), ZN => n1176);
   U1791 : AOI22_X1 port map( A1 => n113, A2 => regs(2519), B1 => n66, B2 => 
                           regs(2007), ZN => n1175);
   U1792 : NAND3_X1 port map( A1 => n1177, A2 => n1176, A3 => n1175, ZN => 
                           curr_proc_regs(471));
   U1793 : NAND2_X1 port map( A1 => regs(1496), A2 => n95, ZN => n1180);
   U1794 : AOI22_X1 port map( A1 => n55, A2 => regs(984), B1 => n19, B2 => 
                           regs(472), ZN => n1179);
   U1795 : AOI22_X1 port map( A1 => n110, A2 => regs(2520), B1 => n5, B2 => 
                           regs(2008), ZN => n1178);
   U1796 : NAND3_X1 port map( A1 => n1180, A2 => n1179, A3 => n1178, ZN => 
                           curr_proc_regs(472));
   U1797 : NAND2_X1 port map( A1 => regs(985), A2 => n55, ZN => n1183);
   U1798 : AOI22_X1 port map( A1 => n81, A2 => regs(1497), B1 => n19, B2 => 
                           regs(473), ZN => n1182);
   U1799 : AOI22_X1 port map( A1 => n111, A2 => regs(2521), B1 => n74, B2 => 
                           regs(2009), ZN => n1181);
   U1800 : NAND3_X1 port map( A1 => n1183, A2 => n1182, A3 => n1181, ZN => 
                           curr_proc_regs(473));
   U1801 : NAND2_X1 port map( A1 => regs(986), A2 => n41, ZN => n1186);
   U1802 : AOI22_X1 port map( A1 => n82, A2 => regs(1498), B1 => n19, B2 => 
                           regs(474), ZN => n1185);
   U1803 : AOI22_X1 port map( A1 => n112, A2 => regs(2522), B1 => n74, B2 => 
                           regs(2010), ZN => n1184);
   U1804 : NAND3_X1 port map( A1 => n1186, A2 => n1185, A3 => n1184, ZN => 
                           curr_proc_regs(474));
   U1805 : NAND2_X1 port map( A1 => regs(1499), A2 => n91, ZN => n1189);
   U1806 : AOI22_X1 port map( A1 => n55, A2 => regs(987), B1 => n19, B2 => 
                           regs(475), ZN => n1188);
   U1807 : AOI22_X1 port map( A1 => n113, A2 => regs(2523), B1 => n5, B2 => 
                           regs(2011), ZN => n1187);
   U1808 : NAND3_X1 port map( A1 => n1189, A2 => n1188, A3 => n1187, ZN => 
                           curr_proc_regs(475));
   U1809 : NAND2_X1 port map( A1 => regs(1500), A2 => n93, ZN => n1192);
   U1810 : AOI22_X1 port map( A1 => n54, A2 => regs(988), B1 => n19, B2 => 
                           regs(476), ZN => n1191);
   U1811 : AOI22_X1 port map( A1 => n110, A2 => regs(2524), B1 => n68, B2 => 
                           regs(2012), ZN => n1190);
   U1812 : NAND3_X1 port map( A1 => n1192, A2 => n1191, A3 => n1190, ZN => 
                           curr_proc_regs(476));
   U1813 : NAND2_X1 port map( A1 => regs(989), A2 => n56, ZN => n1195);
   U1814 : AOI22_X1 port map( A1 => n81, A2 => regs(1501), B1 => n19, B2 => 
                           regs(477), ZN => n1194);
   U1815 : AOI22_X1 port map( A1 => n111, A2 => regs(2525), B1 => n5, B2 => 
                           regs(2013), ZN => n1193);
   U1816 : NAND3_X1 port map( A1 => n1195, A2 => n1194, A3 => n1193, ZN => 
                           curr_proc_regs(477));
   U1817 : NAND2_X1 port map( A1 => regs(990), A2 => n8, ZN => n1198);
   U1818 : AOI22_X1 port map( A1 => n80, A2 => regs(1502), B1 => n19, B2 => 
                           regs(478), ZN => n1197);
   U1819 : AOI22_X1 port map( A1 => n112, A2 => regs(2526), B1 => n74, B2 => 
                           regs(2014), ZN => n1196);
   U1820 : NAND3_X1 port map( A1 => n1198, A2 => n1197, A3 => n1196, ZN => 
                           curr_proc_regs(478));
   U1821 : NAND2_X1 port map( A1 => regs(991), A2 => n1, ZN => n1201);
   U1822 : AOI22_X1 port map( A1 => n85, A2 => regs(1503), B1 => n20, B2 => 
                           regs(479), ZN => n1200);
   U1823 : AOI22_X1 port map( A1 => n113, A2 => regs(2527), B1 => n72, B2 => 
                           regs(2015), ZN => n1199);
   U1824 : NAND3_X1 port map( A1 => n1201, A2 => n1200, A3 => n1199, ZN => 
                           curr_proc_regs(479));
   U1825 : INV_X1 port map( A => regs(559), ZN => n1456);
   U1826 : AOI22_X1 port map( A1 => n113, A2 => regs(2095), B1 => n71, B2 => 
                           regs(1583), ZN => n1203);
   U1827 : AOI22_X1 port map( A1 => n86, A2 => regs(1071), B1 => n20, B2 => 
                           regs(47), ZN => n1202);
   U1828 : OAI211_X1 port map( C1 => n57, C2 => n1456, A => n1203, B => n1202, 
                           ZN => curr_proc_regs(47));
   U1829 : NAND2_X1 port map( A1 => regs(992), A2 => n3, ZN => n1206);
   U1830 : AOI22_X1 port map( A1 => n87, A2 => regs(1504), B1 => n20, B2 => 
                           regs(480), ZN => n1205);
   U1831 : AOI22_X1 port map( A1 => n113, A2 => regs(2528), B1 => n63, B2 => 
                           regs(2016), ZN => n1204);
   U1832 : NAND3_X1 port map( A1 => n1206, A2 => n1205, A3 => n1204, ZN => 
                           curr_proc_regs(480));
   U1833 : NAND2_X1 port map( A1 => regs(1505), A2 => n93, ZN => n1209);
   U1834 : AOI22_X1 port map( A1 => n8, A2 => regs(993), B1 => n20, B2 => 
                           regs(481), ZN => n1208);
   U1835 : AOI22_X1 port map( A1 => n113, A2 => regs(2529), B1 => n70, B2 => 
                           regs(2017), ZN => n1207);
   U1836 : NAND3_X1 port map( A1 => n1209, A2 => n1208, A3 => n1207, ZN => 
                           curr_proc_regs(481));
   U1837 : NAND2_X1 port map( A1 => regs(1506), A2 => n93, ZN => n1212);
   U1838 : AOI22_X1 port map( A1 => n1, A2 => regs(994), B1 => n20, B2 => 
                           regs(482), ZN => n1211);
   U1839 : AOI22_X1 port map( A1 => n113, A2 => regs(2530), B1 => n65, B2 => 
                           regs(2018), ZN => n1210);
   U1840 : NAND3_X1 port map( A1 => n1212, A2 => n1211, A3 => n1210, ZN => 
                           curr_proc_regs(482));
   U1841 : NAND2_X1 port map( A1 => regs(995), A2 => n3, ZN => n1215);
   U1842 : AOI22_X1 port map( A1 => n86, A2 => regs(1507), B1 => n20, B2 => 
                           regs(483), ZN => n1214);
   U1843 : AOI22_X1 port map( A1 => n113, A2 => regs(2531), B1 => n73, B2 => 
                           regs(2019), ZN => n1213);
   U1844 : NAND3_X1 port map( A1 => n1215, A2 => n1214, A3 => n1213, ZN => 
                           curr_proc_regs(483));
   U1845 : NAND2_X1 port map( A1 => regs(996), A2 => n8, ZN => n1218);
   U1846 : AOI22_X1 port map( A1 => n80, A2 => regs(1508), B1 => n20, B2 => 
                           regs(484), ZN => n1217);
   U1847 : AOI22_X1 port map( A1 => n113, A2 => regs(2532), B1 => n66, B2 => 
                           regs(2020), ZN => n1216);
   U1848 : NAND3_X1 port map( A1 => n1218, A2 => n1217, A3 => n1216, ZN => 
                           curr_proc_regs(484));
   U1849 : NAND2_X1 port map( A1 => regs(997), A2 => n3, ZN => n1221);
   U1850 : AOI22_X1 port map( A1 => n85, A2 => regs(1509), B1 => n20, B2 => 
                           regs(485), ZN => n1220);
   U1851 : AOI22_X1 port map( A1 => n113, A2 => regs(2533), B1 => n68, B2 => 
                           regs(2021), ZN => n1219);
   U1852 : NAND3_X1 port map( A1 => n1221, A2 => n1220, A3 => n1219, ZN => 
                           curr_proc_regs(485));
   U1853 : NAND2_X1 port map( A1 => regs(998), A2 => n8, ZN => n1224);
   U1854 : AOI22_X1 port map( A1 => n86, A2 => regs(1510), B1 => n20, B2 => 
                           regs(486), ZN => n1223);
   U1855 : AOI22_X1 port map( A1 => n113, A2 => regs(2534), B1 => n72, B2 => 
                           regs(2022), ZN => n1222);
   U1856 : NAND3_X1 port map( A1 => n1224, A2 => n1223, A3 => n1222, ZN => 
                           curr_proc_regs(486));
   U1857 : NAND2_X1 port map( A1 => regs(1511), A2 => n93, ZN => n1227);
   U1858 : AOI22_X1 port map( A1 => n53, A2 => regs(999), B1 => n20, B2 => 
                           regs(487), ZN => n1226);
   U1859 : AOI22_X1 port map( A1 => n113, A2 => regs(2535), B1 => n73, B2 => 
                           regs(2023), ZN => n1225);
   U1860 : NAND3_X1 port map( A1 => n1227, A2 => n1226, A3 => n1225, ZN => 
                           curr_proc_regs(487));
   U1861 : NAND2_X1 port map( A1 => regs(1000), A2 => n1, ZN => n1230);
   U1862 : AOI22_X1 port map( A1 => n87, A2 => regs(1512), B1 => n20, B2 => 
                           regs(488), ZN => n1229);
   U1863 : AOI22_X1 port map( A1 => n113, A2 => regs(2536), B1 => n66, B2 => 
                           regs(2024), ZN => n1228);
   U1864 : NAND3_X1 port map( A1 => n1230, A2 => n1229, A3 => n1228, ZN => 
                           curr_proc_regs(488));
   U1865 : NAND2_X1 port map( A1 => regs(1513), A2 => n94, ZN => n1233);
   U1866 : AOI22_X1 port map( A1 => n1, A2 => regs(1001), B1 => n20, B2 => 
                           regs(489), ZN => n1232);
   U1867 : AOI22_X1 port map( A1 => n113, A2 => regs(2537), B1 => n5, B2 => 
                           regs(2025), ZN => n1231);
   U1868 : NAND3_X1 port map( A1 => n1233, A2 => n1232, A3 => n1231, ZN => 
                           curr_proc_regs(489));
   U1869 : INV_X1 port map( A => regs(560), ZN => n1461);
   U1870 : AOI22_X1 port map( A1 => n113, A2 => regs(2096), B1 => n68, B2 => 
                           regs(1584), ZN => n1235);
   U1871 : AOI22_X1 port map( A1 => n87, A2 => regs(1072), B1 => n24, B2 => 
                           regs(48), ZN => n1234);
   U1872 : OAI211_X1 port map( C1 => n57, C2 => n1461, A => n1235, B => n1234, 
                           ZN => curr_proc_regs(48));
   U1873 : NAND2_X1 port map( A1 => regs(1002), A2 => n1, ZN => n1238);
   U1874 : AOI22_X1 port map( A1 => n80, A2 => regs(1514), B1 => n17, B2 => 
                           regs(490), ZN => n1237);
   U1875 : AOI22_X1 port map( A1 => n112, A2 => regs(2538), B1 => n68, B2 => 
                           regs(2026), ZN => n1236);
   U1876 : NAND3_X1 port map( A1 => n1238, A2 => n1237, A3 => n1236, ZN => 
                           curr_proc_regs(490));
   U1877 : NAND2_X1 port map( A1 => regs(1003), A2 => n1, ZN => n1241);
   U1878 : AOI22_X1 port map( A1 => n82, A2 => regs(1515), B1 => n18, B2 => 
                           regs(491), ZN => n1240);
   U1879 : AOI22_X1 port map( A1 => n112, A2 => regs(2539), B1 => n68, B2 => 
                           regs(2027), ZN => n1239);
   U1880 : NAND3_X1 port map( A1 => n1241, A2 => n1240, A3 => n1239, ZN => 
                           curr_proc_regs(491));
   U1881 : NAND2_X1 port map( A1 => regs(1516), A2 => n94, ZN => n1244);
   U1882 : AOI22_X1 port map( A1 => n55, A2 => regs(1004), B1 => n19, B2 => 
                           regs(492), ZN => n1243);
   U1883 : AOI22_X1 port map( A1 => n112, A2 => regs(2540), B1 => n68, B2 => 
                           regs(2028), ZN => n1242);
   U1884 : NAND3_X1 port map( A1 => n1244, A2 => n1243, A3 => n1242, ZN => 
                           curr_proc_regs(492));
   U1885 : NAND2_X1 port map( A1 => regs(1517), A2 => n94, ZN => n1247);
   U1886 : AOI22_X1 port map( A1 => n55, A2 => regs(1005), B1 => n27, B2 => 
                           regs(493), ZN => n1246);
   U1887 : AOI22_X1 port map( A1 => n112, A2 => regs(2541), B1 => n68, B2 => 
                           regs(2029), ZN => n1245);
   U1888 : NAND3_X1 port map( A1 => n1247, A2 => n1246, A3 => n1245, ZN => 
                           curr_proc_regs(493));
   U1889 : NAND2_X1 port map( A1 => regs(1518), A2 => n94, ZN => n1250);
   U1890 : AOI22_X1 port map( A1 => n43, A2 => regs(1006), B1 => n26, B2 => 
                           regs(494), ZN => n1249);
   U1891 : AOI22_X1 port map( A1 => n112, A2 => regs(2542), B1 => n68, B2 => 
                           regs(2030), ZN => n1248);
   U1892 : NAND3_X1 port map( A1 => n1250, A2 => n1249, A3 => n1248, ZN => 
                           curr_proc_regs(494));
   U1893 : NAND2_X1 port map( A1 => regs(1519), A2 => n94, ZN => n1253);
   U1894 : AOI22_X1 port map( A1 => n45, A2 => regs(1007), B1 => n25, B2 => 
                           regs(495), ZN => n1252);
   U1895 : AOI22_X1 port map( A1 => n112, A2 => regs(2543), B1 => n68, B2 => 
                           regs(2031), ZN => n1251);
   U1896 : NAND3_X1 port map( A1 => n1253, A2 => n1252, A3 => n1251, ZN => 
                           curr_proc_regs(495));
   U1897 : NAND2_X1 port map( A1 => regs(1008), A2 => n54, ZN => n1256);
   U1898 : AOI22_X1 port map( A1 => n84, A2 => regs(1520), B1 => n38, B2 => 
                           regs(496), ZN => n1255);
   U1899 : AOI22_X1 port map( A1 => n112, A2 => regs(2544), B1 => n68, B2 => 
                           regs(2032), ZN => n1254);
   U1900 : NAND3_X1 port map( A1 => n1256, A2 => n1255, A3 => n1254, ZN => 
                           curr_proc_regs(496));
   U1901 : NAND2_X1 port map( A1 => regs(1009), A2 => n41, ZN => n1259);
   U1902 : AOI22_X1 port map( A1 => n81, A2 => regs(1521), B1 => n38, B2 => 
                           regs(497), ZN => n1258);
   U1903 : AOI22_X1 port map( A1 => n112, A2 => regs(2545), B1 => n68, B2 => 
                           regs(2033), ZN => n1257);
   U1904 : NAND3_X1 port map( A1 => n1259, A2 => n1258, A3 => n1257, ZN => 
                           curr_proc_regs(497));
   U1905 : NAND2_X1 port map( A1 => regs(1010), A2 => n1, ZN => n1262);
   U1906 : AOI22_X1 port map( A1 => n80, A2 => regs(1522), B1 => n36, B2 => 
                           regs(498), ZN => n1261);
   U1907 : AOI22_X1 port map( A1 => n112, A2 => regs(2546), B1 => n68, B2 => 
                           regs(2034), ZN => n1260);
   U1908 : NAND3_X1 port map( A1 => n1262, A2 => n1261, A3 => n1260, ZN => 
                           curr_proc_regs(498));
   U1909 : NAND2_X1 port map( A1 => regs(1523), A2 => n95, ZN => n1265);
   U1910 : AOI22_X1 port map( A1 => n44, A2 => regs(1011), B1 => n33, B2 => 
                           regs(499), ZN => n1264);
   U1911 : AOI22_X1 port map( A1 => n112, A2 => regs(2547), B1 => n68, B2 => 
                           regs(2035), ZN => n1263);
   U1912 : NAND3_X1 port map( A1 => n1265, A2 => n1264, A3 => n1263, ZN => 
                           curr_proc_regs(499));
   U1913 : INV_X1 port map( A => regs(1073), ZN => n1464);
   U1914 : AOI22_X1 port map( A1 => n112, A2 => regs(2097), B1 => n68, B2 => 
                           regs(1585), ZN => n1267);
   U1915 : AOI22_X1 port map( A1 => n45, A2 => regs(561), B1 => n20, B2 => 
                           regs(49), ZN => n1266);
   U1916 : OAI211_X1 port map( C1 => n2215, C2 => n1464, A => n1267, B => n1266
                           , ZN => curr_proc_regs(49));
   U1917 : INV_X1 port map( A => regs(1028), ZN => n1322);
   U1918 : AOI22_X1 port map( A1 => n112, A2 => regs(2052), B1 => n67, B2 => 
                           regs(1540), ZN => n1269);
   U1919 : AOI22_X1 port map( A1 => n3, A2 => regs(516), B1 => n23, B2 => 
                           regs(4), ZN => n1268);
   U1920 : OAI211_X1 port map( C1 => n2215, C2 => n1322, A => n1269, B => n1268
                           , ZN => curr_proc_regs(4));
   U1921 : NAND2_X1 port map( A1 => regs(1012), A2 => n1, ZN => n1272);
   U1922 : AOI22_X1 port map( A1 => n85, A2 => regs(1524), B1 => n26, B2 => 
                           regs(500), ZN => n1271);
   U1923 : AOI22_X1 port map( A1 => n111, A2 => regs(2548), B1 => n71, B2 => 
                           regs(2036), ZN => n1270);
   U1924 : NAND3_X1 port map( A1 => n1272, A2 => n1271, A3 => n1270, ZN => 
                           curr_proc_regs(500));
   U1925 : NAND2_X1 port map( A1 => regs(1525), A2 => n95, ZN => n1275);
   U1926 : AOI22_X1 port map( A1 => n47, A2 => regs(1013), B1 => n28, B2 => 
                           regs(501), ZN => n1274);
   U1927 : AOI22_X1 port map( A1 => n111, A2 => regs(2549), B1 => n67, B2 => 
                           regs(2037), ZN => n1273);
   U1928 : NAND3_X1 port map( A1 => n1275, A2 => n1274, A3 => n1273, ZN => 
                           curr_proc_regs(501));
   U1929 : NAND2_X1 port map( A1 => regs(1526), A2 => n96, ZN => n1278);
   U1930 : AOI22_X1 port map( A1 => n8, A2 => regs(1014), B1 => n20, B2 => 
                           regs(502), ZN => n1277);
   U1931 : AOI22_X1 port map( A1 => n111, A2 => regs(2550), B1 => n5, B2 => 
                           regs(2038), ZN => n1276);
   U1932 : NAND3_X1 port map( A1 => n1278, A2 => n1277, A3 => n1276, ZN => 
                           curr_proc_regs(502));
   U1933 : NAND2_X1 port map( A1 => regs(1527), A2 => n96, ZN => n1281);
   U1934 : AOI22_X1 port map( A1 => n8, A2 => regs(1015), B1 => n28, B2 => 
                           regs(503), ZN => n1280);
   U1935 : AOI22_X1 port map( A1 => n111, A2 => regs(2551), B1 => n67, B2 => 
                           regs(2039), ZN => n1279);
   U1936 : NAND3_X1 port map( A1 => n1281, A2 => n1280, A3 => n1279, ZN => 
                           curr_proc_regs(503));
   U1937 : NAND2_X1 port map( A1 => regs(1528), A2 => n96, ZN => n1284);
   U1938 : AOI22_X1 port map( A1 => n8, A2 => regs(1016), B1 => n29, B2 => 
                           regs(504), ZN => n1283);
   U1939 : AOI22_X1 port map( A1 => n111, A2 => regs(2552), B1 => n72, B2 => 
                           regs(2040), ZN => n1282);
   U1940 : NAND3_X1 port map( A1 => n1284, A2 => n1283, A3 => n1282, ZN => 
                           curr_proc_regs(504));
   U1941 : NAND2_X1 port map( A1 => regs(1017), A2 => n8, ZN => n1287);
   U1942 : AOI22_X1 port map( A1 => n86, A2 => regs(1529), B1 => n30, B2 => 
                           regs(505), ZN => n1286);
   U1943 : AOI22_X1 port map( A1 => n111, A2 => regs(2553), B1 => n67, B2 => 
                           regs(2041), ZN => n1285);
   U1944 : NAND3_X1 port map( A1 => n1287, A2 => n1286, A3 => n1285, ZN => 
                           curr_proc_regs(505));
   U1945 : NAND2_X1 port map( A1 => regs(1018), A2 => n55, ZN => n1290);
   U1946 : AOI22_X1 port map( A1 => n85, A2 => regs(1530), B1 => n32, B2 => 
                           regs(506), ZN => n1289);
   U1947 : AOI22_X1 port map( A1 => n111, A2 => regs(2554), B1 => n69, B2 => 
                           regs(2042), ZN => n1288);
   U1948 : NAND3_X1 port map( A1 => n1290, A2 => n1289, A3 => n1288, ZN => 
                           curr_proc_regs(506));
   U1949 : NAND2_X1 port map( A1 => regs(1531), A2 => n96, ZN => n1293);
   U1950 : AOI22_X1 port map( A1 => n8, A2 => regs(1019), B1 => n35, B2 => 
                           regs(507), ZN => n1292);
   U1951 : AOI22_X1 port map( A1 => n111, A2 => regs(2555), B1 => n67, B2 => 
                           regs(2043), ZN => n1291);
   U1952 : NAND3_X1 port map( A1 => n1293, A2 => n1292, A3 => n1291, ZN => 
                           curr_proc_regs(507));
   U1953 : NAND2_X1 port map( A1 => regs(1020), A2 => n43, ZN => n1296);
   U1954 : AOI22_X1 port map( A1 => n86, A2 => regs(1532), B1 => n39, B2 => 
                           regs(508), ZN => n1295);
   U1955 : AOI22_X1 port map( A1 => n111, A2 => regs(2556), B1 => n73, B2 => 
                           regs(2044), ZN => n1294);
   U1956 : NAND3_X1 port map( A1 => n1296, A2 => n1295, A3 => n1294, ZN => 
                           curr_proc_regs(508));
   U1957 : NAND2_X1 port map( A1 => regs(1021), A2 => n55, ZN => n1299);
   U1958 : AOI22_X1 port map( A1 => n87, A2 => regs(1533), B1 => n38, B2 => 
                           regs(509), ZN => n1298);
   U1959 : AOI22_X1 port map( A1 => n111, A2 => regs(2557), B1 => n67, B2 => 
                           regs(2045), ZN => n1297);
   U1960 : NAND3_X1 port map( A1 => n1299, A2 => n1298, A3 => n1297, ZN => 
                           curr_proc_regs(509));
   U1961 : INV_X1 port map( A => regs(562), ZN => n1467);
   U1962 : AOI22_X1 port map( A1 => n111, A2 => regs(2098), B1 => n67, B2 => 
                           regs(1586), ZN => n1301);
   U1963 : AOI22_X1 port map( A1 => n82, A2 => regs(1074), B1 => n37, B2 => 
                           regs(50), ZN => n1300);
   U1964 : OAI211_X1 port map( C1 => n10, C2 => n1467, A => n1301, B => n1300, 
                           ZN => curr_proc_regs(50));
   U1965 : NAND2_X1 port map( A1 => regs(1022), A2 => n43, ZN => n1304);
   U1966 : AOI22_X1 port map( A1 => n82, A2 => regs(1534), B1 => n33, B2 => 
                           regs(510), ZN => n1303);
   U1967 : AOI22_X1 port map( A1 => n111, A2 => regs(2558), B1 => n63, B2 => 
                           regs(2046), ZN => n1302);
   U1968 : NAND3_X1 port map( A1 => n1304, A2 => n1303, A3 => n1302, ZN => 
                           curr_proc_regs(510));
   U1969 : NAND2_X1 port map( A1 => regs(1535), A2 => n96, ZN => n1307);
   U1970 : AOI22_X1 port map( A1 => n8, A2 => regs(1023), B1 => n31, B2 => 
                           regs(511), ZN => n1306);
   U1971 : AOI22_X1 port map( A1 => n110, A2 => regs(2559), B1 => n72, B2 => 
                           regs(2047), ZN => n1305);
   U1972 : NAND3_X1 port map( A1 => n1307, A2 => n1306, A3 => n1305, ZN => 
                           curr_proc_regs(511));
   U1973 : AOI22_X1 port map( A1 => n110, A2 => regs(0), B1 => n68, B2 => 
                           regs(2048), ZN => n1309);
   U1974 : AOI22_X1 port map( A1 => n43, A2 => regs(1024), B1 => n102, B2 => 
                           regs(1536), ZN => n1308);
   U1975 : OAI211_X1 port map( C1 => n1310, C2 => n2128, A => n1309, B => n1308
                           , ZN => curr_proc_regs(512));
   U1976 : AOI22_X1 port map( A1 => n110, A2 => regs(1), B1 => n68, B2 => 
                           regs(2049), ZN => n1312);
   U1977 : AOI22_X1 port map( A1 => n56, A2 => regs(1025), B1 => n101, B2 => 
                           regs(1537), ZN => n1311);
   U1978 : OAI211_X1 port map( C1 => n14, C2 => n1313, A => n1312, B => n1311, 
                           ZN => curr_proc_regs(513));
   U1979 : AOI22_X1 port map( A1 => n110, A2 => regs(2), B1 => n63, B2 => 
                           regs(2050), ZN => n1315);
   U1980 : AOI22_X1 port map( A1 => n8, A2 => regs(1026), B1 => n102, B2 => 
                           regs(1538), ZN => n1314);
   U1981 : OAI211_X1 port map( C1 => n2128, C2 => n1316, A => n1315, B => n1314
                           , ZN => curr_proc_regs(514));
   U1982 : AOI22_X1 port map( A1 => n110, A2 => regs(3), B1 => n63, B2 => 
                           regs(2051), ZN => n1318);
   U1983 : AOI22_X1 port map( A1 => n41, A2 => regs(1027), B1 => n102, B2 => 
                           regs(1539), ZN => n1317);
   U1984 : OAI211_X1 port map( C1 => n14, C2 => n1319, A => n1318, B => n1317, 
                           ZN => curr_proc_regs(515));
   U1985 : AOI22_X1 port map( A1 => n110, A2 => regs(4), B1 => n72, B2 => 
                           regs(2052), ZN => n1321);
   U1986 : AOI22_X1 port map( A1 => n84, A2 => regs(1540), B1 => n21, B2 => 
                           regs(516), ZN => n1320);
   U1987 : OAI211_X1 port map( C1 => n2201, C2 => n1322, A => n1321, B => n1320
                           , ZN => curr_proc_regs(516));
   U1988 : INV_X1 port map( A => regs(1541), ZN => n1325);
   U1989 : AOI22_X1 port map( A1 => n110, A2 => regs(5), B1 => n63, B2 => 
                           regs(2053), ZN => n1324);
   U1990 : AOI22_X1 port map( A1 => n42, A2 => regs(1029), B1 => n22, B2 => 
                           regs(517), ZN => n1323);
   U1991 : OAI211_X1 port map( C1 => n2215, C2 => n1325, A => n1324, B => n1323
                           , ZN => curr_proc_regs(517));
   U1992 : INV_X1 port map( A => regs(1030), ZN => n1908);
   U1993 : AOI22_X1 port map( A1 => n110, A2 => regs(6), B1 => n68, B2 => 
                           regs(2054), ZN => n1327);
   U1994 : AOI22_X1 port map( A1 => n81, A2 => regs(1542), B1 => n23, B2 => 
                           regs(518), ZN => n1326);
   U1995 : OAI211_X1 port map( C1 => n57, C2 => n1908, A => n1327, B => n1326, 
                           ZN => curr_proc_regs(518));
   U1996 : INV_X1 port map( A => regs(1031), ZN => n2146);
   U1997 : AOI22_X1 port map( A1 => n110, A2 => regs(7), B1 => n68, B2 => 
                           regs(2055), ZN => n1329);
   U1998 : AOI22_X1 port map( A1 => n80, A2 => regs(1543), B1 => n24, B2 => 
                           regs(519), ZN => n1328);
   U1999 : OAI211_X1 port map( C1 => n2201, C2 => n2146, A => n1329, B => n1328
                           , ZN => curr_proc_regs(519));
   U2000 : INV_X1 port map( A => regs(563), ZN => n1470);
   U2001 : AOI22_X1 port map( A1 => n110, A2 => regs(2099), B1 => n72, B2 => 
                           regs(1587), ZN => n1331);
   U2002 : AOI22_X1 port map( A1 => n85, A2 => regs(1075), B1 => n17, B2 => 
                           regs(51), ZN => n1330);
   U2003 : OAI211_X1 port map( C1 => n10, C2 => n1470, A => n1331, B => n1330, 
                           ZN => curr_proc_regs(51));
   U2004 : INV_X1 port map( A => regs(1032), ZN => n2179);
   U2005 : AOI22_X1 port map( A1 => n110, A2 => regs(8), B1 => n72, B2 => 
                           regs(2056), ZN => n1333);
   U2006 : AOI22_X1 port map( A1 => n86, A2 => regs(1544), B1 => n18, B2 => 
                           regs(520), ZN => n1332);
   U2007 : OAI211_X1 port map( C1 => n10, C2 => n2179, A => n1333, B => n1332, 
                           ZN => curr_proc_regs(520));
   U2008 : INV_X1 port map( A => regs(1545), ZN => n1336);
   U2009 : AOI22_X1 port map( A1 => n110, A2 => regs(9), B1 => n5, B2 => 
                           regs(2057), ZN => n1335);
   U2010 : AOI22_X1 port map( A1 => n56, A2 => regs(1033), B1 => n19, B2 => 
                           regs(521), ZN => n1334);
   U2011 : OAI211_X1 port map( C1 => n78, C2 => n1336, A => n1335, B => n1334, 
                           ZN => curr_proc_regs(521));
   U2012 : AOI22_X1 port map( A1 => n109, A2 => regs(10), B1 => n5, B2 => 
                           regs(2058), ZN => n1338);
   U2013 : AOI22_X1 port map( A1 => n52, A2 => regs(1034), B1 => n102, B2 => 
                           regs(1546), ZN => n1337);
   U2014 : OAI211_X1 port map( C1 => n2128, C2 => n1339, A => n1338, B => n1337
                           , ZN => curr_proc_regs(522));
   U2015 : AOI22_X1 port map( A1 => n109, A2 => regs(11), B1 => n5, B2 => 
                           regs(2059), ZN => n1341);
   U2016 : AOI22_X1 port map( A1 => n44, A2 => regs(1035), B1 => n102, B2 => 
                           regs(1547), ZN => n1340);
   U2017 : OAI211_X1 port map( C1 => n14, C2 => n1342, A => n1341, B => n1340, 
                           ZN => curr_proc_regs(523));
   U2018 : AOI22_X1 port map( A1 => n109, A2 => regs(12), B1 => n5, B2 => 
                           regs(2060), ZN => n1344);
   U2019 : AOI22_X1 port map( A1 => n53, A2 => regs(1036), B1 => n102, B2 => 
                           regs(1548), ZN => n1343);
   U2020 : OAI211_X1 port map( C1 => n14, C2 => n1345, A => n1344, B => n1343, 
                           ZN => curr_proc_regs(524));
   U2021 : AOI22_X1 port map( A1 => n109, A2 => regs(13), B1 => n5, B2 => 
                           regs(2061), ZN => n1347);
   U2022 : AOI22_X1 port map( A1 => n55, A2 => regs(1037), B1 => n102, B2 => 
                           regs(1549), ZN => n1346);
   U2023 : OAI211_X1 port map( C1 => n12, C2 => n1348, A => n1347, B => n1346, 
                           ZN => curr_proc_regs(525));
   U2024 : AOI22_X1 port map( A1 => n109, A2 => regs(14), B1 => n5, B2 => 
                           regs(2062), ZN => n1350);
   U2025 : AOI22_X1 port map( A1 => n87, A2 => regs(1550), B1 => n36, B2 => 
                           regs(526), ZN => n1349);
   U2026 : OAI211_X1 port map( C1 => n58, C2 => n1351, A => n1350, B => n1349, 
                           ZN => curr_proc_regs(526));
   U2027 : AOI22_X1 port map( A1 => n109, A2 => regs(15), B1 => n5, B2 => 
                           regs(2063), ZN => n1353);
   U2028 : AOI22_X1 port map( A1 => n84, A2 => regs(1551), B1 => n27, B2 => 
                           regs(527), ZN => n1352);
   U2029 : OAI211_X1 port map( C1 => n10, C2 => n1354, A => n1353, B => n1352, 
                           ZN => curr_proc_regs(527));
   U2030 : AOI22_X1 port map( A1 => n109, A2 => regs(16), B1 => n5, B2 => 
                           regs(2064), ZN => n1356);
   U2031 : AOI22_X1 port map( A1 => n79, A2 => regs(1552), B1 => n26, B2 => 
                           regs(528), ZN => n1355);
   U2032 : OAI211_X1 port map( C1 => n9, C2 => n1357, A => n1356, B => n1355, 
                           ZN => curr_proc_regs(528));
   U2033 : AOI22_X1 port map( A1 => n109, A2 => regs(17), B1 => n5, B2 => 
                           regs(2065), ZN => n1359);
   U2034 : AOI22_X1 port map( A1 => n79, A2 => regs(1553), B1 => n20, B2 => 
                           regs(529), ZN => n1358);
   U2035 : OAI211_X1 port map( C1 => n10, C2 => n1360, A => n1359, B => n1358, 
                           ZN => curr_proc_regs(529));
   U2036 : INV_X1 port map( A => regs(1076), ZN => n1473);
   U2037 : AOI22_X1 port map( A1 => n109, A2 => regs(2100), B1 => n5, B2 => 
                           regs(1588), ZN => n1362);
   U2038 : AOI22_X1 port map( A1 => n41, A2 => regs(564), B1 => n35, B2 => 
                           regs(52), ZN => n1361);
   U2039 : OAI211_X1 port map( C1 => n2215, C2 => n1473, A => n1362, B => n1361
                           , ZN => curr_proc_regs(52));
   U2040 : AOI22_X1 port map( A1 => n109, A2 => regs(18), B1 => n5, B2 => 
                           regs(2066), ZN => n1364);
   U2041 : AOI22_X1 port map( A1 => n79, A2 => regs(1554), B1 => n25, B2 => 
                           regs(530), ZN => n1363);
   U2042 : OAI211_X1 port map( C1 => n9, C2 => n1365, A => n1364, B => n1363, 
                           ZN => curr_proc_regs(530));
   U2043 : AOI22_X1 port map( A1 => n109, A2 => regs(19), B1 => n5, B2 => 
                           regs(2067), ZN => n1367);
   U2044 : AOI22_X1 port map( A1 => n43, A2 => regs(1043), B1 => n102, B2 => 
                           regs(1555), ZN => n1366);
   U2045 : OAI211_X1 port map( C1 => n2128, C2 => n1368, A => n1367, B => n1366
                           , ZN => curr_proc_regs(531));
   U2046 : AOI22_X1 port map( A1 => n109, A2 => regs(20), B1 => n71, B2 => 
                           regs(2068), ZN => n1370);
   U2047 : AOI22_X1 port map( A1 => n79, A2 => regs(1556), B1 => n20, B2 => 
                           regs(532), ZN => n1369);
   U2048 : OAI211_X1 port map( C1 => n10, C2 => n1371, A => n1370, B => n1369, 
                           ZN => curr_proc_regs(532));
   U2049 : AOI22_X1 port map( A1 => n106, A2 => regs(21), B1 => n69, B2 => 
                           regs(2069), ZN => n1373);
   U2050 : AOI22_X1 port map( A1 => n54, A2 => regs(1045), B1 => n102, B2 => 
                           regs(1557), ZN => n1372);
   U2051 : OAI211_X1 port map( C1 => n14, C2 => n1374, A => n1373, B => n1372, 
                           ZN => curr_proc_regs(533));
   U2052 : AOI22_X1 port map( A1 => n107, A2 => regs(22), B1 => n74, B2 => 
                           regs(2070), ZN => n1376);
   U2053 : AOI22_X1 port map( A1 => n53, A2 => regs(1046), B1 => n102, B2 => 
                           regs(1558), ZN => n1375);
   U2054 : OAI211_X1 port map( C1 => n12, C2 => n1377, A => n1376, B => n1375, 
                           ZN => curr_proc_regs(534));
   U2055 : AOI22_X1 port map( A1 => n108, A2 => regs(23), B1 => n74, B2 => 
                           regs(2071), ZN => n1379);
   U2056 : AOI22_X1 port map( A1 => n79, A2 => regs(1559), B1 => n24, B2 => 
                           regs(535), ZN => n1378);
   U2057 : OAI211_X1 port map( C1 => n9, C2 => n1380, A => n1379, B => n1378, 
                           ZN => curr_proc_regs(535));
   U2058 : AOI22_X1 port map( A1 => n109, A2 => regs(24), B1 => n69, B2 => 
                           regs(2072), ZN => n1382);
   U2059 : AOI22_X1 port map( A1 => n42, A2 => regs(1048), B1 => n102, B2 => 
                           regs(1560), ZN => n1381);
   U2060 : OAI211_X1 port map( C1 => n2128, C2 => n1383, A => n1382, B => n1381
                           , ZN => curr_proc_regs(536));
   U2061 : AOI22_X1 port map( A1 => n109, A2 => regs(25), B1 => n66, B2 => 
                           regs(2073), ZN => n1385);
   U2062 : AOI22_X1 port map( A1 => n79, A2 => regs(1561), B1 => n25, B2 => 
                           regs(537), ZN => n1384);
   U2063 : OAI211_X1 port map( C1 => n10, C2 => n1386, A => n1385, B => n1384, 
                           ZN => curr_proc_regs(537));
   U2064 : AOI22_X1 port map( A1 => n109, A2 => regs(26), B1 => n5, B2 => 
                           regs(2074), ZN => n1388);
   U2065 : AOI22_X1 port map( A1 => n79, A2 => regs(1562), B1 => n29, B2 => 
                           regs(538), ZN => n1387);
   U2066 : OAI211_X1 port map( C1 => n10, C2 => n1389, A => n1388, B => n1387, 
                           ZN => curr_proc_regs(538));
   U2067 : AOI22_X1 port map( A1 => n106, A2 => regs(27), B1 => n66, B2 => 
                           regs(2075), ZN => n1391);
   U2068 : AOI22_X1 port map( A1 => n79, A2 => regs(1563), B1 => n19, B2 => 
                           regs(539), ZN => n1390);
   U2069 : OAI211_X1 port map( C1 => n10, C2 => n1392, A => n1391, B => n1390, 
                           ZN => curr_proc_regs(539));
   U2070 : INV_X1 port map( A => regs(565), ZN => n1476);
   U2071 : AOI22_X1 port map( A1 => n107, A2 => regs(2101), B1 => n5, B2 => 
                           regs(1589), ZN => n1394);
   U2072 : AOI22_X1 port map( A1 => n79, A2 => regs(1077), B1 => n28, B2 => 
                           regs(53), ZN => n1393);
   U2073 : OAI211_X1 port map( C1 => n40, C2 => n1476, A => n1394, B => n1393, 
                           ZN => curr_proc_regs(53));
   U2074 : AOI22_X1 port map( A1 => n108, A2 => regs(28), B1 => n68, B2 => 
                           regs(2076), ZN => n1396);
   U2075 : AOI22_X1 port map( A1 => n41, A2 => regs(1052), B1 => n102, B2 => 
                           regs(1564), ZN => n1395);
   U2076 : OAI211_X1 port map( C1 => n14, C2 => n1397, A => n1396, B => n1395, 
                           ZN => curr_proc_regs(540));
   U2077 : AOI22_X1 port map( A1 => n106, A2 => regs(29), B1 => n74, B2 => 
                           regs(2077), ZN => n1399);
   U2078 : AOI22_X1 port map( A1 => n79, A2 => regs(1565), B1 => n29, B2 => 
                           regs(541), ZN => n1398);
   U2079 : OAI211_X1 port map( C1 => n40, C2 => n1400, A => n1399, B => n1398, 
                           ZN => curr_proc_regs(541));
   U2080 : AOI22_X1 port map( A1 => n106, A2 => regs(30), B1 => n69, B2 => 
                           regs(2078), ZN => n1402);
   U2081 : AOI22_X1 port map( A1 => n79, A2 => regs(1566), B1 => n30, B2 => 
                           regs(542), ZN => n1401);
   U2082 : OAI211_X1 port map( C1 => n40, C2 => n1403, A => n1402, B => n1401, 
                           ZN => curr_proc_regs(542));
   U2083 : AOI22_X1 port map( A1 => n107, A2 => regs(31), B1 => n69, B2 => 
                           regs(2079), ZN => n1405);
   U2084 : AOI22_X1 port map( A1 => n56, A2 => regs(1055), B1 => n83, B2 => 
                           regs(1567), ZN => n1404);
   U2085 : OAI211_X1 port map( C1 => n14, C2 => n1406, A => n1405, B => n1404, 
                           ZN => curr_proc_regs(543));
   U2086 : AOI22_X1 port map( A1 => n108, A2 => regs(32), B1 => n63, B2 => 
                           regs(2080), ZN => n1408);
   U2087 : AOI22_X1 port map( A1 => n52, A2 => regs(1056), B1 => n97, B2 => 
                           regs(1568), ZN => n1407);
   U2088 : OAI211_X1 port map( C1 => n14, C2 => n1409, A => n1408, B => n1407, 
                           ZN => curr_proc_regs(544));
   U2089 : AOI22_X1 port map( A1 => n107, A2 => regs(33), B1 => n71, B2 => 
                           regs(2081), ZN => n1411);
   U2090 : AOI22_X1 port map( A1 => n79, A2 => regs(1569), B1 => n32, B2 => 
                           regs(545), ZN => n1410);
   U2091 : OAI211_X1 port map( C1 => n40, C2 => n1412, A => n1411, B => n1410, 
                           ZN => curr_proc_regs(545));
   U2092 : AOI22_X1 port map( A1 => n109, A2 => regs(34), B1 => n68, B2 => 
                           regs(2082), ZN => n1414);
   U2093 : AOI22_X1 port map( A1 => n52, A2 => regs(1058), B1 => n99, B2 => 
                           regs(1570), ZN => n1413);
   U2094 : OAI211_X1 port map( C1 => n14, C2 => n1415, A => n1414, B => n1413, 
                           ZN => curr_proc_regs(546));
   U2095 : AOI22_X1 port map( A1 => n106, A2 => regs(35), B1 => n70, B2 => 
                           regs(2083), ZN => n1417);
   U2096 : AOI22_X1 port map( A1 => n79, A2 => regs(1571), B1 => n34, B2 => 
                           regs(547), ZN => n1416);
   U2097 : OAI211_X1 port map( C1 => n40, C2 => n1418, A => n1417, B => n1416, 
                           ZN => curr_proc_regs(547));
   U2098 : AOI22_X1 port map( A1 => n107, A2 => regs(36), B1 => n65, B2 => 
                           regs(2084), ZN => n1420);
   U2099 : AOI22_X1 port map( A1 => n79, A2 => regs(1572), B1 => n33, B2 => 
                           regs(548), ZN => n1419);
   U2100 : OAI211_X1 port map( C1 => n40, C2 => n1421, A => n1420, B => n1419, 
                           ZN => curr_proc_regs(548));
   U2101 : AOI22_X1 port map( A1 => n108, A2 => regs(37), B1 => n74, B2 => 
                           regs(2085), ZN => n1423);
   U2102 : AOI22_X1 port map( A1 => n52, A2 => regs(1061), B1 => n83, B2 => 
                           regs(1573), ZN => n1422);
   U2103 : OAI211_X1 port map( C1 => n2128, C2 => n1424, A => n1423, B => n1422
                           , ZN => curr_proc_regs(549));
   U2104 : INV_X1 port map( A => regs(1078), ZN => n1479);
   U2105 : AOI22_X1 port map( A1 => n108, A2 => regs(2102), B1 => n72, B2 => 
                           regs(1590), ZN => n1426);
   U2106 : AOI22_X1 port map( A1 => n52, A2 => regs(566), B1 => n31, B2 => 
                           regs(54), ZN => n1425);
   U2107 : OAI211_X1 port map( C1 => n6, C2 => n1479, A => n1426, B => n1425, 
                           ZN => curr_proc_regs(54));
   U2108 : AOI22_X1 port map( A1 => n109, A2 => regs(38), B1 => n73, B2 => 
                           regs(2086), ZN => n1428);
   U2109 : AOI22_X1 port map( A1 => n52, A2 => regs(1062), B1 => n102, B2 => 
                           regs(1574), ZN => n1427);
   U2110 : OAI211_X1 port map( C1 => n14, C2 => n1429, A => n1428, B => n1427, 
                           ZN => curr_proc_regs(550));
   U2111 : AOI22_X1 port map( A1 => n106, A2 => regs(39), B1 => n66, B2 => 
                           regs(2087), ZN => n1431);
   U2112 : AOI22_X1 port map( A1 => n52, A2 => regs(1063), B1 => n102, B2 => 
                           regs(1575), ZN => n1430);
   U2113 : OAI211_X1 port map( C1 => n2128, C2 => n1432, A => n1431, B => n1430
                           , ZN => curr_proc_regs(551));
   U2114 : AOI22_X1 port map( A1 => n107, A2 => regs(40), B1 => n5, B2 => 
                           regs(2088), ZN => n1434);
   U2115 : AOI22_X1 port map( A1 => n52, A2 => regs(1064), B1 => n100, B2 => 
                           regs(1576), ZN => n1433);
   U2116 : OAI211_X1 port map( C1 => n14, C2 => n1435, A => n1434, B => n1433, 
                           ZN => curr_proc_regs(552));
   U2117 : AOI22_X1 port map( A1 => n108, A2 => regs(41), B1 => n67, B2 => 
                           regs(2089), ZN => n1437);
   U2118 : AOI22_X1 port map( A1 => n79, A2 => regs(1577), B1 => n21, B2 => 
                           regs(553), ZN => n1436);
   U2119 : OAI211_X1 port map( C1 => n2201, C2 => n1438, A => n1437, B => n1436
                           , ZN => curr_proc_regs(553));
   U2120 : AOI22_X1 port map( A1 => n109, A2 => regs(42), B1 => n70, B2 => 
                           regs(2090), ZN => n1440);
   U2121 : AOI22_X1 port map( A1 => n79, A2 => regs(1578), B1 => n22, B2 => 
                           regs(554), ZN => n1439);
   U2122 : OAI211_X1 port map( C1 => n40, C2 => n1441, A => n1440, B => n1439, 
                           ZN => curr_proc_regs(554));
   U2123 : AOI22_X1 port map( A1 => n106, A2 => regs(43), B1 => n68, B2 => 
                           regs(2091), ZN => n1443);
   U2124 : AOI22_X1 port map( A1 => n79, A2 => regs(1579), B1 => n23, B2 => 
                           regs(555), ZN => n1442);
   U2125 : OAI211_X1 port map( C1 => n40, C2 => n1444, A => n1443, B => n1442, 
                           ZN => curr_proc_regs(555));
   U2126 : AOI22_X1 port map( A1 => n107, A2 => regs(44), B1 => n5, B2 => 
                           regs(2092), ZN => n1446);
   U2127 : AOI22_X1 port map( A1 => n52, A2 => regs(1068), B1 => n99, B2 => 
                           regs(1580), ZN => n1445);
   U2128 : OAI211_X1 port map( C1 => n14, C2 => n1447, A => n1446, B => n1445, 
                           ZN => curr_proc_regs(556));
   U2129 : AOI22_X1 port map( A1 => n108, A2 => regs(45), B1 => n74, B2 => 
                           regs(2093), ZN => n1449);
   U2130 : AOI22_X1 port map( A1 => n52, A2 => regs(1069), B1 => n99, B2 => 
                           regs(1581), ZN => n1448);
   U2131 : OAI211_X1 port map( C1 => n14, C2 => n1450, A => n1449, B => n1448, 
                           ZN => curr_proc_regs(557));
   U2132 : AOI22_X1 port map( A1 => n109, A2 => regs(46), B1 => n69, B2 => 
                           regs(2094), ZN => n1452);
   U2133 : AOI22_X1 port map( A1 => n52, A2 => regs(1070), B1 => n97, B2 => 
                           regs(1582), ZN => n1451);
   U2134 : OAI211_X1 port map( C1 => n14, C2 => n1453, A => n1452, B => n1451, 
                           ZN => curr_proc_regs(558));
   U2135 : AOI22_X1 port map( A1 => n106, A2 => regs(47), B1 => n68, B2 => 
                           regs(2095), ZN => n1455);
   U2136 : AOI22_X1 port map( A1 => n52, A2 => regs(1071), B1 => n90, B2 => 
                           regs(1583), ZN => n1454);
   U2137 : OAI211_X1 port map( C1 => n2128, C2 => n1456, A => n1455, B => n1454
                           , ZN => curr_proc_regs(559));
   U2138 : INV_X1 port map( A => regs(1079), ZN => n1482);
   U2139 : AOI22_X1 port map( A1 => n107, A2 => regs(2103), B1 => n71, B2 => 
                           regs(1591), ZN => n1458);
   U2140 : AOI22_X1 port map( A1 => n44, A2 => regs(567), B1 => n24, B2 => 
                           regs(55), ZN => n1457);
   U2141 : OAI211_X1 port map( C1 => n6, C2 => n1482, A => n1458, B => n1457, 
                           ZN => curr_proc_regs(55));
   U2142 : AOI22_X1 port map( A1 => n108, A2 => regs(48), B1 => n68, B2 => 
                           regs(2096), ZN => n1460);
   U2143 : AOI22_X1 port map( A1 => n1, A2 => regs(1072), B1 => n93, B2 => 
                           regs(1584), ZN => n1459);
   U2144 : OAI211_X1 port map( C1 => n14, C2 => n1461, A => n1460, B => n1459, 
                           ZN => curr_proc_regs(560));
   U2145 : AOI22_X1 port map( A1 => n109, A2 => regs(49), B1 => n70, B2 => 
                           regs(2097), ZN => n1463);
   U2146 : AOI22_X1 port map( A1 => n79, A2 => regs(1585), B1 => n17, B2 => 
                           regs(561), ZN => n1462);
   U2147 : OAI211_X1 port map( C1 => n40, C2 => n1464, A => n1463, B => n1462, 
                           ZN => curr_proc_regs(561));
   U2148 : AOI22_X1 port map( A1 => n106, A2 => regs(50), B1 => n65, B2 => 
                           regs(2098), ZN => n1466);
   U2149 : AOI22_X1 port map( A1 => n54, A2 => regs(1074), B1 => n85, B2 => 
                           regs(1586), ZN => n1465);
   U2150 : OAI211_X1 port map( C1 => n2128, C2 => n1467, A => n1466, B => n1465
                           , ZN => curr_proc_regs(562));
   U2151 : AOI22_X1 port map( A1 => n107, A2 => regs(51), B1 => n74, B2 => 
                           regs(2099), ZN => n1469);
   U2152 : AOI22_X1 port map( A1 => n3, A2 => regs(1075), B1 => n89, B2 => 
                           regs(1587), ZN => n1468);
   U2153 : OAI211_X1 port map( C1 => n14, C2 => n1470, A => n1469, B => n1468, 
                           ZN => curr_proc_regs(563));
   U2154 : AOI22_X1 port map( A1 => n108, A2 => regs(52), B1 => n5, B2 => 
                           regs(2100), ZN => n1472);
   U2155 : AOI22_X1 port map( A1 => n79, A2 => regs(1588), B1 => n18, B2 => 
                           regs(564), ZN => n1471);
   U2156 : OAI211_X1 port map( C1 => n40, C2 => n1473, A => n1472, B => n1471, 
                           ZN => curr_proc_regs(564));
   U2157 : AOI22_X1 port map( A1 => n108, A2 => regs(53), B1 => n69, B2 => 
                           regs(2101), ZN => n1475);
   U2158 : AOI22_X1 port map( A1 => n48, A2 => regs(1077), B1 => n93, B2 => 
                           regs(1589), ZN => n1474);
   U2159 : OAI211_X1 port map( C1 => n12, C2 => n1476, A => n1475, B => n1474, 
                           ZN => curr_proc_regs(565));
   U2160 : AOI22_X1 port map( A1 => n108, A2 => regs(54), B1 => n69, B2 => 
                           regs(2102), ZN => n1478);
   U2161 : AOI22_X1 port map( A1 => n79, A2 => regs(1590), B1 => n19, B2 => 
                           regs(566), ZN => n1477);
   U2162 : OAI211_X1 port map( C1 => n40, C2 => n1479, A => n1478, B => n1477, 
                           ZN => curr_proc_regs(566));
   U2163 : AOI22_X1 port map( A1 => n108, A2 => regs(55), B1 => n69, B2 => 
                           regs(2103), ZN => n1481);
   U2164 : AOI22_X1 port map( A1 => n79, A2 => regs(1591), B1 => n34, B2 => 
                           regs(567), ZN => n1480);
   U2165 : OAI211_X1 port map( C1 => n40, C2 => n1482, A => n1481, B => n1480, 
                           ZN => curr_proc_regs(567));
   U2166 : INV_X1 port map( A => regs(1592), ZN => n1485);
   U2167 : AOI22_X1 port map( A1 => n108, A2 => regs(56), B1 => n69, B2 => 
                           regs(2104), ZN => n1484);
   U2168 : AOI22_X1 port map( A1 => n56, A2 => regs(1080), B1 => n27, B2 => 
                           regs(568), ZN => n1483);
   U2169 : OAI211_X1 port map( C1 => n11, C2 => n1485, A => n1484, B => n1483, 
                           ZN => curr_proc_regs(568));
   U2170 : INV_X1 port map( A => regs(1593), ZN => n1488);
   U2171 : AOI22_X1 port map( A1 => n108, A2 => regs(57), B1 => n69, B2 => 
                           regs(2105), ZN => n1487);
   U2172 : AOI22_X1 port map( A1 => n8, A2 => regs(1081), B1 => n26, B2 => 
                           regs(569), ZN => n1486);
   U2173 : OAI211_X1 port map( C1 => n78, C2 => n1488, A => n1487, B => n1486, 
                           ZN => curr_proc_regs(569));
   U2174 : INV_X1 port map( A => regs(1080), ZN => n1491);
   U2175 : AOI22_X1 port map( A1 => n108, A2 => regs(2104), B1 => n69, B2 => 
                           regs(1592), ZN => n1490);
   U2176 : AOI22_X1 port map( A1 => n3, A2 => regs(568), B1 => n39, B2 => 
                           regs(56), ZN => n1489);
   U2177 : OAI211_X1 port map( C1 => n6, C2 => n1491, A => n1490, B => n1489, 
                           ZN => curr_proc_regs(56));
   U2178 : INV_X1 port map( A => regs(1594), ZN => n1494);
   U2179 : AOI22_X1 port map( A1 => n108, A2 => regs(58), B1 => n69, B2 => 
                           regs(2106), ZN => n1493);
   U2180 : AOI22_X1 port map( A1 => n1, A2 => regs(1082), B1 => n37, B2 => 
                           regs(570), ZN => n1492);
   U2181 : OAI211_X1 port map( C1 => n11, C2 => n1494, A => n1493, B => n1492, 
                           ZN => curr_proc_regs(570));
   U2182 : INV_X1 port map( A => regs(1595), ZN => n1497);
   U2183 : AOI22_X1 port map( A1 => n108, A2 => regs(59), B1 => n69, B2 => 
                           regs(2107), ZN => n1496);
   U2184 : AOI22_X1 port map( A1 => n8, A2 => regs(1083), B1 => n20, B2 => 
                           regs(571), ZN => n1495);
   U2185 : OAI211_X1 port map( C1 => n11, C2 => n1497, A => n1496, B => n1495, 
                           ZN => curr_proc_regs(571));
   U2186 : INV_X1 port map( A => regs(1084), ZN => n1609);
   U2187 : AOI22_X1 port map( A1 => n108, A2 => regs(60), B1 => n69, B2 => 
                           regs(2108), ZN => n1499);
   U2188 : AOI22_X1 port map( A1 => n79, A2 => regs(1596), B1 => n17, B2 => 
                           regs(572), ZN => n1498);
   U2189 : OAI211_X1 port map( C1 => n40, C2 => n1609, A => n1499, B => n1498, 
                           ZN => curr_proc_regs(572));
   U2190 : INV_X1 port map( A => regs(1597), ZN => n1502);
   U2191 : AOI22_X1 port map( A1 => n108, A2 => regs(61), B1 => n69, B2 => 
                           regs(2109), ZN => n1501);
   U2192 : AOI22_X1 port map( A1 => n3, A2 => regs(1085), B1 => n29, B2 => 
                           regs(573), ZN => n1500);
   U2193 : OAI211_X1 port map( C1 => n6, C2 => n1502, A => n1501, B => n1500, 
                           ZN => curr_proc_regs(573));
   U2194 : INV_X1 port map( A => regs(1598), ZN => n1505);
   U2195 : AOI22_X1 port map( A1 => n108, A2 => regs(62), B1 => n69, B2 => 
                           regs(2110), ZN => n1504);
   U2196 : AOI22_X1 port map( A1 => n1, A2 => regs(1086), B1 => n30, B2 => 
                           regs(574), ZN => n1503);
   U2197 : OAI211_X1 port map( C1 => n2215, C2 => n1505, A => n1504, B => n1503
                           , ZN => curr_proc_regs(574));
   U2198 : INV_X1 port map( A => regs(1599), ZN => n1508);
   U2199 : AOI22_X1 port map( A1 => n108, A2 => regs(63), B1 => n69, B2 => 
                           regs(2111), ZN => n1507);
   U2200 : AOI22_X1 port map( A1 => n8, A2 => regs(1087), B1 => n27, B2 => 
                           regs(575), ZN => n1506);
   U2201 : OAI211_X1 port map( C1 => n6, C2 => n1508, A => n1507, B => n1506, 
                           ZN => curr_proc_regs(575));
   U2202 : INV_X1 port map( A => regs(1088), ZN => n1740);
   U2203 : AOI22_X1 port map( A1 => n107, A2 => regs(64), B1 => n69, B2 => 
                           regs(2112), ZN => n1510);
   U2204 : AOI22_X1 port map( A1 => n79, A2 => regs(1600), B1 => n28, B2 => 
                           regs(576), ZN => n1509);
   U2205 : OAI211_X1 port map( C1 => n58, C2 => n1740, A => n1510, B => n1509, 
                           ZN => curr_proc_regs(576));
   U2206 : INV_X1 port map( A => regs(1601), ZN => n1513);
   U2207 : AOI22_X1 port map( A1 => n107, A2 => regs(65), B1 => n69, B2 => 
                           regs(2113), ZN => n1512);
   U2208 : AOI22_X1 port map( A1 => n54, A2 => regs(1089), B1 => n29, B2 => 
                           regs(577), ZN => n1511);
   U2209 : OAI211_X1 port map( C1 => n2215, C2 => n1513, A => n1512, B => n1511
                           , ZN => curr_proc_regs(577));
   U2210 : INV_X1 port map( A => regs(1090), ZN => n1806);
   U2211 : AOI22_X1 port map( A1 => n107, A2 => regs(66), B1 => n69, B2 => 
                           regs(2114), ZN => n1515);
   U2212 : AOI22_X1 port map( A1 => n84, A2 => regs(1602), B1 => n30, B2 => 
                           regs(578), ZN => n1514);
   U2213 : OAI211_X1 port map( C1 => n59, C2 => n1806, A => n1515, B => n1514, 
                           ZN => curr_proc_regs(578));
   U2214 : INV_X1 port map( A => regs(1603), ZN => n1518);
   U2215 : AOI22_X1 port map( A1 => n107, A2 => regs(67), B1 => n69, B2 => 
                           regs(2115), ZN => n1517);
   U2216 : AOI22_X1 port map( A1 => n54, A2 => regs(1091), B1 => n32, B2 => 
                           regs(579), ZN => n1516);
   U2217 : OAI211_X1 port map( C1 => n11, C2 => n1518, A => n1517, B => n1516, 
                           ZN => curr_proc_regs(579));
   U2218 : INV_X1 port map( A => regs(569), ZN => n1521);
   U2219 : AOI22_X1 port map( A1 => n107, A2 => regs(2105), B1 => n69, B2 => 
                           regs(1593), ZN => n1520);
   U2220 : AOI22_X1 port map( A1 => n86, A2 => regs(1081), B1 => n21, B2 => 
                           regs(57), ZN => n1519);
   U2221 : OAI211_X1 port map( C1 => n58, C2 => n1521, A => n1520, B => n1519, 
                           ZN => curr_proc_regs(57));
   U2222 : INV_X1 port map( A => regs(1604), ZN => n1524);
   U2223 : AOI22_X1 port map( A1 => n107, A2 => regs(68), B1 => n69, B2 => 
                           regs(2116), ZN => n1523);
   U2224 : AOI22_X1 port map( A1 => n54, A2 => regs(1092), B1 => n22, B2 => 
                           regs(580), ZN => n1522);
   U2225 : OAI211_X1 port map( C1 => n11, C2 => n1524, A => n1523, B => n1522, 
                           ZN => curr_proc_regs(580));
   U2226 : INV_X1 port map( A => regs(1605), ZN => n1527);
   U2227 : AOI22_X1 port map( A1 => n107, A2 => regs(69), B1 => n69, B2 => 
                           regs(2117), ZN => n1526);
   U2228 : AOI22_X1 port map( A1 => n54, A2 => regs(1093), B1 => n23, B2 => 
                           regs(581), ZN => n1525);
   U2229 : OAI211_X1 port map( C1 => n6, C2 => n1527, A => n1526, B => n1525, 
                           ZN => curr_proc_regs(581));
   U2230 : INV_X1 port map( A => regs(1094), ZN => n1941);
   U2231 : AOI22_X1 port map( A1 => n107, A2 => regs(70), B1 => n69, B2 => 
                           regs(2118), ZN => n1529);
   U2232 : AOI22_X1 port map( A1 => n97, A2 => regs(1606), B1 => n24, B2 => 
                           regs(582), ZN => n1528);
   U2233 : OAI211_X1 port map( C1 => n57, C2 => n1941, A => n1529, B => n1528, 
                           ZN => curr_proc_regs(582));
   U2234 : INV_X1 port map( A => regs(1607), ZN => n1532);
   U2235 : AOI22_X1 port map( A1 => n107, A2 => regs(71), B1 => n69, B2 => 
                           regs(2119), ZN => n1531);
   U2236 : AOI22_X1 port map( A1 => n54, A2 => regs(1095), B1 => n17, B2 => 
                           regs(583), ZN => n1530);
   U2237 : OAI211_X1 port map( C1 => n13, C2 => n1532, A => n1531, B => n1530, 
                           ZN => curr_proc_regs(583));
   U2238 : INV_X1 port map( A => regs(1096), ZN => n2007);
   U2239 : AOI22_X1 port map( A1 => n107, A2 => regs(72), B1 => n69, B2 => 
                           regs(2120), ZN => n1534);
   U2240 : AOI22_X1 port map( A1 => n90, A2 => regs(1608), B1 => n18, B2 => 
                           regs(584), ZN => n1533);
   U2241 : OAI211_X1 port map( C1 => n57, C2 => n2007, A => n1534, B => n1533, 
                           ZN => curr_proc_regs(584));
   U2242 : INV_X1 port map( A => regs(1097), ZN => n2040);
   U2243 : AOI22_X1 port map( A1 => n107, A2 => regs(73), B1 => n69, B2 => 
                           regs(2121), ZN => n1536);
   U2244 : AOI22_X1 port map( A1 => n83, A2 => regs(1609), B1 => n19, B2 => 
                           regs(585), ZN => n1535);
   U2245 : OAI211_X1 port map( C1 => n59, C2 => n2040, A => n1536, B => n1535, 
                           ZN => curr_proc_regs(585));
   U2246 : INV_X1 port map( A => regs(1098), ZN => n2073);
   U2247 : AOI22_X1 port map( A1 => n107, A2 => regs(74), B1 => n69, B2 => 
                           regs(2122), ZN => n1538);
   U2248 : AOI22_X1 port map( A1 => n94, A2 => regs(1610), B1 => n33, B2 => 
                           regs(586), ZN => n1537);
   U2249 : OAI211_X1 port map( C1 => n59, C2 => n2073, A => n1538, B => n1537, 
                           ZN => curr_proc_regs(586));
   U2250 : INV_X1 port map( A => regs(1611), ZN => n1541);
   U2251 : AOI22_X1 port map( A1 => n106, A2 => regs(75), B1 => n70, B2 => 
                           regs(2123), ZN => n1540);
   U2252 : AOI22_X1 port map( A1 => n3, A2 => regs(1099), B1 => n35, B2 => 
                           regs(587), ZN => n1539);
   U2253 : OAI211_X1 port map( C1 => n13, C2 => n1541, A => n1540, B => n1539, 
                           ZN => curr_proc_regs(587));
   U2254 : INV_X1 port map( A => regs(1100), ZN => n2134);
   U2255 : AOI22_X1 port map( A1 => n106, A2 => regs(76), B1 => n70, B2 => 
                           regs(2124), ZN => n1543);
   U2256 : AOI22_X1 port map( A1 => n88, A2 => regs(1612), B1 => n25, B2 => 
                           regs(588), ZN => n1542);
   U2257 : OAI211_X1 port map( C1 => n40, C2 => n2134, A => n1543, B => n1542, 
                           ZN => curr_proc_regs(588));
   U2258 : INV_X1 port map( A => regs(1613), ZN => n1546);
   U2259 : AOI22_X1 port map( A1 => n106, A2 => regs(77), B1 => n70, B2 => 
                           regs(2125), ZN => n1545);
   U2260 : AOI22_X1 port map( A1 => n41, A2 => regs(1101), B1 => n27, B2 => 
                           regs(589), ZN => n1544);
   U2261 : OAI211_X1 port map( C1 => n13, C2 => n1546, A => n1545, B => n1544, 
                           ZN => curr_proc_regs(589));
   U2262 : INV_X1 port map( A => regs(570), ZN => n1549);
   U2263 : AOI22_X1 port map( A1 => n106, A2 => regs(2106), B1 => n70, B2 => 
                           regs(1594), ZN => n1548);
   U2264 : AOI22_X1 port map( A1 => n99, A2 => regs(1082), B1 => n26, B2 => 
                           regs(58), ZN => n1547);
   U2265 : OAI211_X1 port map( C1 => n40, C2 => n1549, A => n1548, B => n1547, 
                           ZN => curr_proc_regs(58));
   U2266 : INV_X1 port map( A => regs(1102), ZN => n2140);
   U2267 : AOI22_X1 port map( A1 => n106, A2 => regs(78), B1 => n70, B2 => 
                           regs(2126), ZN => n1551);
   U2268 : AOI22_X1 port map( A1 => n93, A2 => regs(1614), B1 => n18, B2 => 
                           regs(590), ZN => n1550);
   U2269 : OAI211_X1 port map( C1 => n2201, C2 => n2140, A => n1551, B => n1550
                           , ZN => curr_proc_regs(590));
   U2270 : INV_X1 port map( A => regs(1103), ZN => n2143);
   U2271 : AOI22_X1 port map( A1 => n106, A2 => regs(79), B1 => n70, B2 => 
                           regs(2127), ZN => n1553);
   U2272 : AOI22_X1 port map( A1 => n97, A2 => regs(1615), B1 => n30, B2 => 
                           regs(591), ZN => n1552);
   U2273 : OAI211_X1 port map( C1 => n40, C2 => n2143, A => n1553, B => n1552, 
                           ZN => curr_proc_regs(591));
   U2274 : INV_X1 port map( A => regs(1104), ZN => n2149);
   U2275 : AOI22_X1 port map( A1 => n106, A2 => regs(80), B1 => n70, B2 => 
                           regs(2128), ZN => n1555);
   U2276 : AOI22_X1 port map( A1 => n90, A2 => regs(1616), B1 => n32, B2 => 
                           regs(592), ZN => n1554);
   U2277 : OAI211_X1 port map( C1 => n40, C2 => n2149, A => n1555, B => n1554, 
                           ZN => curr_proc_regs(592));
   U2278 : INV_X1 port map( A => regs(1105), ZN => n2152);
   U2279 : AOI22_X1 port map( A1 => n106, A2 => regs(81), B1 => n70, B2 => 
                           regs(2129), ZN => n1557);
   U2280 : AOI22_X1 port map( A1 => n83, A2 => regs(1617), B1 => n20, B2 => 
                           regs(593), ZN => n1556);
   U2281 : OAI211_X1 port map( C1 => n40, C2 => n2152, A => n1557, B => n1556, 
                           ZN => curr_proc_regs(593));
   U2282 : INV_X1 port map( A => regs(1618), ZN => n1560);
   U2283 : AOI22_X1 port map( A1 => n106, A2 => regs(82), B1 => n70, B2 => 
                           regs(2130), ZN => n1559);
   U2284 : AOI22_X1 port map( A1 => n42, A2 => regs(1106), B1 => n28, B2 => 
                           regs(594), ZN => n1558);
   U2285 : OAI211_X1 port map( C1 => n13, C2 => n1560, A => n1559, B => n1558, 
                           ZN => curr_proc_regs(594));
   U2286 : INV_X1 port map( A => regs(1619), ZN => n1563);
   U2287 : AOI22_X1 port map( A1 => n106, A2 => regs(83), B1 => n70, B2 => 
                           regs(2131), ZN => n1562);
   U2288 : AOI22_X1 port map( A1 => n53, A2 => regs(1107), B1 => n29, B2 => 
                           regs(595), ZN => n1561);
   U2289 : OAI211_X1 port map( C1 => n13, C2 => n1563, A => n1562, B => n1561, 
                           ZN => curr_proc_regs(595));
   U2290 : INV_X1 port map( A => regs(1620), ZN => n1566);
   U2291 : AOI22_X1 port map( A1 => n106, A2 => regs(84), B1 => n70, B2 => 
                           regs(2132), ZN => n1565);
   U2292 : AOI22_X1 port map( A1 => n54, A2 => regs(1108), B1 => n30, B2 => 
                           regs(596), ZN => n1564);
   U2293 : OAI211_X1 port map( C1 => n13, C2 => n1566, A => n1565, B => n1564, 
                           ZN => curr_proc_regs(596));
   U2294 : INV_X1 port map( A => regs(1621), ZN => n1569);
   U2295 : AOI22_X1 port map( A1 => n106, A2 => regs(85), B1 => n70, B2 => 
                           regs(2133), ZN => n1568);
   U2296 : AOI22_X1 port map( A1 => n43, A2 => regs(1109), B1 => n32, B2 => 
                           regs(597), ZN => n1567);
   U2297 : OAI211_X1 port map( C1 => n13, C2 => n1569, A => n1568, B => n1567, 
                           ZN => curr_proc_regs(597));
   U2298 : INV_X1 port map( A => regs(1110), ZN => n2167);
   U2299 : AOI22_X1 port map( A1 => n105, A2 => regs(86), B1 => n5, B2 => 
                           regs(2134), ZN => n1571);
   U2300 : AOI22_X1 port map( A1 => n95, A2 => regs(1622), B1 => n35, B2 => 
                           regs(598), ZN => n1570);
   U2301 : OAI211_X1 port map( C1 => n40, C2 => n2167, A => n1571, B => n1570, 
                           ZN => curr_proc_regs(598));
   U2302 : INV_X1 port map( A => regs(1111), ZN => n2170);
   U2303 : AOI22_X1 port map( A1 => n105, A2 => regs(87), B1 => n72, B2 => 
                           regs(2135), ZN => n1573);
   U2304 : AOI22_X1 port map( A1 => n99, A2 => regs(1623), B1 => n39, B2 => 
                           regs(599), ZN => n1572);
   U2305 : OAI211_X1 port map( C1 => n40, C2 => n2170, A => n1573, B => n1572, 
                           ZN => curr_proc_regs(599));
   U2306 : INV_X1 port map( A => regs(571), ZN => n1576);
   U2307 : AOI22_X1 port map( A1 => n105, A2 => regs(2107), B1 => n73, B2 => 
                           regs(1595), ZN => n1575);
   U2308 : AOI22_X1 port map( A1 => n85, A2 => regs(1083), B1 => n38, B2 => 
                           regs(59), ZN => n1574);
   U2309 : OAI211_X1 port map( C1 => n40, C2 => n1576, A => n1575, B => n1574, 
                           ZN => curr_proc_regs(59));
   U2310 : INV_X1 port map( A => regs(517), ZN => n1579);
   U2311 : AOI22_X1 port map( A1 => n105, A2 => regs(2053), B1 => n2211, B2 => 
                           regs(1541), ZN => n1578);
   U2312 : AOI22_X1 port map( A1 => n85, A2 => regs(1029), B1 => n37, B2 => 
                           regs(5), ZN => n1577);
   U2313 : OAI211_X1 port map( C1 => n40, C2 => n1579, A => n1578, B => n1577, 
                           ZN => curr_proc_regs(5));
   U2314 : INV_X1 port map( A => regs(1112), ZN => n2173);
   U2315 : AOI22_X1 port map( A1 => n105, A2 => regs(88), B1 => n5, B2 => 
                           regs(2136), ZN => n1581);
   U2316 : AOI22_X1 port map( A1 => n85, A2 => regs(1624), B1 => n31, B2 => 
                           regs(600), ZN => n1580);
   U2317 : OAI211_X1 port map( C1 => n40, C2 => n2173, A => n1581, B => n1580, 
                           ZN => curr_proc_regs(600));
   U2318 : INV_X1 port map( A => regs(1625), ZN => n1584);
   U2319 : AOI22_X1 port map( A1 => n105, A2 => regs(89), B1 => n68, B2 => 
                           regs(2137), ZN => n1583);
   U2320 : AOI22_X1 port map( A1 => n53, A2 => regs(1113), B1 => n39, B2 => 
                           regs(601), ZN => n1582);
   U2321 : OAI211_X1 port map( C1 => n11, C2 => n1584, A => n1583, B => n1582, 
                           ZN => curr_proc_regs(601));
   U2322 : INV_X1 port map( A => regs(1626), ZN => n1587);
   U2323 : AOI22_X1 port map( A1 => n105, A2 => regs(90), B1 => n63, B2 => 
                           regs(2138), ZN => n1586);
   U2324 : AOI22_X1 port map( A1 => n55, A2 => regs(1114), B1 => n34, B2 => 
                           regs(602), ZN => n1585);
   U2325 : OAI211_X1 port map( C1 => n11, C2 => n1587, A => n1586, B => n1585, 
                           ZN => curr_proc_regs(602));
   U2326 : INV_X1 port map( A => regs(1627), ZN => n1590);
   U2327 : AOI22_X1 port map( A1 => n105, A2 => regs(91), B1 => n70, B2 => 
                           regs(2139), ZN => n1589);
   U2328 : AOI22_X1 port map( A1 => n44, A2 => regs(1115), B1 => n36, B2 => 
                           regs(603), ZN => n1588);
   U2329 : OAI211_X1 port map( C1 => n11, C2 => n1590, A => n1589, B => n1588, 
                           ZN => curr_proc_regs(603));
   U2330 : INV_X1 port map( A => regs(1116), ZN => n2188);
   U2331 : AOI22_X1 port map( A1 => n105, A2 => regs(92), B1 => n65, B2 => 
                           regs(2140), ZN => n1592);
   U2332 : AOI22_X1 port map( A1 => n85, A2 => regs(1628), B1 => n27, B2 => 
                           regs(604), ZN => n1591);
   U2333 : OAI211_X1 port map( C1 => n40, C2 => n2188, A => n1592, B => n1591, 
                           ZN => curr_proc_regs(604));
   U2334 : INV_X1 port map( A => regs(1629), ZN => n1595);
   U2335 : AOI22_X1 port map( A1 => n105, A2 => regs(93), B1 => n66, B2 => 
                           regs(2141), ZN => n1594);
   U2336 : AOI22_X1 port map( A1 => n42, A2 => regs(1117), B1 => n26, B2 => 
                           regs(605), ZN => n1593);
   U2337 : OAI211_X1 port map( C1 => n11, C2 => n1595, A => n1594, B => n1593, 
                           ZN => curr_proc_regs(605));
   U2338 : INV_X1 port map( A => regs(1630), ZN => n1598);
   U2339 : AOI22_X1 port map( A1 => n105, A2 => regs(94), B1 => n66, B2 => 
                           regs(2142), ZN => n1597);
   U2340 : AOI22_X1 port map( A1 => n41, A2 => regs(1118), B1 => n25, B2 => 
                           regs(606), ZN => n1596);
   U2341 : OAI211_X1 port map( C1 => n11, C2 => n1598, A => n1597, B => n1596, 
                           ZN => curr_proc_regs(606));
   U2342 : INV_X1 port map( A => regs(1119), ZN => n2197);
   U2343 : AOI22_X1 port map( A1 => n105, A2 => regs(95), B1 => n71, B2 => 
                           regs(2143), ZN => n1600);
   U2344 : AOI22_X1 port map( A1 => n85, A2 => regs(1631), B1 => n33, B2 => 
                           regs(607), ZN => n1599);
   U2345 : OAI211_X1 port map( C1 => n40, C2 => n2197, A => n1600, B => n1599, 
                           ZN => curr_proc_regs(607));
   U2346 : INV_X1 port map( A => regs(1632), ZN => n1603);
   U2347 : AOI22_X1 port map( A1 => n104, A2 => regs(96), B1 => n71, B2 => 
                           regs(2144), ZN => n1602);
   U2348 : AOI22_X1 port map( A1 => n3, A2 => regs(1120), B1 => n33, B2 => 
                           regs(608), ZN => n1601);
   U2349 : OAI211_X1 port map( C1 => n11, C2 => n1603, A => n1602, B => n1601, 
                           ZN => curr_proc_regs(608));
   U2350 : INV_X1 port map( A => regs(1633), ZN => n1606);
   U2351 : AOI22_X1 port map( A1 => n104, A2 => regs(97), B1 => n71, B2 => 
                           regs(2145), ZN => n1605);
   U2352 : AOI22_X1 port map( A1 => n3, A2 => regs(1121), B1 => n20, B2 => 
                           regs(609), ZN => n1604);
   U2353 : OAI211_X1 port map( C1 => n11, C2 => n1606, A => n1605, B => n1604, 
                           ZN => curr_proc_regs(609));
   U2354 : AOI22_X1 port map( A1 => n104, A2 => regs(2108), B1 => n71, B2 => 
                           regs(1596), ZN => n1608);
   U2355 : AOI22_X1 port map( A1 => n3, A2 => regs(572), B1 => n22, B2 => 
                           regs(60), ZN => n1607);
   U2356 : OAI211_X1 port map( C1 => n78, C2 => n1609, A => n1608, B => n1607, 
                           ZN => curr_proc_regs(60));
   U2357 : INV_X1 port map( A => regs(1634), ZN => n1612);
   U2358 : AOI22_X1 port map( A1 => n104, A2 => regs(98), B1 => n71, B2 => 
                           regs(2146), ZN => n1611);
   U2359 : AOI22_X1 port map( A1 => n3, A2 => regs(1122), B1 => n25, B2 => 
                           regs(610), ZN => n1610);
   U2360 : OAI211_X1 port map( C1 => n103, C2 => n1612, A => n1611, B => n1610,
                           ZN => curr_proc_regs(610));
   U2361 : INV_X1 port map( A => regs(1123), ZN => n2210);
   U2362 : AOI22_X1 port map( A1 => n104, A2 => regs(99), B1 => n71, B2 => 
                           regs(2147), ZN => n1614);
   U2363 : AOI22_X1 port map( A1 => n85, A2 => regs(1635), B1 => n35, B2 => 
                           regs(611), ZN => n1613);
   U2364 : OAI211_X1 port map( C1 => n40, C2 => n2210, A => n1614, B => n1613, 
                           ZN => curr_proc_regs(611));
   U2365 : AOI22_X1 port map( A1 => n104, A2 => regs(100), B1 => n71, B2 => 
                           regs(2148), ZN => n1616);
   U2366 : AOI22_X1 port map( A1 => n85, A2 => regs(1636), B1 => n39, B2 => 
                           regs(612), ZN => n1615);
   U2367 : OAI211_X1 port map( C1 => n57, C2 => n1617, A => n1616, B => n1615, 
                           ZN => curr_proc_regs(612));
   U2368 : AOI22_X1 port map( A1 => n104, A2 => regs(101), B1 => n71, B2 => 
                           regs(2149), ZN => n1619);
   U2369 : AOI22_X1 port map( A1 => n3, A2 => regs(1125), B1 => n102, B2 => 
                           regs(1637), ZN => n1618);
   U2370 : OAI211_X1 port map( C1 => n14, C2 => n1620, A => n1619, B => n1618, 
                           ZN => curr_proc_regs(613));
   U2371 : AOI22_X1 port map( A1 => n104, A2 => regs(102), B1 => n71, B2 => 
                           regs(2150), ZN => n1622);
   U2372 : AOI22_X1 port map( A1 => n3, A2 => regs(1126), B1 => n101, B2 => 
                           regs(1638), ZN => n1621);
   U2373 : OAI211_X1 port map( C1 => n12, C2 => n1623, A => n1622, B => n1621, 
                           ZN => curr_proc_regs(614));
   U2374 : AOI22_X1 port map( A1 => n104, A2 => regs(103), B1 => n71, B2 => 
                           regs(2151), ZN => n1625);
   U2375 : AOI22_X1 port map( A1 => n3, A2 => regs(1127), B1 => n101, B2 => 
                           regs(1639), ZN => n1624);
   U2376 : OAI211_X1 port map( C1 => n2128, C2 => n1626, A => n1625, B => n1624
                           , ZN => curr_proc_regs(615));
   U2377 : AOI22_X1 port map( A1 => n104, A2 => regs(104), B1 => n71, B2 => 
                           regs(2152), ZN => n1628);
   U2378 : AOI22_X1 port map( A1 => n3, A2 => regs(1128), B1 => n102, B2 => 
                           regs(1640), ZN => n1627);
   U2379 : OAI211_X1 port map( C1 => n14, C2 => n1629, A => n1628, B => n1627, 
                           ZN => curr_proc_regs(616));
   U2380 : AOI22_X1 port map( A1 => n109, A2 => regs(105), B1 => n71, B2 => 
                           regs(2153), ZN => n1631);
   U2381 : AOI22_X1 port map( A1 => n3, A2 => regs(1129), B1 => n101, B2 => 
                           regs(1641), ZN => n1630);
   U2382 : OAI211_X1 port map( C1 => n12, C2 => n1632, A => n1631, B => n1630, 
                           ZN => curr_proc_regs(617));
   U2383 : AOI22_X1 port map( A1 => n127, A2 => regs(106), B1 => n71, B2 => 
                           regs(2154), ZN => n1634);
   U2384 : AOI22_X1 port map( A1 => n3, A2 => regs(1130), B1 => n102, B2 => 
                           regs(1642), ZN => n1633);
   U2385 : OAI211_X1 port map( C1 => n2128, C2 => n1635, A => n1634, B => n1633
                           , ZN => curr_proc_regs(618));
   U2386 : AOI22_X1 port map( A1 => n120, A2 => regs(107), B1 => n68, B2 => 
                           regs(2155), ZN => n1637);
   U2387 : AOI22_X1 port map( A1 => n85, A2 => regs(1643), B1 => n38, B2 => 
                           regs(619), ZN => n1636);
   U2388 : OAI211_X1 port map( C1 => n57, C2 => n1638, A => n1637, B => n1636, 
                           ZN => curr_proc_regs(619));
   U2389 : INV_X1 port map( A => regs(1085), ZN => n1641);
   U2390 : AOI22_X1 port map( A1 => n120, A2 => regs(2109), B1 => n68, B2 => 
                           regs(1597), ZN => n1640);
   U2391 : AOI22_X1 port map( A1 => n3, A2 => regs(573), B1 => n37, B2 => 
                           regs(61), ZN => n1639);
   U2392 : OAI211_X1 port map( C1 => n78, C2 => n1641, A => n1640, B => n1639, 
                           ZN => curr_proc_regs(61));
   U2393 : AOI22_X1 port map( A1 => n120, A2 => regs(108), B1 => n63, B2 => 
                           regs(2156), ZN => n1643);
   U2394 : AOI22_X1 port map( A1 => n3, A2 => regs(1132), B1 => n102, B2 => 
                           regs(1644), ZN => n1642);
   U2395 : OAI211_X1 port map( C1 => n14, C2 => n1644, A => n1643, B => n1642, 
                           ZN => curr_proc_regs(620));
   U2396 : AOI22_X1 port map( A1 => n120, A2 => regs(109), B1 => n72, B2 => 
                           regs(2157), ZN => n1646);
   U2397 : AOI22_X1 port map( A1 => n85, A2 => regs(1645), B1 => n36, B2 => 
                           regs(621), ZN => n1645);
   U2398 : OAI211_X1 port map( C1 => n57, C2 => n1647, A => n1646, B => n1645, 
                           ZN => curr_proc_regs(621));
   U2399 : AOI22_X1 port map( A1 => n120, A2 => regs(110), B1 => n63, B2 => 
                           regs(2158), ZN => n1649);
   U2400 : AOI22_X1 port map( A1 => n3, A2 => regs(1134), B1 => n101, B2 => 
                           regs(1646), ZN => n1648);
   U2401 : OAI211_X1 port map( C1 => n14, C2 => n1650, A => n1649, B => n1648, 
                           ZN => curr_proc_regs(622));
   U2402 : AOI22_X1 port map( A1 => n120, A2 => regs(111), B1 => n68, B2 => 
                           regs(2159), ZN => n1652);
   U2403 : AOI22_X1 port map( A1 => n45, A2 => regs(1135), B1 => n101, B2 => 
                           regs(1647), ZN => n1651);
   U2404 : OAI211_X1 port map( C1 => n2128, C2 => n1653, A => n1652, B => n1651
                           , ZN => curr_proc_regs(623));
   U2405 : AOI22_X1 port map( A1 => n120, A2 => regs(112), B1 => n63, B2 => 
                           regs(2160), ZN => n1655);
   U2406 : AOI22_X1 port map( A1 => n3, A2 => regs(1136), B1 => n101, B2 => 
                           regs(1648), ZN => n1654);
   U2407 : OAI211_X1 port map( C1 => n2128, C2 => n1656, A => n1655, B => n1654
                           , ZN => curr_proc_regs(624));
   U2408 : AOI22_X1 port map( A1 => n120, A2 => regs(113), B1 => n72, B2 => 
                           regs(2161), ZN => n1658);
   U2409 : AOI22_X1 port map( A1 => n3, A2 => regs(1137), B1 => n102, B2 => 
                           regs(1649), ZN => n1657);
   U2410 : OAI211_X1 port map( C1 => n14, C2 => n1659, A => n1658, B => n1657, 
                           ZN => curr_proc_regs(625));
   U2411 : AOI22_X1 port map( A1 => n120, A2 => regs(114), B1 => n72, B2 => 
                           regs(2162), ZN => n1661);
   U2412 : AOI22_X1 port map( A1 => n3, A2 => regs(1138), B1 => n101, B2 => 
                           regs(1650), ZN => n1660);
   U2413 : OAI211_X1 port map( C1 => n2128, C2 => n1662, A => n1661, B => n1660
                           , ZN => curr_proc_regs(626));
   U2414 : AOI22_X1 port map( A1 => n120, A2 => regs(115), B1 => n68, B2 => 
                           regs(2163), ZN => n1664);
   U2415 : AOI22_X1 port map( A1 => n3, A2 => regs(1139), B1 => n93, B2 => 
                           regs(1651), ZN => n1663);
   U2416 : OAI211_X1 port map( C1 => n14, C2 => n1665, A => n1664, B => n1663, 
                           ZN => curr_proc_regs(627));
   U2417 : AOI22_X1 port map( A1 => n120, A2 => regs(116), B1 => n63, B2 => 
                           regs(2164), ZN => n1667);
   U2418 : AOI22_X1 port map( A1 => n3, A2 => regs(1140), B1 => n97, B2 => 
                           regs(1652), ZN => n1666);
   U2419 : OAI211_X1 port map( C1 => n14, C2 => n1668, A => n1667, B => n1666, 
                           ZN => curr_proc_regs(628));
   U2420 : AOI22_X1 port map( A1 => n120, A2 => regs(117), B1 => n72, B2 => 
                           regs(2165), ZN => n1670);
   U2421 : AOI22_X1 port map( A1 => n3, A2 => regs(1141), B1 => n90, B2 => 
                           regs(1653), ZN => n1669);
   U2422 : OAI211_X1 port map( C1 => n2128, C2 => n1671, A => n1670, B => n1669
                           , ZN => curr_proc_regs(629));
   U2423 : INV_X1 port map( A => regs(1086), ZN => n1674);
   U2424 : AOI22_X1 port map( A1 => n119, A2 => regs(2110), B1 => n74, B2 => 
                           regs(1598), ZN => n1673);
   U2425 : AOI22_X1 port map( A1 => n3, A2 => regs(574), B1 => n34, B2 => 
                           regs(62), ZN => n1672);
   U2426 : OAI211_X1 port map( C1 => n103, C2 => n1674, A => n1673, B => n1672,
                           ZN => curr_proc_regs(62));
   U2427 : AOI22_X1 port map( A1 => n119, A2 => regs(118), B1 => n74, B2 => 
                           regs(2166), ZN => n1676);
   U2428 : AOI22_X1 port map( A1 => n3, A2 => regs(1142), B1 => n83, B2 => 
                           regs(1654), ZN => n1675);
   U2429 : OAI211_X1 port map( C1 => n14, C2 => n1677, A => n1676, B => n1675, 
                           ZN => curr_proc_regs(630));
   U2430 : AOI22_X1 port map( A1 => n119, A2 => regs(119), B1 => n74, B2 => 
                           regs(2167), ZN => n1679);
   U2431 : AOI22_X1 port map( A1 => n85, A2 => regs(1655), B1 => n33, B2 => 
                           regs(631), ZN => n1678);
   U2432 : OAI211_X1 port map( C1 => n58, C2 => n1680, A => n1679, B => n1678, 
                           ZN => curr_proc_regs(631));
   U2433 : AOI22_X1 port map( A1 => n119, A2 => regs(120), B1 => n74, B2 => 
                           regs(2168), ZN => n1682);
   U2434 : AOI22_X1 port map( A1 => n85, A2 => regs(1656), B1 => n31, B2 => 
                           regs(632), ZN => n1681);
   U2435 : OAI211_X1 port map( C1 => n57, C2 => n1683, A => n1682, B => n1681, 
                           ZN => curr_proc_regs(632));
   U2436 : AOI22_X1 port map( A1 => n119, A2 => regs(121), B1 => n74, B2 => 
                           regs(2169), ZN => n1685);
   U2437 : AOI22_X1 port map( A1 => n3, A2 => regs(1145), B1 => n86, B2 => 
                           regs(1657), ZN => n1684);
   U2438 : OAI211_X1 port map( C1 => n2128, C2 => n1686, A => n1685, B => n1684
                           , ZN => curr_proc_regs(633));
   U2439 : AOI22_X1 port map( A1 => n119, A2 => regs(122), B1 => n74, B2 => 
                           regs(2170), ZN => n1688);
   U2440 : AOI22_X1 port map( A1 => n85, A2 => regs(1658), B1 => n21, B2 => 
                           regs(634), ZN => n1687);
   U2441 : OAI211_X1 port map( C1 => n59, C2 => n1689, A => n1688, B => n1687, 
                           ZN => curr_proc_regs(634));
   U2442 : AOI22_X1 port map( A1 => n119, A2 => regs(123), B1 => n74, B2 => 
                           regs(2171), ZN => n1691);
   U2443 : AOI22_X1 port map( A1 => n3, A2 => regs(1147), B1 => n88, B2 => 
                           regs(1659), ZN => n1690);
   U2444 : OAI211_X1 port map( C1 => n14, C2 => n1692, A => n1691, B => n1690, 
                           ZN => curr_proc_regs(635));
   U2445 : AOI22_X1 port map( A1 => n119, A2 => regs(124), B1 => n74, B2 => 
                           regs(2172), ZN => n1694);
   U2446 : AOI22_X1 port map( A1 => n84, A2 => regs(1660), B1 => n22, B2 => 
                           regs(636), ZN => n1693);
   U2447 : OAI211_X1 port map( C1 => n59, C2 => n1695, A => n1694, B => n1693, 
                           ZN => curr_proc_regs(636));
   U2448 : AOI22_X1 port map( A1 => n119, A2 => regs(125), B1 => n74, B2 => 
                           regs(2173), ZN => n1697);
   U2449 : AOI22_X1 port map( A1 => n84, A2 => regs(1661), B1 => n23, B2 => 
                           regs(637), ZN => n1696);
   U2450 : OAI211_X1 port map( C1 => n59, C2 => n1698, A => n1697, B => n1696, 
                           ZN => curr_proc_regs(637));
   U2451 : AOI22_X1 port map( A1 => n119, A2 => regs(126), B1 => n74, B2 => 
                           regs(2174), ZN => n1700);
   U2452 : AOI22_X1 port map( A1 => n84, A2 => regs(1662), B1 => n24, B2 => 
                           regs(638), ZN => n1699);
   U2453 : OAI211_X1 port map( C1 => n59, C2 => n1701, A => n1700, B => n1699, 
                           ZN => curr_proc_regs(638));
   U2454 : AOI22_X1 port map( A1 => n119, A2 => regs(127), B1 => n74, B2 => 
                           regs(2175), ZN => n1703);
   U2455 : AOI22_X1 port map( A1 => n84, A2 => regs(1663), B1 => n23, B2 => 
                           regs(639), ZN => n1702);
   U2456 : OAI211_X1 port map( C1 => n59, C2 => n1704, A => n1703, B => n1702, 
                           ZN => curr_proc_regs(639));
   U2457 : INV_X1 port map( A => regs(1087), ZN => n1707);
   U2458 : AOI22_X1 port map( A1 => n119, A2 => regs(2111), B1 => n74, B2 => 
                           regs(1599), ZN => n1706);
   U2459 : AOI22_X1 port map( A1 => n3, A2 => regs(575), B1 => n29, B2 => 
                           regs(63), ZN => n1705);
   U2460 : OAI211_X1 port map( C1 => n103, C2 => n1707, A => n1706, B => n1705,
                           ZN => curr_proc_regs(63));
   U2461 : AOI22_X1 port map( A1 => n108, A2 => regs(128), B1 => n71, B2 => 
                           regs(2176), ZN => n1709);
   U2462 : AOI22_X1 port map( A1 => n84, A2 => regs(1664), B1 => n38, B2 => 
                           regs(640), ZN => n1708);
   U2463 : OAI211_X1 port map( C1 => n59, C2 => n1710, A => n1709, B => n1708, 
                           ZN => curr_proc_regs(640));
   U2464 : AOI22_X1 port map( A1 => n116, A2 => regs(129), B1 => n71, B2 => 
                           regs(2177), ZN => n1712);
   U2465 : AOI22_X1 port map( A1 => n44, A2 => regs(1153), B1 => n93, B2 => 
                           regs(1665), ZN => n1711);
   U2466 : OAI211_X1 port map( C1 => n2128, C2 => n1713, A => n1712, B => n1711
                           , ZN => curr_proc_regs(641));
   U2467 : AOI22_X1 port map( A1 => n117, A2 => regs(130), B1 => n71, B2 => 
                           regs(2178), ZN => n1715);
   U2468 : AOI22_X1 port map( A1 => n84, A2 => regs(1666), B1 => n36, B2 => 
                           regs(642), ZN => n1714);
   U2469 : OAI211_X1 port map( C1 => n59, C2 => n1716, A => n1715, B => n1714, 
                           ZN => curr_proc_regs(642));
   U2470 : AOI22_X1 port map( A1 => n118, A2 => regs(131), B1 => n71, B2 => 
                           regs(2179), ZN => n1718);
   U2471 : AOI22_X1 port map( A1 => n84, A2 => regs(1667), B1 => n37, B2 => 
                           regs(643), ZN => n1717);
   U2472 : OAI211_X1 port map( C1 => n59, C2 => n1719, A => n1718, B => n1717, 
                           ZN => curr_proc_regs(643));
   U2473 : AOI22_X1 port map( A1 => n122, A2 => regs(132), B1 => n71, B2 => 
                           regs(2180), ZN => n1721);
   U2474 : AOI22_X1 port map( A1 => n84, A2 => regs(1668), B1 => n34, B2 => 
                           regs(644), ZN => n1720);
   U2475 : OAI211_X1 port map( C1 => n59, C2 => n1722, A => n1721, B => n1720, 
                           ZN => curr_proc_regs(644));
   U2476 : AOI22_X1 port map( A1 => n108, A2 => regs(133), B1 => n71, B2 => 
                           regs(2181), ZN => n1724);
   U2477 : AOI22_X1 port map( A1 => n84, A2 => regs(1669), B1 => n20, B2 => 
                           regs(645), ZN => n1723);
   U2478 : OAI211_X1 port map( C1 => n59, C2 => n1725, A => n1724, B => n1723, 
                           ZN => curr_proc_regs(645));
   U2479 : AOI22_X1 port map( A1 => n116, A2 => regs(134), B1 => n71, B2 => 
                           regs(2182), ZN => n1727);
   U2480 : AOI22_X1 port map( A1 => n84, A2 => regs(1670), B1 => n19, B2 => 
                           regs(646), ZN => n1726);
   U2481 : OAI211_X1 port map( C1 => n59, C2 => n1728, A => n1727, B => n1726, 
                           ZN => curr_proc_regs(646));
   U2482 : AOI22_X1 port map( A1 => n116, A2 => regs(135), B1 => n71, B2 => 
                           regs(2183), ZN => n1730);
   U2483 : AOI22_X1 port map( A1 => n45, A2 => regs(1159), B1 => n90, B2 => 
                           regs(1671), ZN => n1729);
   U2484 : OAI211_X1 port map( C1 => n2128, C2 => n1731, A => n1730, B => n1729
                           , ZN => curr_proc_regs(647));
   U2485 : AOI22_X1 port map( A1 => n117, A2 => regs(136), B1 => n71, B2 => 
                           regs(2184), ZN => n1733);
   U2486 : AOI22_X1 port map( A1 => n45, A2 => regs(1160), B1 => n93, B2 => 
                           regs(1672), ZN => n1732);
   U2487 : OAI211_X1 port map( C1 => n12, C2 => n1734, A => n1733, B => n1732, 
                           ZN => curr_proc_regs(648));
   U2488 : AOI22_X1 port map( A1 => n118, A2 => regs(137), B1 => n71, B2 => 
                           regs(2185), ZN => n1736);
   U2489 : AOI22_X1 port map( A1 => n84, A2 => regs(1673), B1 => n39, B2 => 
                           regs(649), ZN => n1735);
   U2490 : OAI211_X1 port map( C1 => n59, C2 => n1737, A => n1736, B => n1735, 
                           ZN => curr_proc_regs(649));
   U2491 : AOI22_X1 port map( A1 => n116, A2 => regs(2112), B1 => n71, B2 => 
                           regs(1600), ZN => n1739);
   U2492 : AOI22_X1 port map( A1 => n45, A2 => regs(576), B1 => n35, B2 => 
                           regs(64), ZN => n1738);
   U2493 : OAI211_X1 port map( C1 => n78, C2 => n1740, A => n1739, B => n1738, 
                           ZN => curr_proc_regs(64));
   U2494 : AOI22_X1 port map( A1 => n116, A2 => regs(138), B1 => n71, B2 => 
                           regs(2186), ZN => n1742);
   U2495 : AOI22_X1 port map( A1 => n45, A2 => regs(1162), B1 => n87, B2 => 
                           regs(1674), ZN => n1741);
   U2496 : OAI211_X1 port map( C1 => n12, C2 => n1743, A => n1742, B => n1741, 
                           ZN => curr_proc_regs(650));
   U2497 : AOI22_X1 port map( A1 => n117, A2 => regs(139), B1 => n5, B2 => 
                           regs(2187), ZN => n1745);
   U2498 : AOI22_X1 port map( A1 => n84, A2 => regs(1675), B1 => n21, B2 => 
                           regs(651), ZN => n1744);
   U2499 : OAI211_X1 port map( C1 => n59, C2 => n1746, A => n1745, B => n1744, 
                           ZN => curr_proc_regs(651));
   U2500 : AOI22_X1 port map( A1 => n118, A2 => regs(140), B1 => n74, B2 => 
                           regs(2188), ZN => n1748);
   U2501 : AOI22_X1 port map( A1 => n45, A2 => regs(1164), B1 => n99, B2 => 
                           regs(1676), ZN => n1747);
   U2502 : OAI211_X1 port map( C1 => n12, C2 => n1749, A => n1748, B => n1747, 
                           ZN => curr_proc_regs(652));
   U2503 : AOI22_X1 port map( A1 => n117, A2 => regs(141), B1 => n5, B2 => 
                           regs(2189), ZN => n1751);
   U2504 : AOI22_X1 port map( A1 => n83, A2 => regs(1677), B1 => n28, B2 => 
                           regs(653), ZN => n1750);
   U2505 : OAI211_X1 port map( C1 => n59, C2 => n1752, A => n1751, B => n1750, 
                           ZN => curr_proc_regs(653));
   U2506 : AOI22_X1 port map( A1 => n106, A2 => regs(142), B1 => n74, B2 => 
                           regs(2190), ZN => n1754);
   U2507 : AOI22_X1 port map( A1 => n45, A2 => regs(1166), B1 => n97, B2 => 
                           regs(1678), ZN => n1753);
   U2508 : OAI211_X1 port map( C1 => n12, C2 => n1755, A => n1754, B => n1753, 
                           ZN => curr_proc_regs(654));
   U2509 : AOI22_X1 port map( A1 => n116, A2 => regs(143), B1 => n5, B2 => 
                           regs(2191), ZN => n1757);
   U2510 : AOI22_X1 port map( A1 => n83, A2 => regs(1679), B1 => n17, B2 => 
                           regs(655), ZN => n1756);
   U2511 : OAI211_X1 port map( C1 => n59, C2 => n1758, A => n1757, B => n1756, 
                           ZN => curr_proc_regs(655));
   U2512 : AOI22_X1 port map( A1 => n117, A2 => regs(144), B1 => n74, B2 => 
                           regs(2192), ZN => n1760);
   U2513 : AOI22_X1 port map( A1 => n83, A2 => regs(1680), B1 => n18, B2 => 
                           regs(656), ZN => n1759);
   U2514 : OAI211_X1 port map( C1 => n59, C2 => n1761, A => n1760, B => n1759, 
                           ZN => curr_proc_regs(656));
   U2515 : AOI22_X1 port map( A1 => n118, A2 => regs(145), B1 => n5, B2 => 
                           regs(2193), ZN => n1763);
   U2516 : AOI22_X1 port map( A1 => n45, A2 => regs(1169), B1 => n102, B2 => 
                           regs(1681), ZN => n1762);
   U2517 : OAI211_X1 port map( C1 => n12, C2 => n1764, A => n1763, B => n1762, 
                           ZN => curr_proc_regs(657));
   U2518 : AOI22_X1 port map( A1 => n118, A2 => regs(146), B1 => n74, B2 => 
                           regs(2194), ZN => n1766);
   U2519 : AOI22_X1 port map( A1 => n83, A2 => regs(1682), B1 => n19, B2 => 
                           regs(658), ZN => n1765);
   U2520 : OAI211_X1 port map( C1 => n2201, C2 => n1767, A => n1766, B => n1765
                           , ZN => curr_proc_regs(658));
   U2521 : AOI22_X1 port map( A1 => n107, A2 => regs(147), B1 => n5, B2 => 
                           regs(2195), ZN => n1769);
   U2522 : AOI22_X1 port map( A1 => n83, A2 => regs(1683), B1 => n21, B2 => 
                           regs(659), ZN => n1768);
   U2523 : OAI211_X1 port map( C1 => n59, C2 => n1770, A => n1769, B => n1768, 
                           ZN => curr_proc_regs(659));
   U2524 : INV_X1 port map( A => regs(577), ZN => n1773);
   U2525 : AOI22_X1 port map( A1 => n116, A2 => regs(2113), B1 => n74, B2 => 
                           regs(1601), ZN => n1772);
   U2526 : AOI22_X1 port map( A1 => n83, A2 => regs(1089), B1 => n38, B2 => 
                           regs(65), ZN => n1771);
   U2527 : OAI211_X1 port map( C1 => n2201, C2 => n1773, A => n1772, B => n1771
                           , ZN => curr_proc_regs(65));
   U2528 : AOI22_X1 port map( A1 => n117, A2 => regs(148), B1 => n5, B2 => 
                           regs(2196), ZN => n1775);
   U2529 : AOI22_X1 port map( A1 => n45, A2 => regs(1172), B1 => n101, B2 => 
                           regs(1684), ZN => n1774);
   U2530 : OAI211_X1 port map( C1 => n12, C2 => n1776, A => n1775, B => n1774, 
                           ZN => curr_proc_regs(660));
   U2531 : AOI22_X1 port map( A1 => n118, A2 => regs(149), B1 => n74, B2 => 
                           regs(2197), ZN => n1778);
   U2532 : AOI22_X1 port map( A1 => n83, A2 => regs(1685), B1 => n34, B2 => 
                           regs(661), ZN => n1777);
   U2533 : OAI211_X1 port map( C1 => n59, C2 => n1779, A => n1778, B => n1777, 
                           ZN => curr_proc_regs(661));
   U2534 : AOI22_X1 port map( A1 => n129, A2 => regs(150), B1 => n63, B2 => 
                           regs(2198), ZN => n1781);
   U2535 : AOI22_X1 port map( A1 => n83, A2 => regs(1686), B1 => n34, B2 => 
                           regs(662), ZN => n1780);
   U2536 : OAI211_X1 port map( C1 => n2201, C2 => n1782, A => n1781, B => n1780
                           , ZN => curr_proc_regs(662));
   U2537 : AOI22_X1 port map( A1 => n116, A2 => regs(151), B1 => n72, B2 => 
                           regs(2199), ZN => n1784);
   U2538 : AOI22_X1 port map( A1 => n83, A2 => regs(1687), B1 => n17, B2 => 
                           regs(663), ZN => n1783);
   U2539 : OAI211_X1 port map( C1 => n59, C2 => n1785, A => n1784, B => n1783, 
                           ZN => curr_proc_regs(663));
   U2540 : AOI22_X1 port map( A1 => n117, A2 => regs(152), B1 => n72, B2 => 
                           regs(2200), ZN => n1787);
   U2541 : AOI22_X1 port map( A1 => n45, A2 => regs(1176), B1 => n102, B2 => 
                           regs(1688), ZN => n1786);
   U2542 : OAI211_X1 port map( C1 => n15, C2 => n1788, A => n1787, B => n1786, 
                           ZN => curr_proc_regs(664));
   U2543 : AOI22_X1 port map( A1 => n118, A2 => regs(153), B1 => n70, B2 => 
                           regs(2201), ZN => n1790);
   U2544 : AOI22_X1 port map( A1 => n45, A2 => regs(1177), B1 => n101, B2 => 
                           regs(1689), ZN => n1789);
   U2545 : OAI211_X1 port map( C1 => n2128, C2 => n1791, A => n1790, B => n1789
                           , ZN => curr_proc_regs(665));
   U2546 : AOI22_X1 port map( A1 => n111, A2 => regs(154), B1 => n74, B2 => 
                           regs(2202), ZN => n1793);
   U2547 : AOI22_X1 port map( A1 => n45, A2 => regs(1178), B1 => n102, B2 => 
                           regs(1690), ZN => n1792);
   U2548 : OAI211_X1 port map( C1 => n15, C2 => n1794, A => n1793, B => n1792, 
                           ZN => curr_proc_regs(666));
   U2549 : AOI22_X1 port map( A1 => n116, A2 => regs(155), B1 => n65, B2 => 
                           regs(2203), ZN => n1796);
   U2550 : AOI22_X1 port map( A1 => n45, A2 => regs(1179), B1 => n101, B2 => 
                           regs(1691), ZN => n1795);
   U2551 : OAI211_X1 port map( C1 => n15, C2 => n1797, A => n1796, B => n1795, 
                           ZN => curr_proc_regs(667));
   U2552 : AOI22_X1 port map( A1 => n117, A2 => regs(156), B1 => n69, B2 => 
                           regs(2204), ZN => n1799);
   U2553 : AOI22_X1 port map( A1 => n44, A2 => regs(1180), B1 => n102, B2 => 
                           regs(1692), ZN => n1798);
   U2554 : OAI211_X1 port map( C1 => n15, C2 => n1800, A => n1799, B => n1798, 
                           ZN => curr_proc_regs(668));
   U2555 : AOI22_X1 port map( A1 => n118, A2 => regs(157), B1 => n63, B2 => 
                           regs(2205), ZN => n1802);
   U2556 : AOI22_X1 port map( A1 => n44, A2 => regs(1181), B1 => n101, B2 => 
                           regs(1693), ZN => n1801);
   U2557 : OAI211_X1 port map( C1 => n15, C2 => n1803, A => n1802, B => n1801, 
                           ZN => curr_proc_regs(669));
   U2558 : AOI22_X1 port map( A1 => n110, A2 => regs(2114), B1 => n66, B2 => 
                           regs(1602), ZN => n1805);
   U2559 : AOI22_X1 port map( A1 => n44, A2 => regs(578), B1 => n27, B2 => 
                           regs(66), ZN => n1804);
   U2560 : OAI211_X1 port map( C1 => n103, C2 => n1806, A => n1805, B => n1804,
                           ZN => curr_proc_regs(66));
   U2561 : AOI22_X1 port map( A1 => n116, A2 => regs(158), B1 => n66, B2 => 
                           regs(2206), ZN => n1808);
   U2562 : AOI22_X1 port map( A1 => n83, A2 => regs(1694), B1 => n26, B2 => 
                           regs(670), ZN => n1807);
   U2563 : OAI211_X1 port map( C1 => n2201, C2 => n1809, A => n1808, B => n1807
                           , ZN => curr_proc_regs(670));
   U2564 : AOI22_X1 port map( A1 => n117, A2 => regs(159), B1 => n5, B2 => 
                           regs(2207), ZN => n1811);
   U2565 : AOI22_X1 port map( A1 => n83, A2 => regs(1695), B1 => n25, B2 => 
                           regs(671), ZN => n1810);
   U2566 : OAI211_X1 port map( C1 => n40, C2 => n1812, A => n1811, B => n1810, 
                           ZN => curr_proc_regs(671));
   U2567 : AOI22_X1 port map( A1 => n118, A2 => regs(160), B1 => n74, B2 => 
                           regs(2208), ZN => n1814);
   U2568 : AOI22_X1 port map( A1 => n83, A2 => regs(1696), B1 => n31, B2 => 
                           regs(672), ZN => n1813);
   U2569 : OAI211_X1 port map( C1 => n40, C2 => n1815, A => n1814, B => n1813, 
                           ZN => curr_proc_regs(672));
   U2570 : AOI22_X1 port map( A1 => n118, A2 => regs(161), B1 => n73, B2 => 
                           regs(2209), ZN => n1817);
   U2571 : AOI22_X1 port map( A1 => n44, A2 => regs(1185), B1 => n102, B2 => 
                           regs(1697), ZN => n1816);
   U2572 : OAI211_X1 port map( C1 => n15, C2 => n1818, A => n1817, B => n1816, 
                           ZN => curr_proc_regs(673));
   U2573 : AOI22_X1 port map( A1 => n118, A2 => regs(162), B1 => n73, B2 => 
                           regs(2210), ZN => n1820);
   U2574 : AOI22_X1 port map( A1 => n82, A2 => regs(1698), B1 => n30, B2 => 
                           regs(674), ZN => n1819);
   U2575 : OAI211_X1 port map( C1 => n40, C2 => n1821, A => n1820, B => n1819, 
                           ZN => curr_proc_regs(674));
   U2576 : AOI22_X1 port map( A1 => n118, A2 => regs(163), B1 => n73, B2 => 
                           regs(2211), ZN => n1823);
   U2577 : AOI22_X1 port map( A1 => n82, A2 => regs(1699), B1 => n32, B2 => 
                           regs(675), ZN => n1822);
   U2578 : OAI211_X1 port map( C1 => n40, C2 => n1824, A => n1823, B => n1822, 
                           ZN => curr_proc_regs(675));
   U2579 : AOI22_X1 port map( A1 => n118, A2 => regs(164), B1 => n73, B2 => 
                           regs(2212), ZN => n1826);
   U2580 : AOI22_X1 port map( A1 => n44, A2 => regs(1188), B1 => n101, B2 => 
                           regs(1700), ZN => n1825);
   U2581 : OAI211_X1 port map( C1 => n12, C2 => n1827, A => n1826, B => n1825, 
                           ZN => curr_proc_regs(676));
   U2582 : AOI22_X1 port map( A1 => n118, A2 => regs(165), B1 => n73, B2 => 
                           regs(2213), ZN => n1829);
   U2583 : AOI22_X1 port map( A1 => n82, A2 => regs(1701), B1 => n35, B2 => 
                           regs(677), ZN => n1828);
   U2584 : OAI211_X1 port map( C1 => n2201, C2 => n1830, A => n1829, B => n1828
                           , ZN => curr_proc_regs(677));
   U2585 : AOI22_X1 port map( A1 => n118, A2 => regs(166), B1 => n73, B2 => 
                           regs(2214), ZN => n1832);
   U2586 : AOI22_X1 port map( A1 => n44, A2 => regs(1190), B1 => n102, B2 => 
                           regs(1702), ZN => n1831);
   U2587 : OAI211_X1 port map( C1 => n12, C2 => n1833, A => n1832, B => n1831, 
                           ZN => curr_proc_regs(678));
   U2588 : AOI22_X1 port map( A1 => n118, A2 => regs(167), B1 => n73, B2 => 
                           regs(2215), ZN => n1835);
   U2589 : AOI22_X1 port map( A1 => n44, A2 => regs(1191), B1 => n101, B2 => 
                           regs(1703), ZN => n1834);
   U2590 : OAI211_X1 port map( C1 => n12, C2 => n1836, A => n1835, B => n1834, 
                           ZN => curr_proc_regs(679));
   U2591 : INV_X1 port map( A => regs(579), ZN => n1839);
   U2592 : AOI22_X1 port map( A1 => n118, A2 => regs(2115), B1 => n5, B2 => 
                           regs(1603), ZN => n1838);
   U2593 : AOI22_X1 port map( A1 => n82, A2 => regs(1091), B1 => n39, B2 => 
                           regs(67), ZN => n1837);
   U2594 : OAI211_X1 port map( C1 => n40, C2 => n1839, A => n1838, B => n1837, 
                           ZN => curr_proc_regs(67));
   U2595 : AOI22_X1 port map( A1 => n118, A2 => regs(168), B1 => n74, B2 => 
                           regs(2216), ZN => n1841);
   U2596 : AOI22_X1 port map( A1 => n44, A2 => regs(1192), B1 => n101, B2 => 
                           regs(1704), ZN => n1840);
   U2597 : OAI211_X1 port map( C1 => n12, C2 => n1842, A => n1841, B => n1840, 
                           ZN => curr_proc_regs(680));
   U2598 : AOI22_X1 port map( A1 => n118, A2 => regs(169), B1 => n5, B2 => 
                           regs(2217), ZN => n1844);
   U2599 : AOI22_X1 port map( A1 => n82, A2 => regs(1705), B1 => n38, B2 => 
                           regs(681), ZN => n1843);
   U2600 : OAI211_X1 port map( C1 => n40, C2 => n1845, A => n1844, B => n1843, 
                           ZN => curr_proc_regs(681));
   U2601 : AOI22_X1 port map( A1 => n118, A2 => regs(170), B1 => n74, B2 => 
                           regs(2218), ZN => n1847);
   U2602 : AOI22_X1 port map( A1 => n82, A2 => regs(1706), B1 => n37, B2 => 
                           regs(682), ZN => n1846);
   U2603 : OAI211_X1 port map( C1 => n40, C2 => n1848, A => n1847, B => n1846, 
                           ZN => curr_proc_regs(682));
   U2604 : AOI22_X1 port map( A1 => n118, A2 => regs(171), B1 => n5, B2 => 
                           regs(2219), ZN => n1850);
   U2605 : AOI22_X1 port map( A1 => n82, A2 => regs(1707), B1 => n36, B2 => 
                           regs(683), ZN => n1849);
   U2606 : OAI211_X1 port map( C1 => n40, C2 => n1851, A => n1850, B => n1849, 
                           ZN => curr_proc_regs(683));
   U2607 : AOI22_X1 port map( A1 => n117, A2 => regs(172), B1 => n72, B2 => 
                           regs(2220), ZN => n1853);
   U2608 : AOI22_X1 port map( A1 => n82, A2 => regs(1708), B1 => n34, B2 => 
                           regs(684), ZN => n1852);
   U2609 : OAI211_X1 port map( C1 => n2201, C2 => n1854, A => n1853, B => n1852
                           , ZN => curr_proc_regs(684));
   U2610 : AOI22_X1 port map( A1 => n117, A2 => regs(173), B1 => n72, B2 => 
                           regs(2221), ZN => n1856);
   U2611 : AOI22_X1 port map( A1 => n82, A2 => regs(1709), B1 => n33, B2 => 
                           regs(685), ZN => n1855);
   U2612 : OAI211_X1 port map( C1 => n40, C2 => n1857, A => n1856, B => n1855, 
                           ZN => curr_proc_regs(685));
   U2613 : AOI22_X1 port map( A1 => n117, A2 => regs(174), B1 => n72, B2 => 
                           regs(2222), ZN => n1859);
   U2614 : AOI22_X1 port map( A1 => n44, A2 => regs(1198), B1 => n101, B2 => 
                           regs(1710), ZN => n1858);
   U2615 : OAI211_X1 port map( C1 => n12, C2 => n1860, A => n1859, B => n1858, 
                           ZN => curr_proc_regs(686));
   U2616 : AOI22_X1 port map( A1 => n117, A2 => regs(175), B1 => n72, B2 => 
                           regs(2223), ZN => n1862);
   U2617 : AOI22_X1 port map( A1 => n44, A2 => regs(1199), B1 => n101, B2 => 
                           regs(1711), ZN => n1861);
   U2618 : OAI211_X1 port map( C1 => n12, C2 => n1863, A => n1862, B => n1861, 
                           ZN => curr_proc_regs(687));
   U2619 : AOI22_X1 port map( A1 => n117, A2 => regs(176), B1 => n72, B2 => 
                           regs(2224), ZN => n1865);
   U2620 : AOI22_X1 port map( A1 => n82, A2 => regs(1712), B1 => n31, B2 => 
                           regs(688), ZN => n1864);
   U2621 : OAI211_X1 port map( C1 => n2201, C2 => n1866, A => n1865, B => n1864
                           , ZN => curr_proc_regs(688));
   U2622 : AOI22_X1 port map( A1 => n117, A2 => regs(177), B1 => n72, B2 => 
                           regs(2225), ZN => n1868);
   U2623 : AOI22_X1 port map( A1 => n44, A2 => regs(1201), B1 => n101, B2 => 
                           regs(1713), ZN => n1867);
   U2624 : OAI211_X1 port map( C1 => n12, C2 => n1869, A => n1868, B => n1867, 
                           ZN => curr_proc_regs(689));
   U2625 : INV_X1 port map( A => regs(580), ZN => n1872);
   U2626 : AOI22_X1 port map( A1 => n117, A2 => regs(2116), B1 => n72, B2 => 
                           regs(1604), ZN => n1871);
   U2627 : AOI22_X1 port map( A1 => n82, A2 => regs(1092), B1 => n21, B2 => 
                           regs(68), ZN => n1870);
   U2628 : OAI211_X1 port map( C1 => n40, C2 => n1872, A => n1871, B => n1870, 
                           ZN => curr_proc_regs(68));
   U2629 : AOI22_X1 port map( A1 => n117, A2 => regs(178), B1 => n72, B2 => 
                           regs(2226), ZN => n1874);
   U2630 : AOI22_X1 port map( A1 => n92, A2 => regs(1714), B1 => n22, B2 => 
                           regs(690), ZN => n1873);
   U2631 : OAI211_X1 port map( C1 => n40, C2 => n1875, A => n1874, B => n1873, 
                           ZN => curr_proc_regs(690));
   U2632 : AOI22_X1 port map( A1 => n117, A2 => regs(179), B1 => n72, B2 => 
                           regs(2227), ZN => n1877);
   U2633 : AOI22_X1 port map( A1 => n43, A2 => regs(1203), B1 => n101, B2 => 
                           regs(1715), ZN => n1876);
   U2634 : OAI211_X1 port map( C1 => n15, C2 => n1878, A => n1877, B => n1876, 
                           ZN => curr_proc_regs(691));
   U2635 : AOI22_X1 port map( A1 => n117, A2 => regs(180), B1 => n72, B2 => 
                           regs(2228), ZN => n1880);
   U2636 : AOI22_X1 port map( A1 => n45, A2 => regs(1204), B1 => n101, B2 => 
                           regs(1716), ZN => n1879);
   U2637 : OAI211_X1 port map( C1 => n15, C2 => n1881, A => n1880, B => n1879, 
                           ZN => curr_proc_regs(692));
   U2638 : AOI22_X1 port map( A1 => n117, A2 => regs(181), B1 => n72, B2 => 
                           regs(2229), ZN => n1883);
   U2639 : AOI22_X1 port map( A1 => n45, A2 => regs(1205), B1 => n101, B2 => 
                           regs(1717), ZN => n1882);
   U2640 : OAI211_X1 port map( C1 => n15, C2 => n1884, A => n1883, B => n1882, 
                           ZN => curr_proc_regs(693));
   U2641 : AOI22_X1 port map( A1 => n117, A2 => regs(182), B1 => n72, B2 => 
                           regs(2230), ZN => n1886);
   U2642 : AOI22_X1 port map( A1 => n42, A2 => regs(1206), B1 => n101, B2 => 
                           regs(1718), ZN => n1885);
   U2643 : OAI211_X1 port map( C1 => n15, C2 => n1887, A => n1886, B => n1885, 
                           ZN => curr_proc_regs(694));
   U2644 : AOI22_X1 port map( A1 => n118, A2 => regs(183), B1 => n73, B2 => 
                           regs(2231), ZN => n1889);
   U2645 : AOI22_X1 port map( A1 => n41, A2 => regs(1207), B1 => n101, B2 => 
                           regs(1719), ZN => n1888);
   U2646 : OAI211_X1 port map( C1 => n15, C2 => n1890, A => n1889, B => n1888, 
                           ZN => curr_proc_regs(695));
   U2647 : AOI22_X1 port map( A1 => n119, A2 => regs(184), B1 => n73, B2 => 
                           regs(2232), ZN => n1892);
   U2648 : AOI22_X1 port map( A1 => n53, A2 => regs(1208), B1 => n101, B2 => 
                           regs(1720), ZN => n1891);
   U2649 : OAI211_X1 port map( C1 => n15, C2 => n1893, A => n1892, B => n1891, 
                           ZN => curr_proc_regs(696));
   U2650 : AOI22_X1 port map( A1 => n121, A2 => regs(185), B1 => n73, B2 => 
                           regs(2233), ZN => n1895);
   U2651 : AOI22_X1 port map( A1 => n56, A2 => regs(1209), B1 => n101, B2 => 
                           regs(1721), ZN => n1894);
   U2652 : OAI211_X1 port map( C1 => n15, C2 => n1896, A => n1895, B => n1894, 
                           ZN => curr_proc_regs(697));
   U2653 : AOI22_X1 port map( A1 => n123, A2 => regs(186), B1 => n73, B2 => 
                           regs(2234), ZN => n1898);
   U2654 : AOI22_X1 port map( A1 => n83, A2 => regs(1722), B1 => n24, B2 => 
                           regs(698), ZN => n1897);
   U2655 : OAI211_X1 port map( C1 => n40, C2 => n1899, A => n1898, B => n1897, 
                           ZN => curr_proc_regs(698));
   U2656 : AOI22_X1 port map( A1 => win(4), A2 => regs(187), B1 => n73, B2 => 
                           regs(2235), ZN => n1901);
   U2657 : AOI22_X1 port map( A1 => n86, A2 => regs(1723), B1 => n31, B2 => 
                           regs(699), ZN => n1900);
   U2658 : OAI211_X1 port map( C1 => n40, C2 => n1902, A => n1901, B => n1900, 
                           ZN => curr_proc_regs(699));
   U2659 : INV_X1 port map( A => regs(581), ZN => n1905);
   U2660 : AOI22_X1 port map( A1 => n126, A2 => regs(2117), B1 => n73, B2 => 
                           regs(1605), ZN => n1904);
   U2661 : AOI22_X1 port map( A1 => n89, A2 => regs(1093), B1 => n30, B2 => 
                           regs(69), ZN => n1903);
   U2662 : OAI211_X1 port map( C1 => n2201, C2 => n1905, A => n1904, B => n1903
                           , ZN => curr_proc_regs(69));
   U2663 : AOI22_X1 port map( A1 => n127, A2 => regs(2054), B1 => n73, B2 => 
                           regs(1542), ZN => n1907);
   U2664 : AOI22_X1 port map( A1 => n46, A2 => regs(518), B1 => n37, B2 => 
                           regs(6), ZN => n1906);
   U2665 : OAI211_X1 port map( C1 => n6, C2 => n1908, A => n1907, B => n1906, 
                           ZN => curr_proc_regs(6));
   U2666 : AOI22_X1 port map( A1 => n129, A2 => regs(188), B1 => n73, B2 => 
                           regs(2236), ZN => n1910);
   U2667 : AOI22_X1 port map( A1 => n54, A2 => regs(1212), B1 => n100, B2 => 
                           regs(1724), ZN => n1909);
   U2668 : OAI211_X1 port map( C1 => n15, C2 => n1911, A => n1910, B => n1909, 
                           ZN => curr_proc_regs(700));
   U2669 : AOI22_X1 port map( A1 => n111, A2 => regs(189), B1 => n73, B2 => 
                           regs(2237), ZN => n1913);
   U2670 : AOI22_X1 port map( A1 => n55, A2 => regs(1213), B1 => n100, B2 => 
                           regs(1725), ZN => n1912);
   U2671 : OAI211_X1 port map( C1 => n15, C2 => n1914, A => n1913, B => n1912, 
                           ZN => curr_proc_regs(701));
   U2672 : AOI22_X1 port map( A1 => n110, A2 => regs(190), B1 => n73, B2 => 
                           regs(2238), ZN => n1916);
   U2673 : AOI22_X1 port map( A1 => n42, A2 => regs(1214), B1 => n100, B2 => 
                           regs(1726), ZN => n1915);
   U2674 : OAI211_X1 port map( C1 => n15, C2 => n1917, A => n1916, B => n1915, 
                           ZN => curr_proc_regs(702));
   U2675 : AOI22_X1 port map( A1 => n107, A2 => regs(191), B1 => n73, B2 => 
                           regs(2239), ZN => n1919);
   U2676 : AOI22_X1 port map( A1 => n51, A2 => regs(1215), B1 => n100, B2 => 
                           regs(1727), ZN => n1918);
   U2677 : OAI211_X1 port map( C1 => n15, C2 => n1920, A => n1919, B => n1918, 
                           ZN => curr_proc_regs(703));
   U2678 : AOI22_X1 port map( A1 => n116, A2 => regs(192), B1 => n73, B2 => 
                           regs(2240), ZN => n1922);
   U2679 : AOI22_X1 port map( A1 => n88, A2 => regs(1728), B1 => n36, B2 => 
                           regs(704), ZN => n1921);
   U2680 : OAI211_X1 port map( C1 => n40, C2 => n1923, A => n1922, B => n1921, 
                           ZN => curr_proc_regs(704));
   U2681 : AOI22_X1 port map( A1 => n116, A2 => regs(193), B1 => n66, B2 => 
                           regs(2241), ZN => n1925);
   U2682 : AOI22_X1 port map( A1 => n101, A2 => regs(1729), B1 => n36, B2 => 
                           regs(705), ZN => n1924);
   U2683 : OAI211_X1 port map( C1 => n40, C2 => n1926, A => n1925, B => n1924, 
                           ZN => curr_proc_regs(705));
   U2684 : AOI22_X1 port map( A1 => n116, A2 => regs(194), B1 => n66, B2 => 
                           regs(2242), ZN => n1928);
   U2685 : AOI22_X1 port map( A1 => n102, A2 => regs(1730), B1 => n31, B2 => 
                           regs(706), ZN => n1927);
   U2686 : OAI211_X1 port map( C1 => n2201, C2 => n1929, A => n1928, B => n1927
                           , ZN => curr_proc_regs(706));
   U2687 : AOI22_X1 port map( A1 => n116, A2 => regs(195), B1 => n66, B2 => 
                           regs(2243), ZN => n1931);
   U2688 : AOI22_X1 port map( A1 => n79, A2 => regs(1731), B1 => n20, B2 => 
                           regs(707), ZN => n1930);
   U2689 : OAI211_X1 port map( C1 => n40, C2 => n1932, A => n1931, B => n1930, 
                           ZN => curr_proc_regs(707));
   U2690 : AOI22_X1 port map( A1 => n116, A2 => regs(196), B1 => n66, B2 => 
                           regs(2244), ZN => n1934);
   U2691 : AOI22_X1 port map( A1 => n51, A2 => regs(1220), B1 => n100, B2 => 
                           regs(1732), ZN => n1933);
   U2692 : OAI211_X1 port map( C1 => n15, C2 => n1935, A => n1934, B => n1933, 
                           ZN => curr_proc_regs(708));
   U2693 : AOI22_X1 port map( A1 => n116, A2 => regs(197), B1 => n66, B2 => 
                           regs(2245), ZN => n1937);
   U2694 : AOI22_X1 port map( A1 => n84, A2 => regs(1733), B1 => n27, B2 => 
                           regs(709), ZN => n1936);
   U2695 : OAI211_X1 port map( C1 => n2201, C2 => n1938, A => n1937, B => n1936
                           , ZN => curr_proc_regs(709));
   U2696 : AOI22_X1 port map( A1 => n116, A2 => regs(2118), B1 => n66, B2 => 
                           regs(1606), ZN => n1940);
   U2697 : AOI22_X1 port map( A1 => n51, A2 => regs(582), B1 => n36, B2 => 
                           regs(70), ZN => n1939);
   U2698 : OAI211_X1 port map( C1 => n6, C2 => n1941, A => n1940, B => n1939, 
                           ZN => curr_proc_regs(70));
   U2699 : AOI22_X1 port map( A1 => n116, A2 => regs(198), B1 => n66, B2 => 
                           regs(2246), ZN => n1943);
   U2700 : AOI22_X1 port map( A1 => n82, A2 => regs(1734), B1 => n39, B2 => 
                           regs(710), ZN => n1942);
   U2701 : OAI211_X1 port map( C1 => n2201, C2 => n1944, A => n1943, B => n1942
                           , ZN => curr_proc_regs(710));
   U2702 : AOI22_X1 port map( A1 => n116, A2 => regs(199), B1 => n66, B2 => 
                           regs(2247), ZN => n1946);
   U2703 : AOI22_X1 port map( A1 => n51, A2 => regs(1223), B1 => n99, B2 => 
                           regs(1735), ZN => n1945);
   U2704 : OAI211_X1 port map( C1 => n15, C2 => n1947, A => n1946, B => n1945, 
                           ZN => curr_proc_regs(711));
   U2705 : AOI22_X1 port map( A1 => n116, A2 => regs(200), B1 => n66, B2 => 
                           regs(2248), ZN => n1949);
   U2706 : AOI22_X1 port map( A1 => n81, A2 => regs(1736), B1 => n22, B2 => 
                           regs(712), ZN => n1948);
   U2707 : OAI211_X1 port map( C1 => n10, C2 => n1950, A => n1949, B => n1948, 
                           ZN => curr_proc_regs(712));
   U2708 : AOI22_X1 port map( A1 => n116, A2 => regs(201), B1 => n66, B2 => 
                           regs(2249), ZN => n1952);
   U2709 : AOI22_X1 port map( A1 => n80, A2 => regs(1737), B1 => n22, B2 => 
                           regs(713), ZN => n1951);
   U2710 : OAI211_X1 port map( C1 => n2201, C2 => n1953, A => n1952, B => n1951
                           , ZN => curr_proc_regs(713));
   U2711 : AOI22_X1 port map( A1 => n116, A2 => regs(202), B1 => n66, B2 => 
                           regs(2250), ZN => n1955);
   U2712 : AOI22_X1 port map( A1 => n51, A2 => regs(1226), B1 => n99, B2 => 
                           regs(1738), ZN => n1954);
   U2713 : OAI211_X1 port map( C1 => n2128, C2 => n1956, A => n1955, B => n1954
                           , ZN => curr_proc_regs(714));
   U2714 : AOI22_X1 port map( A1 => n123, A2 => regs(203), B1 => n66, B2 => 
                           regs(2251), ZN => n1958);
   U2715 : AOI22_X1 port map( A1 => n51, A2 => regs(1227), B1 => n98, B2 => 
                           regs(1739), ZN => n1957);
   U2716 : OAI211_X1 port map( C1 => n12, C2 => n1959, A => n1958, B => n1957, 
                           ZN => curr_proc_regs(715));
   U2717 : AOI22_X1 port map( A1 => n126, A2 => regs(204), B1 => n74, B2 => 
                           regs(2252), ZN => n1961);
   U2718 : AOI22_X1 port map( A1 => n81, A2 => regs(1740), B1 => n37, B2 => 
                           regs(716), ZN => n1960);
   U2719 : OAI211_X1 port map( C1 => n2201, C2 => n1962, A => n1961, B => n1960
                           , ZN => curr_proc_regs(716));
   U2720 : AOI22_X1 port map( A1 => n114, A2 => regs(205), B1 => n74, B2 => 
                           regs(2253), ZN => n1964);
   U2721 : AOI22_X1 port map( A1 => n81, A2 => regs(1741), B1 => n31, B2 => 
                           regs(717), ZN => n1963);
   U2722 : OAI211_X1 port map( C1 => n2201, C2 => n1965, A => n1964, B => n1963
                           , ZN => curr_proc_regs(717));
   U2723 : AOI22_X1 port map( A1 => n115, A2 => regs(206), B1 => n74, B2 => 
                           regs(2254), ZN => n1967);
   U2724 : AOI22_X1 port map( A1 => n51, A2 => regs(1230), B1 => n99, B2 => 
                           regs(1742), ZN => n1966);
   U2725 : OAI211_X1 port map( C1 => n12, C2 => n1968, A => n1967, B => n1966, 
                           ZN => curr_proc_regs(718));
   U2726 : AOI22_X1 port map( A1 => win(4), A2 => regs(207), B1 => n74, B2 => 
                           regs(2255), ZN => n1970);
   U2727 : AOI22_X1 port map( A1 => n51, A2 => regs(1231), B1 => n98, B2 => 
                           regs(1743), ZN => n1969);
   U2728 : OAI211_X1 port map( C1 => n12, C2 => n1971, A => n1970, B => n1969, 
                           ZN => curr_proc_regs(719));
   U2729 : INV_X1 port map( A => regs(583), ZN => n1974);
   U2730 : AOI22_X1 port map( A1 => n126, A2 => regs(2119), B1 => n74, B2 => 
                           regs(1607), ZN => n1973);
   U2731 : AOI22_X1 port map( A1 => n81, A2 => regs(1095), B1 => n33, B2 => 
                           regs(71), ZN => n1972);
   U2732 : OAI211_X1 port map( C1 => n2201, C2 => n1974, A => n1973, B => n1972
                           , ZN => curr_proc_regs(71));
   U2733 : AOI22_X1 port map( A1 => n127, A2 => regs(208), B1 => n74, B2 => 
                           regs(2256), ZN => n1976);
   U2734 : AOI22_X1 port map( A1 => n81, A2 => regs(1744), B1 => n18, B2 => 
                           regs(720), ZN => n1975);
   U2735 : OAI211_X1 port map( C1 => n9, C2 => n1977, A => n1976, B => n1975, 
                           ZN => curr_proc_regs(720));
   U2736 : AOI22_X1 port map( A1 => n127, A2 => regs(209), B1 => n74, B2 => 
                           regs(2257), ZN => n1979);
   U2737 : AOI22_X1 port map( A1 => n81, A2 => regs(1745), B1 => n27, B2 => 
                           regs(721), ZN => n1978);
   U2738 : OAI211_X1 port map( C1 => n2201, C2 => n1980, A => n1979, B => n1978
                           , ZN => curr_proc_regs(721));
   U2739 : AOI22_X1 port map( A1 => n114, A2 => regs(210), B1 => n74, B2 => 
                           regs(2258), ZN => n1982);
   U2740 : AOI22_X1 port map( A1 => n81, A2 => regs(1746), B1 => n26, B2 => 
                           regs(722), ZN => n1981);
   U2741 : OAI211_X1 port map( C1 => n10, C2 => n1983, A => n1982, B => n1981, 
                           ZN => curr_proc_regs(722));
   U2742 : AOI22_X1 port map( A1 => n115, A2 => regs(211), B1 => n74, B2 => 
                           regs(2259), ZN => n1985);
   U2743 : AOI22_X1 port map( A1 => n81, A2 => regs(1747), B1 => n25, B2 => 
                           regs(723), ZN => n1984);
   U2744 : OAI211_X1 port map( C1 => n9, C2 => n1986, A => n1985, B => n1984, 
                           ZN => curr_proc_regs(723));
   U2745 : AOI22_X1 port map( A1 => n129, A2 => regs(212), B1 => n74, B2 => 
                           regs(2260), ZN => n1988);
   U2746 : AOI22_X1 port map( A1 => n51, A2 => regs(1236), B1 => n98, B2 => 
                           regs(1748), ZN => n1987);
   U2747 : OAI211_X1 port map( C1 => n12, C2 => n1989, A => n1988, B => n1987, 
                           ZN => curr_proc_regs(724));
   U2748 : AOI22_X1 port map( A1 => n111, A2 => regs(213), B1 => n74, B2 => 
                           regs(2261), ZN => n1991);
   U2749 : AOI22_X1 port map( A1 => n81, A2 => regs(1749), B1 => n23, B2 => 
                           regs(725), ZN => n1990);
   U2750 : OAI211_X1 port map( C1 => n2201, C2 => n1992, A => n1991, B => n1990
                           , ZN => curr_proc_regs(725));
   U2751 : AOI22_X1 port map( A1 => n114, A2 => regs(214), B1 => n74, B2 => 
                           regs(2262), ZN => n1994);
   U2752 : AOI22_X1 port map( A1 => n81, A2 => regs(1750), B1 => n20, B2 => 
                           regs(726), ZN => n1993);
   U2753 : OAI211_X1 port map( C1 => n10, C2 => n1995, A => n1994, B => n1993, 
                           ZN => curr_proc_regs(726));
   U2754 : AOI22_X1 port map( A1 => n115, A2 => regs(215), B1 => n75, B2 => 
                           regs(2263), ZN => n1997);
   U2755 : AOI22_X1 port map( A1 => n81, A2 => regs(1751), B1 => n28, B2 => 
                           regs(727), ZN => n1996);
   U2756 : OAI211_X1 port map( C1 => n9, C2 => n1998, A => n1997, B => n1996, 
                           ZN => curr_proc_regs(727));
   U2757 : AOI22_X1 port map( A1 => n114, A2 => regs(216), B1 => n75, B2 => 
                           regs(2264), ZN => n2000);
   U2758 : AOI22_X1 port map( A1 => n81, A2 => regs(1752), B1 => n4, B2 => 
                           regs(728), ZN => n1999);
   U2759 : OAI211_X1 port map( C1 => n2201, C2 => n2001, A => n2000, B => n1999
                           , ZN => curr_proc_regs(728));
   U2760 : AOI22_X1 port map( A1 => n119, A2 => regs(217), B1 => n75, B2 => 
                           regs(2265), ZN => n2003);
   U2761 : AOI22_X1 port map( A1 => n81, A2 => regs(1753), B1 => n38, B2 => 
                           regs(729), ZN => n2002);
   U2762 : OAI211_X1 port map( C1 => n2201, C2 => n2004, A => n2003, B => n2002
                           , ZN => curr_proc_regs(729));
   U2763 : AOI22_X1 port map( A1 => n114, A2 => regs(2120), B1 => n75, B2 => 
                           regs(1608), ZN => n2006);
   U2764 : AOI22_X1 port map( A1 => n51, A2 => regs(584), B1 => n37, B2 => 
                           regs(72), ZN => n2005);
   U2765 : OAI211_X1 port map( C1 => n6, C2 => n2007, A => n2006, B => n2005, 
                           ZN => curr_proc_regs(72));
   U2766 : AOI22_X1 port map( A1 => n114, A2 => regs(218), B1 => n75, B2 => 
                           regs(2266), ZN => n2009);
   U2767 : AOI22_X1 port map( A1 => n100, A2 => regs(1754), B1 => n36, B2 => 
                           regs(730), ZN => n2008);
   U2768 : OAI211_X1 port map( C1 => n2201, C2 => n2010, A => n2009, B => n2008
                           , ZN => curr_proc_regs(730));
   U2769 : AOI22_X1 port map( A1 => n115, A2 => regs(219), B1 => n75, B2 => 
                           regs(2267), ZN => n2012);
   U2770 : AOI22_X1 port map( A1 => n51, A2 => regs(1243), B1 => n98, B2 => 
                           regs(1755), ZN => n2011);
   U2771 : OAI211_X1 port map( C1 => n12, C2 => n2013, A => n2012, B => n2011, 
                           ZN => curr_proc_regs(731));
   U2772 : AOI22_X1 port map( A1 => n115, A2 => regs(220), B1 => n75, B2 => 
                           regs(2268), ZN => n2015);
   U2773 : AOI22_X1 port map( A1 => n52, A2 => regs(1244), B1 => n99, B2 => 
                           regs(1756), ZN => n2014);
   U2774 : OAI211_X1 port map( C1 => n12, C2 => n2016, A => n2015, B => n2014, 
                           ZN => curr_proc_regs(732));
   U2775 : AOI22_X1 port map( A1 => n121, A2 => regs(221), B1 => n75, B2 => 
                           regs(2269), ZN => n2018);
   U2776 : AOI22_X1 port map( A1 => n93, A2 => regs(1757), B1 => n34, B2 => 
                           regs(733), ZN => n2017);
   U2777 : OAI211_X1 port map( C1 => n2201, C2 => n2019, A => n2018, B => n2017
                           , ZN => curr_proc_regs(733));
   U2778 : AOI22_X1 port map( A1 => n115, A2 => regs(222), B1 => n75, B2 => 
                           regs(2270), ZN => n2021);
   U2779 : AOI22_X1 port map( A1 => n50, A2 => regs(1246), B1 => n99, B2 => 
                           regs(1758), ZN => n2020);
   U2780 : OAI211_X1 port map( C1 => n12, C2 => n2022, A => n2021, B => n2020, 
                           ZN => curr_proc_regs(734));
   U2781 : AOI22_X1 port map( A1 => n114, A2 => regs(223), B1 => n75, B2 => 
                           regs(2271), ZN => n2024);
   U2782 : AOI22_X1 port map( A1 => n50, A2 => regs(1247), B1 => n98, B2 => 
                           regs(1759), ZN => n2023);
   U2783 : OAI211_X1 port map( C1 => n15, C2 => n2025, A => n2024, B => n2023, 
                           ZN => curr_proc_regs(735));
   U2784 : AOI22_X1 port map( A1 => n115, A2 => regs(224), B1 => n75, B2 => 
                           regs(2272), ZN => n2027);
   U2785 : AOI22_X1 port map( A1 => n98, A2 => regs(1760), B1 => n33, B2 => 
                           regs(736), ZN => n2026);
   U2786 : OAI211_X1 port map( C1 => n2201, C2 => n2028, A => n2027, B => n2026
                           , ZN => curr_proc_regs(736));
   U2787 : AOI22_X1 port map( A1 => win(4), A2 => regs(225), B1 => n75, B2 => 
                           regs(2273), ZN => n2030);
   U2788 : AOI22_X1 port map( A1 => n97, A2 => regs(1761), B1 => n31, B2 => 
                           regs(737), ZN => n2029);
   U2789 : OAI211_X1 port map( C1 => n59, C2 => n2031, A => n2030, B => n2029, 
                           ZN => curr_proc_regs(737));
   U2790 : AOI22_X1 port map( A1 => n105, A2 => regs(226), B1 => n76, B2 => 
                           regs(2274), ZN => n2033);
   U2791 : AOI22_X1 port map( A1 => n50, A2 => regs(1250), B1 => n99, B2 => 
                           regs(1762), ZN => n2032);
   U2792 : OAI211_X1 port map( C1 => n15, C2 => n2034, A => n2033, B => n2032, 
                           ZN => curr_proc_regs(738));
   U2793 : AOI22_X1 port map( A1 => n114, A2 => regs(227), B1 => n76, B2 => 
                           regs(2275), ZN => n2036);
   U2794 : AOI22_X1 port map( A1 => n90, A2 => regs(1763), B1 => n21, B2 => 
                           regs(739), ZN => n2035);
   U2795 : OAI211_X1 port map( C1 => n2201, C2 => n2037, A => n2036, B => n2035
                           , ZN => curr_proc_regs(739));
   U2796 : AOI22_X1 port map( A1 => n115, A2 => regs(2121), B1 => n76, B2 => 
                           regs(1609), ZN => n2039);
   U2797 : AOI22_X1 port map( A1 => n50, A2 => regs(585), B1 => n22, B2 => 
                           regs(73), ZN => n2038);
   U2798 : OAI211_X1 port map( C1 => n6, C2 => n2040, A => n2039, B => n2038, 
                           ZN => curr_proc_regs(73));
   U2799 : AOI22_X1 port map( A1 => n116, A2 => regs(228), B1 => n76, B2 => 
                           regs(2276), ZN => n2042);
   U2800 : AOI22_X1 port map( A1 => n94, A2 => regs(1764), B1 => n23, B2 => 
                           regs(740), ZN => n2041);
   U2801 : OAI211_X1 port map( C1 => n58, C2 => n2043, A => n2042, B => n2041, 
                           ZN => curr_proc_regs(740));
   U2802 : AOI22_X1 port map( A1 => n120, A2 => regs(229), B1 => n76, B2 => 
                           regs(2277), ZN => n2045);
   U2803 : AOI22_X1 port map( A1 => n95, A2 => regs(1765), B1 => n24, B2 => 
                           regs(741), ZN => n2044);
   U2804 : OAI211_X1 port map( C1 => n58, C2 => n2046, A => n2045, B => n2044, 
                           ZN => curr_proc_regs(741));
   U2805 : AOI22_X1 port map( A1 => n114, A2 => regs(230), B1 => n76, B2 => 
                           regs(2278), ZN => n2048);
   U2806 : AOI22_X1 port map( A1 => n91, A2 => regs(1766), B1 => n17, B2 => 
                           regs(742), ZN => n2047);
   U2807 : OAI211_X1 port map( C1 => n58, C2 => n2049, A => n2048, B => n2047, 
                           ZN => curr_proc_regs(742));
   U2808 : AOI22_X1 port map( A1 => n115, A2 => regs(231), B1 => n76, B2 => 
                           regs(2279), ZN => n2051);
   U2809 : AOI22_X1 port map( A1 => n92, A2 => regs(1767), B1 => n18, B2 => 
                           regs(743), ZN => n2050);
   U2810 : OAI211_X1 port map( C1 => n57, C2 => n2052, A => n2051, B => n2050, 
                           ZN => curr_proc_regs(743));
   U2811 : AOI22_X1 port map( A1 => n118, A2 => regs(232), B1 => n76, B2 => 
                           regs(2280), ZN => n2054);
   U2812 : AOI22_X1 port map( A1 => n83, A2 => regs(1768), B1 => n34, B2 => 
                           regs(744), ZN => n2053);
   U2813 : OAI211_X1 port map( C1 => n58, C2 => n2055, A => n2054, B => n2053, 
                           ZN => curr_proc_regs(744));
   U2814 : AOI22_X1 port map( A1 => n117, A2 => regs(233), B1 => n76, B2 => 
                           regs(2281), ZN => n2057);
   U2815 : AOI22_X1 port map( A1 => n91, A2 => regs(1769), B1 => n20, B2 => 
                           regs(745), ZN => n2056);
   U2816 : OAI211_X1 port map( C1 => n57, C2 => n2058, A => n2057, B => n2056, 
                           ZN => curr_proc_regs(745));
   U2817 : AOI22_X1 port map( A1 => n114, A2 => regs(234), B1 => n76, B2 => 
                           regs(2282), ZN => n2060);
   U2818 : AOI22_X1 port map( A1 => n96, A2 => regs(1770), B1 => n20, B2 => 
                           regs(746), ZN => n2059);
   U2819 : OAI211_X1 port map( C1 => n58, C2 => n2061, A => n2060, B => n2059, 
                           ZN => curr_proc_regs(746));
   U2820 : AOI22_X1 port map( A1 => n115, A2 => regs(235), B1 => n76, B2 => 
                           regs(2283), ZN => n2063);
   U2821 : AOI22_X1 port map( A1 => n50, A2 => regs(1259), B1 => n98, B2 => 
                           regs(1771), ZN => n2062);
   U2822 : OAI211_X1 port map( C1 => n2128, C2 => n2064, A => n2063, B => n2062
                           , ZN => curr_proc_regs(747));
   U2823 : AOI22_X1 port map( A1 => n115, A2 => regs(236), B1 => n76, B2 => 
                           regs(2284), ZN => n2066);
   U2824 : AOI22_X1 port map( A1 => n50, A2 => regs(1260), B1 => n99, B2 => 
                           regs(1772), ZN => n2065);
   U2825 : OAI211_X1 port map( C1 => n15, C2 => n2067, A => n2066, B => n2065, 
                           ZN => curr_proc_regs(748));
   U2826 : AOI22_X1 port map( A1 => n115, A2 => regs(237), B1 => n76, B2 => 
                           regs(2285), ZN => n2069);
   U2827 : AOI22_X1 port map( A1 => n80, A2 => regs(1773), B1 => n26, B2 => 
                           regs(749), ZN => n2068);
   U2828 : OAI211_X1 port map( C1 => n40, C2 => n2070, A => n2069, B => n2068, 
                           ZN => curr_proc_regs(749));
   U2829 : AOI22_X1 port map( A1 => n115, A2 => regs(2122), B1 => n2211, B2 => 
                           regs(1610), ZN => n2072);
   U2830 : AOI22_X1 port map( A1 => n50, A2 => regs(586), B1 => n22, B2 => 
                           regs(74), ZN => n2071);
   U2831 : OAI211_X1 port map( C1 => n6, C2 => n2073, A => n2072, B => n2071, 
                           ZN => curr_proc_regs(74));
   U2832 : AOI22_X1 port map( A1 => n115, A2 => regs(238), B1 => n75, B2 => 
                           regs(2286), ZN => n2075);
   U2833 : AOI22_X1 port map( A1 => n50, A2 => regs(1262), B1 => n99, B2 => 
                           regs(1774), ZN => n2074);
   U2834 : OAI211_X1 port map( C1 => n15, C2 => n2076, A => n2075, B => n2074, 
                           ZN => curr_proc_regs(750));
   U2835 : AOI22_X1 port map( A1 => n115, A2 => regs(239), B1 => n76, B2 => 
                           regs(2287), ZN => n2078);
   U2836 : AOI22_X1 port map( A1 => n50, A2 => regs(1263), B1 => n99, B2 => 
                           regs(1775), ZN => n2077);
   U2837 : OAI211_X1 port map( C1 => n15, C2 => n2079, A => n2078, B => n2077, 
                           ZN => curr_proc_regs(751));
   U2838 : AOI22_X1 port map( A1 => n115, A2 => regs(240), B1 => n67, B2 => 
                           regs(2288), ZN => n2081);
   U2839 : AOI22_X1 port map( A1 => n80, A2 => regs(1776), B1 => n38, B2 => 
                           regs(752), ZN => n2080);
   U2840 : OAI211_X1 port map( C1 => n40, C2 => n2082, A => n2081, B => n2080, 
                           ZN => curr_proc_regs(752));
   U2841 : AOI22_X1 port map( A1 => n115, A2 => regs(241), B1 => n75, B2 => 
                           regs(2289), ZN => n2084);
   U2842 : AOI22_X1 port map( A1 => n50, A2 => regs(1265), B1 => n99, B2 => 
                           regs(1777), ZN => n2083);
   U2843 : OAI211_X1 port map( C1 => n15, C2 => n2085, A => n2084, B => n2083, 
                           ZN => curr_proc_regs(753));
   U2844 : AOI22_X1 port map( A1 => n115, A2 => regs(242), B1 => n76, B2 => 
                           regs(2290), ZN => n2087);
   U2845 : AOI22_X1 port map( A1 => n80, A2 => regs(1778), B1 => n23, B2 => 
                           regs(754), ZN => n2086);
   U2846 : OAI211_X1 port map( C1 => n40, C2 => n2088, A => n2087, B => n2086, 
                           ZN => curr_proc_regs(754));
   U2847 : AOI22_X1 port map( A1 => n115, A2 => regs(243), B1 => n5, B2 => 
                           regs(2291), ZN => n2090);
   U2848 : AOI22_X1 port map( A1 => n50, A2 => regs(1267), B1 => n99, B2 => 
                           regs(1779), ZN => n2089);
   U2849 : OAI211_X1 port map( C1 => n15, C2 => n2091, A => n2090, B => n2089, 
                           ZN => curr_proc_regs(755));
   U2850 : AOI22_X1 port map( A1 => n115, A2 => regs(244), B1 => n75, B2 => 
                           regs(2292), ZN => n2093);
   U2851 : AOI22_X1 port map( A1 => n51, A2 => regs(1268), B1 => n100, B2 => 
                           regs(1780), ZN => n2092);
   U2852 : OAI211_X1 port map( C1 => n15, C2 => n2094, A => n2093, B => n2092, 
                           ZN => curr_proc_regs(756));
   U2853 : AOI22_X1 port map( A1 => n115, A2 => regs(245), B1 => n76, B2 => 
                           regs(2293), ZN => n2096);
   U2854 : AOI22_X1 port map( A1 => n80, A2 => regs(1781), B1 => n28, B2 => 
                           regs(757), ZN => n2095);
   U2855 : OAI211_X1 port map( C1 => n40, C2 => n2097, A => n2096, B => n2095, 
                           ZN => curr_proc_regs(757));
   U2856 : AOI22_X1 port map( A1 => n115, A2 => regs(246), B1 => n73, B2 => 
                           regs(2294), ZN => n2099);
   U2857 : AOI22_X1 port map( A1 => n80, A2 => regs(1782), B1 => n29, B2 => 
                           regs(758), ZN => n2098);
   U2858 : OAI211_X1 port map( C1 => n40, C2 => n2100, A => n2099, B => n2098, 
                           ZN => curr_proc_regs(758));
   U2859 : AOI22_X1 port map( A1 => n114, A2 => regs(247), B1 => n75, B2 => 
                           regs(2295), ZN => n2102);
   U2860 : AOI22_X1 port map( A1 => n49, A2 => regs(1271), B1 => n100, B2 => 
                           regs(1783), ZN => n2101);
   U2861 : OAI211_X1 port map( C1 => n15, C2 => n2103, A => n2102, B => n2101, 
                           ZN => curr_proc_regs(759));
   U2862 : INV_X1 port map( A => regs(1099), ZN => n2106);
   U2863 : AOI22_X1 port map( A1 => n114, A2 => regs(2123), B1 => n75, B2 => 
                           regs(1611), ZN => n2105);
   U2864 : AOI22_X1 port map( A1 => n49, A2 => regs(587), B1 => n30, B2 => 
                           regs(75), ZN => n2104);
   U2865 : OAI211_X1 port map( C1 => n6, C2 => n2106, A => n2105, B => n2104, 
                           ZN => curr_proc_regs(75));
   U2866 : AOI22_X1 port map( A1 => n114, A2 => regs(248), B1 => n76, B2 => 
                           regs(2296), ZN => n2108);
   U2867 : AOI22_X1 port map( A1 => n49, A2 => regs(1272), B1 => n99, B2 => 
                           regs(1784), ZN => n2107);
   U2868 : OAI211_X1 port map( C1 => n15, C2 => n2109, A => n2108, B => n2107, 
                           ZN => curr_proc_regs(760));
   U2869 : AOI22_X1 port map( A1 => n114, A2 => regs(249), B1 => n72, B2 => 
                           regs(2297), ZN => n2111);
   U2870 : AOI22_X1 port map( A1 => n49, A2 => regs(1273), B1 => n100, B2 => 
                           regs(1785), ZN => n2110);
   U2871 : OAI211_X1 port map( C1 => n15, C2 => n2112, A => n2111, B => n2110, 
                           ZN => curr_proc_regs(761));
   U2872 : AOI22_X1 port map( A1 => n114, A2 => regs(250), B1 => n76, B2 => 
                           regs(2298), ZN => n2114);
   U2873 : AOI22_X1 port map( A1 => n49, A2 => regs(1274), B1 => n100, B2 => 
                           regs(1786), ZN => n2113);
   U2874 : OAI211_X1 port map( C1 => n15, C2 => n2115, A => n2114, B => n2113, 
                           ZN => curr_proc_regs(762));
   U2875 : AOI22_X1 port map( A1 => n114, A2 => regs(251), B1 => n75, B2 => 
                           regs(2299), ZN => n2117);
   U2876 : AOI22_X1 port map( A1 => n80, A2 => regs(1787), B1 => n32, B2 => 
                           regs(763), ZN => n2116);
   U2877 : OAI211_X1 port map( C1 => n40, C2 => n2118, A => n2117, B => n2116, 
                           ZN => curr_proc_regs(763));
   U2878 : AOI22_X1 port map( A1 => n114, A2 => regs(252), B1 => n76, B2 => 
                           regs(2300), ZN => n2120);
   U2879 : AOI22_X1 port map( A1 => n80, A2 => regs(1788), B1 => n35, B2 => 
                           regs(764), ZN => n2119);
   U2880 : OAI211_X1 port map( C1 => n40, C2 => n2121, A => n2120, B => n2119, 
                           ZN => curr_proc_regs(764));
   U2881 : AOI22_X1 port map( A1 => n114, A2 => regs(253), B1 => n69, B2 => 
                           regs(2301), ZN => n2123);
   U2882 : AOI22_X1 port map( A1 => n49, A2 => regs(1277), B1 => n100, B2 => 
                           regs(1789), ZN => n2122);
   U2883 : OAI211_X1 port map( C1 => n15, C2 => n2124, A => n2123, B => n2122, 
                           ZN => curr_proc_regs(765));
   U2884 : AOI22_X1 port map( A1 => n114, A2 => regs(254), B1 => n71, B2 => 
                           regs(2302), ZN => n2126);
   U2885 : AOI22_X1 port map( A1 => n49, A2 => regs(1278), B1 => n100, B2 => 
                           regs(1790), ZN => n2125);
   U2886 : OAI211_X1 port map( C1 => n12, C2 => n2127, A => n2126, B => n2125, 
                           ZN => curr_proc_regs(766));
   U2887 : AOI22_X1 port map( A1 => n114, A2 => regs(255), B1 => n75, B2 => 
                           regs(2303), ZN => n2130);
   U2888 : AOI22_X1 port map( A1 => n80, A2 => regs(1791), B1 => n21, B2 => 
                           regs(767), ZN => n2129);
   U2889 : OAI211_X1 port map( C1 => n2201, C2 => n2131, A => n2130, B => n2129
                           , ZN => curr_proc_regs(767));
   U2890 : AOI22_X1 port map( A1 => n114, A2 => regs(2124), B1 => n76, B2 => 
                           regs(1612), ZN => n2133);
   U2891 : AOI22_X1 port map( A1 => n49, A2 => regs(588), B1 => n39, B2 => 
                           regs(76), ZN => n2132);
   U2892 : OAI211_X1 port map( C1 => n6, C2 => n2134, A => n2133, B => n2132, 
                           ZN => curr_proc_regs(76));
   U2893 : INV_X1 port map( A => regs(589), ZN => n2137);
   U2894 : AOI22_X1 port map( A1 => n114, A2 => regs(2125), B1 => n68, B2 => 
                           regs(1613), ZN => n2136);
   U2895 : AOI22_X1 port map( A1 => n80, A2 => regs(1101), B1 => n33, B2 => 
                           regs(77), ZN => n2135);
   U2896 : OAI211_X1 port map( C1 => n2201, C2 => n2137, A => n2136, B => n2135
                           , ZN => curr_proc_regs(77));
   U2897 : AOI22_X1 port map( A1 => n110, A2 => regs(2126), B1 => n75, B2 => 
                           regs(1614), ZN => n2139);
   U2898 : AOI22_X1 port map( A1 => n49, A2 => regs(590), B1 => n19, B2 => 
                           regs(78), ZN => n2138);
   U2899 : OAI211_X1 port map( C1 => n103, C2 => n2140, A => n2139, B => n2138,
                           ZN => curr_proc_regs(78));
   U2900 : AOI22_X1 port map( A1 => n106, A2 => regs(2127), B1 => n66, B2 => 
                           regs(1615), ZN => n2142);
   U2901 : AOI22_X1 port map( A1 => n49, A2 => regs(591), B1 => n29, B2 => 
                           regs(79), ZN => n2141);
   U2902 : OAI211_X1 port map( C1 => n78, C2 => n2143, A => n2142, B => n2141, 
                           ZN => curr_proc_regs(79));
   U2903 : AOI22_X1 port map( A1 => n107, A2 => regs(2055), B1 => n75, B2 => 
                           regs(1543), ZN => n2145);
   U2904 : AOI22_X1 port map( A1 => n49, A2 => regs(519), B1 => n4, B2 => 
                           regs(7), ZN => n2144);
   U2905 : OAI211_X1 port map( C1 => n103, C2 => n2146, A => n2145, B => n2144,
                           ZN => curr_proc_regs(7));
   U2906 : AOI22_X1 port map( A1 => n108, A2 => regs(2128), B1 => n76, B2 => 
                           regs(1616), ZN => n2148);
   U2907 : AOI22_X1 port map( A1 => n50, A2 => regs(592), B1 => n2, B2 => 
                           regs(80), ZN => n2147);
   U2908 : OAI211_X1 port map( C1 => n78, C2 => n2149, A => n2148, B => n2147, 
                           ZN => curr_proc_regs(80));
   U2909 : AOI22_X1 port map( A1 => n116, A2 => regs(2129), B1 => n75, B2 => 
                           regs(1617), ZN => n2151);
   U2910 : AOI22_X1 port map( A1 => n48, A2 => regs(593), B1 => n22, B2 => 
                           regs(81), ZN => n2150);
   U2911 : OAI211_X1 port map( C1 => n103, C2 => n2152, A => n2151, B => n2150,
                           ZN => curr_proc_regs(81));
   U2912 : INV_X1 port map( A => regs(1106), ZN => n2155);
   U2913 : AOI22_X1 port map( A1 => n118, A2 => regs(2130), B1 => n76, B2 => 
                           regs(1618), ZN => n2154);
   U2914 : AOI22_X1 port map( A1 => n48, A2 => regs(594), B1 => n17, B2 => 
                           regs(82), ZN => n2153);
   U2915 : OAI211_X1 port map( C1 => n103, C2 => n2155, A => n2154, B => n2153,
                           ZN => curr_proc_regs(82));
   U2916 : INV_X1 port map( A => regs(1107), ZN => n2158);
   U2917 : AOI22_X1 port map( A1 => n119, A2 => regs(2131), B1 => n5, B2 => 
                           regs(1619), ZN => n2157);
   U2918 : AOI22_X1 port map( A1 => n48, A2 => regs(595), B1 => n2, B2 => 
                           regs(83), ZN => n2156);
   U2919 : OAI211_X1 port map( C1 => n103, C2 => n2158, A => n2157, B => n2156,
                           ZN => curr_proc_regs(83));
   U2920 : INV_X1 port map( A => regs(1108), ZN => n2161);
   U2921 : AOI22_X1 port map( A1 => n121, A2 => regs(2132), B1 => n76, B2 => 
                           regs(1620), ZN => n2160);
   U2922 : AOI22_X1 port map( A1 => n48, A2 => regs(596), B1 => n32, B2 => 
                           regs(84), ZN => n2159);
   U2923 : OAI211_X1 port map( C1 => n103, C2 => n2161, A => n2160, B => n2159,
                           ZN => curr_proc_regs(84));
   U2924 : INV_X1 port map( A => regs(597), ZN => n2164);
   U2925 : AOI22_X1 port map( A1 => n123, A2 => regs(2133), B1 => n74, B2 => 
                           regs(1621), ZN => n2163);
   U2926 : AOI22_X1 port map( A1 => n80, A2 => regs(1109), B1 => n20, B2 => 
                           regs(85), ZN => n2162);
   U2927 : OAI211_X1 port map( C1 => n2201, C2 => n2164, A => n2163, B => n2162
                           , ZN => curr_proc_regs(85));
   U2928 : AOI22_X1 port map( A1 => n104, A2 => regs(2134), B1 => n75, B2 => 
                           regs(1622), ZN => n2166);
   U2929 : AOI22_X1 port map( A1 => n48, A2 => regs(598), B1 => n17, B2 => 
                           regs(86), ZN => n2165);
   U2930 : OAI211_X1 port map( C1 => n78, C2 => n2167, A => n2166, B => n2165, 
                           ZN => curr_proc_regs(86));
   U2931 : AOI22_X1 port map( A1 => n7, A2 => regs(2135), B1 => n76, B2 => 
                           regs(1623), ZN => n2169);
   U2932 : AOI22_X1 port map( A1 => n48, A2 => regs(599), B1 => n18, B2 => 
                           regs(87), ZN => n2168);
   U2933 : OAI211_X1 port map( C1 => n103, C2 => n2170, A => n2169, B => n2168,
                           ZN => curr_proc_regs(87));
   U2934 : AOI22_X1 port map( A1 => n7, A2 => regs(2136), B1 => n71, B2 => 
                           regs(1624), ZN => n2172);
   U2935 : AOI22_X1 port map( A1 => n48, A2 => regs(600), B1 => n19, B2 => 
                           regs(88), ZN => n2171);
   U2936 : OAI211_X1 port map( C1 => n103, C2 => n2173, A => n2172, B => n2171,
                           ZN => curr_proc_regs(88));
   U2937 : INV_X1 port map( A => regs(1113), ZN => n2176);
   U2938 : AOI22_X1 port map( A1 => n129, A2 => regs(2137), B1 => n5, B2 => 
                           regs(1625), ZN => n2175);
   U2939 : AOI22_X1 port map( A1 => n48, A2 => regs(601), B1 => n23, B2 => 
                           regs(89), ZN => n2174);
   U2940 : OAI211_X1 port map( C1 => n78, C2 => n2176, A => n2175, B => n2174, 
                           ZN => curr_proc_regs(89));
   U2941 : AOI22_X1 port map( A1 => n111, A2 => regs(2056), B1 => n72, B2 => 
                           regs(1544), ZN => n2178);
   U2942 : AOI22_X1 port map( A1 => n48, A2 => regs(520), B1 => n36, B2 => 
                           regs(8), ZN => n2177);
   U2943 : OAI211_X1 port map( C1 => n103, C2 => n2179, A => n2178, B => n2177,
                           ZN => curr_proc_regs(8));
   U2944 : INV_X1 port map( A => regs(602), ZN => n2182);
   U2945 : AOI22_X1 port map( A1 => n110, A2 => regs(2138), B1 => n68, B2 => 
                           regs(1626), ZN => n2181);
   U2946 : AOI22_X1 port map( A1 => n80, A2 => regs(1114), B1 => n21, B2 => 
                           regs(90), ZN => n2180);
   U2947 : OAI211_X1 port map( C1 => n2201, C2 => n2182, A => n2181, B => n2180
                           , ZN => curr_proc_regs(90));
   U2948 : INV_X1 port map( A => regs(603), ZN => n2185);
   U2949 : AOI22_X1 port map( A1 => n106, A2 => regs(2139), B1 => n68, B2 => 
                           regs(1627), ZN => n2184);
   U2950 : AOI22_X1 port map( A1 => n82, A2 => regs(1115), B1 => n31, B2 => 
                           regs(91), ZN => n2183);
   U2951 : OAI211_X1 port map( C1 => n2201, C2 => n2185, A => n2184, B => n2183
                           , ZN => curr_proc_regs(91));
   U2952 : AOI22_X1 port map( A1 => n107, A2 => regs(2140), B1 => n70, B2 => 
                           regs(1628), ZN => n2187);
   U2953 : AOI22_X1 port map( A1 => n48, A2 => regs(604), B1 => n19, B2 => 
                           regs(92), ZN => n2186);
   U2954 : OAI211_X1 port map( C1 => n103, C2 => n2188, A => n2187, B => n2186,
                           ZN => curr_proc_regs(92));
   U2955 : INV_X1 port map( A => regs(1117), ZN => n2191);
   U2956 : AOI22_X1 port map( A1 => n108, A2 => regs(2141), B1 => n75, B2 => 
                           regs(1629), ZN => n2190);
   U2957 : AOI22_X1 port map( A1 => n48, A2 => regs(605), B1 => n27, B2 => 
                           regs(93), ZN => n2189);
   U2958 : OAI211_X1 port map( C1 => n78, C2 => n2191, A => n2190, B => n2189, 
                           ZN => curr_proc_regs(93));
   U2959 : INV_X1 port map( A => regs(1118), ZN => n2194);
   U2960 : AOI22_X1 port map( A1 => n124, A2 => regs(2142), B1 => n76, B2 => 
                           regs(1630), ZN => n2193);
   U2961 : AOI22_X1 port map( A1 => n49, A2 => regs(606), B1 => n26, B2 => 
                           regs(94), ZN => n2192);
   U2962 : OAI211_X1 port map( C1 => n103, C2 => n2194, A => n2193, B => n2192,
                           ZN => curr_proc_regs(94));
   U2963 : AOI22_X1 port map( A1 => n116, A2 => regs(2143), B1 => n74, B2 => 
                           regs(1631), ZN => n2196);
   U2964 : AOI22_X1 port map( A1 => n47, A2 => regs(607), B1 => n25, B2 => 
                           regs(95), ZN => n2195);
   U2965 : OAI211_X1 port map( C1 => n78, C2 => n2197, A => n2196, B => n2195, 
                           ZN => curr_proc_regs(95));
   U2966 : INV_X1 port map( A => regs(608), ZN => n2200);
   U2967 : AOI22_X1 port map( A1 => n118, A2 => regs(2144), B1 => n65, B2 => 
                           regs(1632), ZN => n2199);
   U2968 : AOI22_X1 port map( A1 => n96, A2 => regs(1120), B1 => n24, B2 => 
                           regs(96), ZN => n2198);
   U2969 : OAI211_X1 port map( C1 => n2201, C2 => n2200, A => n2199, B => n2198
                           , ZN => curr_proc_regs(96));
   U2970 : INV_X1 port map( A => regs(1121), ZN => n2204);
   U2971 : AOI22_X1 port map( A1 => n119, A2 => regs(2145), B1 => n69, B2 => 
                           regs(1633), ZN => n2203);
   U2972 : AOI22_X1 port map( A1 => n47, A2 => regs(609), B1 => n24, B2 => 
                           regs(97), ZN => n2202);
   U2973 : OAI211_X1 port map( C1 => n103, C2 => n2204, A => n2203, B => n2202,
                           ZN => curr_proc_regs(97));
   U2974 : INV_X1 port map( A => regs(1122), ZN => n2207);
   U2975 : AOI22_X1 port map( A1 => n106, A2 => regs(2146), B1 => n67, B2 => 
                           regs(1634), ZN => n2206);
   U2976 : AOI22_X1 port map( A1 => n47, A2 => regs(610), B1 => n21, B2 => 
                           regs(98), ZN => n2205);
   U2977 : OAI211_X1 port map( C1 => n78, C2 => n2207, A => n2206, B => n2205, 
                           ZN => curr_proc_regs(98));
   U2978 : AOI22_X1 port map( A1 => n104, A2 => regs(2147), B1 => n68, B2 => 
                           regs(1635), ZN => n2209);
   U2979 : AOI22_X1 port map( A1 => n8, A2 => regs(611), B1 => n22, B2 => 
                           regs(99), ZN => n2208);
   U2980 : OAI211_X1 port map( C1 => n103, C2 => n2210, A => n2209, B => n2208,
                           ZN => curr_proc_regs(99));
   U2981 : INV_X1 port map( A => regs(1033), ZN => n2214);
   U2982 : AOI22_X1 port map( A1 => n126, A2 => regs(2057), B1 => n66, B2 => 
                           regs(1545), ZN => n2213);
   U2983 : AOI22_X1 port map( A1 => n55, A2 => regs(521), B1 => n23, B2 => 
                           regs(9), ZN => n2212);
   U2984 : OAI211_X1 port map( C1 => n78, C2 => n2214, A => n2213, B => n2212, 
                           ZN => curr_proc_regs(9));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32.all;

entity mux_N32_M5_1 is

   port( S : in std_logic_vector (4 downto 0);  Q : in std_logic_vector (1023 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end mux_N32_M5_1;

architecture SYN_behav of mux_N32_M5_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705 : std_logic;

begin
   
   U2 : AOI22_X1 port map( A1 => n255, A2 => Q(501), B1 => n254, B2 => Q(565), 
                           ZN => n1);
   U3 : AOI22_X1 port map( A1 => n257, A2 => Q(661), B1 => n256, B2 => Q(469), 
                           ZN => n2);
   U4 : AOI22_X1 port map( A1 => n259, A2 => Q(373), B1 => n258, B2 => Q(309), 
                           ZN => n3);
   U5 : AOI22_X1 port map( A1 => n261, A2 => Q(405), B1 => n260, B2 => Q(277), 
                           ZN => n4);
   U6 : NAND4_X1 port map( A1 => n1, A2 => n2, A3 => n3, A4 => n4, ZN => n5);
   U7 : AOI22_X1 port map( A1 => n263, A2 => Q(341), B1 => n262, B2 => Q(437), 
                           ZN => n6);
   U8 : AOI22_X1 port map( A1 => n265, A2 => Q(245), B1 => n264, B2 => Q(149), 
                           ZN => n7);
   U9 : AOI22_X1 port map( A1 => n267, A2 => Q(85), B1 => n266, B2 => Q(181), 
                           ZN => n8);
   U10 : AOI22_X1 port map( A1 => n269, A2 => Q(213), B1 => n268, B2 => Q(53), 
                           ZN => n9);
   U11 : NAND4_X1 port map( A1 => n6, A2 => n7, A3 => n8, A4 => n9, ZN => n10);
   U12 : AOI22_X1 port map( A1 => n240, A2 => Q(1013), B1 => n239, B2 => Q(949)
                           , ZN => n11);
   U13 : AOI22_X1 port map( A1 => n242, A2 => Q(981), B1 => n241, B2 => Q(917),
                           ZN => n12);
   U14 : AOI222_X1 port map( A1 => n244, A2 => Q(821), B1 => n245, B2 => Q(117)
                           , C1 => n243, C2 => Q(757), ZN => n13);
   U15 : NAND3_X1 port map( A1 => n11, A2 => n12, A3 => n13, ZN => n14);
   U16 : AOI22_X1 port map( A1 => n247, A2 => Q(853), B1 => n246, B2 => Q(725),
                           ZN => n15);
   U17 : AOI22_X1 port map( A1 => n249, A2 => Q(789), B1 => n248, B2 => Q(885),
                           ZN => n16);
   U18 : NAND4_X1 port map( A1 => n457, A2 => n458, A3 => n15, A4 => n16, ZN =>
                           n17);
   U19 : OR4_X1 port map( A1 => n5, A2 => n10, A3 => n14, A4 => n17, ZN => 
                           Y(21));
   U20 : AOI22_X1 port map( A1 => n255, A2 => Q(500), B1 => n254, B2 => Q(564),
                           ZN => n18);
   U21 : AOI22_X1 port map( A1 => n257, A2 => Q(660), B1 => n256, B2 => Q(468),
                           ZN => n19);
   U22 : AOI22_X1 port map( A1 => n259, A2 => Q(372), B1 => n258, B2 => Q(308),
                           ZN => n20);
   U23 : AOI22_X1 port map( A1 => n261, A2 => Q(404), B1 => n260, B2 => Q(276),
                           ZN => n21);
   U24 : NAND4_X1 port map( A1 => n18, A2 => n19, A3 => n20, A4 => n21, ZN => 
                           n22);
   U25 : AOI22_X1 port map( A1 => n263, A2 => Q(340), B1 => n262, B2 => Q(436),
                           ZN => n23);
   U26 : AOI22_X1 port map( A1 => n265, A2 => Q(244), B1 => n264, B2 => Q(148),
                           ZN => n24);
   U27 : AOI22_X1 port map( A1 => n267, A2 => Q(84), B1 => n266, B2 => Q(180), 
                           ZN => n25);
   U28 : AOI22_X1 port map( A1 => n269, A2 => Q(212), B1 => n268, B2 => Q(52), 
                           ZN => n26);
   U29 : NAND4_X1 port map( A1 => n23, A2 => n24, A3 => n25, A4 => n26, ZN => 
                           n27);
   U30 : AOI22_X1 port map( A1 => n240, A2 => Q(1012), B1 => n239, B2 => Q(948)
                           , ZN => n28);
   U31 : AOI22_X1 port map( A1 => n242, A2 => Q(980), B1 => n241, B2 => Q(916),
                           ZN => n29);
   U32 : AOI222_X1 port map( A1 => n244, A2 => Q(820), B1 => n245, B2 => Q(116)
                           , C1 => n243, C2 => Q(756), ZN => n30);
   U33 : NAND3_X1 port map( A1 => n28, A2 => n29, A3 => n30, ZN => n31);
   U34 : AOI22_X1 port map( A1 => n247, A2 => Q(852), B1 => n246, B2 => Q(724),
                           ZN => n32);
   U35 : AOI22_X1 port map( A1 => n249, A2 => Q(788), B1 => n248, B2 => Q(884),
                           ZN => n33);
   U36 : NAND4_X1 port map( A1 => n455, A2 => n456, A3 => n32, A4 => n33, ZN =>
                           n34);
   U37 : OR4_X1 port map( A1 => n22, A2 => n27, A3 => n31, A4 => n34, ZN => 
                           Y(20));
   U38 : AOI22_X1 port map( A1 => n255, A2 => Q(493), B1 => n254, B2 => Q(557),
                           ZN => n35);
   U39 : AOI22_X1 port map( A1 => n257, A2 => Q(653), B1 => n256, B2 => Q(461),
                           ZN => n36);
   U40 : AOI22_X1 port map( A1 => n259, A2 => Q(365), B1 => n258, B2 => Q(301),
                           ZN => n37);
   U41 : AOI22_X1 port map( A1 => n261, A2 => Q(397), B1 => n260, B2 => Q(269),
                           ZN => n38);
   U42 : NAND4_X1 port map( A1 => n35, A2 => n36, A3 => n37, A4 => n38, ZN => 
                           n39);
   U43 : AOI22_X1 port map( A1 => n263, A2 => Q(333), B1 => n262, B2 => Q(429),
                           ZN => n40);
   U44 : AOI22_X1 port map( A1 => n265, A2 => Q(237), B1 => n264, B2 => Q(141),
                           ZN => n41);
   U45 : AOI22_X1 port map( A1 => n267, A2 => Q(77), B1 => n266, B2 => Q(173), 
                           ZN => n42);
   U46 : AOI22_X1 port map( A1 => n269, A2 => Q(205), B1 => n268, B2 => Q(45), 
                           ZN => n43);
   U47 : NAND4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n44);
   U48 : AOI22_X1 port map( A1 => n240, A2 => Q(1005), B1 => n239, B2 => Q(941)
                           , ZN => n45);
   U49 : AOI22_X1 port map( A1 => n242, A2 => Q(973), B1 => n241, B2 => Q(909),
                           ZN => n46);
   U50 : AOI222_X1 port map( A1 => n244, A2 => Q(813), B1 => n245, B2 => Q(109)
                           , C1 => n243, C2 => Q(749), ZN => n47);
   U51 : NAND3_X1 port map( A1 => n45, A2 => n46, A3 => n47, ZN => n48);
   U52 : AOI22_X1 port map( A1 => n247, A2 => Q(845), B1 => n246, B2 => Q(717),
                           ZN => n49);
   U53 : AOI22_X1 port map( A1 => n249, A2 => Q(781), B1 => n248, B2 => Q(877),
                           ZN => n50);
   U54 : NAND4_X1 port map( A1 => n331, A2 => n332, A3 => n49, A4 => n50, ZN =>
                           n51);
   U55 : OR4_X1 port map( A1 => n39, A2 => n44, A3 => n48, A4 => n51, ZN => 
                           Y(13));
   U56 : AOI22_X1 port map( A1 => n255, A2 => Q(491), B1 => n254, B2 => Q(555),
                           ZN => n52);
   U57 : AOI22_X1 port map( A1 => n257, A2 => Q(651), B1 => n256, B2 => Q(459),
                           ZN => n53);
   U58 : AOI22_X1 port map( A1 => n259, A2 => Q(363), B1 => n258, B2 => Q(299),
                           ZN => n54);
   U59 : AOI22_X1 port map( A1 => n261, A2 => Q(395), B1 => n260, B2 => Q(267),
                           ZN => n55);
   U60 : NAND4_X1 port map( A1 => n52, A2 => n53, A3 => n54, A4 => n55, ZN => 
                           n56);
   U61 : AOI22_X1 port map( A1 => n263, A2 => Q(331), B1 => n262, B2 => Q(427),
                           ZN => n57);
   U62 : AOI22_X1 port map( A1 => n265, A2 => Q(235), B1 => n264, B2 => Q(139),
                           ZN => n58);
   U63 : AOI22_X1 port map( A1 => n267, A2 => Q(75), B1 => n266, B2 => Q(171), 
                           ZN => n59);
   U64 : AOI22_X1 port map( A1 => n269, A2 => Q(203), B1 => n268, B2 => Q(43), 
                           ZN => n60);
   U65 : NAND4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           n61);
   U66 : AOI22_X1 port map( A1 => n240, A2 => Q(1003), B1 => n239, B2 => Q(939)
                           , ZN => n62);
   U67 : AOI22_X1 port map( A1 => n242, A2 => Q(971), B1 => n241, B2 => Q(907),
                           ZN => n63);
   U68 : AOI222_X1 port map( A1 => n244, A2 => Q(811), B1 => n245, B2 => Q(107)
                           , C1 => n243, C2 => Q(747), ZN => n64);
   U69 : NAND3_X1 port map( A1 => n62, A2 => n63, A3 => n64, ZN => n65);
   U70 : AOI22_X1 port map( A1 => n247, A2 => Q(843), B1 => n246, B2 => Q(715),
                           ZN => n66);
   U71 : AOI22_X1 port map( A1 => n249, A2 => Q(779), B1 => n248, B2 => Q(875),
                           ZN => n67);
   U72 : NAND4_X1 port map( A1 => n309, A2 => n310, A3 => n66, A4 => n67, ZN =>
                           n68);
   U73 : OR4_X1 port map( A1 => n56, A2 => n61, A3 => n65, A4 => n68, ZN => 
                           Y(11));
   U74 : AOI22_X1 port map( A1 => n255, A2 => Q(489), B1 => n254, B2 => Q(553),
                           ZN => n69);
   U75 : AOI22_X1 port map( A1 => n257, A2 => Q(649), B1 => n256, B2 => Q(457),
                           ZN => n70);
   U76 : AOI22_X1 port map( A1 => n259, A2 => Q(361), B1 => n258, B2 => Q(297),
                           ZN => n71);
   U77 : AOI22_X1 port map( A1 => n261, A2 => Q(393), B1 => n260, B2 => Q(265),
                           ZN => n72);
   U78 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           n73);
   U79 : AOI22_X1 port map( A1 => n263, A2 => Q(329), B1 => n262, B2 => Q(425),
                           ZN => n74);
   U80 : AOI22_X1 port map( A1 => n265, A2 => Q(233), B1 => n264, B2 => Q(137),
                           ZN => n75);
   U81 : AOI22_X1 port map( A1 => n267, A2 => Q(73), B1 => n266, B2 => Q(169), 
                           ZN => n76);
   U82 : AOI22_X1 port map( A1 => n269, A2 => Q(201), B1 => n268, B2 => Q(41), 
                           ZN => n77);
   U83 : NAND4_X1 port map( A1 => n74, A2 => n75, A3 => n76, A4 => n77, ZN => 
                           n78);
   U84 : AOI22_X1 port map( A1 => n240, A2 => Q(1001), B1 => n239, B2 => Q(937)
                           , ZN => n79);
   U85 : AOI22_X1 port map( A1 => n242, A2 => Q(969), B1 => n241, B2 => Q(905),
                           ZN => n80);
   U86 : AOI222_X1 port map( A1 => n244, A2 => Q(809), B1 => n245, B2 => Q(105)
                           , C1 => n243, C2 => Q(745), ZN => n81);
   U87 : NAND3_X1 port map( A1 => n79, A2 => n80, A3 => n81, ZN => n82);
   U88 : AOI22_X1 port map( A1 => n247, A2 => Q(841), B1 => n246, B2 => Q(713),
                           ZN => n83);
   U89 : AOI22_X1 port map( A1 => n249, A2 => Q(777), B1 => n248, B2 => Q(873),
                           ZN => n84);
   U90 : NAND4_X1 port map( A1 => n688, A2 => n689, A3 => n83, A4 => n84, ZN =>
                           n85);
   U91 : OR4_X1 port map( A1 => n73, A2 => n78, A3 => n82, A4 => n85, ZN => 
                           Y(9));
   U92 : AOI22_X1 port map( A1 => n255, A2 => Q(488), B1 => n254, B2 => Q(552),
                           ZN => n86);
   U93 : AOI22_X1 port map( A1 => n257, A2 => Q(648), B1 => n256, B2 => Q(456),
                           ZN => n87);
   U94 : AOI22_X1 port map( A1 => n259, A2 => Q(360), B1 => n258, B2 => Q(296),
                           ZN => n88);
   U95 : AOI22_X1 port map( A1 => n261, A2 => Q(392), B1 => n260, B2 => Q(264),
                           ZN => n89);
   U96 : NAND4_X1 port map( A1 => n86, A2 => n87, A3 => n88, A4 => n89, ZN => 
                           n90);
   U97 : AOI22_X1 port map( A1 => n263, A2 => Q(328), B1 => n262, B2 => Q(424),
                           ZN => n91);
   U98 : AOI22_X1 port map( A1 => n265, A2 => Q(232), B1 => n264, B2 => Q(136),
                           ZN => n92);
   U99 : AOI22_X1 port map( A1 => n267, A2 => Q(72), B1 => n266, B2 => Q(168), 
                           ZN => n93);
   U100 : AOI22_X1 port map( A1 => n269, A2 => Q(200), B1 => n268, B2 => Q(40),
                           ZN => n94);
   U101 : NAND4_X1 port map( A1 => n91, A2 => n92, A3 => n93, A4 => n94, ZN => 
                           n95);
   U102 : AOI22_X1 port map( A1 => n240, A2 => Q(1000), B1 => n239, B2 => 
                           Q(936), ZN => n96);
   U103 : AOI22_X1 port map( A1 => n242, A2 => Q(968), B1 => n241, B2 => Q(904)
                           , ZN => n97);
   U104 : AOI222_X1 port map( A1 => n244, A2 => Q(808), B1 => n245, B2 => 
                           Q(104), C1 => n243, C2 => Q(744), ZN => n98);
   U105 : NAND3_X1 port map( A1 => n96, A2 => n97, A3 => n98, ZN => n99);
   U106 : AOI22_X1 port map( A1 => n247, A2 => Q(840), B1 => n246, B2 => Q(712)
                           , ZN => n100);
   U107 : AOI22_X1 port map( A1 => n249, A2 => Q(776), B1 => n248, B2 => Q(872)
                           , ZN => n101);
   U108 : NAND4_X1 port map( A1 => n671, A2 => n672, A3 => n100, A4 => n101, ZN
                           => n102);
   U109 : OR4_X1 port map( A1 => n90, A2 => n95, A3 => n99, A4 => n102, ZN => 
                           Y(8));
   U110 : AOI22_X1 port map( A1 => n255, A2 => Q(487), B1 => n254, B2 => Q(551)
                           , ZN => n103);
   U111 : AOI22_X1 port map( A1 => n257, A2 => Q(647), B1 => n256, B2 => Q(455)
                           , ZN => n104);
   U112 : AOI22_X1 port map( A1 => n259, A2 => Q(359), B1 => n258, B2 => Q(295)
                           , ZN => n105);
   U113 : AOI22_X1 port map( A1 => n261, A2 => Q(391), B1 => n260, B2 => Q(263)
                           , ZN => n106);
   U114 : NAND4_X1 port map( A1 => n103, A2 => n104, A3 => n105, A4 => n106, ZN
                           => n107);
   U115 : AOI22_X1 port map( A1 => n263, A2 => Q(327), B1 => n262, B2 => Q(423)
                           , ZN => n108);
   U116 : AOI22_X1 port map( A1 => n265, A2 => Q(231), B1 => n264, B2 => Q(135)
                           , ZN => n109);
   U117 : AOI22_X1 port map( A1 => n267, A2 => Q(71), B1 => n266, B2 => Q(167),
                           ZN => n110);
   U118 : AOI22_X1 port map( A1 => n269, A2 => Q(199), B1 => n268, B2 => Q(39),
                           ZN => n111);
   U119 : NAND4_X1 port map( A1 => n108, A2 => n109, A3 => n110, A4 => n111, ZN
                           => n112);
   U120 : AOI22_X1 port map( A1 => n240, A2 => Q(999), B1 => n239, B2 => Q(935)
                           , ZN => n113);
   U121 : AOI22_X1 port map( A1 => n242, A2 => Q(967), B1 => n241, B2 => Q(903)
                           , ZN => n114);
   U122 : AOI222_X1 port map( A1 => n244, A2 => Q(807), B1 => n245, B2 => 
                           Q(103), C1 => n243, C2 => Q(743), ZN => n115);
   U123 : NAND3_X1 port map( A1 => n113, A2 => n114, A3 => n115, ZN => n116);
   U124 : AOI22_X1 port map( A1 => n247, A2 => Q(839), B1 => n246, B2 => Q(711)
                           , ZN => n117);
   U125 : AOI22_X1 port map( A1 => n249, A2 => Q(775), B1 => n248, B2 => Q(871)
                           , ZN => n118);
   U126 : NAND4_X1 port map( A1 => n669, A2 => n670, A3 => n117, A4 => n118, ZN
                           => n119);
   U127 : OR4_X1 port map( A1 => n107, A2 => n112, A3 => n116, A4 => n119, ZN 
                           => Y(7));
   U128 : AOI22_X1 port map( A1 => n255, A2 => Q(486), B1 => n254, B2 => Q(550)
                           , ZN => n120);
   U129 : AOI22_X1 port map( A1 => n257, A2 => Q(646), B1 => n256, B2 => Q(454)
                           , ZN => n121);
   U130 : AOI22_X1 port map( A1 => n259, A2 => Q(358), B1 => n258, B2 => Q(294)
                           , ZN => n122);
   U131 : AOI22_X1 port map( A1 => n261, A2 => Q(390), B1 => n260, B2 => Q(262)
                           , ZN => n123);
   U132 : NAND4_X1 port map( A1 => n120, A2 => n121, A3 => n122, A4 => n123, ZN
                           => n124);
   U133 : AOI22_X1 port map( A1 => n263, A2 => Q(326), B1 => n262, B2 => Q(422)
                           , ZN => n125);
   U134 : AOI22_X1 port map( A1 => n265, A2 => Q(230), B1 => n264, B2 => Q(134)
                           , ZN => n126);
   U135 : AOI22_X1 port map( A1 => n267, A2 => Q(70), B1 => n266, B2 => Q(166),
                           ZN => n127);
   U136 : AOI22_X1 port map( A1 => n269, A2 => Q(198), B1 => n268, B2 => Q(38),
                           ZN => n128);
   U137 : NAND4_X1 port map( A1 => n125, A2 => n126, A3 => n127, A4 => n128, ZN
                           => n129);
   U138 : AOI22_X1 port map( A1 => n240, A2 => Q(998), B1 => n239, B2 => Q(934)
                           , ZN => n130);
   U139 : AOI22_X1 port map( A1 => n242, A2 => Q(966), B1 => n241, B2 => Q(902)
                           , ZN => n131);
   U140 : AOI222_X1 port map( A1 => n244, A2 => Q(806), B1 => n245, B2 => 
                           Q(102), C1 => n243, C2 => Q(742), ZN => n132);
   U141 : NAND3_X1 port map( A1 => n130, A2 => n131, A3 => n132, ZN => n133);
   U142 : AOI22_X1 port map( A1 => n247, A2 => Q(838), B1 => n246, B2 => Q(710)
                           , ZN => n134);
   U143 : AOI22_X1 port map( A1 => n249, A2 => Q(774), B1 => n248, B2 => Q(870)
                           , ZN => n135);
   U144 : NAND4_X1 port map( A1 => n667, A2 => n668, A3 => n134, A4 => n135, ZN
                           => n136);
   U145 : OR4_X1 port map( A1 => n124, A2 => n129, A3 => n133, A4 => n136, ZN 
                           => Y(6));
   U146 : AOI22_X1 port map( A1 => n255, A2 => Q(485), B1 => n254, B2 => Q(549)
                           , ZN => n137);
   U147 : AOI22_X1 port map( A1 => n257, A2 => Q(645), B1 => n256, B2 => Q(453)
                           , ZN => n138);
   U148 : AOI22_X1 port map( A1 => n259, A2 => Q(357), B1 => n258, B2 => Q(293)
                           , ZN => n139);
   U149 : AOI22_X1 port map( A1 => n261, A2 => Q(389), B1 => n260, B2 => Q(261)
                           , ZN => n140);
   U150 : NAND4_X1 port map( A1 => n137, A2 => n138, A3 => n139, A4 => n140, ZN
                           => n141);
   U151 : AOI22_X1 port map( A1 => n263, A2 => Q(325), B1 => n262, B2 => Q(421)
                           , ZN => n142);
   U152 : AOI22_X1 port map( A1 => n265, A2 => Q(229), B1 => n264, B2 => Q(133)
                           , ZN => n143);
   U153 : AOI22_X1 port map( A1 => n267, A2 => Q(69), B1 => n266, B2 => Q(165),
                           ZN => n144);
   U154 : AOI22_X1 port map( A1 => n269, A2 => Q(197), B1 => n268, B2 => Q(37),
                           ZN => n145);
   U155 : NAND4_X1 port map( A1 => n142, A2 => n143, A3 => n144, A4 => n145, ZN
                           => n146);
   U156 : AOI22_X1 port map( A1 => n240, A2 => Q(997), B1 => n239, B2 => Q(933)
                           , ZN => n147);
   U157 : AOI22_X1 port map( A1 => n242, A2 => Q(965), B1 => n241, B2 => Q(901)
                           , ZN => n148);
   U158 : AOI222_X1 port map( A1 => n244, A2 => Q(805), B1 => n245, B2 => 
                           Q(101), C1 => n243, C2 => Q(741), ZN => n149);
   U159 : NAND3_X1 port map( A1 => n147, A2 => n148, A3 => n149, ZN => n150);
   U160 : AOI22_X1 port map( A1 => n247, A2 => Q(837), B1 => n246, B2 => Q(709)
                           , ZN => n151);
   U161 : AOI22_X1 port map( A1 => n249, A2 => Q(773), B1 => n248, B2 => Q(869)
                           , ZN => n152);
   U162 : NAND4_X1 port map( A1 => n665, A2 => n666, A3 => n151, A4 => n152, ZN
                           => n153);
   U163 : OR4_X1 port map( A1 => n141, A2 => n146, A3 => n150, A4 => n153, ZN 
                           => Y(5));
   U164 : AOI22_X1 port map( A1 => n255, A2 => Q(484), B1 => n254, B2 => Q(548)
                           , ZN => n154);
   U165 : AOI22_X1 port map( A1 => n257, A2 => Q(644), B1 => n256, B2 => Q(452)
                           , ZN => n155);
   U166 : AOI22_X1 port map( A1 => n259, A2 => Q(356), B1 => n258, B2 => Q(292)
                           , ZN => n156);
   U167 : AOI22_X1 port map( A1 => n261, A2 => Q(388), B1 => n260, B2 => Q(260)
                           , ZN => n157);
   U168 : NAND4_X1 port map( A1 => n154, A2 => n155, A3 => n156, A4 => n157, ZN
                           => n158);
   U169 : AOI22_X1 port map( A1 => n263, A2 => Q(324), B1 => n262, B2 => Q(420)
                           , ZN => n159);
   U170 : AOI22_X1 port map( A1 => n265, A2 => Q(228), B1 => n264, B2 => Q(132)
                           , ZN => n160);
   U171 : AOI22_X1 port map( A1 => n267, A2 => Q(68), B1 => n266, B2 => Q(164),
                           ZN => n161);
   U172 : AOI22_X1 port map( A1 => n269, A2 => Q(196), B1 => n268, B2 => Q(36),
                           ZN => n162);
   U173 : NAND4_X1 port map( A1 => n159, A2 => n160, A3 => n161, A4 => n162, ZN
                           => n163);
   U174 : AOI22_X1 port map( A1 => n240, A2 => Q(996), B1 => n239, B2 => Q(932)
                           , ZN => n164);
   U175 : AOI22_X1 port map( A1 => n242, A2 => Q(964), B1 => n241, B2 => Q(900)
                           , ZN => n165);
   U176 : AOI222_X1 port map( A1 => n244, A2 => Q(804), B1 => n245, B2 => 
                           Q(100), C1 => n243, C2 => Q(740), ZN => n166);
   U177 : NAND3_X1 port map( A1 => n164, A2 => n165, A3 => n166, ZN => n167);
   U178 : AOI22_X1 port map( A1 => n247, A2 => Q(836), B1 => n246, B2 => Q(708)
                           , ZN => n168);
   U179 : AOI22_X1 port map( A1 => n249, A2 => Q(772), B1 => n248, B2 => Q(868)
                           , ZN => n169);
   U180 : NAND4_X1 port map( A1 => n663, A2 => n664, A3 => n168, A4 => n169, ZN
                           => n170);
   U181 : OR4_X1 port map( A1 => n158, A2 => n163, A3 => n167, A4 => n170, ZN 
                           => Y(4));
   U182 : AOI22_X1 port map( A1 => n255, A2 => Q(483), B1 => n254, B2 => Q(547)
                           , ZN => n171);
   U183 : AOI22_X1 port map( A1 => n257, A2 => Q(643), B1 => n256, B2 => Q(451)
                           , ZN => n172);
   U184 : AOI22_X1 port map( A1 => n259, A2 => Q(355), B1 => n258, B2 => Q(291)
                           , ZN => n173);
   U185 : AOI22_X1 port map( A1 => n261, A2 => Q(387), B1 => n260, B2 => Q(259)
                           , ZN => n174);
   U186 : NAND4_X1 port map( A1 => n171, A2 => n172, A3 => n173, A4 => n174, ZN
                           => n175);
   U187 : AOI22_X1 port map( A1 => n263, A2 => Q(323), B1 => n262, B2 => Q(419)
                           , ZN => n176);
   U188 : AOI22_X1 port map( A1 => n265, A2 => Q(227), B1 => n264, B2 => Q(131)
                           , ZN => n177);
   U189 : AOI22_X1 port map( A1 => n267, A2 => Q(67), B1 => n266, B2 => Q(163),
                           ZN => n178);
   U190 : AOI22_X1 port map( A1 => n269, A2 => Q(195), B1 => n268, B2 => Q(35),
                           ZN => n179);
   U191 : NAND4_X1 port map( A1 => n176, A2 => n177, A3 => n178, A4 => n179, ZN
                           => n180);
   U192 : AOI22_X1 port map( A1 => n240, A2 => Q(995), B1 => n239, B2 => Q(931)
                           , ZN => n181);
   U193 : AOI22_X1 port map( A1 => n242, A2 => Q(963), B1 => n241, B2 => Q(899)
                           , ZN => n182);
   U194 : AOI222_X1 port map( A1 => n244, A2 => Q(803), B1 => n245, B2 => Q(99)
                           , C1 => n243, C2 => Q(739), ZN => n183);
   U195 : NAND3_X1 port map( A1 => n181, A2 => n182, A3 => n183, ZN => n184);
   U196 : AOI22_X1 port map( A1 => n247, A2 => Q(835), B1 => n246, B2 => Q(707)
                           , ZN => n185);
   U197 : AOI22_X1 port map( A1 => n249, A2 => Q(771), B1 => n248, B2 => Q(867)
                           , ZN => n186);
   U198 : NAND4_X1 port map( A1 => n661, A2 => n662, A3 => n185, A4 => n186, ZN
                           => n187);
   U199 : OR4_X1 port map( A1 => n175, A2 => n180, A3 => n184, A4 => n187, ZN 
                           => Y(3));
   U200 : AOI22_X1 port map( A1 => n690, A2 => Q(545), B1 => n691, B2 => Q(481)
                           , ZN => n188);
   U201 : AOI22_X1 port map( A1 => n692, A2 => Q(449), B1 => n693, B2 => Q(641)
                           , ZN => n189);
   U202 : AOI22_X1 port map( A1 => n694, A2 => Q(289), B1 => n695, B2 => Q(353)
                           , ZN => n190);
   U203 : AOI22_X1 port map( A1 => n696, A2 => Q(257), B1 => n697, B2 => Q(385)
                           , ZN => n191);
   U204 : NAND4_X1 port map( A1 => n188, A2 => n189, A3 => n190, A4 => n191, ZN
                           => n192);
   U205 : AOI22_X1 port map( A1 => n698, A2 => Q(417), B1 => n699, B2 => Q(321)
                           , ZN => n193);
   U206 : AOI22_X1 port map( A1 => n700, A2 => Q(129), B1 => n701, B2 => Q(225)
                           , ZN => n194);
   U207 : AOI22_X1 port map( A1 => n702, A2 => Q(161), B1 => n703, B2 => Q(65),
                           ZN => n195);
   U208 : AOI22_X1 port map( A1 => n704, A2 => Q(33), B1 => n705, B2 => Q(193),
                           ZN => n196);
   U209 : NAND4_X1 port map( A1 => n193, A2 => n194, A3 => n195, A4 => n196, ZN
                           => n197);
   U210 : AOI22_X1 port map( A1 => n673, A2 => Q(929), B1 => n674, B2 => Q(993)
                           , ZN => n198);
   U211 : AOI22_X1 port map( A1 => n675, A2 => Q(897), B1 => n676, B2 => Q(961)
                           , ZN => n199);
   U212 : AOI222_X1 port map( A1 => n677, A2 => Q(737), B1 => n678, B2 => 
                           Q(801), C1 => n679, C2 => Q(97), ZN => n200);
   U213 : NAND3_X1 port map( A1 => n198, A2 => n199, A3 => n200, ZN => n201);
   U214 : AOI22_X1 port map( A1 => n680, A2 => Q(705), B1 => n681, B2 => Q(833)
                           , ZN => n202);
   U215 : AOI22_X1 port map( A1 => n682, A2 => Q(865), B1 => n683, B2 => Q(769)
                           , ZN => n203);
   U216 : NAND4_X1 port map( A1 => n453, A2 => n454, A3 => n202, A4 => n203, ZN
                           => n204);
   U217 : OR4_X1 port map( A1 => n192, A2 => n197, A3 => n201, A4 => n204, ZN 
                           => Y(1));
   U218 : AOI22_X1 port map( A1 => n255, A2 => Q(480), B1 => n254, B2 => Q(544)
                           , ZN => n205);
   U219 : AOI22_X1 port map( A1 => n257, A2 => Q(640), B1 => n256, B2 => Q(448)
                           , ZN => n206);
   U220 : AOI22_X1 port map( A1 => n259, A2 => Q(352), B1 => n258, B2 => Q(288)
                           , ZN => n207);
   U221 : AOI22_X1 port map( A1 => n261, A2 => Q(384), B1 => n260, B2 => Q(256)
                           , ZN => n208);
   U222 : NAND4_X1 port map( A1 => n205, A2 => n206, A3 => n207, A4 => n208, ZN
                           => n209);
   U223 : AOI22_X1 port map( A1 => n263, A2 => Q(320), B1 => n262, B2 => Q(416)
                           , ZN => n210);
   U224 : AOI22_X1 port map( A1 => n265, A2 => Q(224), B1 => n264, B2 => Q(128)
                           , ZN => n211);
   U225 : AOI22_X1 port map( A1 => n267, A2 => Q(64), B1 => n266, B2 => Q(160),
                           ZN => n212);
   U226 : AOI22_X1 port map( A1 => n269, A2 => Q(192), B1 => n268, B2 => Q(32),
                           ZN => n213);
   U227 : NAND4_X1 port map( A1 => n210, A2 => n211, A3 => n212, A4 => n213, ZN
                           => n214);
   U228 : AOI22_X1 port map( A1 => n240, A2 => Q(992), B1 => n239, B2 => Q(928)
                           , ZN => n215);
   U229 : AOI22_X1 port map( A1 => n242, A2 => Q(960), B1 => n241, B2 => Q(896)
                           , ZN => n216);
   U230 : AOI222_X1 port map( A1 => n244, A2 => Q(800), B1 => n245, B2 => Q(96)
                           , C1 => n243, C2 => Q(736), ZN => n217);
   U231 : NAND3_X1 port map( A1 => n215, A2 => n216, A3 => n217, ZN => n218);
   U232 : AOI22_X1 port map( A1 => n247, A2 => Q(832), B1 => n246, B2 => Q(704)
                           , ZN => n219);
   U233 : AOI22_X1 port map( A1 => n249, A2 => Q(768), B1 => n248, B2 => Q(864)
                           , ZN => n220);
   U234 : NAND4_X1 port map( A1 => n274, A2 => n275, A3 => n219, A4 => n220, ZN
                           => n221);
   U235 : OR4_X1 port map( A1 => n209, A2 => n214, A3 => n218, A4 => n221, ZN 
                           => Y(0));
   U236 : AOI22_X1 port map( A1 => n255, A2 => Q(511), B1 => n254, B2 => Q(575)
                           , ZN => n222);
   U237 : AOI22_X1 port map( A1 => n257, A2 => Q(671), B1 => n256, B2 => Q(479)
                           , ZN => n223);
   U238 : AOI22_X1 port map( A1 => n259, A2 => Q(383), B1 => n258, B2 => Q(319)
                           , ZN => n224);
   U239 : AOI22_X1 port map( A1 => n261, A2 => Q(415), B1 => n260, B2 => Q(287)
                           , ZN => n225);
   U240 : NAND4_X1 port map( A1 => n222, A2 => n223, A3 => n224, A4 => n225, ZN
                           => n226);
   U241 : AOI22_X1 port map( A1 => n263, A2 => Q(351), B1 => n262, B2 => Q(447)
                           , ZN => n227);
   U242 : AOI22_X1 port map( A1 => n265, A2 => Q(255), B1 => n264, B2 => Q(159)
                           , ZN => n228);
   U243 : AOI22_X1 port map( A1 => n267, A2 => Q(95), B1 => n266, B2 => Q(191),
                           ZN => n229);
   U244 : AOI22_X1 port map( A1 => n269, A2 => Q(223), B1 => n268, B2 => Q(63),
                           ZN => n230);
   U245 : NAND4_X1 port map( A1 => n227, A2 => n228, A3 => n229, A4 => n230, ZN
                           => n231);
   U246 : AOI22_X1 port map( A1 => n240, A2 => Q(1023), B1 => n239, B2 => 
                           Q(959), ZN => n232);
   U247 : AOI22_X1 port map( A1 => n242, A2 => Q(991), B1 => n241, B2 => Q(927)
                           , ZN => n233);
   U248 : AOI222_X1 port map( A1 => n244, A2 => Q(831), B1 => n245, B2 => 
                           Q(127), C1 => n243, C2 => Q(767), ZN => n234);
   U249 : NAND3_X1 port map( A1 => n232, A2 => n233, A3 => n234, ZN => n235);
   U250 : AOI22_X1 port map( A1 => n247, A2 => Q(863), B1 => n246, B2 => Q(735)
                           , ZN => n236);
   U251 : AOI22_X1 port map( A1 => n249, A2 => Q(799), B1 => n248, B2 => Q(895)
                           , ZN => n237);
   U252 : NAND4_X1 port map( A1 => n659, A2 => n660, A3 => n236, A4 => n237, ZN
                           => n238);
   U253 : OR4_X1 port map( A1 => n226, A2 => n231, A3 => n235, A4 => n238, ZN 
                           => Y(31));
   U254 : OR4_X1 port map( A1 => n658, A2 => n657, A3 => n656, A4 => n655, ZN 
                           => Y(30));
   U255 : OR4_X1 port map( A1 => n432, A2 => n431, A3 => n430, A4 => n429, ZN 
                           => Y(18));
   U256 : OR4_X1 port map( A1 => n452, A2 => n451, A3 => n450, A4 => n449, ZN 
                           => Y(19));
   U257 : OR4_X1 port map( A1 => n412, A2 => n411, A3 => n410, A4 => n409, ZN 
                           => Y(17));
   U258 : OR4_X1 port map( A1 => n598, A2 => n597, A3 => n596, A4 => n595, ZN 
                           => Y(28));
   U259 : OR4_X1 port map( A1 => n392, A2 => n391, A3 => n390, A4 => n389, ZN 
                           => Y(16));
   U260 : OR4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN 
                           => Y(12));
   U261 : OR4_X1 port map( A1 => n558, A2 => n557, A3 => n556, A4 => n555, ZN 
                           => Y(26));
   U262 : OR4_X1 port map( A1 => n372, A2 => n371, A3 => n370, A4 => n369, ZN 
                           => Y(15));
   U263 : OR4_X1 port map( A1 => n538, A2 => n537, A3 => n536, A4 => n535, ZN 
                           => Y(25));
   U264 : OR4_X1 port map( A1 => n308, A2 => n307, A3 => n306, A4 => n305, ZN 
                           => Y(10));
   U265 : OR4_X1 port map( A1 => n518, A2 => n517, A3 => n516, A4 => n515, ZN 
                           => Y(24));
   U266 : OR4_X1 port map( A1 => n352, A2 => n351, A3 => n350, A4 => n349, ZN 
                           => Y(14));
   U267 : OR4_X1 port map( A1 => n618, A2 => n617, A3 => n616, A4 => n615, ZN 
                           => Y(29));
   U268 : OR4_X1 port map( A1 => n498, A2 => n497, A3 => n496, A4 => n495, ZN 
                           => Y(23));
   U269 : OR4_X1 port map( A1 => n478, A2 => n477, A3 => n476, A4 => n475, ZN 
                           => Y(22));
   U270 : OR4_X1 port map( A1 => n638, A2 => n637, A3 => n636, A4 => n635, ZN 
                           => Y(2));
   U271 : OR4_X1 port map( A1 => n578, A2 => n577, A3 => n576, A4 => n575, ZN 
                           => Y(27));
   U272 : BUF_X1 port map( A => n704, Z => n268);
   U273 : BUF_X1 port map( A => n705, Z => n269);
   U274 : BUF_X1 port map( A => n702, Z => n266);
   U275 : BUF_X1 port map( A => n703, Z => n267);
   U276 : BUF_X1 port map( A => n700, Z => n264);
   U277 : BUF_X1 port map( A => n701, Z => n265);
   U278 : BUF_X1 port map( A => n698, Z => n262);
   U279 : BUF_X1 port map( A => n699, Z => n263);
   U280 : BUF_X1 port map( A => n696, Z => n260);
   U281 : BUF_X1 port map( A => n697, Z => n261);
   U282 : BUF_X1 port map( A => n694, Z => n258);
   U283 : BUF_X1 port map( A => n695, Z => n259);
   U284 : BUF_X1 port map( A => n692, Z => n256);
   U285 : BUF_X1 port map( A => n693, Z => n257);
   U286 : BUF_X1 port map( A => n690, Z => n254);
   U287 : BUF_X1 port map( A => n691, Z => n255);
   U288 : BUF_X1 port map( A => n686, Z => n252);
   U289 : BUF_X1 port map( A => n687, Z => n253);
   U290 : BUF_X1 port map( A => n684, Z => n250);
   U291 : BUF_X1 port map( A => n685, Z => n251);
   U292 : BUF_X1 port map( A => n682, Z => n248);
   U293 : BUF_X1 port map( A => n683, Z => n249);
   U294 : BUF_X1 port map( A => n680, Z => n246);
   U295 : BUF_X1 port map( A => n681, Z => n247);
   U296 : BUF_X1 port map( A => n679, Z => n245);
   U297 : BUF_X1 port map( A => n677, Z => n243);
   U298 : BUF_X1 port map( A => n678, Z => n244);
   U299 : BUF_X1 port map( A => n675, Z => n241);
   U300 : BUF_X1 port map( A => n676, Z => n242);
   U301 : BUF_X1 port map( A => n673, Z => n239);
   U302 : OR2_X1 port map( A1 => n270, A2 => S(1), ZN => n284);
   U303 : BUF_X1 port map( A => n674, Z => n240);
   U304 : NAND2_X1 port map( A1 => S(1), A2 => S(2), ZN => n286);
   U305 : NAND3_X1 port map( A1 => S(3), A2 => S(4), A3 => S(0), ZN => n273);
   U306 : NOR2_X1 port map( A1 => n286, A2 => n273, ZN => n674);
   U307 : INV_X1 port map( A => S(2), ZN => n270);
   U308 : NOR2_X1 port map( A1 => n273, A2 => n284, ZN => n673);
   U309 : INV_X1 port map( A => S(0), ZN => n271);
   U310 : NAND3_X1 port map( A1 => S(4), A2 => S(3), A3 => n271, ZN => n272);
   U311 : NOR2_X1 port map( A1 => n286, A2 => n272, ZN => n676);
   U312 : NOR2_X1 port map( A1 => n284, A2 => n272, ZN => n675);
   U313 : OR2_X1 port map( A1 => S(1), A2 => S(2), ZN => n287);
   U314 : NOR2_X1 port map( A1 => n273, A2 => n287, ZN => n678);
   U315 : INV_X1 port map( A => S(3), ZN => n281);
   U316 : NAND3_X1 port map( A1 => S(4), A2 => S(0), A3 => n281, ZN => n277);
   U317 : NOR2_X1 port map( A1 => n286, A2 => n277, ZN => n677);
   U318 : NAND2_X1 port map( A1 => S(1), A2 => n270, ZN => n283);
   U319 : INV_X1 port map( A => S(4), ZN => n276);
   U320 : NAND3_X1 port map( A1 => S(0), A2 => n281, A3 => n276, ZN => n288);
   U321 : NOR2_X1 port map( A1 => n283, A2 => n288, ZN => n679);
   U322 : NOR2_X1 port map( A1 => n283, A2 => n272, ZN => n681);
   U323 : NAND3_X1 port map( A1 => S(4), A2 => n281, A3 => n271, ZN => n278);
   U324 : NOR2_X1 port map( A1 => n286, A2 => n278, ZN => n680);
   U325 : NOR2_X1 port map( A1 => n272, A2 => n287, ZN => n683);
   U326 : NOR2_X1 port map( A1 => n283, A2 => n273, ZN => n682);
   U327 : NOR2_X1 port map( A1 => n284, A2 => n277, ZN => n685);
   U328 : NOR2_X1 port map( A1 => n283, A2 => n278, ZN => n684);
   U329 : AOI22_X1 port map( A1 => n251, A2 => Q(672), B1 => n250, B2 => Q(576)
                           , ZN => n275);
   U330 : NOR2_X1 port map( A1 => n287, A2 => n278, ZN => n687);
   U331 : NOR2_X1 port map( A1 => n283, A2 => n277, ZN => n686);
   U332 : AOI22_X1 port map( A1 => n253, A2 => Q(512), B1 => n252, B2 => Q(608)
                           , ZN => n274);
   U333 : NAND3_X1 port map( A1 => S(3), A2 => S(0), A3 => n276, ZN => n280);
   U334 : NOR2_X1 port map( A1 => n286, A2 => n280, ZN => n691);
   U335 : NOR2_X1 port map( A1 => n287, A2 => n277, ZN => n690);
   U336 : NOR2_X1 port map( A1 => n284, A2 => n278, ZN => n693);
   U337 : NOR2_X1 port map( A1 => S(4), A2 => S(0), ZN => n282);
   U338 : NAND2_X1 port map( A1 => S(3), A2 => n282, ZN => n279);
   U339 : NOR2_X1 port map( A1 => n286, A2 => n279, ZN => n692);
   U340 : NOR2_X1 port map( A1 => n283, A2 => n280, ZN => n695);
   U341 : NOR2_X1 port map( A1 => n287, A2 => n280, ZN => n694);
   U342 : NOR2_X1 port map( A1 => n284, A2 => n279, ZN => n697);
   U343 : NOR2_X1 port map( A1 => n287, A2 => n279, ZN => n696);
   U344 : NOR2_X1 port map( A1 => n283, A2 => n279, ZN => n699);
   U345 : NOR2_X1 port map( A1 => n284, A2 => n280, ZN => n698);
   U346 : NOR2_X1 port map( A1 => n288, A2 => n286, ZN => n701);
   U347 : NAND2_X1 port map( A1 => n282, A2 => n281, ZN => n285);
   U348 : NOR2_X1 port map( A1 => n284, A2 => n285, ZN => n700);
   U349 : NOR2_X1 port map( A1 => n283, A2 => n285, ZN => n703);
   U350 : NOR2_X1 port map( A1 => n288, A2 => n284, ZN => n702);
   U351 : NOR2_X1 port map( A1 => n286, A2 => n285, ZN => n705);
   U352 : NOR2_X1 port map( A1 => n288, A2 => n287, ZN => n704);
   U353 : AOI22_X1 port map( A1 => n674, A2 => Q(1002), B1 => n673, B2 => 
                           Q(938), ZN => n292);
   U354 : AOI22_X1 port map( A1 => n676, A2 => Q(970), B1 => n675, B2 => Q(906)
                           , ZN => n291);
   U355 : AOI22_X1 port map( A1 => n678, A2 => Q(810), B1 => n677, B2 => Q(746)
                           , ZN => n290);
   U356 : NAND2_X1 port map( A1 => n679, A2 => Q(106), ZN => n289);
   U357 : NAND4_X1 port map( A1 => n292, A2 => n291, A3 => n290, A4 => n289, ZN
                           => n308);
   U358 : AOI22_X1 port map( A1 => n681, A2 => Q(842), B1 => n680, B2 => Q(714)
                           , ZN => n296);
   U359 : AOI22_X1 port map( A1 => n683, A2 => Q(778), B1 => n682, B2 => Q(874)
                           , ZN => n295);
   U360 : AOI22_X1 port map( A1 => n685, A2 => Q(682), B1 => n684, B2 => Q(586)
                           , ZN => n294);
   U361 : AOI22_X1 port map( A1 => n687, A2 => Q(522), B1 => n686, B2 => Q(618)
                           , ZN => n293);
   U362 : NAND4_X1 port map( A1 => n296, A2 => n295, A3 => n294, A4 => n293, ZN
                           => n307);
   U363 : AOI22_X1 port map( A1 => n691, A2 => Q(490), B1 => n690, B2 => Q(554)
                           , ZN => n300);
   U364 : AOI22_X1 port map( A1 => n693, A2 => Q(650), B1 => n692, B2 => Q(458)
                           , ZN => n299);
   U365 : AOI22_X1 port map( A1 => n695, A2 => Q(362), B1 => n694, B2 => Q(298)
                           , ZN => n298);
   U366 : AOI22_X1 port map( A1 => n697, A2 => Q(394), B1 => n696, B2 => Q(266)
                           , ZN => n297);
   U367 : NAND4_X1 port map( A1 => n300, A2 => n299, A3 => n298, A4 => n297, ZN
                           => n306);
   U368 : AOI22_X1 port map( A1 => n699, A2 => Q(330), B1 => n698, B2 => Q(426)
                           , ZN => n304);
   U369 : AOI22_X1 port map( A1 => n701, A2 => Q(234), B1 => n700, B2 => Q(138)
                           , ZN => n303);
   U370 : AOI22_X1 port map( A1 => n703, A2 => Q(74), B1 => n702, B2 => Q(170),
                           ZN => n302);
   U371 : AOI22_X1 port map( A1 => n705, A2 => Q(202), B1 => n704, B2 => Q(42),
                           ZN => n301);
   U372 : NAND4_X1 port map( A1 => n304, A2 => n303, A3 => n302, A4 => n301, ZN
                           => n305);
   U373 : AOI22_X1 port map( A1 => n251, A2 => Q(683), B1 => n250, B2 => Q(587)
                           , ZN => n310);
   U374 : AOI22_X1 port map( A1 => n253, A2 => Q(523), B1 => n252, B2 => Q(619)
                           , ZN => n309);
   U375 : AOI22_X1 port map( A1 => n674, A2 => Q(1004), B1 => n673, B2 => 
                           Q(940), ZN => n314);
   U376 : AOI22_X1 port map( A1 => n676, A2 => Q(972), B1 => n675, B2 => Q(908)
                           , ZN => n313);
   U377 : AOI22_X1 port map( A1 => n678, A2 => Q(812), B1 => n677, B2 => Q(748)
                           , ZN => n312);
   U378 : NAND2_X1 port map( A1 => n679, A2 => Q(108), ZN => n311);
   U379 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => n330);
   U380 : AOI22_X1 port map( A1 => n681, A2 => Q(844), B1 => n680, B2 => Q(716)
                           , ZN => n318);
   U381 : AOI22_X1 port map( A1 => n683, A2 => Q(780), B1 => n682, B2 => Q(876)
                           , ZN => n317);
   U382 : AOI22_X1 port map( A1 => n685, A2 => Q(684), B1 => n684, B2 => Q(588)
                           , ZN => n316);
   U383 : AOI22_X1 port map( A1 => n687, A2 => Q(524), B1 => n686, B2 => Q(620)
                           , ZN => n315);
   U384 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => n329);
   U385 : AOI22_X1 port map( A1 => n691, A2 => Q(492), B1 => n690, B2 => Q(556)
                           , ZN => n322);
   U386 : AOI22_X1 port map( A1 => n693, A2 => Q(652), B1 => n692, B2 => Q(460)
                           , ZN => n321);
   U387 : AOI22_X1 port map( A1 => n695, A2 => Q(364), B1 => n694, B2 => Q(300)
                           , ZN => n320);
   U388 : AOI22_X1 port map( A1 => n697, A2 => Q(396), B1 => n696, B2 => Q(268)
                           , ZN => n319);
   U389 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => n328);
   U390 : AOI22_X1 port map( A1 => n699, A2 => Q(332), B1 => n698, B2 => Q(428)
                           , ZN => n326);
   U391 : AOI22_X1 port map( A1 => n701, A2 => Q(236), B1 => n700, B2 => Q(140)
                           , ZN => n325);
   U392 : AOI22_X1 port map( A1 => n703, A2 => Q(76), B1 => n702, B2 => Q(172),
                           ZN => n324);
   U393 : AOI22_X1 port map( A1 => n705, A2 => Q(204), B1 => n704, B2 => Q(44),
                           ZN => n323);
   U394 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => n327);
   U395 : AOI22_X1 port map( A1 => n251, A2 => Q(685), B1 => n250, B2 => Q(589)
                           , ZN => n332);
   U396 : AOI22_X1 port map( A1 => n253, A2 => Q(525), B1 => n252, B2 => Q(621)
                           , ZN => n331);
   U397 : AOI22_X1 port map( A1 => n674, A2 => Q(1006), B1 => n673, B2 => 
                           Q(942), ZN => n336);
   U398 : AOI22_X1 port map( A1 => n676, A2 => Q(974), B1 => n675, B2 => Q(910)
                           , ZN => n335);
   U399 : AOI22_X1 port map( A1 => n678, A2 => Q(814), B1 => n677, B2 => Q(750)
                           , ZN => n334);
   U400 : NAND2_X1 port map( A1 => n679, A2 => Q(110), ZN => n333);
   U401 : NAND4_X1 port map( A1 => n336, A2 => n335, A3 => n334, A4 => n333, ZN
                           => n352);
   U402 : AOI22_X1 port map( A1 => n681, A2 => Q(846), B1 => n680, B2 => Q(718)
                           , ZN => n340);
   U403 : AOI22_X1 port map( A1 => n683, A2 => Q(782), B1 => n682, B2 => Q(878)
                           , ZN => n339);
   U404 : AOI22_X1 port map( A1 => n685, A2 => Q(686), B1 => n684, B2 => Q(590)
                           , ZN => n338);
   U405 : AOI22_X1 port map( A1 => n687, A2 => Q(526), B1 => n686, B2 => Q(622)
                           , ZN => n337);
   U406 : NAND4_X1 port map( A1 => n340, A2 => n339, A3 => n338, A4 => n337, ZN
                           => n351);
   U407 : AOI22_X1 port map( A1 => n691, A2 => Q(494), B1 => n690, B2 => Q(558)
                           , ZN => n344);
   U408 : AOI22_X1 port map( A1 => n693, A2 => Q(654), B1 => n692, B2 => Q(462)
                           , ZN => n343);
   U409 : AOI22_X1 port map( A1 => n695, A2 => Q(366), B1 => n694, B2 => Q(302)
                           , ZN => n342);
   U410 : AOI22_X1 port map( A1 => n697, A2 => Q(398), B1 => n696, B2 => Q(270)
                           , ZN => n341);
   U411 : NAND4_X1 port map( A1 => n344, A2 => n343, A3 => n342, A4 => n341, ZN
                           => n350);
   U412 : AOI22_X1 port map( A1 => n699, A2 => Q(334), B1 => n698, B2 => Q(430)
                           , ZN => n348);
   U413 : AOI22_X1 port map( A1 => n701, A2 => Q(238), B1 => n700, B2 => Q(142)
                           , ZN => n347);
   U414 : AOI22_X1 port map( A1 => n703, A2 => Q(78), B1 => n702, B2 => Q(174),
                           ZN => n346);
   U415 : AOI22_X1 port map( A1 => n705, A2 => Q(206), B1 => n704, B2 => Q(46),
                           ZN => n345);
   U416 : NAND4_X1 port map( A1 => n348, A2 => n347, A3 => n346, A4 => n345, ZN
                           => n349);
   U417 : AOI22_X1 port map( A1 => n674, A2 => Q(1007), B1 => n673, B2 => 
                           Q(943), ZN => n356);
   U418 : AOI22_X1 port map( A1 => n676, A2 => Q(975), B1 => n675, B2 => Q(911)
                           , ZN => n355);
   U419 : AOI22_X1 port map( A1 => n678, A2 => Q(815), B1 => n677, B2 => Q(751)
                           , ZN => n354);
   U420 : NAND2_X1 port map( A1 => n679, A2 => Q(111), ZN => n353);
   U421 : NAND4_X1 port map( A1 => n356, A2 => n355, A3 => n354, A4 => n353, ZN
                           => n372);
   U422 : AOI22_X1 port map( A1 => n681, A2 => Q(847), B1 => n680, B2 => Q(719)
                           , ZN => n360);
   U423 : AOI22_X1 port map( A1 => n683, A2 => Q(783), B1 => n682, B2 => Q(879)
                           , ZN => n359);
   U424 : AOI22_X1 port map( A1 => n685, A2 => Q(687), B1 => n684, B2 => Q(591)
                           , ZN => n358);
   U425 : AOI22_X1 port map( A1 => n687, A2 => Q(527), B1 => n686, B2 => Q(623)
                           , ZN => n357);
   U426 : NAND4_X1 port map( A1 => n360, A2 => n359, A3 => n358, A4 => n357, ZN
                           => n371);
   U427 : AOI22_X1 port map( A1 => n691, A2 => Q(495), B1 => n690, B2 => Q(559)
                           , ZN => n364);
   U428 : AOI22_X1 port map( A1 => n693, A2 => Q(655), B1 => n692, B2 => Q(463)
                           , ZN => n363);
   U429 : AOI22_X1 port map( A1 => n695, A2 => Q(367), B1 => n694, B2 => Q(303)
                           , ZN => n362);
   U430 : AOI22_X1 port map( A1 => n697, A2 => Q(399), B1 => n696, B2 => Q(271)
                           , ZN => n361);
   U431 : NAND4_X1 port map( A1 => n364, A2 => n363, A3 => n362, A4 => n361, ZN
                           => n370);
   U432 : AOI22_X1 port map( A1 => n699, A2 => Q(335), B1 => n698, B2 => Q(431)
                           , ZN => n368);
   U433 : AOI22_X1 port map( A1 => n701, A2 => Q(239), B1 => n700, B2 => Q(143)
                           , ZN => n367);
   U434 : AOI22_X1 port map( A1 => n703, A2 => Q(79), B1 => n702, B2 => Q(175),
                           ZN => n366);
   U435 : AOI22_X1 port map( A1 => n705, A2 => Q(207), B1 => n704, B2 => Q(47),
                           ZN => n365);
   U436 : NAND4_X1 port map( A1 => n368, A2 => n367, A3 => n366, A4 => n365, ZN
                           => n369);
   U437 : AOI22_X1 port map( A1 => n674, A2 => Q(1008), B1 => n673, B2 => 
                           Q(944), ZN => n376);
   U438 : AOI22_X1 port map( A1 => n676, A2 => Q(976), B1 => n675, B2 => Q(912)
                           , ZN => n375);
   U439 : AOI22_X1 port map( A1 => n678, A2 => Q(816), B1 => n677, B2 => Q(752)
                           , ZN => n374);
   U440 : NAND2_X1 port map( A1 => n679, A2 => Q(112), ZN => n373);
   U441 : NAND4_X1 port map( A1 => n376, A2 => n375, A3 => n374, A4 => n373, ZN
                           => n392);
   U442 : AOI22_X1 port map( A1 => n681, A2 => Q(848), B1 => n680, B2 => Q(720)
                           , ZN => n380);
   U443 : AOI22_X1 port map( A1 => n683, A2 => Q(784), B1 => n682, B2 => Q(880)
                           , ZN => n379);
   U444 : AOI22_X1 port map( A1 => n685, A2 => Q(688), B1 => n684, B2 => Q(592)
                           , ZN => n378);
   U445 : AOI22_X1 port map( A1 => n687, A2 => Q(528), B1 => n686, B2 => Q(624)
                           , ZN => n377);
   U446 : NAND4_X1 port map( A1 => n380, A2 => n379, A3 => n378, A4 => n377, ZN
                           => n391);
   U447 : AOI22_X1 port map( A1 => n691, A2 => Q(496), B1 => n690, B2 => Q(560)
                           , ZN => n384);
   U448 : AOI22_X1 port map( A1 => n693, A2 => Q(656), B1 => n692, B2 => Q(464)
                           , ZN => n383);
   U449 : AOI22_X1 port map( A1 => n695, A2 => Q(368), B1 => n694, B2 => Q(304)
                           , ZN => n382);
   U450 : AOI22_X1 port map( A1 => n697, A2 => Q(400), B1 => n696, B2 => Q(272)
                           , ZN => n381);
   U451 : NAND4_X1 port map( A1 => n384, A2 => n383, A3 => n382, A4 => n381, ZN
                           => n390);
   U452 : AOI22_X1 port map( A1 => n699, A2 => Q(336), B1 => n698, B2 => Q(432)
                           , ZN => n388);
   U453 : AOI22_X1 port map( A1 => n701, A2 => Q(240), B1 => n700, B2 => Q(144)
                           , ZN => n387);
   U454 : AOI22_X1 port map( A1 => n703, A2 => Q(80), B1 => n702, B2 => Q(176),
                           ZN => n386);
   U455 : AOI22_X1 port map( A1 => n705, A2 => Q(208), B1 => n704, B2 => Q(48),
                           ZN => n385);
   U456 : NAND4_X1 port map( A1 => n388, A2 => n387, A3 => n386, A4 => n385, ZN
                           => n389);
   U457 : AOI22_X1 port map( A1 => n674, A2 => Q(1009), B1 => n673, B2 => 
                           Q(945), ZN => n396);
   U458 : AOI22_X1 port map( A1 => n676, A2 => Q(977), B1 => n675, B2 => Q(913)
                           , ZN => n395);
   U459 : AOI22_X1 port map( A1 => n678, A2 => Q(817), B1 => n677, B2 => Q(753)
                           , ZN => n394);
   U460 : NAND2_X1 port map( A1 => n679, A2 => Q(113), ZN => n393);
   U461 : NAND4_X1 port map( A1 => n396, A2 => n395, A3 => n394, A4 => n393, ZN
                           => n412);
   U462 : AOI22_X1 port map( A1 => n681, A2 => Q(849), B1 => n680, B2 => Q(721)
                           , ZN => n400);
   U463 : AOI22_X1 port map( A1 => n683, A2 => Q(785), B1 => n682, B2 => Q(881)
                           , ZN => n399);
   U464 : AOI22_X1 port map( A1 => n685, A2 => Q(689), B1 => n684, B2 => Q(593)
                           , ZN => n398);
   U465 : AOI22_X1 port map( A1 => n687, A2 => Q(529), B1 => n686, B2 => Q(625)
                           , ZN => n397);
   U466 : NAND4_X1 port map( A1 => n400, A2 => n399, A3 => n398, A4 => n397, ZN
                           => n411);
   U467 : AOI22_X1 port map( A1 => n691, A2 => Q(497), B1 => n690, B2 => Q(561)
                           , ZN => n404);
   U468 : AOI22_X1 port map( A1 => n693, A2 => Q(657), B1 => n692, B2 => Q(465)
                           , ZN => n403);
   U469 : AOI22_X1 port map( A1 => n695, A2 => Q(369), B1 => n694, B2 => Q(305)
                           , ZN => n402);
   U470 : AOI22_X1 port map( A1 => n697, A2 => Q(401), B1 => n696, B2 => Q(273)
                           , ZN => n401);
   U471 : NAND4_X1 port map( A1 => n404, A2 => n403, A3 => n402, A4 => n401, ZN
                           => n410);
   U472 : AOI22_X1 port map( A1 => n699, A2 => Q(337), B1 => n698, B2 => Q(433)
                           , ZN => n408);
   U473 : AOI22_X1 port map( A1 => n701, A2 => Q(241), B1 => n700, B2 => Q(145)
                           , ZN => n407);
   U474 : AOI22_X1 port map( A1 => n703, A2 => Q(81), B1 => n702, B2 => Q(177),
                           ZN => n406);
   U475 : AOI22_X1 port map( A1 => n705, A2 => Q(209), B1 => n704, B2 => Q(49),
                           ZN => n405);
   U476 : NAND4_X1 port map( A1 => n408, A2 => n407, A3 => n406, A4 => n405, ZN
                           => n409);
   U477 : AOI22_X1 port map( A1 => n674, A2 => Q(1010), B1 => n673, B2 => 
                           Q(946), ZN => n416);
   U478 : AOI22_X1 port map( A1 => n676, A2 => Q(978), B1 => n675, B2 => Q(914)
                           , ZN => n415);
   U479 : AOI22_X1 port map( A1 => n678, A2 => Q(818), B1 => n677, B2 => Q(754)
                           , ZN => n414);
   U480 : NAND2_X1 port map( A1 => n679, A2 => Q(114), ZN => n413);
   U481 : NAND4_X1 port map( A1 => n416, A2 => n415, A3 => n414, A4 => n413, ZN
                           => n432);
   U482 : AOI22_X1 port map( A1 => n681, A2 => Q(850), B1 => n680, B2 => Q(722)
                           , ZN => n420);
   U483 : AOI22_X1 port map( A1 => n683, A2 => Q(786), B1 => n682, B2 => Q(882)
                           , ZN => n419);
   U484 : AOI22_X1 port map( A1 => n685, A2 => Q(690), B1 => n684, B2 => Q(594)
                           , ZN => n418);
   U485 : AOI22_X1 port map( A1 => n687, A2 => Q(530), B1 => n686, B2 => Q(626)
                           , ZN => n417);
   U486 : NAND4_X1 port map( A1 => n420, A2 => n419, A3 => n418, A4 => n417, ZN
                           => n431);
   U487 : AOI22_X1 port map( A1 => n691, A2 => Q(498), B1 => n690, B2 => Q(562)
                           , ZN => n424);
   U488 : AOI22_X1 port map( A1 => n693, A2 => Q(658), B1 => n692, B2 => Q(466)
                           , ZN => n423);
   U489 : AOI22_X1 port map( A1 => n695, A2 => Q(370), B1 => n694, B2 => Q(306)
                           , ZN => n422);
   U490 : AOI22_X1 port map( A1 => n697, A2 => Q(402), B1 => n696, B2 => Q(274)
                           , ZN => n421);
   U491 : NAND4_X1 port map( A1 => n424, A2 => n423, A3 => n422, A4 => n421, ZN
                           => n430);
   U492 : AOI22_X1 port map( A1 => n699, A2 => Q(338), B1 => n698, B2 => Q(434)
                           , ZN => n428);
   U493 : AOI22_X1 port map( A1 => n701, A2 => Q(242), B1 => n700, B2 => Q(146)
                           , ZN => n427);
   U494 : AOI22_X1 port map( A1 => n703, A2 => Q(82), B1 => n702, B2 => Q(178),
                           ZN => n426);
   U495 : AOI22_X1 port map( A1 => n705, A2 => Q(210), B1 => n704, B2 => Q(50),
                           ZN => n425);
   U496 : NAND4_X1 port map( A1 => n428, A2 => n427, A3 => n426, A4 => n425, ZN
                           => n429);
   U497 : AOI22_X1 port map( A1 => n674, A2 => Q(1011), B1 => n673, B2 => 
                           Q(947), ZN => n436);
   U498 : AOI22_X1 port map( A1 => n676, A2 => Q(979), B1 => n675, B2 => Q(915)
                           , ZN => n435);
   U499 : AOI22_X1 port map( A1 => n678, A2 => Q(819), B1 => n677, B2 => Q(755)
                           , ZN => n434);
   U500 : NAND2_X1 port map( A1 => n679, A2 => Q(115), ZN => n433);
   U501 : NAND4_X1 port map( A1 => n436, A2 => n435, A3 => n434, A4 => n433, ZN
                           => n452);
   U502 : AOI22_X1 port map( A1 => n681, A2 => Q(851), B1 => n680, B2 => Q(723)
                           , ZN => n440);
   U503 : AOI22_X1 port map( A1 => n683, A2 => Q(787), B1 => n682, B2 => Q(883)
                           , ZN => n439);
   U504 : AOI22_X1 port map( A1 => n685, A2 => Q(691), B1 => n684, B2 => Q(595)
                           , ZN => n438);
   U505 : AOI22_X1 port map( A1 => n687, A2 => Q(531), B1 => n686, B2 => Q(627)
                           , ZN => n437);
   U506 : NAND4_X1 port map( A1 => n440, A2 => n439, A3 => n438, A4 => n437, ZN
                           => n451);
   U507 : AOI22_X1 port map( A1 => n691, A2 => Q(499), B1 => n690, B2 => Q(563)
                           , ZN => n444);
   U508 : AOI22_X1 port map( A1 => n693, A2 => Q(659), B1 => n692, B2 => Q(467)
                           , ZN => n443);
   U509 : AOI22_X1 port map( A1 => n695, A2 => Q(371), B1 => n694, B2 => Q(307)
                           , ZN => n442);
   U510 : AOI22_X1 port map( A1 => n697, A2 => Q(403), B1 => n696, B2 => Q(275)
                           , ZN => n441);
   U511 : NAND4_X1 port map( A1 => n444, A2 => n443, A3 => n442, A4 => n441, ZN
                           => n450);
   U512 : AOI22_X1 port map( A1 => n699, A2 => Q(339), B1 => n698, B2 => Q(435)
                           , ZN => n448);
   U513 : AOI22_X1 port map( A1 => n701, A2 => Q(243), B1 => n700, B2 => Q(147)
                           , ZN => n447);
   U514 : AOI22_X1 port map( A1 => n703, A2 => Q(83), B1 => n702, B2 => Q(179),
                           ZN => n446);
   U515 : AOI22_X1 port map( A1 => n705, A2 => Q(211), B1 => n704, B2 => Q(51),
                           ZN => n445);
   U516 : NAND4_X1 port map( A1 => n448, A2 => n447, A3 => n446, A4 => n445, ZN
                           => n449);
   U517 : AOI22_X1 port map( A1 => n685, A2 => Q(673), B1 => n684, B2 => Q(577)
                           , ZN => n454);
   U518 : AOI22_X1 port map( A1 => n687, A2 => Q(513), B1 => n686, B2 => Q(609)
                           , ZN => n453);
   U519 : AOI22_X1 port map( A1 => n251, A2 => Q(692), B1 => n250, B2 => Q(596)
                           , ZN => n456);
   U520 : AOI22_X1 port map( A1 => n253, A2 => Q(532), B1 => n252, B2 => Q(628)
                           , ZN => n455);
   U521 : AOI22_X1 port map( A1 => n251, A2 => Q(693), B1 => n250, B2 => Q(597)
                           , ZN => n458);
   U522 : AOI22_X1 port map( A1 => n253, A2 => Q(533), B1 => n252, B2 => Q(629)
                           , ZN => n457);
   U523 : AOI22_X1 port map( A1 => n240, A2 => Q(1014), B1 => n239, B2 => 
                           Q(950), ZN => n462);
   U524 : AOI22_X1 port map( A1 => n242, A2 => Q(982), B1 => n241, B2 => Q(918)
                           , ZN => n461);
   U525 : AOI22_X1 port map( A1 => n244, A2 => Q(822), B1 => n243, B2 => Q(758)
                           , ZN => n460);
   U526 : NAND2_X1 port map( A1 => n245, A2 => Q(118), ZN => n459);
   U527 : NAND4_X1 port map( A1 => n462, A2 => n461, A3 => n460, A4 => n459, ZN
                           => n478);
   U528 : AOI22_X1 port map( A1 => n247, A2 => Q(854), B1 => n246, B2 => Q(726)
                           , ZN => n466);
   U529 : AOI22_X1 port map( A1 => n249, A2 => Q(790), B1 => n248, B2 => Q(886)
                           , ZN => n465);
   U530 : AOI22_X1 port map( A1 => n251, A2 => Q(694), B1 => n250, B2 => Q(598)
                           , ZN => n464);
   U531 : AOI22_X1 port map( A1 => n253, A2 => Q(534), B1 => n252, B2 => Q(630)
                           , ZN => n463);
   U532 : NAND4_X1 port map( A1 => n466, A2 => n465, A3 => n464, A4 => n463, ZN
                           => n477);
   U533 : AOI22_X1 port map( A1 => n255, A2 => Q(502), B1 => n254, B2 => Q(566)
                           , ZN => n470);
   U534 : AOI22_X1 port map( A1 => n257, A2 => Q(662), B1 => n256, B2 => Q(470)
                           , ZN => n469);
   U535 : AOI22_X1 port map( A1 => n259, A2 => Q(374), B1 => n258, B2 => Q(310)
                           , ZN => n468);
   U536 : AOI22_X1 port map( A1 => n261, A2 => Q(406), B1 => n260, B2 => Q(278)
                           , ZN => n467);
   U537 : NAND4_X1 port map( A1 => n470, A2 => n469, A3 => n468, A4 => n467, ZN
                           => n476);
   U538 : AOI22_X1 port map( A1 => n263, A2 => Q(342), B1 => n262, B2 => Q(438)
                           , ZN => n474);
   U539 : AOI22_X1 port map( A1 => n265, A2 => Q(246), B1 => n264, B2 => Q(150)
                           , ZN => n473);
   U540 : AOI22_X1 port map( A1 => n267, A2 => Q(86), B1 => n266, B2 => Q(182),
                           ZN => n472);
   U541 : AOI22_X1 port map( A1 => n269, A2 => Q(214), B1 => n268, B2 => Q(54),
                           ZN => n471);
   U542 : NAND4_X1 port map( A1 => n474, A2 => n473, A3 => n472, A4 => n471, ZN
                           => n475);
   U543 : AOI22_X1 port map( A1 => n240, A2 => Q(1015), B1 => n239, B2 => 
                           Q(951), ZN => n482);
   U544 : AOI22_X1 port map( A1 => n242, A2 => Q(983), B1 => n241, B2 => Q(919)
                           , ZN => n481);
   U545 : AOI22_X1 port map( A1 => n244, A2 => Q(823), B1 => n243, B2 => Q(759)
                           , ZN => n480);
   U546 : NAND2_X1 port map( A1 => n245, A2 => Q(119), ZN => n479);
   U547 : NAND4_X1 port map( A1 => n482, A2 => n481, A3 => n480, A4 => n479, ZN
                           => n498);
   U548 : AOI22_X1 port map( A1 => n247, A2 => Q(855), B1 => n246, B2 => Q(727)
                           , ZN => n486);
   U549 : AOI22_X1 port map( A1 => n249, A2 => Q(791), B1 => n248, B2 => Q(887)
                           , ZN => n485);
   U550 : AOI22_X1 port map( A1 => n251, A2 => Q(695), B1 => n250, B2 => Q(599)
                           , ZN => n484);
   U551 : AOI22_X1 port map( A1 => n253, A2 => Q(535), B1 => n252, B2 => Q(631)
                           , ZN => n483);
   U552 : NAND4_X1 port map( A1 => n486, A2 => n485, A3 => n484, A4 => n483, ZN
                           => n497);
   U553 : AOI22_X1 port map( A1 => n255, A2 => Q(503), B1 => n254, B2 => Q(567)
                           , ZN => n490);
   U554 : AOI22_X1 port map( A1 => n257, A2 => Q(663), B1 => n256, B2 => Q(471)
                           , ZN => n489);
   U555 : AOI22_X1 port map( A1 => n259, A2 => Q(375), B1 => n258, B2 => Q(311)
                           , ZN => n488);
   U556 : AOI22_X1 port map( A1 => n261, A2 => Q(407), B1 => n260, B2 => Q(279)
                           , ZN => n487);
   U557 : NAND4_X1 port map( A1 => n490, A2 => n489, A3 => n488, A4 => n487, ZN
                           => n496);
   U558 : AOI22_X1 port map( A1 => n263, A2 => Q(343), B1 => n262, B2 => Q(439)
                           , ZN => n494);
   U559 : AOI22_X1 port map( A1 => n265, A2 => Q(247), B1 => n264, B2 => Q(151)
                           , ZN => n493);
   U560 : AOI22_X1 port map( A1 => n267, A2 => Q(87), B1 => n266, B2 => Q(183),
                           ZN => n492);
   U561 : AOI22_X1 port map( A1 => n269, A2 => Q(215), B1 => n268, B2 => Q(55),
                           ZN => n491);
   U562 : NAND4_X1 port map( A1 => n494, A2 => n493, A3 => n492, A4 => n491, ZN
                           => n495);
   U563 : AOI22_X1 port map( A1 => n240, A2 => Q(1016), B1 => n239, B2 => 
                           Q(952), ZN => n502);
   U564 : AOI22_X1 port map( A1 => n242, A2 => Q(984), B1 => n241, B2 => Q(920)
                           , ZN => n501);
   U565 : AOI22_X1 port map( A1 => n244, A2 => Q(824), B1 => n243, B2 => Q(760)
                           , ZN => n500);
   U566 : NAND2_X1 port map( A1 => n245, A2 => Q(120), ZN => n499);
   U567 : NAND4_X1 port map( A1 => n502, A2 => n501, A3 => n500, A4 => n499, ZN
                           => n518);
   U568 : AOI22_X1 port map( A1 => n247, A2 => Q(856), B1 => n246, B2 => Q(728)
                           , ZN => n506);
   U569 : AOI22_X1 port map( A1 => n249, A2 => Q(792), B1 => n248, B2 => Q(888)
                           , ZN => n505);
   U570 : AOI22_X1 port map( A1 => n251, A2 => Q(696), B1 => n250, B2 => Q(600)
                           , ZN => n504);
   U571 : AOI22_X1 port map( A1 => n253, A2 => Q(536), B1 => n252, B2 => Q(632)
                           , ZN => n503);
   U572 : NAND4_X1 port map( A1 => n506, A2 => n505, A3 => n504, A4 => n503, ZN
                           => n517);
   U573 : AOI22_X1 port map( A1 => n255, A2 => Q(504), B1 => n254, B2 => Q(568)
                           , ZN => n510);
   U574 : AOI22_X1 port map( A1 => n257, A2 => Q(664), B1 => n256, B2 => Q(472)
                           , ZN => n509);
   U575 : AOI22_X1 port map( A1 => n259, A2 => Q(376), B1 => n258, B2 => Q(312)
                           , ZN => n508);
   U576 : AOI22_X1 port map( A1 => n261, A2 => Q(408), B1 => n260, B2 => Q(280)
                           , ZN => n507);
   U577 : NAND4_X1 port map( A1 => n510, A2 => n509, A3 => n508, A4 => n507, ZN
                           => n516);
   U578 : AOI22_X1 port map( A1 => n263, A2 => Q(344), B1 => n262, B2 => Q(440)
                           , ZN => n514);
   U579 : AOI22_X1 port map( A1 => n265, A2 => Q(248), B1 => n264, B2 => Q(152)
                           , ZN => n513);
   U580 : AOI22_X1 port map( A1 => n267, A2 => Q(88), B1 => n266, B2 => Q(184),
                           ZN => n512);
   U581 : AOI22_X1 port map( A1 => n269, A2 => Q(216), B1 => n268, B2 => Q(56),
                           ZN => n511);
   U582 : NAND4_X1 port map( A1 => n514, A2 => n513, A3 => n512, A4 => n511, ZN
                           => n515);
   U583 : AOI22_X1 port map( A1 => n240, A2 => Q(1017), B1 => n239, B2 => 
                           Q(953), ZN => n522);
   U584 : AOI22_X1 port map( A1 => n242, A2 => Q(985), B1 => n241, B2 => Q(921)
                           , ZN => n521);
   U585 : AOI22_X1 port map( A1 => n244, A2 => Q(825), B1 => n243, B2 => Q(761)
                           , ZN => n520);
   U586 : NAND2_X1 port map( A1 => n245, A2 => Q(121), ZN => n519);
   U587 : NAND4_X1 port map( A1 => n522, A2 => n521, A3 => n520, A4 => n519, ZN
                           => n538);
   U588 : AOI22_X1 port map( A1 => n247, A2 => Q(857), B1 => n246, B2 => Q(729)
                           , ZN => n526);
   U589 : AOI22_X1 port map( A1 => n249, A2 => Q(793), B1 => n248, B2 => Q(889)
                           , ZN => n525);
   U590 : AOI22_X1 port map( A1 => n251, A2 => Q(697), B1 => n250, B2 => Q(601)
                           , ZN => n524);
   U591 : AOI22_X1 port map( A1 => n253, A2 => Q(537), B1 => n252, B2 => Q(633)
                           , ZN => n523);
   U592 : NAND4_X1 port map( A1 => n526, A2 => n525, A3 => n524, A4 => n523, ZN
                           => n537);
   U593 : AOI22_X1 port map( A1 => n255, A2 => Q(505), B1 => n254, B2 => Q(569)
                           , ZN => n530);
   U594 : AOI22_X1 port map( A1 => n257, A2 => Q(665), B1 => n256, B2 => Q(473)
                           , ZN => n529);
   U595 : AOI22_X1 port map( A1 => n259, A2 => Q(377), B1 => n258, B2 => Q(313)
                           , ZN => n528);
   U596 : AOI22_X1 port map( A1 => n261, A2 => Q(409), B1 => n260, B2 => Q(281)
                           , ZN => n527);
   U597 : NAND4_X1 port map( A1 => n530, A2 => n529, A3 => n528, A4 => n527, ZN
                           => n536);
   U598 : AOI22_X1 port map( A1 => n263, A2 => Q(345), B1 => n262, B2 => Q(441)
                           , ZN => n534);
   U599 : AOI22_X1 port map( A1 => n265, A2 => Q(249), B1 => n264, B2 => Q(153)
                           , ZN => n533);
   U600 : AOI22_X1 port map( A1 => n267, A2 => Q(89), B1 => n266, B2 => Q(185),
                           ZN => n532);
   U601 : AOI22_X1 port map( A1 => n269, A2 => Q(217), B1 => n268, B2 => Q(57),
                           ZN => n531);
   U602 : NAND4_X1 port map( A1 => n534, A2 => n533, A3 => n532, A4 => n531, ZN
                           => n535);
   U603 : AOI22_X1 port map( A1 => n240, A2 => Q(1018), B1 => n239, B2 => 
                           Q(954), ZN => n542);
   U604 : AOI22_X1 port map( A1 => n242, A2 => Q(986), B1 => n241, B2 => Q(922)
                           , ZN => n541);
   U605 : AOI22_X1 port map( A1 => n244, A2 => Q(826), B1 => n243, B2 => Q(762)
                           , ZN => n540);
   U606 : NAND2_X1 port map( A1 => n245, A2 => Q(122), ZN => n539);
   U607 : NAND4_X1 port map( A1 => n542, A2 => n541, A3 => n540, A4 => n539, ZN
                           => n558);
   U608 : AOI22_X1 port map( A1 => n247, A2 => Q(858), B1 => n246, B2 => Q(730)
                           , ZN => n546);
   U609 : AOI22_X1 port map( A1 => n249, A2 => Q(794), B1 => n248, B2 => Q(890)
                           , ZN => n545);
   U610 : AOI22_X1 port map( A1 => n251, A2 => Q(698), B1 => n250, B2 => Q(602)
                           , ZN => n544);
   U611 : AOI22_X1 port map( A1 => n253, A2 => Q(538), B1 => n252, B2 => Q(634)
                           , ZN => n543);
   U612 : NAND4_X1 port map( A1 => n546, A2 => n545, A3 => n544, A4 => n543, ZN
                           => n557);
   U613 : AOI22_X1 port map( A1 => n255, A2 => Q(506), B1 => n254, B2 => Q(570)
                           , ZN => n550);
   U614 : AOI22_X1 port map( A1 => n257, A2 => Q(666), B1 => n256, B2 => Q(474)
                           , ZN => n549);
   U615 : AOI22_X1 port map( A1 => n259, A2 => Q(378), B1 => n258, B2 => Q(314)
                           , ZN => n548);
   U616 : AOI22_X1 port map( A1 => n261, A2 => Q(410), B1 => n260, B2 => Q(282)
                           , ZN => n547);
   U617 : NAND4_X1 port map( A1 => n550, A2 => n549, A3 => n548, A4 => n547, ZN
                           => n556);
   U618 : AOI22_X1 port map( A1 => n263, A2 => Q(346), B1 => n262, B2 => Q(442)
                           , ZN => n554);
   U619 : AOI22_X1 port map( A1 => n265, A2 => Q(250), B1 => n264, B2 => Q(154)
                           , ZN => n553);
   U620 : AOI22_X1 port map( A1 => n267, A2 => Q(90), B1 => n266, B2 => Q(186),
                           ZN => n552);
   U621 : AOI22_X1 port map( A1 => n269, A2 => Q(218), B1 => n268, B2 => Q(58),
                           ZN => n551);
   U622 : NAND4_X1 port map( A1 => n554, A2 => n553, A3 => n552, A4 => n551, ZN
                           => n555);
   U623 : AOI22_X1 port map( A1 => n240, A2 => Q(1019), B1 => n239, B2 => 
                           Q(955), ZN => n562);
   U624 : AOI22_X1 port map( A1 => n242, A2 => Q(987), B1 => n241, B2 => Q(923)
                           , ZN => n561);
   U625 : AOI22_X1 port map( A1 => n244, A2 => Q(827), B1 => n243, B2 => Q(763)
                           , ZN => n560);
   U626 : NAND2_X1 port map( A1 => n245, A2 => Q(123), ZN => n559);
   U627 : NAND4_X1 port map( A1 => n562, A2 => n561, A3 => n560, A4 => n559, ZN
                           => n578);
   U628 : AOI22_X1 port map( A1 => n247, A2 => Q(859), B1 => n246, B2 => Q(731)
                           , ZN => n566);
   U629 : AOI22_X1 port map( A1 => n249, A2 => Q(795), B1 => n248, B2 => Q(891)
                           , ZN => n565);
   U630 : AOI22_X1 port map( A1 => n251, A2 => Q(699), B1 => n250, B2 => Q(603)
                           , ZN => n564);
   U631 : AOI22_X1 port map( A1 => n253, A2 => Q(539), B1 => n252, B2 => Q(635)
                           , ZN => n563);
   U632 : NAND4_X1 port map( A1 => n566, A2 => n565, A3 => n564, A4 => n563, ZN
                           => n577);
   U633 : AOI22_X1 port map( A1 => n255, A2 => Q(507), B1 => n254, B2 => Q(571)
                           , ZN => n570);
   U634 : AOI22_X1 port map( A1 => n257, A2 => Q(667), B1 => n256, B2 => Q(475)
                           , ZN => n569);
   U635 : AOI22_X1 port map( A1 => n259, A2 => Q(379), B1 => n258, B2 => Q(315)
                           , ZN => n568);
   U636 : AOI22_X1 port map( A1 => n261, A2 => Q(411), B1 => n260, B2 => Q(283)
                           , ZN => n567);
   U637 : NAND4_X1 port map( A1 => n570, A2 => n569, A3 => n568, A4 => n567, ZN
                           => n576);
   U638 : AOI22_X1 port map( A1 => n263, A2 => Q(347), B1 => n262, B2 => Q(443)
                           , ZN => n574);
   U639 : AOI22_X1 port map( A1 => n265, A2 => Q(251), B1 => n264, B2 => Q(155)
                           , ZN => n573);
   U640 : AOI22_X1 port map( A1 => n267, A2 => Q(91), B1 => n266, B2 => Q(187),
                           ZN => n572);
   U641 : AOI22_X1 port map( A1 => n269, A2 => Q(219), B1 => n268, B2 => Q(59),
                           ZN => n571);
   U642 : NAND4_X1 port map( A1 => n574, A2 => n573, A3 => n572, A4 => n571, ZN
                           => n575);
   U643 : AOI22_X1 port map( A1 => n240, A2 => Q(1020), B1 => n673, B2 => 
                           Q(956), ZN => n582);
   U644 : AOI22_X1 port map( A1 => n242, A2 => Q(988), B1 => n675, B2 => Q(924)
                           , ZN => n581);
   U645 : AOI22_X1 port map( A1 => n244, A2 => Q(828), B1 => n677, B2 => Q(764)
                           , ZN => n580);
   U646 : NAND2_X1 port map( A1 => n245, A2 => Q(124), ZN => n579);
   U647 : NAND4_X1 port map( A1 => n582, A2 => n581, A3 => n580, A4 => n579, ZN
                           => n598);
   U648 : AOI22_X1 port map( A1 => n247, A2 => Q(860), B1 => n680, B2 => Q(732)
                           , ZN => n586);
   U649 : AOI22_X1 port map( A1 => n249, A2 => Q(796), B1 => n682, B2 => Q(892)
                           , ZN => n585);
   U650 : AOI22_X1 port map( A1 => n251, A2 => Q(700), B1 => n684, B2 => Q(604)
                           , ZN => n584);
   U651 : AOI22_X1 port map( A1 => n253, A2 => Q(540), B1 => n686, B2 => Q(636)
                           , ZN => n583);
   U652 : NAND4_X1 port map( A1 => n586, A2 => n585, A3 => n584, A4 => n583, ZN
                           => n597);
   U653 : AOI22_X1 port map( A1 => n255, A2 => Q(508), B1 => n690, B2 => Q(572)
                           , ZN => n590);
   U654 : AOI22_X1 port map( A1 => n257, A2 => Q(668), B1 => n692, B2 => Q(476)
                           , ZN => n589);
   U655 : AOI22_X1 port map( A1 => n259, A2 => Q(380), B1 => n694, B2 => Q(316)
                           , ZN => n588);
   U656 : AOI22_X1 port map( A1 => n261, A2 => Q(412), B1 => n696, B2 => Q(284)
                           , ZN => n587);
   U657 : NAND4_X1 port map( A1 => n590, A2 => n589, A3 => n588, A4 => n587, ZN
                           => n596);
   U658 : AOI22_X1 port map( A1 => n263, A2 => Q(348), B1 => n698, B2 => Q(444)
                           , ZN => n594);
   U659 : AOI22_X1 port map( A1 => n265, A2 => Q(252), B1 => n700, B2 => Q(156)
                           , ZN => n593);
   U660 : AOI22_X1 port map( A1 => n267, A2 => Q(92), B1 => n702, B2 => Q(188),
                           ZN => n592);
   U661 : AOI22_X1 port map( A1 => n269, A2 => Q(220), B1 => n704, B2 => Q(60),
                           ZN => n591);
   U662 : NAND4_X1 port map( A1 => n594, A2 => n593, A3 => n592, A4 => n591, ZN
                           => n595);
   U663 : AOI22_X1 port map( A1 => n240, A2 => Q(1021), B1 => n239, B2 => 
                           Q(957), ZN => n602);
   U664 : AOI22_X1 port map( A1 => n242, A2 => Q(989), B1 => n241, B2 => Q(925)
                           , ZN => n601);
   U665 : AOI22_X1 port map( A1 => n244, A2 => Q(829), B1 => n243, B2 => Q(765)
                           , ZN => n600);
   U666 : NAND2_X1 port map( A1 => n245, A2 => Q(125), ZN => n599);
   U667 : NAND4_X1 port map( A1 => n602, A2 => n601, A3 => n600, A4 => n599, ZN
                           => n618);
   U668 : AOI22_X1 port map( A1 => n247, A2 => Q(861), B1 => n246, B2 => Q(733)
                           , ZN => n606);
   U669 : AOI22_X1 port map( A1 => n249, A2 => Q(797), B1 => n248, B2 => Q(893)
                           , ZN => n605);
   U670 : AOI22_X1 port map( A1 => n251, A2 => Q(701), B1 => n250, B2 => Q(605)
                           , ZN => n604);
   U671 : AOI22_X1 port map( A1 => n253, A2 => Q(541), B1 => n252, B2 => Q(637)
                           , ZN => n603);
   U672 : NAND4_X1 port map( A1 => n606, A2 => n605, A3 => n604, A4 => n603, ZN
                           => n617);
   U673 : AOI22_X1 port map( A1 => n255, A2 => Q(509), B1 => n254, B2 => Q(573)
                           , ZN => n610);
   U674 : AOI22_X1 port map( A1 => n257, A2 => Q(669), B1 => n256, B2 => Q(477)
                           , ZN => n609);
   U675 : AOI22_X1 port map( A1 => n259, A2 => Q(381), B1 => n258, B2 => Q(317)
                           , ZN => n608);
   U676 : AOI22_X1 port map( A1 => n261, A2 => Q(413), B1 => n260, B2 => Q(285)
                           , ZN => n607);
   U677 : NAND4_X1 port map( A1 => n610, A2 => n609, A3 => n608, A4 => n607, ZN
                           => n616);
   U678 : AOI22_X1 port map( A1 => n263, A2 => Q(349), B1 => n262, B2 => Q(445)
                           , ZN => n614);
   U679 : AOI22_X1 port map( A1 => n265, A2 => Q(253), B1 => n264, B2 => Q(157)
                           , ZN => n613);
   U680 : AOI22_X1 port map( A1 => n267, A2 => Q(93), B1 => n266, B2 => Q(189),
                           ZN => n612);
   U681 : AOI22_X1 port map( A1 => n269, A2 => Q(221), B1 => n268, B2 => Q(61),
                           ZN => n611);
   U682 : NAND4_X1 port map( A1 => n614, A2 => n613, A3 => n612, A4 => n611, ZN
                           => n615);
   U683 : AOI22_X1 port map( A1 => n674, A2 => Q(994), B1 => n673, B2 => Q(930)
                           , ZN => n622);
   U684 : AOI22_X1 port map( A1 => n676, A2 => Q(962), B1 => n675, B2 => Q(898)
                           , ZN => n621);
   U685 : AOI22_X1 port map( A1 => n678, A2 => Q(802), B1 => n677, B2 => Q(738)
                           , ZN => n620);
   U686 : NAND2_X1 port map( A1 => n679, A2 => Q(98), ZN => n619);
   U687 : NAND4_X1 port map( A1 => n622, A2 => n621, A3 => n620, A4 => n619, ZN
                           => n638);
   U688 : AOI22_X1 port map( A1 => n681, A2 => Q(834), B1 => n680, B2 => Q(706)
                           , ZN => n626);
   U689 : AOI22_X1 port map( A1 => n683, A2 => Q(770), B1 => n682, B2 => Q(866)
                           , ZN => n625);
   U690 : AOI22_X1 port map( A1 => n685, A2 => Q(674), B1 => n684, B2 => Q(578)
                           , ZN => n624);
   U691 : AOI22_X1 port map( A1 => n687, A2 => Q(514), B1 => n686, B2 => Q(610)
                           , ZN => n623);
   U692 : NAND4_X1 port map( A1 => n626, A2 => n625, A3 => n624, A4 => n623, ZN
                           => n637);
   U693 : AOI22_X1 port map( A1 => n691, A2 => Q(482), B1 => n690, B2 => Q(546)
                           , ZN => n630);
   U694 : AOI22_X1 port map( A1 => n693, A2 => Q(642), B1 => n692, B2 => Q(450)
                           , ZN => n629);
   U695 : AOI22_X1 port map( A1 => n695, A2 => Q(354), B1 => n694, B2 => Q(290)
                           , ZN => n628);
   U696 : AOI22_X1 port map( A1 => n697, A2 => Q(386), B1 => n696, B2 => Q(258)
                           , ZN => n627);
   U697 : NAND4_X1 port map( A1 => n630, A2 => n629, A3 => n628, A4 => n627, ZN
                           => n636);
   U698 : AOI22_X1 port map( A1 => n699, A2 => Q(322), B1 => n698, B2 => Q(418)
                           , ZN => n634);
   U699 : AOI22_X1 port map( A1 => n701, A2 => Q(226), B1 => n700, B2 => Q(130)
                           , ZN => n633);
   U700 : AOI22_X1 port map( A1 => n703, A2 => Q(66), B1 => n702, B2 => Q(162),
                           ZN => n632);
   U701 : AOI22_X1 port map( A1 => n705, A2 => Q(194), B1 => n704, B2 => Q(34),
                           ZN => n631);
   U702 : NAND4_X1 port map( A1 => n634, A2 => n633, A3 => n632, A4 => n631, ZN
                           => n635);
   U703 : AOI22_X1 port map( A1 => n674, A2 => Q(1022), B1 => n673, B2 => 
                           Q(958), ZN => n642);
   U704 : AOI22_X1 port map( A1 => n676, A2 => Q(990), B1 => n675, B2 => Q(926)
                           , ZN => n641);
   U705 : AOI22_X1 port map( A1 => n678, A2 => Q(830), B1 => n677, B2 => Q(766)
                           , ZN => n640);
   U706 : NAND2_X1 port map( A1 => n679, A2 => Q(126), ZN => n639);
   U707 : NAND4_X1 port map( A1 => n642, A2 => n641, A3 => n640, A4 => n639, ZN
                           => n658);
   U708 : AOI22_X1 port map( A1 => n681, A2 => Q(862), B1 => n680, B2 => Q(734)
                           , ZN => n646);
   U709 : AOI22_X1 port map( A1 => n683, A2 => Q(798), B1 => n682, B2 => Q(894)
                           , ZN => n645);
   U710 : AOI22_X1 port map( A1 => n685, A2 => Q(702), B1 => n684, B2 => Q(606)
                           , ZN => n644);
   U711 : AOI22_X1 port map( A1 => n687, A2 => Q(542), B1 => n686, B2 => Q(638)
                           , ZN => n643);
   U712 : NAND4_X1 port map( A1 => n646, A2 => n645, A3 => n644, A4 => n643, ZN
                           => n657);
   U713 : AOI22_X1 port map( A1 => n691, A2 => Q(510), B1 => n690, B2 => Q(574)
                           , ZN => n650);
   U714 : AOI22_X1 port map( A1 => n693, A2 => Q(670), B1 => n692, B2 => Q(478)
                           , ZN => n649);
   U715 : AOI22_X1 port map( A1 => n695, A2 => Q(382), B1 => n694, B2 => Q(318)
                           , ZN => n648);
   U716 : AOI22_X1 port map( A1 => n697, A2 => Q(414), B1 => n696, B2 => Q(286)
                           , ZN => n647);
   U717 : NAND4_X1 port map( A1 => n650, A2 => n649, A3 => n648, A4 => n647, ZN
                           => n656);
   U718 : AOI22_X1 port map( A1 => n699, A2 => Q(350), B1 => n698, B2 => Q(446)
                           , ZN => n654);
   U719 : AOI22_X1 port map( A1 => n701, A2 => Q(254), B1 => n700, B2 => Q(158)
                           , ZN => n653);
   U720 : AOI22_X1 port map( A1 => n703, A2 => Q(94), B1 => n702, B2 => Q(190),
                           ZN => n652);
   U721 : AOI22_X1 port map( A1 => n705, A2 => Q(222), B1 => n704, B2 => Q(62),
                           ZN => n651);
   U722 : NAND4_X1 port map( A1 => n654, A2 => n653, A3 => n652, A4 => n651, ZN
                           => n655);
   U723 : AOI22_X1 port map( A1 => n251, A2 => Q(703), B1 => n250, B2 => Q(607)
                           , ZN => n660);
   U724 : AOI22_X1 port map( A1 => n253, A2 => Q(543), B1 => n252, B2 => Q(639)
                           , ZN => n659);
   U725 : AOI22_X1 port map( A1 => n251, A2 => Q(675), B1 => n250, B2 => Q(579)
                           , ZN => n662);
   U726 : AOI22_X1 port map( A1 => n253, A2 => Q(515), B1 => n252, B2 => Q(611)
                           , ZN => n661);
   U727 : AOI22_X1 port map( A1 => n251, A2 => Q(676), B1 => n250, B2 => Q(580)
                           , ZN => n664);
   U728 : AOI22_X1 port map( A1 => n253, A2 => Q(516), B1 => n252, B2 => Q(612)
                           , ZN => n663);
   U729 : AOI22_X1 port map( A1 => n251, A2 => Q(677), B1 => n250, B2 => Q(581)
                           , ZN => n666);
   U730 : AOI22_X1 port map( A1 => n253, A2 => Q(517), B1 => n252, B2 => Q(613)
                           , ZN => n665);
   U731 : AOI22_X1 port map( A1 => n251, A2 => Q(678), B1 => n250, B2 => Q(582)
                           , ZN => n668);
   U732 : AOI22_X1 port map( A1 => n253, A2 => Q(518), B1 => n252, B2 => Q(614)
                           , ZN => n667);
   U733 : AOI22_X1 port map( A1 => n251, A2 => Q(679), B1 => n250, B2 => Q(583)
                           , ZN => n670);
   U734 : AOI22_X1 port map( A1 => n253, A2 => Q(519), B1 => n252, B2 => Q(615)
                           , ZN => n669);
   U735 : AOI22_X1 port map( A1 => n251, A2 => Q(680), B1 => n250, B2 => Q(584)
                           , ZN => n672);
   U736 : AOI22_X1 port map( A1 => n253, A2 => Q(520), B1 => n252, B2 => Q(616)
                           , ZN => n671);
   U737 : AOI22_X1 port map( A1 => n251, A2 => Q(681), B1 => n250, B2 => Q(585)
                           , ZN => n689);
   U738 : AOI22_X1 port map( A1 => n253, A2 => Q(521), B1 => n252, B2 => Q(617)
                           , ZN => n688);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32.all;

entity in_loc_selblock_NBIT_DATA32_N8_F5 is

   port( regs : in std_logic_vector (2559 downto 0);  win : in std_logic_vector
         (4 downto 0);  curr_proc_regs : out std_logic_vector (511 downto 0));

end in_loc_selblock_NBIT_DATA32_N8_F5;

architecture SYN_behav of in_loc_selblock_NBIT_DATA32_N8_F5 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
      n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, 
      n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, 
      n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
      n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
      n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601 : std_logic
      ;

begin
   
   U2 : CLKBUF_X3 port map( A => n1595, Z => n3);
   U3 : BUF_X4 port map( A => n21, Z => n23);
   U4 : BUF_X4 port map( A => n31, Z => n29);
   U5 : CLKBUF_X3 port map( A => n26, Z => n21);
   U6 : BUF_X4 port map( A => n33, Z => n31);
   U7 : CLKBUF_X3 port map( A => n33, Z => n30);
   U8 : CLKBUF_X3 port map( A => n20, Z => n19);
   U9 : BUF_X4 port map( A => n1595, Z => n16);
   U10 : BUF_X2 port map( A => n4, Z => n1);
   U11 : BUF_X4 port map( A => n35, Z => n42);
   U12 : BUF_X4 port map( A => n1597, Z => n2);
   U13 : BUF_X1 port map( A => n44, Z => n5);
   U14 : BUF_X1 port map( A => n44, Z => n6);
   U15 : BUF_X1 port map( A => n55, Z => n8);
   U16 : BUF_X1 port map( A => n53, Z => n7);
   U17 : CLKBUF_X3 port map( A => n19, Z => n26);
   U18 : BUF_X2 port map( A => n3, Z => n13);
   U19 : BUF_X2 port map( A => n3, Z => n15);
   U20 : CLKBUF_X3 port map( A => n1598, Z => n36);
   U21 : BUF_X2 port map( A => n1595, Z => n14);
   U22 : CLKBUF_X3 port map( A => n1597, Z => n33);
   U23 : CLKBUF_X3 port map( A => n1598, Z => n40);
   U24 : CLKBUF_X3 port map( A => n1598, Z => n35);
   U25 : BUF_X2 port map( A => n1595, Z => n4);
   U26 : BUF_X2 port map( A => n56, Z => n57);
   U27 : CLKBUF_X3 port map( A => n1598, Z => n38);
   U28 : BUF_X1 port map( A => n4, Z => n9);
   U29 : BUF_X1 port map( A => n21, Z => n25);
   U30 : BUF_X1 port map( A => n13, Z => n12);
   U31 : BUF_X1 port map( A => n4, Z => n11);
   U32 : BUF_X1 port map( A => n23, Z => n22);
   U33 : BUF_X1 port map( A => n2, Z => n32);
   U34 : BUF_X1 port map( A => n38, Z => n34);
   U35 : BUF_X1 port map( A => n15, Z => n10);
   U36 : BUF_X1 port map( A => n38, Z => n37);
   U37 : BUF_X1 port map( A => n40, Z => n41);
   U38 : NOR2_X1 port map( A1 => n45, A2 => n61, ZN => n1598);
   U39 : AND2_X1 port map( A1 => n59, A2 => win(1), ZN => n1595);
   U40 : BUF_X2 port map( A => n1597, Z => n27);
   U41 : BUF_X2 port map( A => n1598, Z => n39);
   U42 : BUF_X2 port map( A => n1596, Z => n20);
   U43 : BUF_X1 port map( A => n53, Z => n56);
   U44 : BUF_X1 port map( A => win(4), Z => n55);
   U45 : BUF_X1 port map( A => win(4), Z => n48);
   U46 : BUF_X1 port map( A => n52, Z => n50);
   U47 : BUF_X1 port map( A => n44, Z => n47);
   U48 : BUF_X1 port map( A => n52, Z => n45);
   U49 : BUF_X1 port map( A => n44, Z => n51);
   U50 : BUF_X1 port map( A => n44, Z => n53);
   U51 : BUF_X1 port map( A => win(4), Z => n54);
   U52 : BUF_X1 port map( A => n50, Z => n43);
   U53 : BUF_X1 port map( A => win(4), Z => n44);
   U54 : BUF_X1 port map( A => win(4), Z => n49);
   U55 : BUF_X1 port map( A => n55, Z => n46);
   U56 : BUF_X1 port map( A => win(4), Z => n52);
   U57 : BUF_X1 port map( A => n1596, Z => n17);
   U58 : BUF_X1 port map( A => n1596, Z => n18);
   U59 : BUF_X1 port map( A => n1596, Z => n24);
   U60 : BUF_X1 port map( A => n1597, Z => n28);
   U61 : NOR3_X1 port map( A1 => win(2), A2 => win(3), A3 => n46, ZN => n59);
   U62 : INV_X1 port map( A => win(1), ZN => n58);
   U63 : AND3_X1 port map( A1 => n59, A2 => win(0), A3 => n58, ZN => n1596);
   U64 : NAND2_X1 port map( A1 => regs(0), A2 => n17, ZN => n64);
   U65 : INV_X1 port map( A => win(2), ZN => n60);
   U66 : NOR3_X1 port map( A1 => win(3), A2 => n57, A3 => n60, ZN => n1597);
   U67 : AOI22_X1 port map( A1 => n10, A2 => regs(512), B1 => n33, B2 => 
                           regs(1024), ZN => n63);
   U68 : INV_X1 port map( A => win(3), ZN => n61);
   U69 : AOI22_X1 port map( A1 => win(4), A2 => regs(2048), B1 => n34, B2 => 
                           regs(1536), ZN => n62);
   U70 : NAND3_X1 port map( A1 => n64, A2 => n63, A3 => n62, ZN => 
                           curr_proc_regs(0));
   U71 : NAND2_X1 port map( A1 => regs(612), A2 => n1595, ZN => n67);
   U72 : AOI22_X1 port map( A1 => n27, A2 => regs(1124), B1 => n17, B2 => 
                           regs(100), ZN => n66);
   U73 : AOI22_X1 port map( A1 => n54, A2 => regs(2148), B1 => n34, B2 => 
                           regs(1636), ZN => n65);
   U74 : NAND3_X1 port map( A1 => n67, A2 => n66, A3 => n65, ZN => 
                           curr_proc_regs(100));
   U75 : NAND2_X1 port map( A1 => regs(613), A2 => n10, ZN => n70);
   U76 : AOI22_X1 port map( A1 => n29, A2 => regs(1125), B1 => n17, B2 => 
                           regs(101), ZN => n69);
   U77 : AOI22_X1 port map( A1 => n54, A2 => regs(2149), B1 => n34, B2 => 
                           regs(1637), ZN => n68);
   U78 : NAND3_X1 port map( A1 => n70, A2 => n69, A3 => n68, ZN => 
                           curr_proc_regs(101));
   U79 : NAND2_X1 port map( A1 => regs(614), A2 => n12, ZN => n73);
   U80 : AOI22_X1 port map( A1 => n30, A2 => regs(1126), B1 => n17, B2 => 
                           regs(102), ZN => n72);
   U81 : AOI22_X1 port map( A1 => n54, A2 => regs(2150), B1 => n34, B2 => 
                           regs(1638), ZN => n71);
   U82 : NAND3_X1 port map( A1 => n73, A2 => n72, A3 => n71, ZN => 
                           curr_proc_regs(102));
   U83 : NAND2_X1 port map( A1 => regs(615), A2 => n16, ZN => n76);
   U84 : AOI22_X1 port map( A1 => n33, A2 => regs(1127), B1 => n17, B2 => 
                           regs(103), ZN => n75);
   U85 : AOI22_X1 port map( A1 => n54, A2 => regs(2151), B1 => n34, B2 => 
                           regs(1639), ZN => n74);
   U86 : NAND3_X1 port map( A1 => n76, A2 => n75, A3 => n74, ZN => 
                           curr_proc_regs(103));
   U87 : NAND2_X1 port map( A1 => regs(616), A2 => n9, ZN => n79);
   U88 : AOI22_X1 port map( A1 => n30, A2 => regs(1128), B1 => n17, B2 => 
                           regs(104), ZN => n78);
   U89 : AOI22_X1 port map( A1 => n54, A2 => regs(2152), B1 => n34, B2 => 
                           regs(1640), ZN => n77);
   U90 : NAND3_X1 port map( A1 => n79, A2 => n78, A3 => n77, ZN => 
                           curr_proc_regs(104));
   U91 : NAND2_X1 port map( A1 => regs(617), A2 => n11, ZN => n82);
   U92 : AOI22_X1 port map( A1 => n33, A2 => regs(1129), B1 => n17, B2 => 
                           regs(105), ZN => n81);
   U93 : AOI22_X1 port map( A1 => n54, A2 => regs(2153), B1 => n34, B2 => 
                           regs(1641), ZN => n80);
   U94 : NAND3_X1 port map( A1 => n82, A2 => n81, A3 => n80, ZN => 
                           curr_proc_regs(105));
   U95 : NAND2_X1 port map( A1 => regs(618), A2 => n1595, ZN => n85);
   U96 : AOI22_X1 port map( A1 => n27, A2 => regs(1130), B1 => n17, B2 => 
                           regs(106), ZN => n84);
   U97 : AOI22_X1 port map( A1 => n54, A2 => regs(2154), B1 => n34, B2 => 
                           regs(1642), ZN => n83);
   U98 : NAND3_X1 port map( A1 => n85, A2 => n84, A3 => n83, ZN => 
                           curr_proc_regs(106));
   U99 : NAND2_X1 port map( A1 => regs(619), A2 => n10, ZN => n88);
   U100 : AOI22_X1 port map( A1 => n27, A2 => regs(1131), B1 => n17, B2 => 
                           regs(107), ZN => n87);
   U101 : AOI22_X1 port map( A1 => n54, A2 => regs(2155), B1 => n34, B2 => 
                           regs(1643), ZN => n86);
   U102 : NAND3_X1 port map( A1 => n88, A2 => n87, A3 => n86, ZN => 
                           curr_proc_regs(107));
   U103 : NAND2_X1 port map( A1 => regs(620), A2 => n12, ZN => n91);
   U104 : AOI22_X1 port map( A1 => n33, A2 => regs(1132), B1 => n17, B2 => 
                           regs(108), ZN => n90);
   U105 : AOI22_X1 port map( A1 => n54, A2 => regs(2156), B1 => n34, B2 => 
                           regs(1644), ZN => n89);
   U106 : NAND3_X1 port map( A1 => n91, A2 => n90, A3 => n89, ZN => 
                           curr_proc_regs(108));
   U107 : NAND2_X1 port map( A1 => regs(621), A2 => n16, ZN => n94);
   U108 : AOI22_X1 port map( A1 => n30, A2 => regs(1133), B1 => n17, B2 => 
                           regs(109), ZN => n93);
   U109 : AOI22_X1 port map( A1 => n54, A2 => regs(2157), B1 => n34, B2 => 
                           regs(1645), ZN => n92);
   U110 : NAND3_X1 port map( A1 => n94, A2 => n93, A3 => n92, ZN => 
                           curr_proc_regs(109));
   U111 : NAND2_X1 port map( A1 => regs(522), A2 => n9, ZN => n97);
   U112 : AOI22_X1 port map( A1 => n33, A2 => regs(1034), B1 => n17, B2 => 
                           regs(10), ZN => n96);
   U113 : AOI22_X1 port map( A1 => n54, A2 => regs(2058), B1 => n34, B2 => 
                           regs(1546), ZN => n95);
   U114 : NAND3_X1 port map( A1 => n97, A2 => n96, A3 => n95, ZN => 
                           curr_proc_regs(10));
   U115 : NAND2_X1 port map( A1 => regs(622), A2 => n3, ZN => n100);
   U116 : AOI22_X1 port map( A1 => n27, A2 => regs(1134), B1 => n19, B2 => 
                           regs(110), ZN => n99);
   U117 : AOI22_X1 port map( A1 => n54, A2 => regs(2158), B1 => n35, B2 => 
                           regs(1646), ZN => n98);
   U118 : NAND3_X1 port map( A1 => n100, A2 => n99, A3 => n98, ZN => 
                           curr_proc_regs(110));
   U119 : NAND2_X1 port map( A1 => regs(623), A2 => n3, ZN => n103);
   U120 : AOI22_X1 port map( A1 => n33, A2 => regs(1135), B1 => n21, B2 => 
                           regs(111), ZN => n102);
   U121 : AOI22_X1 port map( A1 => n53, A2 => regs(2159), B1 => n35, B2 => 
                           regs(1647), ZN => n101);
   U122 : NAND3_X1 port map( A1 => n103, A2 => n102, A3 => n101, ZN => 
                           curr_proc_regs(111));
   U123 : NAND2_X1 port map( A1 => regs(624), A2 => n3, ZN => n106);
   U124 : AOI22_X1 port map( A1 => n27, A2 => regs(1136), B1 => n19, B2 => 
                           regs(112), ZN => n105);
   U125 : AOI22_X1 port map( A1 => n55, A2 => regs(2160), B1 => n35, B2 => 
                           regs(1648), ZN => n104);
   U126 : NAND3_X1 port map( A1 => n106, A2 => n105, A3 => n104, ZN => 
                           curr_proc_regs(112));
   U127 : NAND2_X1 port map( A1 => regs(625), A2 => n3, ZN => n109);
   U128 : AOI22_X1 port map( A1 => n33, A2 => regs(1137), B1 => n21, B2 => 
                           regs(113), ZN => n108);
   U129 : AOI22_X1 port map( A1 => n52, A2 => regs(2161), B1 => n35, B2 => 
                           regs(1649), ZN => n107);
   U130 : NAND3_X1 port map( A1 => n109, A2 => n108, A3 => n107, ZN => 
                           curr_proc_regs(113));
   U131 : NAND2_X1 port map( A1 => regs(626), A2 => n3, ZN => n112);
   U132 : AOI22_X1 port map( A1 => n33, A2 => regs(1138), B1 => n19, B2 => 
                           regs(114), ZN => n111);
   U133 : AOI22_X1 port map( A1 => win(4), A2 => regs(2162), B1 => n35, B2 => 
                           regs(1650), ZN => n110);
   U134 : NAND3_X1 port map( A1 => n112, A2 => n111, A3 => n110, ZN => 
                           curr_proc_regs(114));
   U135 : NAND2_X1 port map( A1 => regs(627), A2 => n3, ZN => n115);
   U136 : AOI22_X1 port map( A1 => n29, A2 => regs(1139), B1 => n21, B2 => 
                           regs(115), ZN => n114);
   U137 : AOI22_X1 port map( A1 => n56, A2 => regs(2163), B1 => n35, B2 => 
                           regs(1651), ZN => n113);
   U138 : NAND3_X1 port map( A1 => n115, A2 => n114, A3 => n113, ZN => 
                           curr_proc_regs(115));
   U139 : NAND2_X1 port map( A1 => regs(628), A2 => n3, ZN => n118);
   U140 : AOI22_X1 port map( A1 => n30, A2 => regs(1140), B1 => n26, B2 => 
                           regs(116), ZN => n117);
   U141 : AOI22_X1 port map( A1 => n43, A2 => regs(2164), B1 => n35, B2 => 
                           regs(1652), ZN => n116);
   U142 : NAND3_X1 port map( A1 => n118, A2 => n117, A3 => n116, ZN => 
                           curr_proc_regs(116));
   U143 : NAND2_X1 port map( A1 => regs(629), A2 => n3, ZN => n121);
   U144 : AOI22_X1 port map( A1 => n29, A2 => regs(1141), B1 => n19, B2 => 
                           regs(117), ZN => n120);
   U145 : AOI22_X1 port map( A1 => n45, A2 => regs(2165), B1 => n35, B2 => 
                           regs(1653), ZN => n119);
   U146 : NAND3_X1 port map( A1 => n121, A2 => n120, A3 => n119, ZN => 
                           curr_proc_regs(117));
   U147 : NAND2_X1 port map( A1 => regs(630), A2 => n3, ZN => n124);
   U148 : AOI22_X1 port map( A1 => n33, A2 => regs(1142), B1 => n1596, B2 => 
                           regs(118), ZN => n123);
   U149 : AOI22_X1 port map( A1 => n49, A2 => regs(2166), B1 => n35, B2 => 
                           regs(1654), ZN => n122);
   U150 : NAND3_X1 port map( A1 => n124, A2 => n123, A3 => n122, ZN => 
                           curr_proc_regs(118));
   U151 : NAND2_X1 port map( A1 => regs(631), A2 => n3, ZN => n127);
   U152 : AOI22_X1 port map( A1 => n33, A2 => regs(1143), B1 => n21, B2 => 
                           regs(119), ZN => n126);
   U153 : AOI22_X1 port map( A1 => n48, A2 => regs(2167), B1 => n35, B2 => 
                           regs(1655), ZN => n125);
   U154 : NAND3_X1 port map( A1 => n127, A2 => n126, A3 => n125, ZN => 
                           curr_proc_regs(119));
   U155 : NAND2_X1 port map( A1 => regs(523), A2 => n3, ZN => n130);
   U156 : AOI22_X1 port map( A1 => n33, A2 => regs(1035), B1 => n17, B2 => 
                           regs(11), ZN => n129);
   U157 : AOI22_X1 port map( A1 => n54, A2 => regs(2059), B1 => n35, B2 => 
                           regs(1547), ZN => n128);
   U158 : NAND3_X1 port map( A1 => n130, A2 => n129, A3 => n128, ZN => 
                           curr_proc_regs(11));
   U159 : NAND2_X1 port map( A1 => regs(632), A2 => n3, ZN => n133);
   U160 : AOI22_X1 port map( A1 => n33, A2 => regs(1144), B1 => n26, B2 => 
                           regs(120), ZN => n132);
   U161 : AOI22_X1 port map( A1 => n51, A2 => regs(2168), B1 => n35, B2 => 
                           regs(1656), ZN => n131);
   U162 : NAND3_X1 port map( A1 => n133, A2 => n132, A3 => n131, ZN => 
                           curr_proc_regs(120));
   U163 : NAND2_X1 port map( A1 => regs(633), A2 => n16, ZN => n136);
   U164 : AOI22_X1 port map( A1 => n27, A2 => regs(1145), B1 => n23, B2 => 
                           regs(121), ZN => n135);
   U165 : AOI22_X1 port map( A1 => win(4), A2 => regs(2169), B1 => n35, B2 => 
                           regs(1657), ZN => n134);
   U166 : NAND3_X1 port map( A1 => n136, A2 => n135, A3 => n134, ZN => 
                           curr_proc_regs(121));
   U167 : NAND2_X1 port map( A1 => regs(634), A2 => n9, ZN => n139);
   U168 : AOI22_X1 port map( A1 => n27, A2 => regs(1146), B1 => n23, B2 => 
                           regs(122), ZN => n138);
   U169 : AOI22_X1 port map( A1 => n6, A2 => regs(2170), B1 => n40, B2 => 
                           regs(1658), ZN => n137);
   U170 : NAND3_X1 port map( A1 => n139, A2 => n138, A3 => n137, ZN => 
                           curr_proc_regs(122));
   U171 : NAND2_X1 port map( A1 => regs(635), A2 => n11, ZN => n142);
   U172 : AOI22_X1 port map( A1 => n33, A2 => regs(1147), B1 => n23, B2 => 
                           regs(123), ZN => n141);
   U173 : AOI22_X1 port map( A1 => n6, A2 => regs(2171), B1 => n36, B2 => 
                           regs(1659), ZN => n140);
   U174 : NAND3_X1 port map( A1 => n142, A2 => n141, A3 => n140, ZN => 
                           curr_proc_regs(123));
   U175 : NAND2_X1 port map( A1 => regs(636), A2 => n11, ZN => n145);
   U176 : AOI22_X1 port map( A1 => n33, A2 => regs(1148), B1 => n23, B2 => 
                           regs(124), ZN => n144);
   U177 : AOI22_X1 port map( A1 => n6, A2 => regs(2172), B1 => n35, B2 => 
                           regs(1660), ZN => n143);
   U178 : NAND3_X1 port map( A1 => n145, A2 => n144, A3 => n143, ZN => 
                           curr_proc_regs(124));
   U179 : NAND2_X1 port map( A1 => regs(637), A2 => n1595, ZN => n148);
   U180 : AOI22_X1 port map( A1 => n29, A2 => regs(1149), B1 => n23, B2 => 
                           regs(125), ZN => n147);
   U181 : AOI22_X1 port map( A1 => n6, A2 => regs(2173), B1 => n40, B2 => 
                           regs(1661), ZN => n146);
   U182 : NAND3_X1 port map( A1 => n148, A2 => n147, A3 => n146, ZN => 
                           curr_proc_regs(125));
   U183 : NAND2_X1 port map( A1 => regs(638), A2 => n10, ZN => n151);
   U184 : AOI22_X1 port map( A1 => n27, A2 => regs(1150), B1 => n23, B2 => 
                           regs(126), ZN => n150);
   U185 : AOI22_X1 port map( A1 => n6, A2 => regs(2174), B1 => n36, B2 => 
                           regs(1662), ZN => n149);
   U186 : NAND3_X1 port map( A1 => n151, A2 => n150, A3 => n149, ZN => 
                           curr_proc_regs(126));
   U187 : NAND2_X1 port map( A1 => regs(639), A2 => n12, ZN => n154);
   U188 : AOI22_X1 port map( A1 => n30, A2 => regs(1151), B1 => n23, B2 => 
                           regs(127), ZN => n153);
   U189 : AOI22_X1 port map( A1 => n6, A2 => regs(2175), B1 => n35, B2 => 
                           regs(1663), ZN => n152);
   U190 : NAND3_X1 port map( A1 => n154, A2 => n153, A3 => n152, ZN => 
                           curr_proc_regs(127));
   U191 : NAND2_X1 port map( A1 => regs(640), A2 => n16, ZN => n157);
   U192 : AOI22_X1 port map( A1 => n33, A2 => regs(1152), B1 => n23, B2 => 
                           regs(128), ZN => n156);
   U193 : AOI22_X1 port map( A1 => n6, A2 => regs(2176), B1 => n40, B2 => 
                           regs(1664), ZN => n155);
   U194 : NAND3_X1 port map( A1 => n157, A2 => n156, A3 => n155, ZN => 
                           curr_proc_regs(128));
   U195 : NAND2_X1 port map( A1 => regs(641), A2 => n9, ZN => n160);
   U196 : AOI22_X1 port map( A1 => n31, A2 => regs(1153), B1 => n23, B2 => 
                           regs(129), ZN => n159);
   U197 : AOI22_X1 port map( A1 => n6, A2 => regs(2177), B1 => n36, B2 => 
                           regs(1665), ZN => n158);
   U198 : NAND3_X1 port map( A1 => n160, A2 => n159, A3 => n158, ZN => 
                           curr_proc_regs(129));
   U199 : NAND2_X1 port map( A1 => regs(524), A2 => n11, ZN => n163);
   U200 : AOI22_X1 port map( A1 => n33, A2 => regs(1036), B1 => n23, B2 => 
                           regs(12), ZN => n162);
   U201 : AOI22_X1 port map( A1 => n6, A2 => regs(2060), B1 => n35, B2 => 
                           regs(1548), ZN => n161);
   U202 : NAND3_X1 port map( A1 => n163, A2 => n162, A3 => n161, ZN => 
                           curr_proc_regs(12));
   U203 : NAND2_X1 port map( A1 => regs(642), A2 => n1595, ZN => n166);
   U204 : AOI22_X1 port map( A1 => n31, A2 => regs(1154), B1 => n23, B2 => 
                           regs(130), ZN => n165);
   U205 : AOI22_X1 port map( A1 => n6, A2 => regs(2178), B1 => n40, B2 => 
                           regs(1666), ZN => n164);
   U206 : NAND3_X1 port map( A1 => n166, A2 => n165, A3 => n164, ZN => 
                           curr_proc_regs(130));
   U207 : NAND2_X1 port map( A1 => regs(643), A2 => n12, ZN => n169);
   U208 : AOI22_X1 port map( A1 => n2, A2 => regs(1155), B1 => n23, B2 => 
                           regs(131), ZN => n168);
   U209 : AOI22_X1 port map( A1 => n6, A2 => regs(2179), B1 => n36, B2 => 
                           regs(1667), ZN => n167);
   U210 : NAND3_X1 port map( A1 => n169, A2 => n168, A3 => n167, ZN => 
                           curr_proc_regs(131));
   U211 : NAND2_X1 port map( A1 => regs(644), A2 => n16, ZN => n172);
   U212 : AOI22_X1 port map( A1 => n33, A2 => regs(1156), B1 => n18, B2 => 
                           regs(132), ZN => n171);
   U213 : AOI22_X1 port map( A1 => n6, A2 => regs(2180), B1 => n42, B2 => 
                           regs(1668), ZN => n170);
   U214 : NAND3_X1 port map( A1 => n172, A2 => n171, A3 => n170, ZN => 
                           curr_proc_regs(132));
   U215 : NAND2_X1 port map( A1 => regs(645), A2 => n16, ZN => n175);
   U216 : AOI22_X1 port map( A1 => n27, A2 => regs(1157), B1 => n18, B2 => 
                           regs(133), ZN => n174);
   U217 : AOI22_X1 port map( A1 => n48, A2 => regs(2181), B1 => n35, B2 => 
                           regs(1669), ZN => n173);
   U218 : NAND3_X1 port map( A1 => n175, A2 => n174, A3 => n173, ZN => 
                           curr_proc_regs(133));
   U219 : NAND2_X1 port map( A1 => regs(646), A2 => n16, ZN => n178);
   U220 : AOI22_X1 port map( A1 => n29, A2 => regs(1158), B1 => n18, B2 => 
                           regs(134), ZN => n177);
   U221 : AOI22_X1 port map( A1 => n54, A2 => regs(2182), B1 => n34, B2 => 
                           regs(1670), ZN => n176);
   U222 : NAND3_X1 port map( A1 => n178, A2 => n177, A3 => n176, ZN => 
                           curr_proc_regs(134));
   U223 : NAND2_X1 port map( A1 => regs(647), A2 => n16, ZN => n181);
   U224 : AOI22_X1 port map( A1 => n33, A2 => regs(1159), B1 => n18, B2 => 
                           regs(135), ZN => n180);
   U225 : AOI22_X1 port map( A1 => n51, A2 => regs(2183), B1 => n37, B2 => 
                           regs(1671), ZN => n179);
   U226 : NAND3_X1 port map( A1 => n181, A2 => n180, A3 => n179, ZN => 
                           curr_proc_regs(135));
   U227 : NAND2_X1 port map( A1 => regs(648), A2 => n16, ZN => n184);
   U228 : AOI22_X1 port map( A1 => n27, A2 => regs(1160), B1 => n18, B2 => 
                           regs(136), ZN => n183);
   U229 : AOI22_X1 port map( A1 => n47, A2 => regs(2184), B1 => n42, B2 => 
                           regs(1672), ZN => n182);
   U230 : NAND3_X1 port map( A1 => n184, A2 => n183, A3 => n182, ZN => 
                           curr_proc_regs(136));
   U231 : NAND2_X1 port map( A1 => regs(649), A2 => n16, ZN => n187);
   U232 : AOI22_X1 port map( A1 => n30, A2 => regs(1161), B1 => n18, B2 => 
                           regs(137), ZN => n186);
   U233 : AOI22_X1 port map( A1 => n46, A2 => regs(2185), B1 => n40, B2 => 
                           regs(1673), ZN => n185);
   U234 : NAND3_X1 port map( A1 => n187, A2 => n186, A3 => n185, ZN => 
                           curr_proc_regs(137));
   U235 : NAND2_X1 port map( A1 => regs(650), A2 => n16, ZN => n190);
   U236 : AOI22_X1 port map( A1 => n33, A2 => regs(1162), B1 => n18, B2 => 
                           regs(138), ZN => n189);
   U237 : AOI22_X1 port map( A1 => n50, A2 => regs(2186), B1 => n34, B2 => 
                           regs(1674), ZN => n188);
   U238 : NAND3_X1 port map( A1 => n190, A2 => n189, A3 => n188, ZN => 
                           curr_proc_regs(138));
   U239 : NAND2_X1 port map( A1 => regs(651), A2 => n16, ZN => n193);
   U240 : AOI22_X1 port map( A1 => n27, A2 => regs(1163), B1 => n18, B2 => 
                           regs(139), ZN => n192);
   U241 : AOI22_X1 port map( A1 => n53, A2 => regs(2187), B1 => n37, B2 => 
                           regs(1675), ZN => n191);
   U242 : NAND3_X1 port map( A1 => n193, A2 => n192, A3 => n191, ZN => 
                           curr_proc_regs(139));
   U243 : NAND2_X1 port map( A1 => regs(525), A2 => n16, ZN => n196);
   U244 : AOI22_X1 port map( A1 => n33, A2 => regs(1037), B1 => n18, B2 => 
                           regs(13), ZN => n195);
   U245 : AOI22_X1 port map( A1 => n55, A2 => regs(2061), B1 => n42, B2 => 
                           regs(1549), ZN => n194);
   U246 : NAND3_X1 port map( A1 => n196, A2 => n195, A3 => n194, ZN => 
                           curr_proc_regs(13));
   U247 : NAND2_X1 port map( A1 => regs(652), A2 => n16, ZN => n199);
   U248 : AOI22_X1 port map( A1 => n30, A2 => regs(1164), B1 => n18, B2 => 
                           regs(140), ZN => n198);
   U249 : AOI22_X1 port map( A1 => n52, A2 => regs(2188), B1 => n36, B2 => 
                           regs(1676), ZN => n197);
   U250 : NAND3_X1 port map( A1 => n199, A2 => n198, A3 => n197, ZN => 
                           curr_proc_regs(140));
   U251 : NAND2_X1 port map( A1 => regs(653), A2 => n16, ZN => n202);
   U252 : AOI22_X1 port map( A1 => n33, A2 => regs(1165), B1 => n18, B2 => 
                           regs(141), ZN => n201);
   U253 : AOI22_X1 port map( A1 => win(4), A2 => regs(2189), B1 => n34, B2 => 
                           regs(1677), ZN => n200);
   U254 : NAND3_X1 port map( A1 => n202, A2 => n201, A3 => n200, ZN => 
                           curr_proc_regs(141));
   U255 : NAND2_X1 port map( A1 => regs(654), A2 => n16, ZN => n205);
   U256 : AOI22_X1 port map( A1 => n29, A2 => regs(1166), B1 => n18, B2 => 
                           regs(142), ZN => n204);
   U257 : AOI22_X1 port map( A1 => n56, A2 => regs(2190), B1 => n37, B2 => 
                           regs(1678), ZN => n203);
   U258 : NAND3_X1 port map( A1 => n205, A2 => n204, A3 => n203, ZN => 
                           curr_proc_regs(142));
   U259 : NAND2_X1 port map( A1 => regs(655), A2 => n16, ZN => n208);
   U260 : AOI22_X1 port map( A1 => n33, A2 => regs(1167), B1 => n20, B2 => 
                           regs(143), ZN => n207);
   U261 : AOI22_X1 port map( A1 => win(4), A2 => regs(2191), B1 => n34, B2 => 
                           regs(1679), ZN => n206);
   U262 : NAND3_X1 port map( A1 => n208, A2 => n207, A3 => n206, ZN => 
                           curr_proc_regs(143));
   U263 : NAND2_X1 port map( A1 => regs(656), A2 => n16, ZN => n211);
   U264 : AOI22_X1 port map( A1 => n27, A2 => regs(1168), B1 => n20, B2 => 
                           regs(144), ZN => n210);
   U265 : AOI22_X1 port map( A1 => n47, A2 => regs(2192), B1 => n37, B2 => 
                           regs(1680), ZN => n209);
   U266 : NAND3_X1 port map( A1 => n211, A2 => n210, A3 => n209, ZN => 
                           curr_proc_regs(144));
   U267 : NAND2_X1 port map( A1 => regs(657), A2 => n16, ZN => n214);
   U268 : AOI22_X1 port map( A1 => n33, A2 => regs(1169), B1 => n20, B2 => 
                           regs(145), ZN => n213);
   U269 : AOI22_X1 port map( A1 => n51, A2 => regs(2193), B1 => n38, B2 => 
                           regs(1681), ZN => n212);
   U270 : NAND3_X1 port map( A1 => n214, A2 => n213, A3 => n212, ZN => 
                           curr_proc_regs(145));
   U271 : NAND2_X1 port map( A1 => regs(658), A2 => n16, ZN => n217);
   U272 : AOI22_X1 port map( A1 => n28, A2 => regs(1170), B1 => n20, B2 => 
                           regs(146), ZN => n216);
   U273 : AOI22_X1 port map( A1 => n54, A2 => regs(2194), B1 => n38, B2 => 
                           regs(1682), ZN => n215);
   U274 : NAND3_X1 port map( A1 => n217, A2 => n216, A3 => n215, ZN => 
                           curr_proc_regs(146));
   U275 : NAND2_X1 port map( A1 => regs(659), A2 => n16, ZN => n220);
   U276 : AOI22_X1 port map( A1 => n33, A2 => regs(1171), B1 => n20, B2 => 
                           regs(147), ZN => n219);
   U277 : AOI22_X1 port map( A1 => n48, A2 => regs(2195), B1 => n35, B2 => 
                           regs(1683), ZN => n218);
   U278 : NAND3_X1 port map( A1 => n220, A2 => n219, A3 => n218, ZN => 
                           curr_proc_regs(147));
   U279 : NAND2_X1 port map( A1 => regs(660), A2 => n16, ZN => n223);
   U280 : AOI22_X1 port map( A1 => n2, A2 => regs(1172), B1 => n20, B2 => 
                           regs(148), ZN => n222);
   U281 : AOI22_X1 port map( A1 => n49, A2 => regs(2196), B1 => n34, B2 => 
                           regs(1684), ZN => n221);
   U282 : NAND3_X1 port map( A1 => n223, A2 => n222, A3 => n221, ZN => 
                           curr_proc_regs(148));
   U283 : NAND2_X1 port map( A1 => regs(661), A2 => n16, ZN => n226);
   U284 : AOI22_X1 port map( A1 => n33, A2 => regs(1173), B1 => n20, B2 => 
                           regs(149), ZN => n225);
   U285 : AOI22_X1 port map( A1 => n45, A2 => regs(2197), B1 => n37, B2 => 
                           regs(1685), ZN => n224);
   U286 : NAND3_X1 port map( A1 => n226, A2 => n225, A3 => n224, ZN => 
                           curr_proc_regs(149));
   U287 : NAND2_X1 port map( A1 => regs(526), A2 => n16, ZN => n229);
   U288 : AOI22_X1 port map( A1 => n27, A2 => regs(1038), B1 => n20, B2 => 
                           regs(14), ZN => n228);
   U289 : AOI22_X1 port map( A1 => n51, A2 => regs(2062), B1 => n42, B2 => 
                           regs(1550), ZN => n227);
   U290 : NAND3_X1 port map( A1 => n229, A2 => n228, A3 => n227, ZN => 
                           curr_proc_regs(14));
   U291 : NAND2_X1 port map( A1 => regs(662), A2 => n16, ZN => n232);
   U292 : AOI22_X1 port map( A1 => n33, A2 => regs(1174), B1 => n20, B2 => 
                           regs(150), ZN => n231);
   U293 : AOI22_X1 port map( A1 => n52, A2 => regs(2198), B1 => n40, B2 => 
                           regs(1686), ZN => n230);
   U294 : NAND3_X1 port map( A1 => n232, A2 => n231, A3 => n230, ZN => 
                           curr_proc_regs(150));
   U295 : NAND2_X1 port map( A1 => regs(663), A2 => n16, ZN => n235);
   U296 : AOI22_X1 port map( A1 => n33, A2 => regs(1175), B1 => n20, B2 => 
                           regs(151), ZN => n234);
   U297 : AOI22_X1 port map( A1 => n43, A2 => regs(2199), B1 => n36, B2 => 
                           regs(1687), ZN => n233);
   U298 : NAND3_X1 port map( A1 => n235, A2 => n234, A3 => n233, ZN => 
                           curr_proc_regs(151));
   U299 : NAND2_X1 port map( A1 => regs(664), A2 => n16, ZN => n238);
   U300 : AOI22_X1 port map( A1 => n33, A2 => regs(1176), B1 => n20, B2 => 
                           regs(152), ZN => n237);
   U301 : AOI22_X1 port map( A1 => n56, A2 => regs(2200), B1 => n34, B2 => 
                           regs(1688), ZN => n236);
   U302 : NAND3_X1 port map( A1 => n238, A2 => n237, A3 => n236, ZN => 
                           curr_proc_regs(152));
   U303 : NAND2_X1 port map( A1 => regs(665), A2 => n16, ZN => n241);
   U304 : AOI22_X1 port map( A1 => n33, A2 => regs(1177), B1 => n20, B2 => 
                           regs(153), ZN => n240);
   U305 : AOI22_X1 port map( A1 => n52, A2 => regs(2201), B1 => n37, B2 => 
                           regs(1689), ZN => n239);
   U306 : NAND3_X1 port map( A1 => n241, A2 => n240, A3 => n239, ZN => 
                           curr_proc_regs(153));
   U307 : NAND2_X1 port map( A1 => regs(666), A2 => n16, ZN => n244);
   U308 : AOI22_X1 port map( A1 => n33, A2 => regs(1178), B1 => n26, B2 => 
                           regs(154), ZN => n243);
   U309 : AOI22_X1 port map( A1 => n47, A2 => regs(2202), B1 => n36, B2 => 
                           regs(1690), ZN => n242);
   U310 : NAND3_X1 port map( A1 => n244, A2 => n243, A3 => n242, ZN => 
                           curr_proc_regs(154));
   U311 : NAND2_X1 port map( A1 => regs(667), A2 => n16, ZN => n247);
   U312 : AOI22_X1 port map( A1 => n33, A2 => regs(1179), B1 => n19, B2 => 
                           regs(155), ZN => n246);
   U313 : AOI22_X1 port map( A1 => n56, A2 => regs(2203), B1 => n36, B2 => 
                           regs(1691), ZN => n245);
   U314 : NAND3_X1 port map( A1 => n247, A2 => n246, A3 => n245, ZN => 
                           curr_proc_regs(155));
   U315 : NAND2_X1 port map( A1 => regs(668), A2 => n16, ZN => n250);
   U316 : AOI22_X1 port map( A1 => n2, A2 => regs(1180), B1 => n20, B2 => 
                           regs(156), ZN => n249);
   U317 : AOI22_X1 port map( A1 => n49, A2 => regs(2204), B1 => n36, B2 => 
                           regs(1692), ZN => n248);
   U318 : NAND3_X1 port map( A1 => n250, A2 => n249, A3 => n248, ZN => 
                           curr_proc_regs(156));
   U319 : NAND2_X1 port map( A1 => regs(669), A2 => n16, ZN => n253);
   U320 : AOI22_X1 port map( A1 => n33, A2 => regs(1181), B1 => n21, B2 => 
                           regs(157), ZN => n252);
   U321 : AOI22_X1 port map( A1 => n52, A2 => regs(2205), B1 => n36, B2 => 
                           regs(1693), ZN => n251);
   U322 : NAND3_X1 port map( A1 => n253, A2 => n252, A3 => n251, ZN => 
                           curr_proc_regs(157));
   U323 : NAND2_X1 port map( A1 => regs(670), A2 => n16, ZN => n256);
   U324 : AOI22_X1 port map( A1 => n33, A2 => regs(1182), B1 => n21, B2 => 
                           regs(158), ZN => n255);
   U325 : AOI22_X1 port map( A1 => n50, A2 => regs(2206), B1 => n36, B2 => 
                           regs(1694), ZN => n254);
   U326 : NAND3_X1 port map( A1 => n256, A2 => n255, A3 => n254, ZN => 
                           curr_proc_regs(158));
   U327 : NAND2_X1 port map( A1 => regs(671), A2 => n16, ZN => n259);
   U328 : AOI22_X1 port map( A1 => n33, A2 => regs(1183), B1 => n20, B2 => 
                           regs(159), ZN => n258);
   U329 : AOI22_X1 port map( A1 => n53, A2 => regs(2207), B1 => n36, B2 => 
                           regs(1695), ZN => n257);
   U330 : NAND3_X1 port map( A1 => n259, A2 => n258, A3 => n257, ZN => 
                           curr_proc_regs(159));
   U331 : NAND2_X1 port map( A1 => regs(527), A2 => n16, ZN => n262);
   U332 : AOI22_X1 port map( A1 => n27, A2 => regs(1039), B1 => n19, B2 => 
                           regs(15), ZN => n261);
   U333 : AOI22_X1 port map( A1 => n50, A2 => regs(2063), B1 => n36, B2 => 
                           regs(1551), ZN => n260);
   U334 : NAND3_X1 port map( A1 => n262, A2 => n261, A3 => n260, ZN => 
                           curr_proc_regs(15));
   U335 : NAND2_X1 port map( A1 => regs(672), A2 => n16, ZN => n265);
   U336 : AOI22_X1 port map( A1 => n29, A2 => regs(1184), B1 => n26, B2 => 
                           regs(160), ZN => n264);
   U337 : AOI22_X1 port map( A1 => n49, A2 => regs(2208), B1 => n36, B2 => 
                           regs(1696), ZN => n263);
   U338 : NAND3_X1 port map( A1 => n265, A2 => n264, A3 => n263, ZN => 
                           curr_proc_regs(160));
   U339 : NAND2_X1 port map( A1 => regs(673), A2 => n16, ZN => n268);
   U340 : AOI22_X1 port map( A1 => n33, A2 => regs(1185), B1 => n20, B2 => 
                           regs(161), ZN => n267);
   U341 : AOI22_X1 port map( A1 => n53, A2 => regs(2209), B1 => n36, B2 => 
                           regs(1697), ZN => n266);
   U342 : NAND3_X1 port map( A1 => n268, A2 => n267, A3 => n266, ZN => 
                           curr_proc_regs(161));
   U343 : NAND2_X1 port map( A1 => regs(674), A2 => n16, ZN => n271);
   U344 : AOI22_X1 port map( A1 => n33, A2 => regs(1186), B1 => n26, B2 => 
                           regs(162), ZN => n270);
   U345 : AOI22_X1 port map( A1 => n48, A2 => regs(2210), B1 => n36, B2 => 
                           regs(1698), ZN => n269);
   U346 : NAND3_X1 port map( A1 => n271, A2 => n270, A3 => n269, ZN => 
                           curr_proc_regs(162));
   U347 : NAND2_X1 port map( A1 => regs(675), A2 => n16, ZN => n274);
   U348 : AOI22_X1 port map( A1 => n33, A2 => regs(1187), B1 => n19, B2 => 
                           regs(163), ZN => n273);
   U349 : AOI22_X1 port map( A1 => n46, A2 => regs(2211), B1 => n36, B2 => 
                           regs(1699), ZN => n272);
   U350 : NAND3_X1 port map( A1 => n274, A2 => n273, A3 => n272, ZN => 
                           curr_proc_regs(163));
   U351 : NAND2_X1 port map( A1 => regs(676), A2 => n16, ZN => n277);
   U352 : AOI22_X1 port map( A1 => n33, A2 => regs(1188), B1 => n20, B2 => 
                           regs(164), ZN => n276);
   U353 : AOI22_X1 port map( A1 => n54, A2 => regs(2212), B1 => n36, B2 => 
                           regs(1700), ZN => n275);
   U354 : NAND3_X1 port map( A1 => n277, A2 => n276, A3 => n275, ZN => 
                           curr_proc_regs(164));
   U355 : NAND2_X1 port map( A1 => regs(677), A2 => n16, ZN => n280);
   U356 : AOI22_X1 port map( A1 => n33, A2 => regs(1189), B1 => n21, B2 => 
                           regs(165), ZN => n279);
   U357 : AOI22_X1 port map( A1 => n55, A2 => regs(2213), B1 => n40, B2 => 
                           regs(1701), ZN => n278);
   U358 : NAND3_X1 port map( A1 => n280, A2 => n279, A3 => n278, ZN => 
                           curr_proc_regs(165));
   U359 : NAND2_X1 port map( A1 => regs(678), A2 => n16, ZN => n283);
   U360 : AOI22_X1 port map( A1 => n33, A2 => regs(1190), B1 => n21, B2 => 
                           regs(166), ZN => n282);
   U361 : AOI22_X1 port map( A1 => n54, A2 => regs(2214), B1 => n34, B2 => 
                           regs(1702), ZN => n281);
   U362 : NAND3_X1 port map( A1 => n283, A2 => n282, A3 => n281, ZN => 
                           curr_proc_regs(166));
   U363 : NAND2_X1 port map( A1 => regs(679), A2 => n16, ZN => n286);
   U364 : AOI22_X1 port map( A1 => n30, A2 => regs(1191), B1 => n21, B2 => 
                           regs(167), ZN => n285);
   U365 : AOI22_X1 port map( A1 => n48, A2 => regs(2215), B1 => n37, B2 => 
                           regs(1703), ZN => n284);
   U366 : NAND3_X1 port map( A1 => n286, A2 => n285, A3 => n284, ZN => 
                           curr_proc_regs(167));
   U367 : NAND2_X1 port map( A1 => regs(680), A2 => n16, ZN => n289);
   U368 : AOI22_X1 port map( A1 => n29, A2 => regs(1192), B1 => n21, B2 => 
                           regs(168), ZN => n288);
   U369 : AOI22_X1 port map( A1 => n52, A2 => regs(2216), B1 => n38, B2 => 
                           regs(1704), ZN => n287);
   U370 : NAND3_X1 port map( A1 => n289, A2 => n288, A3 => n287, ZN => 
                           curr_proc_regs(168));
   U371 : NAND2_X1 port map( A1 => regs(681), A2 => n16, ZN => n292);
   U372 : AOI22_X1 port map( A1 => n30, A2 => regs(1193), B1 => n21, B2 => 
                           regs(169), ZN => n291);
   U373 : AOI22_X1 port map( A1 => n51, A2 => regs(2217), B1 => n38, B2 => 
                           regs(1705), ZN => n290);
   U374 : NAND3_X1 port map( A1 => n292, A2 => n291, A3 => n290, ZN => 
                           curr_proc_regs(169));
   U375 : NAND2_X1 port map( A1 => regs(528), A2 => n16, ZN => n295);
   U376 : AOI22_X1 port map( A1 => n33, A2 => regs(1040), B1 => n21, B2 => 
                           regs(16), ZN => n294);
   U377 : AOI22_X1 port map( A1 => n49, A2 => regs(2064), B1 => n34, B2 => 
                           regs(1552), ZN => n293);
   U378 : NAND3_X1 port map( A1 => n295, A2 => n294, A3 => n293, ZN => 
                           curr_proc_regs(16));
   U379 : NAND2_X1 port map( A1 => regs(682), A2 => n16, ZN => n298);
   U380 : AOI22_X1 port map( A1 => n29, A2 => regs(1194), B1 => n21, B2 => 
                           regs(170), ZN => n297);
   U381 : AOI22_X1 port map( A1 => n56, A2 => regs(2218), B1 => n36, B2 => 
                           regs(1706), ZN => n296);
   U382 : NAND3_X1 port map( A1 => n298, A2 => n297, A3 => n296, ZN => 
                           curr_proc_regs(170));
   U383 : NAND2_X1 port map( A1 => regs(683), A2 => n16, ZN => n301);
   U384 : AOI22_X1 port map( A1 => n33, A2 => regs(1195), B1 => n21, B2 => 
                           regs(171), ZN => n300);
   U385 : AOI22_X1 port map( A1 => n47, A2 => regs(2219), B1 => n34, B2 => 
                           regs(1707), ZN => n299);
   U386 : NAND3_X1 port map( A1 => n301, A2 => n300, A3 => n299, ZN => 
                           curr_proc_regs(171));
   U387 : NAND2_X1 port map( A1 => regs(684), A2 => n16, ZN => n304);
   U388 : AOI22_X1 port map( A1 => n29, A2 => regs(1196), B1 => n21, B2 => 
                           regs(172), ZN => n303);
   U389 : AOI22_X1 port map( A1 => n45, A2 => regs(2220), B1 => n37, B2 => 
                           regs(1708), ZN => n302);
   U390 : NAND3_X1 port map( A1 => n304, A2 => n303, A3 => n302, ZN => 
                           curr_proc_regs(172));
   U391 : NAND2_X1 port map( A1 => regs(685), A2 => n16, ZN => n307);
   U392 : AOI22_X1 port map( A1 => n33, A2 => regs(1197), B1 => n21, B2 => 
                           regs(173), ZN => n306);
   U393 : AOI22_X1 port map( A1 => n43, A2 => regs(2221), B1 => n38, B2 => 
                           regs(1709), ZN => n305);
   U394 : NAND3_X1 port map( A1 => n307, A2 => n306, A3 => n305, ZN => 
                           curr_proc_regs(173));
   U395 : NAND2_X1 port map( A1 => regs(686), A2 => n16, ZN => n310);
   U396 : AOI22_X1 port map( A1 => n30, A2 => regs(1198), B1 => n21, B2 => 
                           regs(174), ZN => n309);
   U397 : AOI22_X1 port map( A1 => n46, A2 => regs(2222), B1 => n37, B2 => 
                           regs(1710), ZN => n308);
   U398 : NAND3_X1 port map( A1 => n310, A2 => n309, A3 => n308, ZN => 
                           curr_proc_regs(174));
   U399 : NAND2_X1 port map( A1 => regs(687), A2 => n16, ZN => n313);
   U400 : AOI22_X1 port map( A1 => n30, A2 => regs(1199), B1 => n21, B2 => 
                           regs(175), ZN => n312);
   U401 : AOI22_X1 port map( A1 => n43, A2 => regs(2223), B1 => n38, B2 => 
                           regs(1711), ZN => n311);
   U402 : NAND3_X1 port map( A1 => n313, A2 => n312, A3 => n311, ZN => 
                           curr_proc_regs(175));
   U403 : NAND2_X1 port map( A1 => regs(688), A2 => n16, ZN => n316);
   U404 : AOI22_X1 port map( A1 => n33, A2 => regs(1200), B1 => n19, B2 => 
                           regs(176), ZN => n315);
   U405 : AOI22_X1 port map( A1 => n45, A2 => regs(2224), B1 => n34, B2 => 
                           regs(1712), ZN => n314);
   U406 : NAND3_X1 port map( A1 => n316, A2 => n315, A3 => n314, ZN => 
                           curr_proc_regs(176));
   U407 : NAND2_X1 port map( A1 => regs(689), A2 => n16, ZN => n319);
   U408 : AOI22_X1 port map( A1 => n2, A2 => regs(1201), B1 => n19, B2 => 
                           regs(177), ZN => n318);
   U409 : AOI22_X1 port map( A1 => n56, A2 => regs(2225), B1 => n37, B2 => 
                           regs(1713), ZN => n317);
   U410 : NAND3_X1 port map( A1 => n319, A2 => n318, A3 => n317, ZN => 
                           curr_proc_regs(177));
   U411 : NAND2_X1 port map( A1 => regs(690), A2 => n16, ZN => n322);
   U412 : AOI22_X1 port map( A1 => n1597, A2 => regs(1202), B1 => n19, B2 => 
                           regs(178), ZN => n321);
   U413 : AOI22_X1 port map( A1 => n43, A2 => regs(2226), B1 => n38, B2 => 
                           regs(1714), ZN => n320);
   U414 : NAND3_X1 port map( A1 => n322, A2 => n321, A3 => n320, ZN => 
                           curr_proc_regs(178));
   U415 : NAND2_X1 port map( A1 => regs(691), A2 => n16, ZN => n325);
   U416 : AOI22_X1 port map( A1 => n33, A2 => regs(1203), B1 => n19, B2 => 
                           regs(179), ZN => n324);
   U417 : AOI22_X1 port map( A1 => n45, A2 => regs(2227), B1 => n40, B2 => 
                           regs(1715), ZN => n323);
   U418 : NAND3_X1 port map( A1 => n325, A2 => n324, A3 => n323, ZN => 
                           curr_proc_regs(179));
   U419 : NAND2_X1 port map( A1 => regs(529), A2 => n16, ZN => n328);
   U420 : AOI22_X1 port map( A1 => n29, A2 => regs(1041), B1 => n19, B2 => 
                           regs(17), ZN => n327);
   U421 : AOI22_X1 port map( A1 => n49, A2 => regs(2065), B1 => n38, B2 => 
                           regs(1553), ZN => n326);
   U422 : NAND3_X1 port map( A1 => n328, A2 => n327, A3 => n326, ZN => 
                           curr_proc_regs(17));
   U423 : NAND2_X1 port map( A1 => regs(692), A2 => n16, ZN => n331);
   U424 : AOI22_X1 port map( A1 => n33, A2 => regs(1204), B1 => n19, B2 => 
                           regs(180), ZN => n330);
   U425 : AOI22_X1 port map( A1 => n48, A2 => regs(2228), B1 => n36, B2 => 
                           regs(1716), ZN => n329);
   U426 : NAND3_X1 port map( A1 => n331, A2 => n330, A3 => n329, ZN => 
                           curr_proc_regs(180));
   U427 : NAND2_X1 port map( A1 => regs(693), A2 => n16, ZN => n334);
   U428 : AOI22_X1 port map( A1 => n33, A2 => regs(1205), B1 => n19, B2 => 
                           regs(181), ZN => n333);
   U429 : AOI22_X1 port map( A1 => n54, A2 => regs(2229), B1 => n35, B2 => 
                           regs(1717), ZN => n332);
   U430 : NAND3_X1 port map( A1 => n334, A2 => n333, A3 => n332, ZN => 
                           curr_proc_regs(181));
   U431 : NAND2_X1 port map( A1 => regs(694), A2 => n16, ZN => n337);
   U432 : AOI22_X1 port map( A1 => n27, A2 => regs(1206), B1 => n19, B2 => 
                           regs(182), ZN => n336);
   U433 : AOI22_X1 port map( A1 => n51, A2 => regs(2230), B1 => n34, B2 => 
                           regs(1718), ZN => n335);
   U434 : NAND3_X1 port map( A1 => n337, A2 => n336, A3 => n335, ZN => 
                           curr_proc_regs(182));
   U435 : NAND2_X1 port map( A1 => regs(695), A2 => n16, ZN => n340);
   U436 : AOI22_X1 port map( A1 => n29, A2 => regs(1207), B1 => n19, B2 => 
                           regs(183), ZN => n339);
   U437 : AOI22_X1 port map( A1 => n47, A2 => regs(2231), B1 => n37, B2 => 
                           regs(1719), ZN => n338);
   U438 : NAND3_X1 port map( A1 => n340, A2 => n339, A3 => n338, ZN => 
                           curr_proc_regs(183));
   U439 : NAND2_X1 port map( A1 => regs(696), A2 => n16, ZN => n343);
   U440 : AOI22_X1 port map( A1 => n27, A2 => regs(1208), B1 => n19, B2 => 
                           regs(184), ZN => n342);
   U441 : AOI22_X1 port map( A1 => n46, A2 => regs(2232), B1 => n38, B2 => 
                           regs(1720), ZN => n341);
   U442 : NAND3_X1 port map( A1 => n343, A2 => n342, A3 => n341, ZN => 
                           curr_proc_regs(184));
   U443 : NAND2_X1 port map( A1 => regs(697), A2 => n16, ZN => n346);
   U444 : AOI22_X1 port map( A1 => n27, A2 => regs(1209), B1 => n19, B2 => 
                           regs(185), ZN => n345);
   U445 : AOI22_X1 port map( A1 => n50, A2 => regs(2233), B1 => n38, B2 => 
                           regs(1721), ZN => n344);
   U446 : NAND3_X1 port map( A1 => n346, A2 => n345, A3 => n344, ZN => 
                           curr_proc_regs(185));
   U447 : NAND2_X1 port map( A1 => regs(698), A2 => n16, ZN => n349);
   U448 : AOI22_X1 port map( A1 => n27, A2 => regs(1210), B1 => n19, B2 => 
                           regs(186), ZN => n348);
   U449 : AOI22_X1 port map( A1 => n53, A2 => regs(2234), B1 => n38, B2 => 
                           regs(1722), ZN => n347);
   U450 : NAND3_X1 port map( A1 => n349, A2 => n348, A3 => n347, ZN => 
                           curr_proc_regs(186));
   U451 : NAND2_X1 port map( A1 => regs(699), A2 => n1, ZN => n352);
   U452 : AOI22_X1 port map( A1 => n30, A2 => regs(1211), B1 => n23, B2 => 
                           regs(187), ZN => n351);
   U453 : AOI22_X1 port map( A1 => n55, A2 => regs(2235), B1 => n37, B2 => 
                           regs(1723), ZN => n350);
   U454 : NAND3_X1 port map( A1 => n352, A2 => n351, A3 => n350, ZN => 
                           curr_proc_regs(187));
   U455 : NAND2_X1 port map( A1 => regs(700), A2 => n1, ZN => n355);
   U456 : AOI22_X1 port map( A1 => n27, A2 => regs(1212), B1 => n23, B2 => 
                           regs(188), ZN => n354);
   U457 : AOI22_X1 port map( A1 => n46, A2 => regs(2236), B1 => n37, B2 => 
                           regs(1724), ZN => n353);
   U458 : NAND3_X1 port map( A1 => n355, A2 => n354, A3 => n353, ZN => 
                           curr_proc_regs(188));
   U459 : NAND2_X1 port map( A1 => regs(701), A2 => n1, ZN => n358);
   U460 : AOI22_X1 port map( A1 => n29, A2 => regs(1213), B1 => n23, B2 => 
                           regs(189), ZN => n357);
   U461 : AOI22_X1 port map( A1 => n50, A2 => regs(2237), B1 => n37, B2 => 
                           regs(1725), ZN => n356);
   U462 : NAND3_X1 port map( A1 => n358, A2 => n357, A3 => n356, ZN => 
                           curr_proc_regs(189));
   U463 : NAND2_X1 port map( A1 => regs(530), A2 => n1, ZN => n361);
   U464 : AOI22_X1 port map( A1 => n27, A2 => regs(1042), B1 => n23, B2 => 
                           regs(18), ZN => n360);
   U465 : AOI22_X1 port map( A1 => n53, A2 => regs(2066), B1 => n37, B2 => 
                           regs(1554), ZN => n359);
   U466 : NAND3_X1 port map( A1 => n361, A2 => n360, A3 => n359, ZN => 
                           curr_proc_regs(18));
   U467 : NAND2_X1 port map( A1 => regs(702), A2 => n1, ZN => n364);
   U468 : AOI22_X1 port map( A1 => n27, A2 => regs(1214), B1 => n23, B2 => 
                           regs(190), ZN => n363);
   U469 : AOI22_X1 port map( A1 => n55, A2 => regs(2238), B1 => n37, B2 => 
                           regs(1726), ZN => n362);
   U470 : NAND3_X1 port map( A1 => n364, A2 => n363, A3 => n362, ZN => 
                           curr_proc_regs(190));
   U471 : NAND2_X1 port map( A1 => regs(703), A2 => n1, ZN => n367);
   U472 : AOI22_X1 port map( A1 => n27, A2 => regs(1215), B1 => n23, B2 => 
                           regs(191), ZN => n366);
   U473 : AOI22_X1 port map( A1 => n52, A2 => regs(2239), B1 => n37, B2 => 
                           regs(1727), ZN => n365);
   U474 : NAND3_X1 port map( A1 => n367, A2 => n366, A3 => n365, ZN => 
                           curr_proc_regs(191));
   U475 : NAND2_X1 port map( A1 => regs(704), A2 => n1, ZN => n370);
   U476 : AOI22_X1 port map( A1 => n30, A2 => regs(1216), B1 => n23, B2 => 
                           regs(192), ZN => n369);
   U477 : AOI22_X1 port map( A1 => n56, A2 => regs(2240), B1 => n37, B2 => 
                           regs(1728), ZN => n368);
   U478 : NAND3_X1 port map( A1 => n370, A2 => n369, A3 => n368, ZN => 
                           curr_proc_regs(192));
   U479 : NAND2_X1 port map( A1 => regs(705), A2 => n1, ZN => n373);
   U480 : AOI22_X1 port map( A1 => n27, A2 => regs(1217), B1 => n23, B2 => 
                           regs(193), ZN => n372);
   U481 : AOI22_X1 port map( A1 => n43, A2 => regs(2241), B1 => n37, B2 => 
                           regs(1729), ZN => n371);
   U482 : NAND3_X1 port map( A1 => n373, A2 => n372, A3 => n371, ZN => 
                           curr_proc_regs(193));
   U483 : NAND2_X1 port map( A1 => regs(706), A2 => n1, ZN => n376);
   U484 : AOI22_X1 port map( A1 => n29, A2 => regs(1218), B1 => n23, B2 => 
                           regs(194), ZN => n375);
   U485 : AOI22_X1 port map( A1 => n45, A2 => regs(2242), B1 => n37, B2 => 
                           regs(1730), ZN => n374);
   U486 : NAND3_X1 port map( A1 => n376, A2 => n375, A3 => n374, ZN => 
                           curr_proc_regs(194));
   U487 : NAND2_X1 port map( A1 => regs(707), A2 => n1, ZN => n379);
   U488 : AOI22_X1 port map( A1 => n1597, A2 => regs(1219), B1 => n23, B2 => 
                           regs(195), ZN => n378);
   U489 : AOI22_X1 port map( A1 => n49, A2 => regs(2243), B1 => n37, B2 => 
                           regs(1731), ZN => n377);
   U490 : NAND3_X1 port map( A1 => n379, A2 => n378, A3 => n377, ZN => 
                           curr_proc_regs(195));
   U491 : NAND2_X1 port map( A1 => regs(708), A2 => n1, ZN => n382);
   U492 : AOI22_X1 port map( A1 => n27, A2 => regs(1220), B1 => n23, B2 => 
                           regs(196), ZN => n381);
   U493 : AOI22_X1 port map( A1 => n51, A2 => regs(2244), B1 => n37, B2 => 
                           regs(1732), ZN => n380);
   U494 : NAND3_X1 port map( A1 => n382, A2 => n381, A3 => n380, ZN => 
                           curr_proc_regs(196));
   U495 : NAND2_X1 port map( A1 => regs(709), A2 => n1, ZN => n385);
   U496 : AOI22_X1 port map( A1 => n1597, A2 => regs(1221), B1 => n19, B2 => 
                           regs(197), ZN => n384);
   U497 : AOI22_X1 port map( A1 => n43, A2 => regs(2245), B1 => n37, B2 => 
                           regs(1733), ZN => n383);
   U498 : NAND3_X1 port map( A1 => n385, A2 => n384, A3 => n383, ZN => 
                           curr_proc_regs(197));
   U499 : NAND2_X1 port map( A1 => regs(710), A2 => n9, ZN => n388);
   U500 : AOI22_X1 port map( A1 => n27, A2 => regs(1222), B1 => n20, B2 => 
                           regs(198), ZN => n387);
   U501 : AOI22_X1 port map( A1 => n43, A2 => regs(2246), B1 => n38, B2 => 
                           regs(1734), ZN => n386);
   U502 : NAND3_X1 port map( A1 => n388, A2 => n387, A3 => n386, ZN => 
                           curr_proc_regs(198));
   U503 : NAND2_X1 port map( A1 => regs(711), A2 => n4, ZN => n391);
   U504 : AOI22_X1 port map( A1 => n29, A2 => regs(1223), B1 => n26, B2 => 
                           regs(199), ZN => n390);
   U505 : AOI22_X1 port map( A1 => n53, A2 => regs(2247), B1 => n38, B2 => 
                           regs(1735), ZN => n389);
   U506 : NAND3_X1 port map( A1 => n391, A2 => n390, A3 => n389, ZN => 
                           curr_proc_regs(199));
   U507 : NAND2_X1 port map( A1 => regs(531), A2 => n1, ZN => n394);
   U508 : AOI22_X1 port map( A1 => n27, A2 => regs(1043), B1 => n21, B2 => 
                           regs(19), ZN => n393);
   U509 : AOI22_X1 port map( A1 => n53, A2 => regs(2067), B1 => n38, B2 => 
                           regs(1555), ZN => n392);
   U510 : NAND3_X1 port map( A1 => n394, A2 => n393, A3 => n392, ZN => 
                           curr_proc_regs(19));
   U511 : NAND2_X1 port map( A1 => regs(513), A2 => n9, ZN => n397);
   U512 : AOI22_X1 port map( A1 => n30, A2 => regs(1025), B1 => n19, B2 => 
                           regs(1), ZN => n396);
   U513 : AOI22_X1 port map( A1 => n53, A2 => regs(2049), B1 => n38, B2 => 
                           regs(1537), ZN => n395);
   U514 : NAND3_X1 port map( A1 => n397, A2 => n396, A3 => n395, ZN => 
                           curr_proc_regs(1));
   U515 : NAND2_X1 port map( A1 => regs(712), A2 => n4, ZN => n400);
   U516 : AOI22_X1 port map( A1 => n27, A2 => regs(1224), B1 => n21, B2 => 
                           regs(200), ZN => n399);
   U517 : AOI22_X1 port map( A1 => n53, A2 => regs(2248), B1 => n38, B2 => 
                           regs(1736), ZN => n398);
   U518 : NAND3_X1 port map( A1 => n400, A2 => n399, A3 => n398, ZN => 
                           curr_proc_regs(200));
   U519 : NAND2_X1 port map( A1 => regs(713), A2 => n1, ZN => n403);
   U520 : AOI22_X1 port map( A1 => n27, A2 => regs(1225), B1 => n17, B2 => 
                           regs(201), ZN => n402);
   U521 : AOI22_X1 port map( A1 => n53, A2 => regs(2249), B1 => n38, B2 => 
                           regs(1737), ZN => n401);
   U522 : NAND3_X1 port map( A1 => n403, A2 => n402, A3 => n401, ZN => 
                           curr_proc_regs(201));
   U523 : NAND2_X1 port map( A1 => regs(714), A2 => n9, ZN => n406);
   U524 : AOI22_X1 port map( A1 => n27, A2 => regs(1226), B1 => n26, B2 => 
                           regs(202), ZN => n405);
   U525 : AOI22_X1 port map( A1 => n53, A2 => regs(2250), B1 => n38, B2 => 
                           regs(1738), ZN => n404);
   U526 : NAND3_X1 port map( A1 => n406, A2 => n405, A3 => n404, ZN => 
                           curr_proc_regs(202));
   U527 : NAND2_X1 port map( A1 => regs(715), A2 => n4, ZN => n409);
   U528 : AOI22_X1 port map( A1 => n29, A2 => regs(1227), B1 => n21, B2 => 
                           regs(203), ZN => n408);
   U529 : AOI22_X1 port map( A1 => n53, A2 => regs(2251), B1 => n38, B2 => 
                           regs(1739), ZN => n407);
   U530 : NAND3_X1 port map( A1 => n409, A2 => n408, A3 => n407, ZN => 
                           curr_proc_regs(203));
   U531 : NAND2_X1 port map( A1 => regs(716), A2 => n1, ZN => n412);
   U532 : AOI22_X1 port map( A1 => n2, A2 => regs(1228), B1 => n18, B2 => 
                           regs(204), ZN => n411);
   U533 : AOI22_X1 port map( A1 => n53, A2 => regs(2252), B1 => n38, B2 => 
                           regs(1740), ZN => n410);
   U534 : NAND3_X1 port map( A1 => n412, A2 => n411, A3 => n410, ZN => 
                           curr_proc_regs(204));
   U535 : NAND2_X1 port map( A1 => regs(717), A2 => n9, ZN => n415);
   U536 : AOI22_X1 port map( A1 => n2, A2 => regs(1229), B1 => n1596, B2 => 
                           regs(205), ZN => n414);
   U537 : AOI22_X1 port map( A1 => n53, A2 => regs(2253), B1 => n38, B2 => 
                           regs(1741), ZN => n413);
   U538 : NAND3_X1 port map( A1 => n415, A2 => n414, A3 => n413, ZN => 
                           curr_proc_regs(205));
   U539 : NAND2_X1 port map( A1 => regs(718), A2 => n4, ZN => n418);
   U540 : AOI22_X1 port map( A1 => n2, A2 => regs(1230), B1 => n19, B2 => 
                           regs(206), ZN => n417);
   U541 : AOI22_X1 port map( A1 => n53, A2 => regs(2254), B1 => n38, B2 => 
                           regs(1742), ZN => n416);
   U542 : NAND3_X1 port map( A1 => n418, A2 => n417, A3 => n416, ZN => 
                           curr_proc_regs(206));
   U543 : NAND2_X1 port map( A1 => regs(719), A2 => n1, ZN => n421);
   U544 : AOI22_X1 port map( A1 => n2, A2 => regs(1231), B1 => n21, B2 => 
                           regs(207), ZN => n420);
   U545 : AOI22_X1 port map( A1 => n53, A2 => regs(2255), B1 => n38, B2 => 
                           regs(1743), ZN => n419);
   U546 : NAND3_X1 port map( A1 => n421, A2 => n420, A3 => n419, ZN => 
                           curr_proc_regs(207));
   U547 : NAND2_X1 port map( A1 => regs(720), A2 => n9, ZN => n424);
   U548 : AOI22_X1 port map( A1 => n2, A2 => regs(1232), B1 => n20, B2 => 
                           regs(208), ZN => n423);
   U549 : AOI22_X1 port map( A1 => n53, A2 => regs(2256), B1 => n36, B2 => 
                           regs(1744), ZN => n422);
   U550 : NAND3_X1 port map( A1 => n424, A2 => n423, A3 => n422, ZN => 
                           curr_proc_regs(208));
   U551 : NAND2_X1 port map( A1 => regs(721), A2 => n9, ZN => n427);
   U552 : AOI22_X1 port map( A1 => n2, A2 => regs(1233), B1 => n26, B2 => 
                           regs(209), ZN => n426);
   U553 : AOI22_X1 port map( A1 => n6, A2 => regs(2257), B1 => n35, B2 => 
                           regs(1745), ZN => n425);
   U554 : NAND3_X1 port map( A1 => n427, A2 => n426, A3 => n425, ZN => 
                           curr_proc_regs(209));
   U555 : NAND2_X1 port map( A1 => regs(532), A2 => n9, ZN => n430);
   U556 : AOI22_X1 port map( A1 => n32, A2 => regs(1044), B1 => n19, B2 => 
                           regs(20), ZN => n429);
   U557 : AOI22_X1 port map( A1 => n6, A2 => regs(2068), B1 => n40, B2 => 
                           regs(1556), ZN => n428);
   U558 : NAND3_X1 port map( A1 => n430, A2 => n429, A3 => n428, ZN => 
                           curr_proc_regs(20));
   U559 : NAND2_X1 port map( A1 => regs(722), A2 => n9, ZN => n433);
   U560 : AOI22_X1 port map( A1 => n2, A2 => regs(1234), B1 => n21, B2 => 
                           regs(210), ZN => n432);
   U561 : AOI22_X1 port map( A1 => n6, A2 => regs(2258), B1 => n36, B2 => 
                           regs(1746), ZN => n431);
   U562 : NAND3_X1 port map( A1 => n433, A2 => n432, A3 => n431, ZN => 
                           curr_proc_regs(210));
   U563 : NAND2_X1 port map( A1 => regs(723), A2 => n9, ZN => n436);
   U564 : AOI22_X1 port map( A1 => n2, A2 => regs(1235), B1 => n20, B2 => 
                           regs(211), ZN => n435);
   U565 : AOI22_X1 port map( A1 => n6, A2 => regs(2259), B1 => n35, B2 => 
                           regs(1747), ZN => n434);
   U566 : NAND3_X1 port map( A1 => n436, A2 => n435, A3 => n434, ZN => 
                           curr_proc_regs(211));
   U567 : NAND2_X1 port map( A1 => regs(724), A2 => n9, ZN => n439);
   U568 : AOI22_X1 port map( A1 => n2, A2 => regs(1236), B1 => n21, B2 => 
                           regs(212), ZN => n438);
   U569 : AOI22_X1 port map( A1 => n6, A2 => regs(2260), B1 => n40, B2 => 
                           regs(1748), ZN => n437);
   U570 : NAND3_X1 port map( A1 => n439, A2 => n438, A3 => n437, ZN => 
                           curr_proc_regs(212));
   U571 : NAND2_X1 port map( A1 => regs(725), A2 => n9, ZN => n442);
   U572 : AOI22_X1 port map( A1 => n2, A2 => regs(1237), B1 => n19, B2 => 
                           regs(213), ZN => n441);
   U573 : AOI22_X1 port map( A1 => n6, A2 => regs(2261), B1 => n36, B2 => 
                           regs(1749), ZN => n440);
   U574 : NAND3_X1 port map( A1 => n442, A2 => n441, A3 => n440, ZN => 
                           curr_proc_regs(213));
   U575 : NAND2_X1 port map( A1 => regs(726), A2 => n9, ZN => n445);
   U576 : AOI22_X1 port map( A1 => n32, A2 => regs(1238), B1 => n21, B2 => 
                           regs(214), ZN => n444);
   U577 : AOI22_X1 port map( A1 => n55, A2 => regs(2262), B1 => n35, B2 => 
                           regs(1750), ZN => n443);
   U578 : NAND3_X1 port map( A1 => n445, A2 => n444, A3 => n443, ZN => 
                           curr_proc_regs(214));
   U579 : NAND2_X1 port map( A1 => regs(727), A2 => n9, ZN => n448);
   U580 : AOI22_X1 port map( A1 => n2, A2 => regs(1239), B1 => n20, B2 => 
                           regs(215), ZN => n447);
   U581 : AOI22_X1 port map( A1 => n52, A2 => regs(2263), B1 => n40, B2 => 
                           regs(1751), ZN => n446);
   U582 : NAND3_X1 port map( A1 => n448, A2 => n447, A3 => n446, ZN => 
                           curr_proc_regs(215));
   U583 : NAND2_X1 port map( A1 => regs(728), A2 => n9, ZN => n451);
   U584 : AOI22_X1 port map( A1 => n2, A2 => regs(1240), B1 => n19, B2 => 
                           regs(216), ZN => n450);
   U585 : AOI22_X1 port map( A1 => n57, A2 => regs(2264), B1 => n36, B2 => 
                           regs(1752), ZN => n449);
   U586 : NAND3_X1 port map( A1 => n451, A2 => n450, A3 => n449, ZN => 
                           curr_proc_regs(216));
   U587 : NAND2_X1 port map( A1 => regs(729), A2 => n9, ZN => n454);
   U588 : AOI22_X1 port map( A1 => n2, A2 => regs(1241), B1 => n19, B2 => 
                           regs(217), ZN => n453);
   U589 : AOI22_X1 port map( A1 => n57, A2 => regs(2265), B1 => n35, B2 => 
                           regs(1753), ZN => n452);
   U590 : NAND3_X1 port map( A1 => n454, A2 => n453, A3 => n452, ZN => 
                           curr_proc_regs(217));
   U591 : NAND2_X1 port map( A1 => regs(730), A2 => n9, ZN => n457);
   U592 : AOI22_X1 port map( A1 => n2, A2 => regs(1242), B1 => n21, B2 => 
                           regs(218), ZN => n456);
   U593 : AOI22_X1 port map( A1 => n57, A2 => regs(2266), B1 => n40, B2 => 
                           regs(1754), ZN => n455);
   U594 : NAND3_X1 port map( A1 => n457, A2 => n456, A3 => n455, ZN => 
                           curr_proc_regs(218));
   U595 : NAND2_X1 port map( A1 => regs(731), A2 => n1, ZN => n460);
   U596 : AOI22_X1 port map( A1 => n2, A2 => regs(1243), B1 => n20, B2 => 
                           regs(219), ZN => n459);
   U597 : AOI22_X1 port map( A1 => n44, A2 => regs(2267), B1 => n38, B2 => 
                           regs(1755), ZN => n458);
   U598 : NAND3_X1 port map( A1 => n460, A2 => n459, A3 => n458, ZN => 
                           curr_proc_regs(219));
   U599 : NAND2_X1 port map( A1 => regs(533), A2 => n9, ZN => n463);
   U600 : AOI22_X1 port map( A1 => n2, A2 => regs(1045), B1 => n20, B2 => 
                           regs(21), ZN => n462);
   U601 : AOI22_X1 port map( A1 => n47, A2 => regs(2069), B1 => n38, B2 => 
                           regs(1557), ZN => n461);
   U602 : NAND3_X1 port map( A1 => n463, A2 => n462, A3 => n461, ZN => 
                           curr_proc_regs(21));
   U603 : NAND2_X1 port map( A1 => regs(732), A2 => n4, ZN => n466);
   U604 : AOI22_X1 port map( A1 => n32, A2 => regs(1244), B1 => n20, B2 => 
                           regs(220), ZN => n465);
   U605 : AOI22_X1 port map( A1 => n48, A2 => regs(2268), B1 => n38, B2 => 
                           regs(1756), ZN => n464);
   U606 : NAND3_X1 port map( A1 => n466, A2 => n465, A3 => n464, ZN => 
                           curr_proc_regs(220));
   U607 : NAND2_X1 port map( A1 => regs(733), A2 => n9, ZN => n469);
   U608 : AOI22_X1 port map( A1 => n2, A2 => regs(1245), B1 => n20, B2 => 
                           regs(221), ZN => n468);
   U609 : AOI22_X1 port map( A1 => n54, A2 => regs(2269), B1 => n38, B2 => 
                           regs(1757), ZN => n467);
   U610 : NAND3_X1 port map( A1 => n469, A2 => n468, A3 => n467, ZN => 
                           curr_proc_regs(221));
   U611 : NAND2_X1 port map( A1 => regs(734), A2 => n1, ZN => n472);
   U612 : AOI22_X1 port map( A1 => n32, A2 => regs(1246), B1 => n20, B2 => 
                           regs(222), ZN => n471);
   U613 : AOI22_X1 port map( A1 => n57, A2 => regs(2270), B1 => n35, B2 => 
                           regs(1758), ZN => n470);
   U614 : NAND3_X1 port map( A1 => n472, A2 => n471, A3 => n470, ZN => 
                           curr_proc_regs(222));
   U615 : NAND2_X1 port map( A1 => regs(735), A2 => n9, ZN => n475);
   U616 : AOI22_X1 port map( A1 => n2, A2 => regs(1247), B1 => n20, B2 => 
                           regs(223), ZN => n474);
   U617 : AOI22_X1 port map( A1 => n57, A2 => regs(2271), B1 => n34, B2 => 
                           regs(1759), ZN => n473);
   U618 : NAND3_X1 port map( A1 => n475, A2 => n474, A3 => n473, ZN => 
                           curr_proc_regs(223));
   U619 : NAND2_X1 port map( A1 => regs(736), A2 => n4, ZN => n478);
   U620 : AOI22_X1 port map( A1 => n32, A2 => regs(1248), B1 => n20, B2 => 
                           regs(224), ZN => n477);
   U621 : AOI22_X1 port map( A1 => n57, A2 => regs(2272), B1 => n37, B2 => 
                           regs(1760), ZN => n476);
   U622 : NAND3_X1 port map( A1 => n478, A2 => n477, A3 => n476, ZN => 
                           curr_proc_regs(224));
   U623 : NAND2_X1 port map( A1 => regs(737), A2 => n4, ZN => n481);
   U624 : AOI22_X1 port map( A1 => n2, A2 => regs(1249), B1 => n20, B2 => 
                           regs(225), ZN => n480);
   U625 : AOI22_X1 port map( A1 => n57, A2 => regs(2273), B1 => n38, B2 => 
                           regs(1761), ZN => n479);
   U626 : NAND3_X1 port map( A1 => n481, A2 => n480, A3 => n479, ZN => 
                           curr_proc_regs(225));
   U627 : NAND2_X1 port map( A1 => regs(738), A2 => n1, ZN => n484);
   U628 : AOI22_X1 port map( A1 => n2, A2 => regs(1250), B1 => n20, B2 => 
                           regs(226), ZN => n483);
   U629 : AOI22_X1 port map( A1 => n55, A2 => regs(2274), B1 => n1598, B2 => 
                           regs(1762), ZN => n482);
   U630 : NAND3_X1 port map( A1 => n484, A2 => n483, A3 => n482, ZN => 
                           curr_proc_regs(226));
   U631 : NAND2_X1 port map( A1 => regs(739), A2 => n4, ZN => n487);
   U632 : AOI22_X1 port map( A1 => n2, A2 => regs(1251), B1 => n20, B2 => 
                           regs(227), ZN => n486);
   U633 : AOI22_X1 port map( A1 => n57, A2 => regs(2275), B1 => n38, B2 => 
                           regs(1763), ZN => n485);
   U634 : NAND3_X1 port map( A1 => n487, A2 => n486, A3 => n485, ZN => 
                           curr_proc_regs(227));
   U635 : NAND2_X1 port map( A1 => regs(740), A2 => n4, ZN => n490);
   U636 : AOI22_X1 port map( A1 => n32, A2 => regs(1252), B1 => n20, B2 => 
                           regs(228), ZN => n489);
   U637 : AOI22_X1 port map( A1 => n57, A2 => regs(2276), B1 => n1598, B2 => 
                           regs(1764), ZN => n488);
   U638 : NAND3_X1 port map( A1 => n490, A2 => n489, A3 => n488, ZN => 
                           curr_proc_regs(228));
   U639 : NAND2_X1 port map( A1 => regs(741), A2 => n4, ZN => n493);
   U640 : AOI22_X1 port map( A1 => n2, A2 => regs(1253), B1 => n20, B2 => 
                           regs(229), ZN => n492);
   U641 : AOI22_X1 port map( A1 => n53, A2 => regs(2277), B1 => n38, B2 => 
                           regs(1765), ZN => n491);
   U642 : NAND3_X1 port map( A1 => n493, A2 => n492, A3 => n491, ZN => 
                           curr_proc_regs(229));
   U643 : NAND2_X1 port map( A1 => regs(534), A2 => n9, ZN => n496);
   U644 : AOI22_X1 port map( A1 => n2, A2 => regs(1046), B1 => n21, B2 => 
                           regs(22), ZN => n495);
   U645 : AOI22_X1 port map( A1 => n57, A2 => regs(2070), B1 => n39, B2 => 
                           regs(1558), ZN => n494);
   U646 : NAND3_X1 port map( A1 => n496, A2 => n495, A3 => n494, ZN => 
                           curr_proc_regs(22));
   U647 : NAND2_X1 port map( A1 => regs(742), A2 => n4, ZN => n499);
   U648 : AOI22_X1 port map( A1 => n32, A2 => regs(1254), B1 => n18, B2 => 
                           regs(230), ZN => n498);
   U649 : AOI22_X1 port map( A1 => n57, A2 => regs(2278), B1 => n39, B2 => 
                           regs(1766), ZN => n497);
   U650 : NAND3_X1 port map( A1 => n499, A2 => n498, A3 => n497, ZN => 
                           curr_proc_regs(230));
   U651 : NAND2_X1 port map( A1 => regs(743), A2 => n4, ZN => n502);
   U652 : AOI22_X1 port map( A1 => n2, A2 => regs(1255), B1 => n23, B2 => 
                           regs(231), ZN => n501);
   U653 : AOI22_X1 port map( A1 => n57, A2 => regs(2279), B1 => n39, B2 => 
                           regs(1767), ZN => n500);
   U654 : NAND3_X1 port map( A1 => n502, A2 => n501, A3 => n500, ZN => 
                           curr_proc_regs(231));
   U655 : NAND2_X1 port map( A1 => regs(744), A2 => n4, ZN => n505);
   U656 : AOI22_X1 port map( A1 => n2, A2 => regs(1256), B1 => n26, B2 => 
                           regs(232), ZN => n504);
   U657 : AOI22_X1 port map( A1 => n57, A2 => regs(2280), B1 => n39, B2 => 
                           regs(1768), ZN => n503);
   U658 : NAND3_X1 port map( A1 => n505, A2 => n504, A3 => n503, ZN => 
                           curr_proc_regs(232));
   U659 : NAND2_X1 port map( A1 => regs(745), A2 => n1, ZN => n508);
   U660 : AOI22_X1 port map( A1 => n32, A2 => regs(1257), B1 => n26, B2 => 
                           regs(233), ZN => n507);
   U661 : AOI22_X1 port map( A1 => n57, A2 => regs(2281), B1 => n39, B2 => 
                           regs(1769), ZN => n506);
   U662 : NAND3_X1 port map( A1 => n508, A2 => n507, A3 => n506, ZN => 
                           curr_proc_regs(233));
   U663 : NAND2_X1 port map( A1 => regs(746), A2 => n9, ZN => n511);
   U664 : AOI22_X1 port map( A1 => n2, A2 => regs(1258), B1 => n19, B2 => 
                           regs(234), ZN => n510);
   U665 : AOI22_X1 port map( A1 => n57, A2 => regs(2282), B1 => n39, B2 => 
                           regs(1770), ZN => n509);
   U666 : NAND3_X1 port map( A1 => n511, A2 => n510, A3 => n509, ZN => 
                           curr_proc_regs(234));
   U667 : NAND2_X1 port map( A1 => regs(747), A2 => n4, ZN => n514);
   U668 : AOI22_X1 port map( A1 => n2, A2 => regs(1259), B1 => n21, B2 => 
                           regs(235), ZN => n513);
   U669 : AOI22_X1 port map( A1 => n57, A2 => regs(2283), B1 => n39, B2 => 
                           regs(1771), ZN => n512);
   U670 : NAND3_X1 port map( A1 => n514, A2 => n513, A3 => n512, ZN => 
                           curr_proc_regs(235));
   U671 : NAND2_X1 port map( A1 => regs(748), A2 => n4, ZN => n517);
   U672 : AOI22_X1 port map( A1 => n32, A2 => regs(1260), B1 => n17, B2 => 
                           regs(236), ZN => n516);
   U673 : AOI22_X1 port map( A1 => n57, A2 => regs(2284), B1 => n39, B2 => 
                           regs(1772), ZN => n515);
   U674 : NAND3_X1 port map( A1 => n517, A2 => n516, A3 => n515, ZN => 
                           curr_proc_regs(236));
   U675 : NAND2_X1 port map( A1 => regs(749), A2 => n4, ZN => n520);
   U676 : AOI22_X1 port map( A1 => n2, A2 => regs(1261), B1 => n26, B2 => 
                           regs(237), ZN => n519);
   U677 : AOI22_X1 port map( A1 => win(4), A2 => regs(2285), B1 => n39, B2 => 
                           regs(1773), ZN => n518);
   U678 : NAND3_X1 port map( A1 => n520, A2 => n519, A3 => n518, ZN => 
                           curr_proc_regs(237));
   U679 : NAND2_X1 port map( A1 => regs(750), A2 => n4, ZN => n523);
   U680 : AOI22_X1 port map( A1 => n2, A2 => regs(1262), B1 => n20, B2 => 
                           regs(238), ZN => n522);
   U681 : AOI22_X1 port map( A1 => n57, A2 => regs(2286), B1 => n39, B2 => 
                           regs(1774), ZN => n521);
   U682 : NAND3_X1 port map( A1 => n523, A2 => n522, A3 => n521, ZN => 
                           curr_proc_regs(238));
   U683 : NAND2_X1 port map( A1 => regs(751), A2 => n4, ZN => n526);
   U684 : AOI22_X1 port map( A1 => n2, A2 => regs(1263), B1 => n26, B2 => 
                           regs(239), ZN => n525);
   U685 : AOI22_X1 port map( A1 => win(4), A2 => regs(2287), B1 => n39, B2 => 
                           regs(1775), ZN => n524);
   U686 : NAND3_X1 port map( A1 => n526, A2 => n525, A3 => n524, ZN => 
                           curr_proc_regs(239));
   U687 : NAND2_X1 port map( A1 => regs(535), A2 => n4, ZN => n529);
   U688 : AOI22_X1 port map( A1 => n2, A2 => regs(1047), B1 => n18, B2 => 
                           regs(23), ZN => n528);
   U689 : AOI22_X1 port map( A1 => n57, A2 => regs(2071), B1 => n39, B2 => 
                           regs(1559), ZN => n527);
   U690 : NAND3_X1 port map( A1 => n529, A2 => n528, A3 => n527, ZN => 
                           curr_proc_regs(23));
   U691 : NAND2_X1 port map( A1 => regs(752), A2 => n3, ZN => n532);
   U692 : AOI22_X1 port map( A1 => n2, A2 => regs(1264), B1 => n21, B2 => 
                           regs(240), ZN => n531);
   U693 : AOI22_X1 port map( A1 => n56, A2 => regs(2288), B1 => n42, B2 => 
                           regs(1776), ZN => n530);
   U694 : NAND3_X1 port map( A1 => n532, A2 => n531, A3 => n530, ZN => 
                           curr_proc_regs(240));
   U695 : NAND2_X1 port map( A1 => regs(753), A2 => n3, ZN => n535);
   U696 : AOI22_X1 port map( A1 => n2, A2 => regs(1265), B1 => n21, B2 => 
                           regs(241), ZN => n534);
   U697 : AOI22_X1 port map( A1 => n57, A2 => regs(2289), B1 => n42, B2 => 
                           regs(1777), ZN => n533);
   U698 : NAND3_X1 port map( A1 => n535, A2 => n534, A3 => n533, ZN => 
                           curr_proc_regs(241));
   U699 : NAND2_X1 port map( A1 => regs(754), A2 => n3, ZN => n538);
   U700 : AOI22_X1 port map( A1 => n2, A2 => regs(1266), B1 => n21, B2 => 
                           regs(242), ZN => n537);
   U701 : AOI22_X1 port map( A1 => n57, A2 => regs(2290), B1 => n42, B2 => 
                           regs(1778), ZN => n536);
   U702 : NAND3_X1 port map( A1 => n538, A2 => n537, A3 => n536, ZN => 
                           curr_proc_regs(242));
   U703 : NAND2_X1 port map( A1 => regs(755), A2 => n3, ZN => n541);
   U704 : AOI22_X1 port map( A1 => n2, A2 => regs(1267), B1 => n21, B2 => 
                           regs(243), ZN => n540);
   U705 : AOI22_X1 port map( A1 => n57, A2 => regs(2291), B1 => n42, B2 => 
                           regs(1779), ZN => n539);
   U706 : NAND3_X1 port map( A1 => n541, A2 => n540, A3 => n539, ZN => 
                           curr_proc_regs(243));
   U707 : NAND2_X1 port map( A1 => regs(756), A2 => n3, ZN => n544);
   U708 : AOI22_X1 port map( A1 => n2, A2 => regs(1268), B1 => n21, B2 => 
                           regs(244), ZN => n543);
   U709 : AOI22_X1 port map( A1 => n45, A2 => regs(2292), B1 => n42, B2 => 
                           regs(1780), ZN => n542);
   U710 : NAND3_X1 port map( A1 => n544, A2 => n543, A3 => n542, ZN => 
                           curr_proc_regs(244));
   U711 : NAND2_X1 port map( A1 => regs(757), A2 => n3, ZN => n547);
   U712 : AOI22_X1 port map( A1 => n2, A2 => regs(1269), B1 => n21, B2 => 
                           regs(245), ZN => n546);
   U713 : AOI22_X1 port map( A1 => n46, A2 => regs(2293), B1 => n42, B2 => 
                           regs(1781), ZN => n545);
   U714 : NAND3_X1 port map( A1 => n547, A2 => n546, A3 => n545, ZN => 
                           curr_proc_regs(245));
   U715 : NAND2_X1 port map( A1 => regs(758), A2 => n3, ZN => n550);
   U716 : AOI22_X1 port map( A1 => n2, A2 => regs(1270), B1 => n21, B2 => 
                           regs(246), ZN => n549);
   U717 : AOI22_X1 port map( A1 => n57, A2 => regs(2294), B1 => n42, B2 => 
                           regs(1782), ZN => n548);
   U718 : NAND3_X1 port map( A1 => n550, A2 => n549, A3 => n548, ZN => 
                           curr_proc_regs(246));
   U719 : NAND2_X1 port map( A1 => regs(759), A2 => n3, ZN => n553);
   U720 : AOI22_X1 port map( A1 => n2, A2 => regs(1271), B1 => n21, B2 => 
                           regs(247), ZN => n552);
   U721 : AOI22_X1 port map( A1 => n57, A2 => regs(2295), B1 => n42, B2 => 
                           regs(1783), ZN => n551);
   U722 : NAND3_X1 port map( A1 => n553, A2 => n552, A3 => n551, ZN => 
                           curr_proc_regs(247));
   U723 : NAND2_X1 port map( A1 => regs(760), A2 => n3, ZN => n556);
   U724 : AOI22_X1 port map( A1 => n32, A2 => regs(1272), B1 => n21, B2 => 
                           regs(248), ZN => n555);
   U725 : AOI22_X1 port map( A1 => n57, A2 => regs(2296), B1 => n42, B2 => 
                           regs(1784), ZN => n554);
   U726 : NAND3_X1 port map( A1 => n556, A2 => n555, A3 => n554, ZN => 
                           curr_proc_regs(248));
   U727 : NAND2_X1 port map( A1 => regs(761), A2 => n3, ZN => n559);
   U728 : AOI22_X1 port map( A1 => n32, A2 => regs(1273), B1 => n21, B2 => 
                           regs(249), ZN => n558);
   U729 : AOI22_X1 port map( A1 => n57, A2 => regs(2297), B1 => n42, B2 => 
                           regs(1785), ZN => n557);
   U730 : NAND3_X1 port map( A1 => n559, A2 => n558, A3 => n557, ZN => 
                           curr_proc_regs(249));
   U731 : NAND2_X1 port map( A1 => regs(536), A2 => n3, ZN => n562);
   U732 : AOI22_X1 port map( A1 => n32, A2 => regs(1048), B1 => n21, B2 => 
                           regs(24), ZN => n561);
   U733 : AOI22_X1 port map( A1 => n50, A2 => regs(2072), B1 => n42, B2 => 
                           regs(1560), ZN => n560);
   U734 : NAND3_X1 port map( A1 => n562, A2 => n561, A3 => n560, ZN => 
                           curr_proc_regs(24));
   U735 : NAND2_X1 port map( A1 => regs(762), A2 => n3, ZN => n565);
   U736 : AOI22_X1 port map( A1 => n32, A2 => regs(1274), B1 => n21, B2 => 
                           regs(250), ZN => n564);
   U737 : AOI22_X1 port map( A1 => n51, A2 => regs(2298), B1 => n42, B2 => 
                           regs(1786), ZN => n563);
   U738 : NAND3_X1 port map( A1 => n565, A2 => n564, A3 => n563, ZN => 
                           curr_proc_regs(250));
   U739 : NAND2_X1 port map( A1 => regs(763), A2 => n16, ZN => n568);
   U740 : AOI22_X1 port map( A1 => n32, A2 => regs(1275), B1 => n26, B2 => 
                           regs(251), ZN => n567);
   U741 : AOI22_X1 port map( A1 => n57, A2 => regs(2299), B1 => n42, B2 => 
                           regs(1787), ZN => n566);
   U742 : NAND3_X1 port map( A1 => n568, A2 => n567, A3 => n566, ZN => 
                           curr_proc_regs(251));
   U743 : NAND2_X1 port map( A1 => regs(764), A2 => n3, ZN => n571);
   U744 : AOI22_X1 port map( A1 => n32, A2 => regs(1276), B1 => n26, B2 => 
                           regs(252), ZN => n570);
   U745 : AOI22_X1 port map( A1 => n57, A2 => regs(2300), B1 => n42, B2 => 
                           regs(1788), ZN => n569);
   U746 : NAND3_X1 port map( A1 => n571, A2 => n570, A3 => n569, ZN => 
                           curr_proc_regs(252));
   U747 : NAND2_X1 port map( A1 => regs(765), A2 => n3, ZN => n574);
   U748 : AOI22_X1 port map( A1 => n32, A2 => regs(1277), B1 => n21, B2 => 
                           regs(253), ZN => n573);
   U749 : AOI22_X1 port map( A1 => n57, A2 => regs(2301), B1 => n42, B2 => 
                           regs(1789), ZN => n572);
   U750 : NAND3_X1 port map( A1 => n574, A2 => n573, A3 => n572, ZN => 
                           curr_proc_regs(253));
   U751 : NAND2_X1 port map( A1 => regs(766), A2 => n16, ZN => n577);
   U752 : AOI22_X1 port map( A1 => n32, A2 => regs(1278), B1 => n26, B2 => 
                           regs(254), ZN => n576);
   U753 : AOI22_X1 port map( A1 => n57, A2 => regs(2302), B1 => n42, B2 => 
                           regs(1790), ZN => n575);
   U754 : NAND3_X1 port map( A1 => n577, A2 => n576, A3 => n575, ZN => 
                           curr_proc_regs(254));
   U755 : NAND2_X1 port map( A1 => regs(767), A2 => n3, ZN => n580);
   U756 : AOI22_X1 port map( A1 => n32, A2 => regs(1279), B1 => n26, B2 => 
                           regs(255), ZN => n579);
   U757 : AOI22_X1 port map( A1 => n49, A2 => regs(2303), B1 => n42, B2 => 
                           regs(1791), ZN => n578);
   U758 : NAND3_X1 port map( A1 => n580, A2 => n579, A3 => n578, ZN => 
                           curr_proc_regs(255));
   U759 : NAND2_X1 port map( A1 => regs(768), A2 => n3, ZN => n583);
   U760 : AOI22_X1 port map( A1 => n32, A2 => regs(1280), B1 => n21, B2 => 
                           regs(256), ZN => n582);
   U761 : AOI22_X1 port map( A1 => n57, A2 => regs(2304), B1 => n42, B2 => 
                           regs(1792), ZN => n581);
   U762 : NAND3_X1 port map( A1 => n583, A2 => n582, A3 => n581, ZN => 
                           curr_proc_regs(256));
   U763 : NAND2_X1 port map( A1 => regs(769), A2 => n16, ZN => n586);
   U764 : AOI22_X1 port map( A1 => n32, A2 => regs(1281), B1 => n26, B2 => 
                           regs(257), ZN => n585);
   U765 : AOI22_X1 port map( A1 => n57, A2 => regs(2305), B1 => n42, B2 => 
                           regs(1793), ZN => n584);
   U766 : NAND3_X1 port map( A1 => n586, A2 => n585, A3 => n584, ZN => 
                           curr_proc_regs(257));
   U767 : NAND2_X1 port map( A1 => regs(770), A2 => n3, ZN => n589);
   U768 : AOI22_X1 port map( A1 => n32, A2 => regs(1282), B1 => n26, B2 => 
                           regs(258), ZN => n588);
   U769 : AOI22_X1 port map( A1 => n57, A2 => regs(2306), B1 => n42, B2 => 
                           regs(1794), ZN => n587);
   U770 : NAND3_X1 port map( A1 => n589, A2 => n588, A3 => n587, ZN => 
                           curr_proc_regs(258));
   U771 : NAND2_X1 port map( A1 => regs(771), A2 => n3, ZN => n592);
   U772 : AOI22_X1 port map( A1 => n31, A2 => regs(1283), B1 => n21, B2 => 
                           regs(259), ZN => n591);
   U773 : AOI22_X1 port map( A1 => n57, A2 => regs(2307), B1 => n42, B2 => 
                           regs(1795), ZN => n590);
   U774 : NAND3_X1 port map( A1 => n592, A2 => n591, A3 => n590, ZN => 
                           curr_proc_regs(259));
   U775 : NAND2_X1 port map( A1 => regs(537), A2 => n16, ZN => n595);
   U776 : AOI22_X1 port map( A1 => n31, A2 => regs(1049), B1 => n26, B2 => 
                           regs(25), ZN => n594);
   U777 : AOI22_X1 port map( A1 => n57, A2 => regs(2073), B1 => n42, B2 => 
                           regs(1561), ZN => n593);
   U778 : NAND3_X1 port map( A1 => n595, A2 => n594, A3 => n593, ZN => 
                           curr_proc_regs(25));
   U779 : NAND2_X1 port map( A1 => regs(772), A2 => n3, ZN => n598);
   U780 : AOI22_X1 port map( A1 => n31, A2 => regs(1284), B1 => n26, B2 => 
                           regs(260), ZN => n597);
   U781 : AOI22_X1 port map( A1 => n57, A2 => regs(2308), B1 => n42, B2 => 
                           regs(1796), ZN => n596);
   U782 : NAND3_X1 port map( A1 => n598, A2 => n597, A3 => n596, ZN => 
                           curr_proc_regs(260));
   U783 : NAND2_X1 port map( A1 => regs(773), A2 => n3, ZN => n601);
   U784 : AOI22_X1 port map( A1 => n31, A2 => regs(1285), B1 => n21, B2 => 
                           regs(261), ZN => n600);
   U785 : AOI22_X1 port map( A1 => n57, A2 => regs(2309), B1 => n42, B2 => 
                           regs(1797), ZN => n599);
   U786 : NAND3_X1 port map( A1 => n601, A2 => n600, A3 => n599, ZN => 
                           curr_proc_regs(261));
   U787 : NAND2_X1 port map( A1 => regs(774), A2 => n16, ZN => n604);
   U788 : AOI22_X1 port map( A1 => n31, A2 => regs(1286), B1 => n26, B2 => 
                           regs(262), ZN => n603);
   U789 : AOI22_X1 port map( A1 => n57, A2 => regs(2310), B1 => n42, B2 => 
                           regs(1798), ZN => n602);
   U790 : NAND3_X1 port map( A1 => n604, A2 => n603, A3 => n602, ZN => 
                           curr_proc_regs(262));
   U791 : NAND2_X1 port map( A1 => regs(775), A2 => n16, ZN => n607);
   U792 : AOI22_X1 port map( A1 => n31, A2 => regs(1287), B1 => n26, B2 => 
                           regs(263), ZN => n606);
   U793 : AOI22_X1 port map( A1 => n57, A2 => regs(2311), B1 => n42, B2 => 
                           regs(1799), ZN => n605);
   U794 : NAND3_X1 port map( A1 => n607, A2 => n606, A3 => n605, ZN => 
                           curr_proc_regs(263));
   U795 : NAND2_X1 port map( A1 => regs(776), A2 => n16, ZN => n610);
   U796 : AOI22_X1 port map( A1 => n31, A2 => regs(1288), B1 => n26, B2 => 
                           regs(264), ZN => n609);
   U797 : AOI22_X1 port map( A1 => n57, A2 => regs(2312), B1 => n42, B2 => 
                           regs(1800), ZN => n608);
   U798 : NAND3_X1 port map( A1 => n610, A2 => n609, A3 => n608, ZN => 
                           curr_proc_regs(264));
   U799 : NAND2_X1 port map( A1 => regs(777), A2 => n16, ZN => n613);
   U800 : AOI22_X1 port map( A1 => n31, A2 => regs(1289), B1 => n26, B2 => 
                           regs(265), ZN => n612);
   U801 : AOI22_X1 port map( A1 => n57, A2 => regs(2313), B1 => n42, B2 => 
                           regs(1801), ZN => n611);
   U802 : NAND3_X1 port map( A1 => n613, A2 => n612, A3 => n611, ZN => 
                           curr_proc_regs(265));
   U803 : NAND2_X1 port map( A1 => regs(778), A2 => n16, ZN => n616);
   U804 : AOI22_X1 port map( A1 => n31, A2 => regs(1290), B1 => n26, B2 => 
                           regs(266), ZN => n615);
   U805 : AOI22_X1 port map( A1 => n57, A2 => regs(2314), B1 => n42, B2 => 
                           regs(1802), ZN => n614);
   U806 : NAND3_X1 port map( A1 => n616, A2 => n615, A3 => n614, ZN => 
                           curr_proc_regs(266));
   U807 : NAND2_X1 port map( A1 => regs(779), A2 => n16, ZN => n619);
   U808 : AOI22_X1 port map( A1 => n31, A2 => regs(1291), B1 => n26, B2 => 
                           regs(267), ZN => n618);
   U809 : AOI22_X1 port map( A1 => win(4), A2 => regs(2315), B1 => n42, B2 => 
                           regs(1803), ZN => n617);
   U810 : NAND3_X1 port map( A1 => n619, A2 => n618, A3 => n617, ZN => 
                           curr_proc_regs(267));
   U811 : NAND2_X1 port map( A1 => regs(780), A2 => n16, ZN => n622);
   U812 : AOI22_X1 port map( A1 => n31, A2 => regs(1292), B1 => n26, B2 => 
                           regs(268), ZN => n621);
   U813 : AOI22_X1 port map( A1 => win(4), A2 => regs(2316), B1 => n42, B2 => 
                           regs(1804), ZN => n620);
   U814 : NAND3_X1 port map( A1 => n622, A2 => n621, A3 => n620, ZN => 
                           curr_proc_regs(268));
   U815 : NAND2_X1 port map( A1 => regs(781), A2 => n3, ZN => n625);
   U816 : AOI22_X1 port map( A1 => n31, A2 => regs(1293), B1 => n26, B2 => 
                           regs(269), ZN => n624);
   U817 : AOI22_X1 port map( A1 => win(4), A2 => regs(2317), B1 => n42, B2 => 
                           regs(1805), ZN => n623);
   U818 : NAND3_X1 port map( A1 => n625, A2 => n624, A3 => n623, ZN => 
                           curr_proc_regs(269));
   U819 : NAND2_X1 port map( A1 => regs(538), A2 => n16, ZN => n628);
   U820 : AOI22_X1 port map( A1 => n31, A2 => regs(1050), B1 => n26, B2 => 
                           regs(26), ZN => n627);
   U821 : AOI22_X1 port map( A1 => win(4), A2 => regs(2074), B1 => n42, B2 => 
                           regs(1562), ZN => n626);
   U822 : NAND3_X1 port map( A1 => n628, A2 => n627, A3 => n626, ZN => 
                           curr_proc_regs(26));
   U823 : NAND2_X1 port map( A1 => regs(782), A2 => n3, ZN => n631);
   U824 : AOI22_X1 port map( A1 => n31, A2 => regs(1294), B1 => n26, B2 => 
                           regs(270), ZN => n630);
   U825 : AOI22_X1 port map( A1 => win(4), A2 => regs(2318), B1 => n42, B2 => 
                           regs(1806), ZN => n629);
   U826 : NAND3_X1 port map( A1 => n631, A2 => n630, A3 => n629, ZN => 
                           curr_proc_regs(270));
   U827 : NAND2_X1 port map( A1 => regs(783), A2 => n16, ZN => n634);
   U828 : AOI22_X1 port map( A1 => n31, A2 => regs(1295), B1 => n26, B2 => 
                           regs(271), ZN => n633);
   U829 : AOI22_X1 port map( A1 => win(4), A2 => regs(2319), B1 => n42, B2 => 
                           regs(1807), ZN => n632);
   U830 : NAND3_X1 port map( A1 => n634, A2 => n633, A3 => n632, ZN => 
                           curr_proc_regs(271));
   U831 : NAND2_X1 port map( A1 => regs(784), A2 => n3, ZN => n637);
   U832 : AOI22_X1 port map( A1 => n31, A2 => regs(1296), B1 => n26, B2 => 
                           regs(272), ZN => n636);
   U833 : AOI22_X1 port map( A1 => win(4), A2 => regs(2320), B1 => n42, B2 => 
                           regs(1808), ZN => n635);
   U834 : NAND3_X1 port map( A1 => n637, A2 => n636, A3 => n635, ZN => 
                           curr_proc_regs(272));
   U835 : NAND2_X1 port map( A1 => regs(785), A2 => n3, ZN => n640);
   U836 : AOI22_X1 port map( A1 => n31, A2 => regs(1297), B1 => n21, B2 => 
                           regs(273), ZN => n639);
   U837 : AOI22_X1 port map( A1 => win(4), A2 => regs(2321), B1 => n42, B2 => 
                           regs(1809), ZN => n638);
   U838 : NAND3_X1 port map( A1 => n640, A2 => n639, A3 => n638, ZN => 
                           curr_proc_regs(273));
   U839 : NAND2_X1 port map( A1 => regs(786), A2 => n16, ZN => n643);
   U840 : AOI22_X1 port map( A1 => n31, A2 => regs(1298), B1 => n26, B2 => 
                           regs(274), ZN => n642);
   U841 : AOI22_X1 port map( A1 => win(4), A2 => regs(2322), B1 => n42, B2 => 
                           regs(1810), ZN => n641);
   U842 : NAND3_X1 port map( A1 => n643, A2 => n642, A3 => n641, ZN => 
                           curr_proc_regs(274));
   U843 : NAND2_X1 port map( A1 => regs(787), A2 => n3, ZN => n646);
   U844 : AOI22_X1 port map( A1 => n31, A2 => regs(1299), B1 => n26, B2 => 
                           regs(275), ZN => n645);
   U845 : AOI22_X1 port map( A1 => win(4), A2 => regs(2323), B1 => n42, B2 => 
                           regs(1811), ZN => n644);
   U846 : NAND3_X1 port map( A1 => n646, A2 => n645, A3 => n644, ZN => 
                           curr_proc_regs(275));
   U847 : NAND2_X1 port map( A1 => regs(788), A2 => n3, ZN => n649);
   U848 : AOI22_X1 port map( A1 => n31, A2 => regs(1300), B1 => n26, B2 => 
                           regs(276), ZN => n648);
   U849 : AOI22_X1 port map( A1 => win(4), A2 => regs(2324), B1 => n42, B2 => 
                           regs(1812), ZN => n647);
   U850 : NAND3_X1 port map( A1 => n649, A2 => n648, A3 => n647, ZN => 
                           curr_proc_regs(276));
   U851 : NAND2_X1 port map( A1 => regs(789), A2 => n3, ZN => n652);
   U852 : AOI22_X1 port map( A1 => n31, A2 => regs(1301), B1 => n21, B2 => 
                           regs(277), ZN => n651);
   U853 : AOI22_X1 port map( A1 => n56, A2 => regs(2325), B1 => n42, B2 => 
                           regs(1813), ZN => n650);
   U854 : NAND3_X1 port map( A1 => n652, A2 => n651, A3 => n650, ZN => 
                           curr_proc_regs(277));
   U855 : NAND2_X1 port map( A1 => regs(790), A2 => n16, ZN => n655);
   U856 : AOI22_X1 port map( A1 => n31, A2 => regs(1302), B1 => n26, B2 => 
                           regs(278), ZN => n654);
   U857 : AOI22_X1 port map( A1 => n56, A2 => regs(2326), B1 => n42, B2 => 
                           regs(1814), ZN => n653);
   U858 : NAND3_X1 port map( A1 => n655, A2 => n654, A3 => n653, ZN => 
                           curr_proc_regs(278));
   U859 : NAND2_X1 port map( A1 => regs(791), A2 => n3, ZN => n658);
   U860 : AOI22_X1 port map( A1 => n31, A2 => regs(1303), B1 => n26, B2 => 
                           regs(279), ZN => n657);
   U861 : AOI22_X1 port map( A1 => n56, A2 => regs(2327), B1 => n42, B2 => 
                           regs(1815), ZN => n656);
   U862 : NAND3_X1 port map( A1 => n658, A2 => n657, A3 => n656, ZN => 
                           curr_proc_regs(279));
   U863 : NAND2_X1 port map( A1 => regs(539), A2 => n3, ZN => n661);
   U864 : AOI22_X1 port map( A1 => n31, A2 => regs(1051), B1 => n26, B2 => 
                           regs(27), ZN => n660);
   U865 : AOI22_X1 port map( A1 => n56, A2 => regs(2075), B1 => n42, B2 => 
                           regs(1563), ZN => n659);
   U866 : NAND3_X1 port map( A1 => n661, A2 => n660, A3 => n659, ZN => 
                           curr_proc_regs(27));
   U867 : NAND2_X1 port map( A1 => regs(792), A2 => n3, ZN => n664);
   U868 : AOI22_X1 port map( A1 => n29, A2 => regs(1304), B1 => n21, B2 => 
                           regs(280), ZN => n663);
   U869 : AOI22_X1 port map( A1 => n56, A2 => regs(2328), B1 => n42, B2 => 
                           regs(1816), ZN => n662);
   U870 : NAND3_X1 port map( A1 => n664, A2 => n663, A3 => n662, ZN => 
                           curr_proc_regs(280));
   U871 : NAND2_X1 port map( A1 => regs(793), A2 => n3, ZN => n667);
   U872 : AOI22_X1 port map( A1 => n33, A2 => regs(1305), B1 => n26, B2 => 
                           regs(281), ZN => n666);
   U873 : AOI22_X1 port map( A1 => n56, A2 => regs(2329), B1 => n42, B2 => 
                           regs(1817), ZN => n665);
   U874 : NAND3_X1 port map( A1 => n667, A2 => n666, A3 => n665, ZN => 
                           curr_proc_regs(281));
   U875 : NAND2_X1 port map( A1 => regs(794), A2 => n3, ZN => n670);
   U876 : AOI22_X1 port map( A1 => n31, A2 => regs(1306), B1 => n26, B2 => 
                           regs(282), ZN => n669);
   U877 : AOI22_X1 port map( A1 => n56, A2 => regs(2330), B1 => n42, B2 => 
                           regs(1818), ZN => n668);
   U878 : NAND3_X1 port map( A1 => n670, A2 => n669, A3 => n668, ZN => 
                           curr_proc_regs(282));
   U879 : NAND2_X1 port map( A1 => regs(795), A2 => n3, ZN => n673);
   U880 : AOI22_X1 port map( A1 => n31, A2 => regs(1307), B1 => n26, B2 => 
                           regs(283), ZN => n672);
   U881 : AOI22_X1 port map( A1 => n56, A2 => regs(2331), B1 => n42, B2 => 
                           regs(1819), ZN => n671);
   U882 : NAND3_X1 port map( A1 => n673, A2 => n672, A3 => n671, ZN => 
                           curr_proc_regs(283));
   U883 : NAND2_X1 port map( A1 => regs(796), A2 => n16, ZN => n676);
   U884 : AOI22_X1 port map( A1 => n30, A2 => regs(1308), B1 => n26, B2 => 
                           regs(284), ZN => n675);
   U885 : AOI22_X1 port map( A1 => n56, A2 => regs(2332), B1 => n42, B2 => 
                           regs(1820), ZN => n674);
   U886 : NAND3_X1 port map( A1 => n676, A2 => n675, A3 => n674, ZN => 
                           curr_proc_regs(284));
   U887 : NAND2_X1 port map( A1 => regs(797), A2 => n3, ZN => n679);
   U888 : AOI22_X1 port map( A1 => n29, A2 => regs(1309), B1 => n26, B2 => 
                           regs(285), ZN => n678);
   U889 : AOI22_X1 port map( A1 => n56, A2 => regs(2333), B1 => n42, B2 => 
                           regs(1821), ZN => n677);
   U890 : NAND3_X1 port map( A1 => n679, A2 => n678, A3 => n677, ZN => 
                           curr_proc_regs(285));
   U891 : NAND2_X1 port map( A1 => regs(798), A2 => n3, ZN => n682);
   U892 : AOI22_X1 port map( A1 => n31, A2 => regs(1310), B1 => n26, B2 => 
                           regs(286), ZN => n681);
   U893 : AOI22_X1 port map( A1 => n56, A2 => regs(2334), B1 => n42, B2 => 
                           regs(1822), ZN => n680);
   U894 : NAND3_X1 port map( A1 => n682, A2 => n681, A3 => n680, ZN => 
                           curr_proc_regs(286));
   U895 : NAND2_X1 port map( A1 => regs(799), A2 => n3, ZN => n685);
   U896 : AOI22_X1 port map( A1 => n30, A2 => regs(1311), B1 => n26, B2 => 
                           regs(287), ZN => n684);
   U897 : AOI22_X1 port map( A1 => n56, A2 => regs(2335), B1 => n42, B2 => 
                           regs(1823), ZN => n683);
   U898 : NAND3_X1 port map( A1 => n685, A2 => n684, A3 => n683, ZN => 
                           curr_proc_regs(287));
   U899 : NAND2_X1 port map( A1 => regs(800), A2 => n3, ZN => n688);
   U900 : AOI22_X1 port map( A1 => n33, A2 => regs(1312), B1 => n21, B2 => 
                           regs(288), ZN => n687);
   U901 : AOI22_X1 port map( A1 => n5, A2 => regs(2336), B1 => n42, B2 => 
                           regs(1824), ZN => n686);
   U902 : NAND3_X1 port map( A1 => n688, A2 => n687, A3 => n686, ZN => 
                           curr_proc_regs(288));
   U903 : NAND2_X1 port map( A1 => regs(801), A2 => n3, ZN => n691);
   U904 : AOI22_X1 port map( A1 => n31, A2 => regs(1313), B1 => n26, B2 => 
                           regs(289), ZN => n690);
   U905 : AOI22_X1 port map( A1 => n5, A2 => regs(2337), B1 => n42, B2 => 
                           regs(1825), ZN => n689);
   U906 : NAND3_X1 port map( A1 => n691, A2 => n690, A3 => n689, ZN => 
                           curr_proc_regs(289));
   U907 : NAND2_X1 port map( A1 => regs(540), A2 => n3, ZN => n694);
   U908 : AOI22_X1 port map( A1 => n30, A2 => regs(1052), B1 => n26, B2 => 
                           regs(28), ZN => n693);
   U909 : AOI22_X1 port map( A1 => n5, A2 => regs(2076), B1 => n42, B2 => 
                           regs(1564), ZN => n692);
   U910 : NAND3_X1 port map( A1 => n694, A2 => n693, A3 => n692, ZN => 
                           curr_proc_regs(28));
   U911 : NAND2_X1 port map( A1 => regs(802), A2 => n3, ZN => n697);
   U912 : AOI22_X1 port map( A1 => n29, A2 => regs(1314), B1 => n26, B2 => 
                           regs(290), ZN => n696);
   U913 : AOI22_X1 port map( A1 => n5, A2 => regs(2338), B1 => n42, B2 => 
                           regs(1826), ZN => n695);
   U914 : NAND3_X1 port map( A1 => n697, A2 => n696, A3 => n695, ZN => 
                           curr_proc_regs(290));
   U915 : NAND2_X1 port map( A1 => regs(803), A2 => n3, ZN => n700);
   U916 : AOI22_X1 port map( A1 => n33, A2 => regs(1315), B1 => n26, B2 => 
                           regs(291), ZN => n699);
   U917 : AOI22_X1 port map( A1 => n5, A2 => regs(2339), B1 => n42, B2 => 
                           regs(1827), ZN => n698);
   U918 : NAND3_X1 port map( A1 => n700, A2 => n699, A3 => n698, ZN => 
                           curr_proc_regs(291));
   U919 : NAND2_X1 port map( A1 => regs(804), A2 => n3, ZN => n703);
   U920 : AOI22_X1 port map( A1 => n29, A2 => regs(1316), B1 => n26, B2 => 
                           regs(292), ZN => n702);
   U921 : AOI22_X1 port map( A1 => n5, A2 => regs(2340), B1 => n42, B2 => 
                           regs(1828), ZN => n701);
   U922 : NAND3_X1 port map( A1 => n703, A2 => n702, A3 => n701, ZN => 
                           curr_proc_regs(292));
   U923 : NAND2_X1 port map( A1 => regs(805), A2 => n3, ZN => n706);
   U924 : AOI22_X1 port map( A1 => n31, A2 => regs(1317), B1 => n26, B2 => 
                           regs(293), ZN => n705);
   U925 : AOI22_X1 port map( A1 => n5, A2 => regs(2341), B1 => n42, B2 => 
                           regs(1829), ZN => n704);
   U926 : NAND3_X1 port map( A1 => n706, A2 => n705, A3 => n704, ZN => 
                           curr_proc_regs(293));
   U927 : NAND2_X1 port map( A1 => regs(806), A2 => n3, ZN => n709);
   U928 : AOI22_X1 port map( A1 => n31, A2 => regs(1318), B1 => n26, B2 => 
                           regs(294), ZN => n708);
   U929 : AOI22_X1 port map( A1 => n5, A2 => regs(2342), B1 => n42, B2 => 
                           regs(1830), ZN => n707);
   U930 : NAND3_X1 port map( A1 => n709, A2 => n708, A3 => n707, ZN => 
                           curr_proc_regs(294));
   U931 : NAND2_X1 port map( A1 => regs(807), A2 => n15, ZN => n712);
   U932 : AOI22_X1 port map( A1 => n29, A2 => regs(1319), B1 => n20, B2 => 
                           regs(295), ZN => n711);
   U933 : AOI22_X1 port map( A1 => n5, A2 => regs(2343), B1 => n38, B2 => 
                           regs(1831), ZN => n710);
   U934 : NAND3_X1 port map( A1 => n712, A2 => n711, A3 => n710, ZN => 
                           curr_proc_regs(295));
   U935 : NAND2_X1 port map( A1 => regs(808), A2 => n15, ZN => n715);
   U936 : AOI22_X1 port map( A1 => n31, A2 => regs(1320), B1 => n20, B2 => 
                           regs(296), ZN => n714);
   U937 : AOI22_X1 port map( A1 => n5, A2 => regs(2344), B1 => n39, B2 => 
                           regs(1832), ZN => n713);
   U938 : NAND3_X1 port map( A1 => n715, A2 => n714, A3 => n713, ZN => 
                           curr_proc_regs(296));
   U939 : NAND2_X1 port map( A1 => regs(809), A2 => n15, ZN => n718);
   U940 : AOI22_X1 port map( A1 => n30, A2 => regs(1321), B1 => n25, B2 => 
                           regs(297), ZN => n717);
   U941 : AOI22_X1 port map( A1 => n5, A2 => regs(2345), B1 => n36, B2 => 
                           regs(1833), ZN => n716);
   U942 : NAND3_X1 port map( A1 => n718, A2 => n717, A3 => n716, ZN => 
                           curr_proc_regs(297));
   U943 : NAND2_X1 port map( A1 => regs(810), A2 => n15, ZN => n721);
   U944 : AOI22_X1 port map( A1 => n30, A2 => regs(1322), B1 => n21, B2 => 
                           regs(298), ZN => n720);
   U945 : AOI22_X1 port map( A1 => n5, A2 => regs(2346), B1 => n35, B2 => 
                           regs(1834), ZN => n719);
   U946 : NAND3_X1 port map( A1 => n721, A2 => n720, A3 => n719, ZN => 
                           curr_proc_regs(298));
   U947 : NAND2_X1 port map( A1 => regs(811), A2 => n15, ZN => n724);
   U948 : AOI22_X1 port map( A1 => n31, A2 => regs(1323), B1 => n25, B2 => 
                           regs(299), ZN => n723);
   U949 : AOI22_X1 port map( A1 => n48, A2 => regs(2347), B1 => n36, B2 => 
                           regs(1835), ZN => n722);
   U950 : NAND3_X1 port map( A1 => n724, A2 => n723, A3 => n722, ZN => 
                           curr_proc_regs(299));
   U951 : NAND2_X1 port map( A1 => regs(541), A2 => n15, ZN => n727);
   U952 : AOI22_X1 port map( A1 => n29, A2 => regs(1053), B1 => n21, B2 => 
                           regs(29), ZN => n726);
   U953 : AOI22_X1 port map( A1 => n54, A2 => regs(2077), B1 => n34, B2 => 
                           regs(1565), ZN => n725);
   U954 : NAND3_X1 port map( A1 => n727, A2 => n726, A3 => n725, ZN => 
                           curr_proc_regs(29));
   U955 : NAND2_X1 port map( A1 => regs(514), A2 => n15, ZN => n730);
   U956 : AOI22_X1 port map( A1 => n33, A2 => regs(1026), B1 => n25, B2 => 
                           regs(2), ZN => n729);
   U957 : AOI22_X1 port map( A1 => n51, A2 => regs(2050), B1 => n36, B2 => 
                           regs(1538), ZN => n728);
   U958 : NAND3_X1 port map( A1 => n730, A2 => n729, A3 => n728, ZN => 
                           curr_proc_regs(2));
   U959 : NAND2_X1 port map( A1 => regs(812), A2 => n15, ZN => n733);
   U960 : AOI22_X1 port map( A1 => n31, A2 => regs(1324), B1 => n23, B2 => 
                           regs(300), ZN => n732);
   U961 : AOI22_X1 port map( A1 => n5, A2 => regs(2348), B1 => n37, B2 => 
                           regs(1836), ZN => n731);
   U962 : NAND3_X1 port map( A1 => n733, A2 => n732, A3 => n731, ZN => 
                           curr_proc_regs(300));
   U963 : NAND2_X1 port map( A1 => regs(813), A2 => n15, ZN => n736);
   U964 : AOI22_X1 port map( A1 => n33, A2 => regs(1325), B1 => n25, B2 => 
                           regs(301), ZN => n735);
   U965 : AOI22_X1 port map( A1 => n47, A2 => regs(2349), B1 => n36, B2 => 
                           regs(1837), ZN => n734);
   U966 : NAND3_X1 port map( A1 => n736, A2 => n735, A3 => n734, ZN => 
                           curr_proc_regs(301));
   U967 : NAND2_X1 port map( A1 => regs(814), A2 => n15, ZN => n739);
   U968 : AOI22_X1 port map( A1 => n33, A2 => regs(1326), B1 => n25, B2 => 
                           regs(302), ZN => n738);
   U969 : AOI22_X1 port map( A1 => n6, A2 => regs(2350), B1 => n36, B2 => 
                           regs(1838), ZN => n737);
   U970 : NAND3_X1 port map( A1 => n739, A2 => n738, A3 => n737, ZN => 
                           curr_proc_regs(302));
   U971 : NAND2_X1 port map( A1 => regs(815), A2 => n15, ZN => n742);
   U972 : AOI22_X1 port map( A1 => n31, A2 => regs(1327), B1 => n25, B2 => 
                           regs(303), ZN => n741);
   U973 : AOI22_X1 port map( A1 => n7, A2 => regs(2351), B1 => n36, B2 => 
                           regs(1839), ZN => n740);
   U974 : NAND3_X1 port map( A1 => n742, A2 => n741, A3 => n740, ZN => 
                           curr_proc_regs(303));
   U975 : NAND2_X1 port map( A1 => regs(816), A2 => n15, ZN => n745);
   U976 : AOI22_X1 port map( A1 => n31, A2 => regs(1328), B1 => n25, B2 => 
                           regs(304), ZN => n744);
   U977 : AOI22_X1 port map( A1 => n8, A2 => regs(2352), B1 => n36, B2 => 
                           regs(1840), ZN => n743);
   U978 : NAND3_X1 port map( A1 => n745, A2 => n744, A3 => n743, ZN => 
                           curr_proc_regs(304));
   U979 : NAND2_X1 port map( A1 => regs(817), A2 => n10, ZN => n748);
   U980 : AOI22_X1 port map( A1 => n31, A2 => regs(1329), B1 => n26, B2 => 
                           regs(305), ZN => n747);
   U981 : AOI22_X1 port map( A1 => n43, A2 => regs(2353), B1 => n38, B2 => 
                           regs(1841), ZN => n746);
   U982 : NAND3_X1 port map( A1 => n748, A2 => n747, A3 => n746, ZN => 
                           curr_proc_regs(305));
   U983 : NAND2_X1 port map( A1 => regs(818), A2 => n15, ZN => n751);
   U984 : AOI22_X1 port map( A1 => n30, A2 => regs(1330), B1 => n25, B2 => 
                           regs(306), ZN => n750);
   U985 : AOI22_X1 port map( A1 => n46, A2 => regs(2354), B1 => n36, B2 => 
                           regs(1842), ZN => n749);
   U986 : NAND3_X1 port map( A1 => n751, A2 => n750, A3 => n749, ZN => 
                           curr_proc_regs(306));
   U987 : NAND2_X1 port map( A1 => regs(819), A2 => n15, ZN => n754);
   U988 : AOI22_X1 port map( A1 => n33, A2 => regs(1331), B1 => n19, B2 => 
                           regs(307), ZN => n753);
   U989 : AOI22_X1 port map( A1 => n50, A2 => regs(2355), B1 => n39, B2 => 
                           regs(1843), ZN => n752);
   U990 : NAND3_X1 port map( A1 => n754, A2 => n753, A3 => n752, ZN => 
                           curr_proc_regs(307));
   U991 : NAND2_X1 port map( A1 => regs(820), A2 => n10, ZN => n757);
   U992 : AOI22_X1 port map( A1 => n33, A2 => regs(1332), B1 => n21, B2 => 
                           regs(308), ZN => n756);
   U993 : AOI22_X1 port map( A1 => n44, A2 => regs(2356), B1 => n38, B2 => 
                           regs(1844), ZN => n755);
   U994 : NAND3_X1 port map( A1 => n757, A2 => n756, A3 => n755, ZN => 
                           curr_proc_regs(308));
   U995 : NAND2_X1 port map( A1 => regs(821), A2 => n15, ZN => n760);
   U996 : AOI22_X1 port map( A1 => n31, A2 => regs(1333), B1 => n25, B2 => 
                           regs(309), ZN => n759);
   U997 : AOI22_X1 port map( A1 => n55, A2 => regs(2357), B1 => n36, B2 => 
                           regs(1845), ZN => n758);
   U998 : NAND3_X1 port map( A1 => n760, A2 => n759, A3 => n758, ZN => 
                           curr_proc_regs(309));
   U999 : NAND2_X1 port map( A1 => regs(542), A2 => n15, ZN => n763);
   U1000 : AOI22_X1 port map( A1 => n31, A2 => regs(1054), B1 => n1596, B2 => 
                           regs(30), ZN => n762);
   U1001 : AOI22_X1 port map( A1 => n55, A2 => regs(2078), B1 => n39, B2 => 
                           regs(1566), ZN => n761);
   U1002 : NAND3_X1 port map( A1 => n763, A2 => n762, A3 => n761, ZN => 
                           curr_proc_regs(30));
   U1003 : NAND2_X1 port map( A1 => regs(822), A2 => n10, ZN => n766);
   U1004 : AOI22_X1 port map( A1 => n30, A2 => regs(1334), B1 => n17, B2 => 
                           regs(310), ZN => n765);
   U1005 : AOI22_X1 port map( A1 => n55, A2 => regs(2358), B1 => n38, B2 => 
                           regs(1846), ZN => n764);
   U1006 : NAND3_X1 port map( A1 => n766, A2 => n765, A3 => n764, ZN => 
                           curr_proc_regs(310));
   U1007 : NAND2_X1 port map( A1 => regs(823), A2 => n15, ZN => n769);
   U1008 : AOI22_X1 port map( A1 => n31, A2 => regs(1335), B1 => n25, B2 => 
                           regs(311), ZN => n768);
   U1009 : AOI22_X1 port map( A1 => n55, A2 => regs(2359), B1 => n36, B2 => 
                           regs(1847), ZN => n767);
   U1010 : NAND3_X1 port map( A1 => n769, A2 => n768, A3 => n767, ZN => 
                           curr_proc_regs(311));
   U1011 : NAND2_X1 port map( A1 => regs(824), A2 => n15, ZN => n772);
   U1012 : AOI22_X1 port map( A1 => n33, A2 => regs(1336), B1 => n20, B2 => 
                           regs(312), ZN => n771);
   U1013 : AOI22_X1 port map( A1 => n55, A2 => regs(2360), B1 => n39, B2 => 
                           regs(1848), ZN => n770);
   U1014 : NAND3_X1 port map( A1 => n772, A2 => n771, A3 => n770, ZN => 
                           curr_proc_regs(312));
   U1015 : NAND2_X1 port map( A1 => regs(825), A2 => n10, ZN => n775);
   U1016 : AOI22_X1 port map( A1 => n33, A2 => regs(1337), B1 => n26, B2 => 
                           regs(313), ZN => n774);
   U1017 : AOI22_X1 port map( A1 => n55, A2 => regs(2361), B1 => n38, B2 => 
                           regs(1849), ZN => n773);
   U1018 : NAND3_X1 port map( A1 => n775, A2 => n774, A3 => n773, ZN => 
                           curr_proc_regs(313));
   U1019 : NAND2_X1 port map( A1 => regs(826), A2 => n15, ZN => n778);
   U1020 : AOI22_X1 port map( A1 => n33, A2 => regs(1338), B1 => n25, B2 => 
                           regs(314), ZN => n777);
   U1021 : AOI22_X1 port map( A1 => n55, A2 => regs(2362), B1 => n36, B2 => 
                           regs(1850), ZN => n776);
   U1022 : NAND3_X1 port map( A1 => n778, A2 => n777, A3 => n776, ZN => 
                           curr_proc_regs(314));
   U1023 : NAND2_X1 port map( A1 => regs(827), A2 => n15, ZN => n781);
   U1024 : AOI22_X1 port map( A1 => n33, A2 => regs(1339), B1 => n18, B2 => 
                           regs(315), ZN => n780);
   U1025 : AOI22_X1 port map( A1 => n55, A2 => regs(2363), B1 => n42, B2 => 
                           regs(1851), ZN => n779);
   U1026 : NAND3_X1 port map( A1 => n781, A2 => n780, A3 => n779, ZN => 
                           curr_proc_regs(315));
   U1027 : NAND2_X1 port map( A1 => regs(828), A2 => n10, ZN => n784);
   U1028 : AOI22_X1 port map( A1 => n31, A2 => regs(1340), B1 => n21, B2 => 
                           regs(316), ZN => n783);
   U1029 : AOI22_X1 port map( A1 => n55, A2 => regs(2364), B1 => n1598, B2 => 
                           regs(1852), ZN => n782);
   U1030 : NAND3_X1 port map( A1 => n784, A2 => n783, A3 => n782, ZN => 
                           curr_proc_regs(316));
   U1031 : NAND2_X1 port map( A1 => regs(829), A2 => n10, ZN => n787);
   U1032 : AOI22_X1 port map( A1 => n31, A2 => regs(1341), B1 => n1596, B2 => 
                           regs(317), ZN => n786);
   U1033 : AOI22_X1 port map( A1 => n55, A2 => regs(2365), B1 => n36, B2 => 
                           regs(1853), ZN => n785);
   U1034 : NAND3_X1 port map( A1 => n787, A2 => n786, A3 => n785, ZN => 
                           curr_proc_regs(317));
   U1035 : NAND2_X1 port map( A1 => regs(830), A2 => n10, ZN => n790);
   U1036 : AOI22_X1 port map( A1 => n31, A2 => regs(1342), B1 => n19, B2 => 
                           regs(318), ZN => n789);
   U1037 : AOI22_X1 port map( A1 => n55, A2 => regs(2366), B1 => n35, B2 => 
                           regs(1854), ZN => n788);
   U1038 : NAND3_X1 port map( A1 => n790, A2 => n789, A3 => n788, ZN => 
                           curr_proc_regs(318));
   U1039 : NAND2_X1 port map( A1 => regs(831), A2 => n10, ZN => n793);
   U1040 : AOI22_X1 port map( A1 => n29, A2 => regs(1343), B1 => n19, B2 => 
                           regs(319), ZN => n792);
   U1041 : AOI22_X1 port map( A1 => n55, A2 => regs(2367), B1 => n42, B2 => 
                           regs(1855), ZN => n791);
   U1042 : NAND3_X1 port map( A1 => n793, A2 => n792, A3 => n791, ZN => 
                           curr_proc_regs(319));
   U1043 : NAND2_X1 port map( A1 => regs(543), A2 => n10, ZN => n796);
   U1044 : AOI22_X1 port map( A1 => n33, A2 => regs(1055), B1 => n21, B2 => 
                           regs(31), ZN => n795);
   U1045 : AOI22_X1 port map( A1 => n48, A2 => regs(2079), B1 => n37, B2 => 
                           regs(1567), ZN => n794);
   U1046 : NAND3_X1 port map( A1 => n796, A2 => n795, A3 => n794, ZN => 
                           curr_proc_regs(31));
   U1047 : NAND2_X1 port map( A1 => regs(832), A2 => n10, ZN => n799);
   U1048 : AOI22_X1 port map( A1 => n31, A2 => regs(1344), B1 => n17, B2 => 
                           regs(320), ZN => n798);
   U1049 : AOI22_X1 port map( A1 => win(4), A2 => regs(2368), B1 => n34, B2 => 
                           regs(1856), ZN => n797);
   U1050 : NAND3_X1 port map( A1 => n799, A2 => n798, A3 => n797, ZN => 
                           curr_proc_regs(320));
   U1051 : NAND2_X1 port map( A1 => regs(833), A2 => n10, ZN => n802);
   U1052 : AOI22_X1 port map( A1 => n30, A2 => regs(1345), B1 => n17, B2 => 
                           regs(321), ZN => n801);
   U1053 : AOI22_X1 port map( A1 => n44, A2 => regs(2369), B1 => n40, B2 => 
                           regs(1857), ZN => n800);
   U1054 : NAND3_X1 port map( A1 => n802, A2 => n801, A3 => n800, ZN => 
                           curr_proc_regs(321));
   U1055 : NAND2_X1 port map( A1 => regs(834), A2 => n10, ZN => n805);
   U1056 : AOI22_X1 port map( A1 => n33, A2 => regs(1346), B1 => n20, B2 => 
                           regs(322), ZN => n804);
   U1057 : AOI22_X1 port map( A1 => n54, A2 => regs(2370), B1 => n39, B2 => 
                           regs(1858), ZN => n803);
   U1058 : NAND3_X1 port map( A1 => n805, A2 => n804, A3 => n803, ZN => 
                           curr_proc_regs(322));
   U1059 : NAND2_X1 port map( A1 => regs(835), A2 => n10, ZN => n808);
   U1060 : AOI22_X1 port map( A1 => n2, A2 => regs(1347), B1 => n1596, B2 => 
                           regs(323), ZN => n807);
   U1061 : AOI22_X1 port map( A1 => win(4), A2 => regs(2371), B1 => n38, B2 => 
                           regs(1859), ZN => n806);
   U1062 : NAND3_X1 port map( A1 => n808, A2 => n807, A3 => n806, ZN => 
                           curr_proc_regs(323));
   U1063 : NAND2_X1 port map( A1 => regs(836), A2 => n10, ZN => n811);
   U1064 : AOI22_X1 port map( A1 => n2, A2 => regs(1348), B1 => n1596, B2 => 
                           regs(324), ZN => n810);
   U1065 : AOI22_X1 port map( A1 => win(4), A2 => regs(2372), B1 => n1598, B2 
                           => regs(1860), ZN => n809);
   U1066 : NAND3_X1 port map( A1 => n811, A2 => n810, A3 => n809, ZN => 
                           curr_proc_regs(324));
   U1067 : NAND2_X1 port map( A1 => regs(837), A2 => n10, ZN => n814);
   U1068 : AOI22_X1 port map( A1 => n2, A2 => regs(1349), B1 => n1596, B2 => 
                           regs(325), ZN => n813);
   U1069 : AOI22_X1 port map( A1 => win(4), A2 => regs(2373), B1 => n1598, B2 
                           => regs(1861), ZN => n812);
   U1070 : NAND3_X1 port map( A1 => n814, A2 => n813, A3 => n812, ZN => 
                           curr_proc_regs(325));
   U1071 : NAND2_X1 port map( A1 => regs(838), A2 => n10, ZN => n817);
   U1072 : AOI22_X1 port map( A1 => n2, A2 => regs(1350), B1 => n1596, B2 => 
                           regs(326), ZN => n816);
   U1073 : AOI22_X1 port map( A1 => n51, A2 => regs(2374), B1 => n1598, B2 => 
                           regs(1862), ZN => n815);
   U1074 : NAND3_X1 port map( A1 => n817, A2 => n816, A3 => n815, ZN => 
                           curr_proc_regs(326));
   U1075 : NAND2_X1 port map( A1 => regs(839), A2 => n15, ZN => n820);
   U1076 : AOI22_X1 port map( A1 => n2, A2 => regs(1351), B1 => n19, B2 => 
                           regs(327), ZN => n819);
   U1077 : AOI22_X1 port map( A1 => n44, A2 => regs(2375), B1 => n38, B2 => 
                           regs(1863), ZN => n818);
   U1078 : NAND3_X1 port map( A1 => n820, A2 => n819, A3 => n818, ZN => 
                           curr_proc_regs(327));
   U1079 : NAND2_X1 port map( A1 => regs(840), A2 => n10, ZN => n823);
   U1080 : AOI22_X1 port map( A1 => n2, A2 => regs(1352), B1 => n19, B2 => 
                           regs(328), ZN => n822);
   U1081 : AOI22_X1 port map( A1 => win(4), A2 => regs(2376), B1 => n39, B2 => 
                           regs(1864), ZN => n821);
   U1082 : NAND3_X1 port map( A1 => n823, A2 => n822, A3 => n821, ZN => 
                           curr_proc_regs(328));
   U1083 : NAND2_X1 port map( A1 => regs(841), A2 => n15, ZN => n826);
   U1084 : AOI22_X1 port map( A1 => n2, A2 => regs(1353), B1 => n25, B2 => 
                           regs(329), ZN => n825);
   U1085 : AOI22_X1 port map( A1 => win(4), A2 => regs(2377), B1 => n36, B2 => 
                           regs(1865), ZN => n824);
   U1086 : NAND3_X1 port map( A1 => n826, A2 => n825, A3 => n824, ZN => 
                           curr_proc_regs(329));
   U1087 : NAND2_X1 port map( A1 => regs(544), A2 => n10, ZN => n829);
   U1088 : AOI22_X1 port map( A1 => n2, A2 => regs(1056), B1 => n1596, B2 => 
                           regs(32), ZN => n828);
   U1089 : AOI22_X1 port map( A1 => n5, A2 => regs(2080), B1 => n38, B2 => 
                           regs(1568), ZN => n827);
   U1090 : NAND3_X1 port map( A1 => n829, A2 => n828, A3 => n827, ZN => 
                           curr_proc_regs(32));
   U1091 : NAND2_X1 port map( A1 => regs(842), A2 => n15, ZN => n832);
   U1092 : AOI22_X1 port map( A1 => n2, A2 => regs(1354), B1 => n21, B2 => 
                           regs(330), ZN => n831);
   U1093 : AOI22_X1 port map( A1 => n5, A2 => regs(2378), B1 => n39, B2 => 
                           regs(1866), ZN => n830);
   U1094 : NAND3_X1 port map( A1 => n832, A2 => n831, A3 => n830, ZN => 
                           curr_proc_regs(330));
   U1095 : NAND2_X1 port map( A1 => regs(843), A2 => n10, ZN => n835);
   U1096 : AOI22_X1 port map( A1 => n2, A2 => regs(1355), B1 => n20, B2 => 
                           regs(331), ZN => n834);
   U1097 : AOI22_X1 port map( A1 => n5, A2 => regs(2379), B1 => n38, B2 => 
                           regs(1867), ZN => n833);
   U1098 : NAND3_X1 port map( A1 => n835, A2 => n834, A3 => n833, ZN => 
                           curr_proc_regs(331));
   U1099 : NAND2_X1 port map( A1 => regs(844), A2 => n15, ZN => n838);
   U1100 : AOI22_X1 port map( A1 => n2, A2 => regs(1356), B1 => n25, B2 => 
                           regs(332), ZN => n837);
   U1101 : AOI22_X1 port map( A1 => n5, A2 => regs(2380), B1 => n36, B2 => 
                           regs(1868), ZN => n836);
   U1102 : NAND3_X1 port map( A1 => n838, A2 => n837, A3 => n836, ZN => 
                           curr_proc_regs(332));
   U1103 : NAND2_X1 port map( A1 => regs(845), A2 => n15, ZN => n841);
   U1104 : AOI22_X1 port map( A1 => n2, A2 => regs(1357), B1 => n25, B2 => 
                           regs(333), ZN => n840);
   U1105 : AOI22_X1 port map( A1 => n5, A2 => regs(2381), B1 => n36, B2 => 
                           regs(1869), ZN => n839);
   U1106 : NAND3_X1 port map( A1 => n841, A2 => n840, A3 => n839, ZN => 
                           curr_proc_regs(333));
   U1107 : NAND2_X1 port map( A1 => regs(846), A2 => n15, ZN => n844);
   U1108 : AOI22_X1 port map( A1 => n33, A2 => regs(1358), B1 => n1596, B2 => 
                           regs(334), ZN => n843);
   U1109 : AOI22_X1 port map( A1 => n5, A2 => regs(2382), B1 => n39, B2 => 
                           regs(1870), ZN => n842);
   U1110 : NAND3_X1 port map( A1 => n844, A2 => n843, A3 => n842, ZN => 
                           curr_proc_regs(334));
   U1111 : NAND2_X1 port map( A1 => regs(847), A2 => n15, ZN => n847);
   U1112 : AOI22_X1 port map( A1 => n31, A2 => regs(1359), B1 => n25, B2 => 
                           regs(335), ZN => n846);
   U1113 : AOI22_X1 port map( A1 => n5, A2 => regs(2383), B1 => n36, B2 => 
                           regs(1871), ZN => n845);
   U1114 : NAND3_X1 port map( A1 => n847, A2 => n846, A3 => n845, ZN => 
                           curr_proc_regs(335));
   U1115 : NAND2_X1 port map( A1 => regs(848), A2 => n15, ZN => n850);
   U1116 : AOI22_X1 port map( A1 => n29, A2 => regs(1360), B1 => n25, B2 => 
                           regs(336), ZN => n849);
   U1117 : AOI22_X1 port map( A1 => n5, A2 => regs(2384), B1 => n36, B2 => 
                           regs(1872), ZN => n848);
   U1118 : NAND3_X1 port map( A1 => n850, A2 => n849, A3 => n848, ZN => 
                           curr_proc_regs(336));
   U1119 : NAND2_X1 port map( A1 => regs(849), A2 => n15, ZN => n853);
   U1120 : AOI22_X1 port map( A1 => n29, A2 => regs(1361), B1 => n25, B2 => 
                           regs(337), ZN => n852);
   U1121 : AOI22_X1 port map( A1 => n5, A2 => regs(2385), B1 => n36, B2 => 
                           regs(1873), ZN => n851);
   U1122 : NAND3_X1 port map( A1 => n853, A2 => n852, A3 => n851, ZN => 
                           curr_proc_regs(337));
   U1123 : NAND2_X1 port map( A1 => regs(850), A2 => n10, ZN => n856);
   U1124 : AOI22_X1 port map( A1 => n31, A2 => regs(1362), B1 => n21, B2 => 
                           regs(338), ZN => n855);
   U1125 : AOI22_X1 port map( A1 => n5, A2 => regs(2386), B1 => n39, B2 => 
                           regs(1874), ZN => n854);
   U1126 : NAND3_X1 port map( A1 => n856, A2 => n855, A3 => n854, ZN => 
                           curr_proc_regs(338));
   U1127 : NAND2_X1 port map( A1 => regs(851), A2 => n15, ZN => n859);
   U1128 : AOI22_X1 port map( A1 => n31, A2 => regs(1363), B1 => n25, B2 => 
                           regs(339), ZN => n858);
   U1129 : AOI22_X1 port map( A1 => n47, A2 => regs(2387), B1 => n36, B2 => 
                           regs(1875), ZN => n857);
   U1130 : NAND3_X1 port map( A1 => n859, A2 => n858, A3 => n857, ZN => 
                           curr_proc_regs(339));
   U1131 : NAND2_X1 port map( A1 => regs(545), A2 => n15, ZN => n862);
   U1132 : AOI22_X1 port map( A1 => n29, A2 => regs(1057), B1 => n25, B2 => 
                           regs(33), ZN => n861);
   U1133 : AOI22_X1 port map( A1 => n47, A2 => regs(2081), B1 => n36, B2 => 
                           regs(1569), ZN => n860);
   U1134 : NAND3_X1 port map( A1 => n862, A2 => n861, A3 => n860, ZN => 
                           curr_proc_regs(33));
   U1135 : NAND2_X1 port map( A1 => regs(852), A2 => n15, ZN => n865);
   U1136 : AOI22_X1 port map( A1 => n31, A2 => regs(1364), B1 => n25, B2 => 
                           regs(340), ZN => n864);
   U1137 : AOI22_X1 port map( A1 => n47, A2 => regs(2388), B1 => n36, B2 => 
                           regs(1876), ZN => n863);
   U1138 : NAND3_X1 port map( A1 => n865, A2 => n864, A3 => n863, ZN => 
                           curr_proc_regs(340));
   U1139 : NAND2_X1 port map( A1 => regs(853), A2 => n15, ZN => n868);
   U1140 : AOI22_X1 port map( A1 => n31, A2 => regs(1365), B1 => n18, B2 => 
                           regs(341), ZN => n867);
   U1141 : AOI22_X1 port map( A1 => n47, A2 => regs(2389), B1 => n38, B2 => 
                           regs(1877), ZN => n866);
   U1142 : NAND3_X1 port map( A1 => n868, A2 => n867, A3 => n866, ZN => 
                           curr_proc_regs(341));
   U1143 : NAND2_X1 port map( A1 => regs(854), A2 => n10, ZN => n871);
   U1144 : AOI22_X1 port map( A1 => n30, A2 => regs(1366), B1 => n23, B2 => 
                           regs(342), ZN => n870);
   U1145 : AOI22_X1 port map( A1 => n47, A2 => regs(2390), B1 => n39, B2 => 
                           regs(1878), ZN => n869);
   U1146 : NAND3_X1 port map( A1 => n871, A2 => n870, A3 => n869, ZN => 
                           curr_proc_regs(342));
   U1147 : NAND2_X1 port map( A1 => regs(855), A2 => n15, ZN => n874);
   U1148 : AOI22_X1 port map( A1 => n33, A2 => regs(1367), B1 => n25, B2 => 
                           regs(343), ZN => n873);
   U1149 : AOI22_X1 port map( A1 => n47, A2 => regs(2391), B1 => n36, B2 => 
                           regs(1879), ZN => n872);
   U1150 : NAND3_X1 port map( A1 => n874, A2 => n873, A3 => n872, ZN => 
                           curr_proc_regs(343));
   U1151 : NAND2_X1 port map( A1 => regs(856), A2 => n15, ZN => n877);
   U1152 : AOI22_X1 port map( A1 => n31, A2 => regs(1368), B1 => n25, B2 => 
                           regs(344), ZN => n876);
   U1153 : AOI22_X1 port map( A1 => n47, A2 => regs(2392), B1 => n36, B2 => 
                           regs(1880), ZN => n875);
   U1154 : NAND3_X1 port map( A1 => n877, A2 => n876, A3 => n875, ZN => 
                           curr_proc_regs(344));
   U1155 : NAND2_X1 port map( A1 => regs(857), A2 => n15, ZN => n880);
   U1156 : AOI22_X1 port map( A1 => n33, A2 => regs(1369), B1 => n25, B2 => 
                           regs(345), ZN => n879);
   U1157 : AOI22_X1 port map( A1 => n47, A2 => regs(2393), B1 => n36, B2 => 
                           regs(1881), ZN => n878);
   U1158 : NAND3_X1 port map( A1 => n880, A2 => n879, A3 => n878, ZN => 
                           curr_proc_regs(345));
   U1159 : NAND2_X1 port map( A1 => regs(858), A2 => n15, ZN => n883);
   U1160 : AOI22_X1 port map( A1 => n30, A2 => regs(1370), B1 => n25, B2 => 
                           regs(346), ZN => n882);
   U1161 : AOI22_X1 port map( A1 => n47, A2 => regs(2394), B1 => n36, B2 => 
                           regs(1882), ZN => n881);
   U1162 : NAND3_X1 port map( A1 => n883, A2 => n882, A3 => n881, ZN => 
                           curr_proc_regs(346));
   U1163 : NAND2_X1 port map( A1 => regs(859), A2 => n15, ZN => n886);
   U1164 : AOI22_X1 port map( A1 => n29, A2 => regs(1371), B1 => n25, B2 => 
                           regs(347), ZN => n885);
   U1165 : AOI22_X1 port map( A1 => n47, A2 => regs(2395), B1 => n36, B2 => 
                           regs(1883), ZN => n884);
   U1166 : NAND3_X1 port map( A1 => n886, A2 => n885, A3 => n884, ZN => 
                           curr_proc_regs(347));
   U1167 : NAND2_X1 port map( A1 => regs(860), A2 => n15, ZN => n889);
   U1168 : AOI22_X1 port map( A1 => n31, A2 => regs(1372), B1 => n25, B2 => 
                           regs(348), ZN => n888);
   U1169 : AOI22_X1 port map( A1 => n47, A2 => regs(2396), B1 => n36, B2 => 
                           regs(1884), ZN => n887);
   U1170 : NAND3_X1 port map( A1 => n889, A2 => n888, A3 => n887, ZN => 
                           curr_proc_regs(348));
   U1171 : NAND2_X1 port map( A1 => regs(861), A2 => n1, ZN => n892);
   U1172 : AOI22_X1 port map( A1 => n31, A2 => regs(1373), B1 => n24, B2 => 
                           regs(349), ZN => n891);
   U1173 : AOI22_X1 port map( A1 => n47, A2 => regs(2397), B1 => n41, B2 => 
                           regs(1885), ZN => n890);
   U1174 : NAND3_X1 port map( A1 => n892, A2 => n891, A3 => n890, ZN => 
                           curr_proc_regs(349));
   U1175 : NAND2_X1 port map( A1 => regs(546), A2 => n1, ZN => n895);
   U1176 : AOI22_X1 port map( A1 => n31, A2 => regs(1058), B1 => n24, B2 => 
                           regs(34), ZN => n894);
   U1177 : AOI22_X1 port map( A1 => n46, A2 => regs(2082), B1 => n41, B2 => 
                           regs(1570), ZN => n893);
   U1178 : NAND3_X1 port map( A1 => n895, A2 => n894, A3 => n893, ZN => 
                           curr_proc_regs(34));
   U1179 : NAND2_X1 port map( A1 => regs(862), A2 => n1, ZN => n898);
   U1180 : AOI22_X1 port map( A1 => n29, A2 => regs(1374), B1 => n20, B2 => 
                           regs(350), ZN => n897);
   U1181 : AOI22_X1 port map( A1 => n46, A2 => regs(2398), B1 => n39, B2 => 
                           regs(1886), ZN => n896);
   U1182 : NAND3_X1 port map( A1 => n898, A2 => n897, A3 => n896, ZN => 
                           curr_proc_regs(350));
   U1183 : NAND2_X1 port map( A1 => regs(863), A2 => n1, ZN => n901);
   U1184 : AOI22_X1 port map( A1 => n33, A2 => regs(1375), B1 => n26, B2 => 
                           regs(351), ZN => n900);
   U1185 : AOI22_X1 port map( A1 => n46, A2 => regs(2399), B1 => n38, B2 => 
                           regs(1887), ZN => n899);
   U1186 : NAND3_X1 port map( A1 => n901, A2 => n900, A3 => n899, ZN => 
                           curr_proc_regs(351));
   U1187 : NAND2_X1 port map( A1 => regs(864), A2 => n1, ZN => n904);
   U1188 : AOI22_X1 port map( A1 => n30, A2 => regs(1376), B1 => n24, B2 => 
                           regs(352), ZN => n903);
   U1189 : AOI22_X1 port map( A1 => n46, A2 => regs(2400), B1 => n41, B2 => 
                           regs(1888), ZN => n902);
   U1190 : NAND3_X1 port map( A1 => n904, A2 => n903, A3 => n902, ZN => 
                           curr_proc_regs(352));
   U1191 : NAND2_X1 port map( A1 => regs(865), A2 => n1, ZN => n907);
   U1192 : AOI22_X1 port map( A1 => n33, A2 => regs(1377), B1 => n18, B2 => 
                           regs(353), ZN => n906);
   U1193 : AOI22_X1 port map( A1 => n46, A2 => regs(2401), B1 => n39, B2 => 
                           regs(1889), ZN => n905);
   U1194 : NAND3_X1 port map( A1 => n907, A2 => n906, A3 => n905, ZN => 
                           curr_proc_regs(353));
   U1195 : NAND2_X1 port map( A1 => regs(866), A2 => n1, ZN => n910);
   U1196 : AOI22_X1 port map( A1 => n31, A2 => regs(1378), B1 => n24, B2 => 
                           regs(354), ZN => n909);
   U1197 : AOI22_X1 port map( A1 => n46, A2 => regs(2402), B1 => n41, B2 => 
                           regs(1890), ZN => n908);
   U1198 : NAND3_X1 port map( A1 => n910, A2 => n909, A3 => n908, ZN => 
                           curr_proc_regs(354));
   U1199 : NAND2_X1 port map( A1 => regs(867), A2 => n1, ZN => n913);
   U1200 : AOI22_X1 port map( A1 => n33, A2 => regs(1379), B1 => n24, B2 => 
                           regs(355), ZN => n912);
   U1201 : AOI22_X1 port map( A1 => n46, A2 => regs(2403), B1 => n41, B2 => 
                           regs(1891), ZN => n911);
   U1202 : NAND3_X1 port map( A1 => n913, A2 => n912, A3 => n911, ZN => 
                           curr_proc_regs(355));
   U1203 : NAND2_X1 port map( A1 => regs(868), A2 => n1, ZN => n916);
   U1204 : AOI22_X1 port map( A1 => n31, A2 => regs(1380), B1 => n23, B2 => 
                           regs(356), ZN => n915);
   U1205 : AOI22_X1 port map( A1 => n46, A2 => regs(2404), B1 => n38, B2 => 
                           regs(1892), ZN => n914);
   U1206 : NAND3_X1 port map( A1 => n916, A2 => n915, A3 => n914, ZN => 
                           curr_proc_regs(356));
   U1207 : NAND2_X1 port map( A1 => regs(869), A2 => n1, ZN => n919);
   U1208 : AOI22_X1 port map( A1 => n33, A2 => regs(1381), B1 => n24, B2 => 
                           regs(357), ZN => n918);
   U1209 : AOI22_X1 port map( A1 => n46, A2 => regs(2405), B1 => n41, B2 => 
                           regs(1893), ZN => n917);
   U1210 : NAND3_X1 port map( A1 => n919, A2 => n918, A3 => n917, ZN => 
                           curr_proc_regs(357));
   U1211 : NAND2_X1 port map( A1 => regs(870), A2 => n1, ZN => n922);
   U1212 : AOI22_X1 port map( A1 => n31, A2 => regs(1382), B1 => n24, B2 => 
                           regs(358), ZN => n921);
   U1213 : AOI22_X1 port map( A1 => n46, A2 => regs(2406), B1 => n41, B2 => 
                           regs(1894), ZN => n920);
   U1214 : NAND3_X1 port map( A1 => n922, A2 => n921, A3 => n920, ZN => 
                           curr_proc_regs(358));
   U1215 : NAND2_X1 port map( A1 => regs(871), A2 => n1, ZN => n925);
   U1216 : AOI22_X1 port map( A1 => n30, A2 => regs(1383), B1 => n26, B2 => 
                           regs(359), ZN => n924);
   U1217 : AOI22_X1 port map( A1 => n46, A2 => regs(2407), B1 => n39, B2 => 
                           regs(1895), ZN => n923);
   U1218 : NAND3_X1 port map( A1 => n925, A2 => n924, A3 => n923, ZN => 
                           curr_proc_regs(359));
   U1219 : NAND2_X1 port map( A1 => regs(547), A2 => n11, ZN => n928);
   U1220 : AOI22_X1 port map( A1 => n31, A2 => regs(1059), B1 => n24, B2 => 
                           regs(35), ZN => n927);
   U1221 : AOI22_X1 port map( A1 => n46, A2 => regs(2083), B1 => n41, B2 => 
                           regs(1571), ZN => n926);
   U1222 : NAND3_X1 port map( A1 => n928, A2 => n927, A3 => n926, ZN => 
                           curr_proc_regs(35));
   U1223 : NAND2_X1 port map( A1 => regs(872), A2 => n4, ZN => n931);
   U1224 : AOI22_X1 port map( A1 => n31, A2 => regs(1384), B1 => n17, B2 => 
                           regs(360), ZN => n930);
   U1225 : AOI22_X1 port map( A1 => n8, A2 => regs(2408), B1 => n38, B2 => 
                           regs(1896), ZN => n929);
   U1226 : NAND3_X1 port map( A1 => n931, A2 => n930, A3 => n929, ZN => 
                           curr_proc_regs(360));
   U1227 : NAND2_X1 port map( A1 => regs(873), A2 => n1, ZN => n934);
   U1228 : AOI22_X1 port map( A1 => n33, A2 => regs(1385), B1 => n20, B2 => 
                           regs(361), ZN => n933);
   U1229 : AOI22_X1 port map( A1 => n8, A2 => regs(2409), B1 => n39, B2 => 
                           regs(1897), ZN => n932);
   U1230 : NAND3_X1 port map( A1 => n934, A2 => n933, A3 => n932, ZN => 
                           curr_proc_regs(361));
   U1231 : NAND2_X1 port map( A1 => regs(874), A2 => n11, ZN => n937);
   U1232 : AOI22_X1 port map( A1 => n31, A2 => regs(1386), B1 => n21, B2 => 
                           regs(362), ZN => n936);
   U1233 : AOI22_X1 port map( A1 => n8, A2 => regs(2410), B1 => n38, B2 => 
                           regs(1898), ZN => n935);
   U1234 : NAND3_X1 port map( A1 => n937, A2 => n936, A3 => n935, ZN => 
                           curr_proc_regs(362));
   U1235 : NAND2_X1 port map( A1 => regs(875), A2 => n4, ZN => n940);
   U1236 : AOI22_X1 port map( A1 => n30, A2 => regs(1387), B1 => n24, B2 => 
                           regs(363), ZN => n939);
   U1237 : AOI22_X1 port map( A1 => n8, A2 => regs(2411), B1 => n41, B2 => 
                           regs(1899), ZN => n938);
   U1238 : NAND3_X1 port map( A1 => n940, A2 => n939, A3 => n938, ZN => 
                           curr_proc_regs(363));
   U1239 : NAND2_X1 port map( A1 => regs(876), A2 => n1, ZN => n943);
   U1240 : AOI22_X1 port map( A1 => n29, A2 => regs(1388), B1 => n24, B2 => 
                           regs(364), ZN => n942);
   U1241 : AOI22_X1 port map( A1 => n8, A2 => regs(2412), B1 => n41, B2 => 
                           regs(1900), ZN => n941);
   U1242 : NAND3_X1 port map( A1 => n943, A2 => n942, A3 => n941, ZN => 
                           curr_proc_regs(364));
   U1243 : NAND2_X1 port map( A1 => regs(877), A2 => n11, ZN => n946);
   U1244 : AOI22_X1 port map( A1 => n31, A2 => regs(1389), B1 => n19, B2 => 
                           regs(365), ZN => n945);
   U1245 : AOI22_X1 port map( A1 => n8, A2 => regs(2413), B1 => n39, B2 => 
                           regs(1901), ZN => n944);
   U1246 : NAND3_X1 port map( A1 => n946, A2 => n945, A3 => n944, ZN => 
                           curr_proc_regs(365));
   U1247 : NAND2_X1 port map( A1 => regs(878), A2 => n4, ZN => n949);
   U1248 : AOI22_X1 port map( A1 => n33, A2 => regs(1390), B1 => n19, B2 => 
                           regs(366), ZN => n948);
   U1249 : AOI22_X1 port map( A1 => n8, A2 => regs(2414), B1 => n38, B2 => 
                           regs(1902), ZN => n947);
   U1250 : NAND3_X1 port map( A1 => n949, A2 => n948, A3 => n947, ZN => 
                           curr_proc_regs(366));
   U1251 : NAND2_X1 port map( A1 => regs(879), A2 => n1, ZN => n952);
   U1252 : AOI22_X1 port map( A1 => n2, A2 => regs(1391), B1 => n24, B2 => 
                           regs(367), ZN => n951);
   U1253 : AOI22_X1 port map( A1 => n8, A2 => regs(2415), B1 => n41, B2 => 
                           regs(1903), ZN => n950);
   U1254 : NAND3_X1 port map( A1 => n952, A2 => n951, A3 => n950, ZN => 
                           curr_proc_regs(367));
   U1255 : NAND2_X1 port map( A1 => regs(880), A2 => n11, ZN => n955);
   U1256 : AOI22_X1 port map( A1 => n2, A2 => regs(1392), B1 => n24, B2 => 
                           regs(368), ZN => n954);
   U1257 : AOI22_X1 port map( A1 => n8, A2 => regs(2416), B1 => n41, B2 => 
                           regs(1904), ZN => n953);
   U1258 : NAND3_X1 port map( A1 => n955, A2 => n954, A3 => n953, ZN => 
                           curr_proc_regs(368));
   U1259 : NAND2_X1 port map( A1 => regs(881), A2 => n4, ZN => n958);
   U1260 : AOI22_X1 port map( A1 => n2, A2 => regs(1393), B1 => n24, B2 => 
                           regs(369), ZN => n957);
   U1261 : AOI22_X1 port map( A1 => n8, A2 => regs(2417), B1 => n41, B2 => 
                           regs(1905), ZN => n956);
   U1262 : NAND3_X1 port map( A1 => n958, A2 => n957, A3 => n956, ZN => 
                           curr_proc_regs(369));
   U1263 : NAND2_X1 port map( A1 => regs(548), A2 => n1, ZN => n961);
   U1264 : AOI22_X1 port map( A1 => n2, A2 => regs(1060), B1 => n24, B2 => 
                           regs(36), ZN => n960);
   U1265 : AOI22_X1 port map( A1 => n8, A2 => regs(2084), B1 => n41, B2 => 
                           regs(1572), ZN => n959);
   U1266 : NAND3_X1 port map( A1 => n961, A2 => n960, A3 => n959, ZN => 
                           curr_proc_regs(36));
   U1267 : NAND2_X1 port map( A1 => regs(882), A2 => n11, ZN => n964);
   U1268 : AOI22_X1 port map( A1 => n2, A2 => regs(1394), B1 => n20, B2 => 
                           regs(370), ZN => n963);
   U1269 : AOI22_X1 port map( A1 => n8, A2 => regs(2418), B1 => n38, B2 => 
                           regs(1906), ZN => n962);
   U1270 : NAND3_X1 port map( A1 => n964, A2 => n963, A3 => n962, ZN => 
                           curr_proc_regs(370));
   U1271 : NAND2_X1 port map( A1 => regs(883), A2 => n11, ZN => n967);
   U1272 : AOI22_X1 port map( A1 => n2, A2 => regs(1395), B1 => n17, B2 => 
                           regs(371), ZN => n966);
   U1273 : AOI22_X1 port map( A1 => n45, A2 => regs(2419), B1 => n39, B2 => 
                           regs(1907), ZN => n965);
   U1274 : NAND3_X1 port map( A1 => n967, A2 => n966, A3 => n965, ZN => 
                           curr_proc_regs(371));
   U1275 : NAND2_X1 port map( A1 => regs(884), A2 => n11, ZN => n970);
   U1276 : AOI22_X1 port map( A1 => n2, A2 => regs(1396), B1 => n21, B2 => 
                           regs(372), ZN => n969);
   U1277 : AOI22_X1 port map( A1 => n45, A2 => regs(2420), B1 => n38, B2 => 
                           regs(1908), ZN => n968);
   U1278 : NAND3_X1 port map( A1 => n970, A2 => n969, A3 => n968, ZN => 
                           curr_proc_regs(372));
   U1279 : NAND2_X1 port map( A1 => regs(885), A2 => n11, ZN => n973);
   U1280 : AOI22_X1 port map( A1 => n2, A2 => regs(1397), B1 => n21, B2 => 
                           regs(373), ZN => n972);
   U1281 : AOI22_X1 port map( A1 => n45, A2 => regs(2421), B1 => n39, B2 => 
                           regs(1909), ZN => n971);
   U1282 : NAND3_X1 port map( A1 => n973, A2 => n972, A3 => n971, ZN => 
                           curr_proc_regs(373));
   U1283 : NAND2_X1 port map( A1 => regs(886), A2 => n11, ZN => n976);
   U1284 : AOI22_X1 port map( A1 => n2, A2 => regs(1398), B1 => n19, B2 => 
                           regs(374), ZN => n975);
   U1285 : AOI22_X1 port map( A1 => n45, A2 => regs(2422), B1 => n38, B2 => 
                           regs(1910), ZN => n974);
   U1286 : NAND3_X1 port map( A1 => n976, A2 => n975, A3 => n974, ZN => 
                           curr_proc_regs(374));
   U1287 : NAND2_X1 port map( A1 => regs(887), A2 => n11, ZN => n979);
   U1288 : AOI22_X1 port map( A1 => n2, A2 => regs(1399), B1 => n19, B2 => 
                           regs(375), ZN => n978);
   U1289 : AOI22_X1 port map( A1 => n45, A2 => regs(2423), B1 => n39, B2 => 
                           regs(1911), ZN => n977);
   U1290 : NAND3_X1 port map( A1 => n979, A2 => n978, A3 => n977, ZN => 
                           curr_proc_regs(375));
   U1291 : NAND2_X1 port map( A1 => regs(888), A2 => n11, ZN => n982);
   U1292 : AOI22_X1 port map( A1 => n2, A2 => regs(1400), B1 => n1596, B2 => 
                           regs(376), ZN => n981);
   U1293 : AOI22_X1 port map( A1 => n45, A2 => regs(2424), B1 => n38, B2 => 
                           regs(1912), ZN => n980);
   U1294 : NAND3_X1 port map( A1 => n982, A2 => n981, A3 => n980, ZN => 
                           curr_proc_regs(376));
   U1295 : NAND2_X1 port map( A1 => regs(889), A2 => n11, ZN => n985);
   U1296 : AOI22_X1 port map( A1 => n2, A2 => regs(1401), B1 => n19, B2 => 
                           regs(377), ZN => n984);
   U1297 : AOI22_X1 port map( A1 => n45, A2 => regs(2425), B1 => n39, B2 => 
                           regs(1913), ZN => n983);
   U1298 : NAND3_X1 port map( A1 => n985, A2 => n984, A3 => n983, ZN => 
                           curr_proc_regs(377));
   U1299 : NAND2_X1 port map( A1 => regs(890), A2 => n11, ZN => n988);
   U1300 : AOI22_X1 port map( A1 => n30, A2 => regs(1402), B1 => n19, B2 => 
                           regs(378), ZN => n987);
   U1301 : AOI22_X1 port map( A1 => n45, A2 => regs(2426), B1 => n38, B2 => 
                           regs(1914), ZN => n986);
   U1302 : NAND3_X1 port map( A1 => n988, A2 => n987, A3 => n986, ZN => 
                           curr_proc_regs(378));
   U1303 : NAND2_X1 port map( A1 => regs(891), A2 => n11, ZN => n991);
   U1304 : AOI22_X1 port map( A1 => n30, A2 => regs(1403), B1 => n26, B2 => 
                           regs(379), ZN => n990);
   U1305 : AOI22_X1 port map( A1 => n45, A2 => regs(2427), B1 => n39, B2 => 
                           regs(1915), ZN => n989);
   U1306 : NAND3_X1 port map( A1 => n991, A2 => n990, A3 => n989, ZN => 
                           curr_proc_regs(379));
   U1307 : NAND2_X1 port map( A1 => regs(549), A2 => n11, ZN => n994);
   U1308 : AOI22_X1 port map( A1 => n30, A2 => regs(1061), B1 => n21, B2 => 
                           regs(37), ZN => n993);
   U1309 : AOI22_X1 port map( A1 => n45, A2 => regs(2085), B1 => n38, B2 => 
                           regs(1573), ZN => n992);
   U1310 : NAND3_X1 port map( A1 => n994, A2 => n993, A3 => n992, ZN => 
                           curr_proc_regs(37));
   U1311 : NAND2_X1 port map( A1 => regs(892), A2 => n11, ZN => n997);
   U1312 : AOI22_X1 port map( A1 => n30, A2 => regs(1404), B1 => n24, B2 => 
                           regs(380), ZN => n996);
   U1313 : AOI22_X1 port map( A1 => n45, A2 => regs(2428), B1 => n41, B2 => 
                           regs(1916), ZN => n995);
   U1314 : NAND3_X1 port map( A1 => n997, A2 => n996, A3 => n995, ZN => 
                           curr_proc_regs(380));
   U1315 : NAND2_X1 port map( A1 => regs(893), A2 => n1, ZN => n1000);
   U1316 : AOI22_X1 port map( A1 => n30, A2 => regs(1405), B1 => n24, B2 => 
                           regs(381), ZN => n999);
   U1317 : AOI22_X1 port map( A1 => n45, A2 => regs(2429), B1 => n41, B2 => 
                           regs(1917), ZN => n998);
   U1318 : NAND3_X1 port map( A1 => n1000, A2 => n999, A3 => n998, ZN => 
                           curr_proc_regs(381));
   U1319 : NAND2_X1 port map( A1 => regs(894), A2 => n11, ZN => n1003);
   U1320 : AOI22_X1 port map( A1 => n30, A2 => regs(1406), B1 => n24, B2 => 
                           regs(382), ZN => n1002);
   U1321 : AOI22_X1 port map( A1 => n44, A2 => regs(2430), B1 => n41, B2 => 
                           regs(1918), ZN => n1001);
   U1322 : NAND3_X1 port map( A1 => n1003, A2 => n1002, A3 => n1001, ZN => 
                           curr_proc_regs(382));
   U1323 : NAND2_X1 port map( A1 => regs(895), A2 => n4, ZN => n1006);
   U1324 : AOI22_X1 port map( A1 => n30, A2 => regs(1407), B1 => n26, B2 => 
                           regs(383), ZN => n1005);
   U1325 : AOI22_X1 port map( A1 => n44, A2 => regs(2431), B1 => n39, B2 => 
                           regs(1919), ZN => n1004);
   U1326 : NAND3_X1 port map( A1 => n1006, A2 => n1005, A3 => n1004, ZN => 
                           curr_proc_regs(383));
   U1327 : NAND2_X1 port map( A1 => regs(896), A2 => n11, ZN => n1009);
   U1328 : AOI22_X1 port map( A1 => n30, A2 => regs(1408), B1 => n24, B2 => 
                           regs(384), ZN => n1008);
   U1329 : AOI22_X1 port map( A1 => n44, A2 => regs(2432), B1 => n41, B2 => 
                           regs(1920), ZN => n1007);
   U1330 : NAND3_X1 port map( A1 => n1009, A2 => n1008, A3 => n1007, ZN => 
                           curr_proc_regs(384));
   U1331 : NAND2_X1 port map( A1 => regs(897), A2 => n1, ZN => n1012);
   U1332 : AOI22_X1 port map( A1 => n30, A2 => regs(1409), B1 => n24, B2 => 
                           regs(385), ZN => n1011);
   U1333 : AOI22_X1 port map( A1 => n44, A2 => regs(2433), B1 => n41, B2 => 
                           regs(1921), ZN => n1010);
   U1334 : NAND3_X1 port map( A1 => n1012, A2 => n1011, A3 => n1010, ZN => 
                           curr_proc_regs(385));
   U1335 : NAND2_X1 port map( A1 => regs(898), A2 => n11, ZN => n1015);
   U1336 : AOI22_X1 port map( A1 => n30, A2 => regs(1410), B1 => n26, B2 => 
                           regs(386), ZN => n1014);
   U1337 : AOI22_X1 port map( A1 => n44, A2 => regs(2434), B1 => n38, B2 => 
                           regs(1922), ZN => n1013);
   U1338 : NAND3_X1 port map( A1 => n1015, A2 => n1014, A3 => n1013, ZN => 
                           curr_proc_regs(386));
   U1339 : NAND2_X1 port map( A1 => regs(899), A2 => n4, ZN => n1018);
   U1340 : AOI22_X1 port map( A1 => n30, A2 => regs(1411), B1 => n21, B2 => 
                           regs(387), ZN => n1017);
   U1341 : AOI22_X1 port map( A1 => n44, A2 => regs(2435), B1 => n39, B2 => 
                           regs(1923), ZN => n1016);
   U1342 : NAND3_X1 port map( A1 => n1018, A2 => n1017, A3 => n1016, ZN => 
                           curr_proc_regs(387));
   U1343 : NAND2_X1 port map( A1 => regs(900), A2 => n4, ZN => n1021);
   U1344 : AOI22_X1 port map( A1 => n30, A2 => regs(1412), B1 => n21, B2 => 
                           regs(388), ZN => n1020);
   U1345 : AOI22_X1 port map( A1 => n44, A2 => regs(2436), B1 => n38, B2 => 
                           regs(1924), ZN => n1019);
   U1346 : NAND3_X1 port map( A1 => n1021, A2 => n1020, A3 => n1019, ZN => 
                           curr_proc_regs(388));
   U1347 : NAND2_X1 port map( A1 => regs(901), A2 => n1, ZN => n1024);
   U1348 : AOI22_X1 port map( A1 => n31, A2 => regs(1413), B1 => n24, B2 => 
                           regs(389), ZN => n1023);
   U1349 : AOI22_X1 port map( A1 => n44, A2 => regs(2437), B1 => n41, B2 => 
                           regs(1925), ZN => n1022);
   U1350 : NAND3_X1 port map( A1 => n1024, A2 => n1023, A3 => n1022, ZN => 
                           curr_proc_regs(389));
   U1351 : NAND2_X1 port map( A1 => regs(550), A2 => n4, ZN => n1027);
   U1352 : AOI22_X1 port map( A1 => n31, A2 => regs(1062), B1 => n24, B2 => 
                           regs(38), ZN => n1026);
   U1353 : AOI22_X1 port map( A1 => n44, A2 => regs(2086), B1 => n41, B2 => 
                           regs(1574), ZN => n1025);
   U1354 : NAND3_X1 port map( A1 => n1027, A2 => n1026, A3 => n1025, ZN => 
                           curr_proc_regs(38));
   U1355 : NAND2_X1 port map( A1 => regs(902), A2 => n4, ZN => n1030);
   U1356 : AOI22_X1 port map( A1 => n31, A2 => regs(1414), B1 => n1596, B2 => 
                           regs(390), ZN => n1029);
   U1357 : AOI22_X1 port map( A1 => n44, A2 => regs(2438), B1 => n39, B2 => 
                           regs(1926), ZN => n1028);
   U1358 : NAND3_X1 port map( A1 => n1030, A2 => n1029, A3 => n1028, ZN => 
                           curr_proc_regs(390));
   U1359 : NAND2_X1 port map( A1 => regs(903), A2 => n4, ZN => n1033);
   U1360 : AOI22_X1 port map( A1 => n31, A2 => regs(1415), B1 => n24, B2 => 
                           regs(391), ZN => n1032);
   U1361 : AOI22_X1 port map( A1 => n44, A2 => regs(2439), B1 => n41, B2 => 
                           regs(1927), ZN => n1031);
   U1362 : NAND3_X1 port map( A1 => n1033, A2 => n1032, A3 => n1031, ZN => 
                           curr_proc_regs(391));
   U1363 : NAND2_X1 port map( A1 => regs(904), A2 => n11, ZN => n1036);
   U1364 : AOI22_X1 port map( A1 => n31, A2 => regs(1416), B1 => n24, B2 => 
                           regs(392), ZN => n1035);
   U1365 : AOI22_X1 port map( A1 => n8, A2 => regs(2440), B1 => n41, B2 => 
                           regs(1928), ZN => n1034);
   U1366 : NAND3_X1 port map( A1 => n1036, A2 => n1035, A3 => n1034, ZN => 
                           curr_proc_regs(392));
   U1367 : NAND2_X1 port map( A1 => regs(905), A2 => n4, ZN => n1039);
   U1368 : AOI22_X1 port map( A1 => n31, A2 => regs(1417), B1 => n21, B2 => 
                           regs(393), ZN => n1038);
   U1369 : AOI22_X1 port map( A1 => n8, A2 => regs(2441), B1 => n39, B2 => 
                           regs(1929), ZN => n1037);
   U1370 : NAND3_X1 port map( A1 => n1039, A2 => n1038, A3 => n1037, ZN => 
                           curr_proc_regs(393));
   U1371 : NAND2_X1 port map( A1 => regs(906), A2 => n4, ZN => n1042);
   U1372 : AOI22_X1 port map( A1 => n31, A2 => regs(1418), B1 => n24, B2 => 
                           regs(394), ZN => n1041);
   U1373 : AOI22_X1 port map( A1 => n8, A2 => regs(2442), B1 => n41, B2 => 
                           regs(1930), ZN => n1040);
   U1374 : NAND3_X1 port map( A1 => n1042, A2 => n1041, A3 => n1040, ZN => 
                           curr_proc_regs(394));
   U1375 : NAND2_X1 port map( A1 => regs(907), A2 => n4, ZN => n1045);
   U1376 : AOI22_X1 port map( A1 => n31, A2 => regs(1419), B1 => n23, B2 => 
                           regs(395), ZN => n1044);
   U1377 : AOI22_X1 port map( A1 => n8, A2 => regs(2443), B1 => n38, B2 => 
                           regs(1931), ZN => n1043);
   U1378 : NAND3_X1 port map( A1 => n1045, A2 => n1044, A3 => n1043, ZN => 
                           curr_proc_regs(395));
   U1379 : NAND2_X1 port map( A1 => regs(908), A2 => n1, ZN => n1048);
   U1380 : AOI22_X1 port map( A1 => n31, A2 => regs(1420), B1 => n17, B2 => 
                           regs(396), ZN => n1047);
   U1381 : AOI22_X1 port map( A1 => n8, A2 => regs(2444), B1 => n39, B2 => 
                           regs(1932), ZN => n1046);
   U1382 : NAND3_X1 port map( A1 => n1048, A2 => n1047, A3 => n1046, ZN => 
                           curr_proc_regs(396));
   U1383 : NAND2_X1 port map( A1 => regs(909), A2 => n11, ZN => n1051);
   U1384 : AOI22_X1 port map( A1 => n31, A2 => regs(1421), B1 => n24, B2 => 
                           regs(397), ZN => n1050);
   U1385 : AOI22_X1 port map( A1 => n8, A2 => regs(2445), B1 => n41, B2 => 
                           regs(1933), ZN => n1049);
   U1386 : NAND3_X1 port map( A1 => n1051, A2 => n1050, A3 => n1049, ZN => 
                           curr_proc_regs(397));
   U1387 : NAND2_X1 port map( A1 => regs(910), A2 => n4, ZN => n1054);
   U1388 : AOI22_X1 port map( A1 => n31, A2 => regs(1422), B1 => n20, B2 => 
                           regs(398), ZN => n1053);
   U1389 : AOI22_X1 port map( A1 => n8, A2 => regs(2446), B1 => n38, B2 => 
                           regs(1934), ZN => n1052);
   U1390 : NAND3_X1 port map( A1 => n1054, A2 => n1053, A3 => n1052, ZN => 
                           curr_proc_regs(398));
   U1391 : NAND2_X1 port map( A1 => regs(911), A2 => n4, ZN => n1057);
   U1392 : AOI22_X1 port map( A1 => n31, A2 => regs(1423), B1 => n24, B2 => 
                           regs(399), ZN => n1056);
   U1393 : AOI22_X1 port map( A1 => n8, A2 => regs(2447), B1 => n41, B2 => 
                           regs(1935), ZN => n1055);
   U1394 : NAND3_X1 port map( A1 => n1057, A2 => n1056, A3 => n1055, ZN => 
                           curr_proc_regs(399));
   U1395 : NAND2_X1 port map( A1 => regs(551), A2 => n4, ZN => n1060);
   U1396 : AOI22_X1 port map( A1 => n29, A2 => regs(1063), B1 => n26, B2 => 
                           regs(39), ZN => n1059);
   U1397 : AOI22_X1 port map( A1 => n8, A2 => regs(2087), B1 => n39, B2 => 
                           regs(1575), ZN => n1058);
   U1398 : NAND3_X1 port map( A1 => n1060, A2 => n1059, A3 => n1058, ZN => 
                           curr_proc_regs(39));
   U1399 : NAND2_X1 port map( A1 => regs(515), A2 => n4, ZN => n1063);
   U1400 : AOI22_X1 port map( A1 => n29, A2 => regs(1027), B1 => n18, B2 => 
                           regs(3), ZN => n1062);
   U1401 : AOI22_X1 port map( A1 => n8, A2 => regs(2051), B1 => n38, B2 => 
                           regs(1539), ZN => n1061);
   U1402 : NAND3_X1 port map( A1 => n1063, A2 => n1062, A3 => n1061, ZN => 
                           curr_proc_regs(3));
   U1403 : NAND2_X1 port map( A1 => regs(912), A2 => n4, ZN => n1066);
   U1404 : AOI22_X1 port map( A1 => n29, A2 => regs(1424), B1 => n23, B2 => 
                           regs(400), ZN => n1065);
   U1405 : AOI22_X1 port map( A1 => n8, A2 => regs(2448), B1 => n39, B2 => 
                           regs(1936), ZN => n1064);
   U1406 : NAND3_X1 port map( A1 => n1066, A2 => n1065, A3 => n1064, ZN => 
                           curr_proc_regs(400));
   U1407 : NAND2_X1 port map( A1 => regs(913), A2 => n4, ZN => n1069);
   U1408 : AOI22_X1 port map( A1 => n29, A2 => regs(1425), B1 => n26, B2 => 
                           regs(401), ZN => n1068);
   U1409 : AOI22_X1 port map( A1 => n8, A2 => regs(2449), B1 => n38, B2 => 
                           regs(1937), ZN => n1067);
   U1410 : NAND3_X1 port map( A1 => n1069, A2 => n1068, A3 => n1067, ZN => 
                           curr_proc_regs(401));
   U1411 : NAND2_X1 port map( A1 => regs(914), A2 => n15, ZN => n1072);
   U1412 : AOI22_X1 port map( A1 => n29, A2 => regs(1426), B1 => n1596, B2 => 
                           regs(402), ZN => n1071);
   U1413 : AOI22_X1 port map( A1 => n47, A2 => regs(2450), B1 => n1598, B2 => 
                           regs(1938), ZN => n1070);
   U1414 : NAND3_X1 port map( A1 => n1072, A2 => n1071, A3 => n1070, ZN => 
                           curr_proc_regs(402));
   U1415 : NAND2_X1 port map( A1 => regs(915), A2 => n1, ZN => n1075);
   U1416 : AOI22_X1 port map( A1 => n29, A2 => regs(1427), B1 => n23, B2 => 
                           regs(403), ZN => n1074);
   U1417 : AOI22_X1 port map( A1 => n46, A2 => regs(2451), B1 => n40, B2 => 
                           regs(1939), ZN => n1073);
   U1418 : NAND3_X1 port map( A1 => n1075, A2 => n1074, A3 => n1073, ZN => 
                           curr_proc_regs(403));
   U1419 : NAND2_X1 port map( A1 => regs(916), A2 => n4, ZN => n1078);
   U1420 : AOI22_X1 port map( A1 => n29, A2 => regs(1428), B1 => n23, B2 => 
                           regs(404), ZN => n1077);
   U1421 : AOI22_X1 port map( A1 => n50, A2 => regs(2452), B1 => n40, B2 => 
                           regs(1940), ZN => n1076);
   U1422 : NAND3_X1 port map( A1 => n1078, A2 => n1077, A3 => n1076, ZN => 
                           curr_proc_regs(404));
   U1423 : NAND2_X1 port map( A1 => regs(917), A2 => n15, ZN => n1081);
   U1424 : AOI22_X1 port map( A1 => n29, A2 => regs(1429), B1 => n23, B2 => 
                           regs(405), ZN => n1080);
   U1425 : AOI22_X1 port map( A1 => n44, A2 => regs(2453), B1 => n40, B2 => 
                           regs(1941), ZN => n1079);
   U1426 : NAND3_X1 port map( A1 => n1081, A2 => n1080, A3 => n1079, ZN => 
                           curr_proc_regs(405));
   U1427 : NAND2_X1 port map( A1 => regs(918), A2 => n1, ZN => n1084);
   U1428 : AOI22_X1 port map( A1 => n29, A2 => regs(1430), B1 => n23, B2 => 
                           regs(406), ZN => n1083);
   U1429 : AOI22_X1 port map( A1 => n53, A2 => regs(2454), B1 => n40, B2 => 
                           regs(1942), ZN => n1082);
   U1430 : NAND3_X1 port map( A1 => n1084, A2 => n1083, A3 => n1082, ZN => 
                           curr_proc_regs(406));
   U1431 : NAND2_X1 port map( A1 => regs(919), A2 => n13, ZN => n1087);
   U1432 : AOI22_X1 port map( A1 => n29, A2 => regs(1431), B1 => n23, B2 => 
                           regs(407), ZN => n1086);
   U1433 : AOI22_X1 port map( A1 => n55, A2 => regs(2455), B1 => n40, B2 => 
                           regs(1943), ZN => n1085);
   U1434 : NAND3_X1 port map( A1 => n1087, A2 => n1086, A3 => n1085, ZN => 
                           curr_proc_regs(407));
   U1435 : NAND2_X1 port map( A1 => regs(920), A2 => n4, ZN => n1090);
   U1436 : AOI22_X1 port map( A1 => n29, A2 => regs(1432), B1 => n23, B2 => 
                           regs(408), ZN => n1089);
   U1437 : AOI22_X1 port map( A1 => n52, A2 => regs(2456), B1 => n40, B2 => 
                           regs(1944), ZN => n1088);
   U1438 : NAND3_X1 port map( A1 => n1090, A2 => n1089, A3 => n1088, ZN => 
                           curr_proc_regs(408));
   U1439 : NAND2_X1 port map( A1 => regs(921), A2 => n15, ZN => n1093);
   U1440 : AOI22_X1 port map( A1 => n29, A2 => regs(1433), B1 => n23, B2 => 
                           regs(409), ZN => n1092);
   U1441 : AOI22_X1 port map( A1 => win(4), A2 => regs(2457), B1 => n40, B2 => 
                           regs(1945), ZN => n1091);
   U1442 : NAND3_X1 port map( A1 => n1093, A2 => n1092, A3 => n1091, ZN => 
                           curr_proc_regs(409));
   U1443 : NAND2_X1 port map( A1 => regs(552), A2 => n1, ZN => n1096);
   U1444 : AOI22_X1 port map( A1 => n31, A2 => regs(1064), B1 => n23, B2 => 
                           regs(40), ZN => n1095);
   U1445 : AOI22_X1 port map( A1 => n56, A2 => regs(2088), B1 => n40, B2 => 
                           regs(1576), ZN => n1094);
   U1446 : NAND3_X1 port map( A1 => n1096, A2 => n1095, A3 => n1094, ZN => 
                           curr_proc_regs(40));
   U1447 : NAND2_X1 port map( A1 => regs(922), A2 => n13, ZN => n1099);
   U1448 : AOI22_X1 port map( A1 => n29, A2 => regs(1434), B1 => n23, B2 => 
                           regs(410), ZN => n1098);
   U1449 : AOI22_X1 port map( A1 => n43, A2 => regs(2458), B1 => n40, B2 => 
                           regs(1946), ZN => n1097);
   U1450 : NAND3_X1 port map( A1 => n1099, A2 => n1098, A3 => n1097, ZN => 
                           curr_proc_regs(410));
   U1451 : NAND2_X1 port map( A1 => regs(923), A2 => n4, ZN => n1102);
   U1452 : AOI22_X1 port map( A1 => n30, A2 => regs(1435), B1 => n23, B2 => 
                           regs(411), ZN => n1101);
   U1453 : AOI22_X1 port map( A1 => n45, A2 => regs(2459), B1 => n40, B2 => 
                           regs(1947), ZN => n1100);
   U1454 : NAND3_X1 port map( A1 => n1102, A2 => n1101, A3 => n1100, ZN => 
                           curr_proc_regs(411));
   U1455 : NAND2_X1 port map( A1 => regs(924), A2 => n15, ZN => n1105);
   U1456 : AOI22_X1 port map( A1 => n29, A2 => regs(1436), B1 => n23, B2 => 
                           regs(412), ZN => n1104);
   U1457 : AOI22_X1 port map( A1 => n49, A2 => regs(2460), B1 => n40, B2 => 
                           regs(1948), ZN => n1103);
   U1458 : NAND3_X1 port map( A1 => n1105, A2 => n1104, A3 => n1103, ZN => 
                           curr_proc_regs(412));
   U1459 : NAND2_X1 port map( A1 => regs(925), A2 => n12, ZN => n1108);
   U1460 : AOI22_X1 port map( A1 => n30, A2 => regs(1437), B1 => n23, B2 => 
                           regs(413), ZN => n1107);
   U1461 : AOI22_X1 port map( A1 => n43, A2 => regs(2461), B1 => n40, B2 => 
                           regs(1949), ZN => n1106);
   U1462 : NAND3_X1 port map( A1 => n1108, A2 => n1107, A3 => n1106, ZN => 
                           curr_proc_regs(413));
   U1463 : NAND2_X1 port map( A1 => regs(926), A2 => n1, ZN => n1111);
   U1464 : AOI22_X1 port map( A1 => n29, A2 => regs(1438), B1 => n23, B2 => 
                           regs(414), ZN => n1110);
   U1465 : AOI22_X1 port map( A1 => n43, A2 => regs(2462), B1 => n40, B2 => 
                           regs(1950), ZN => n1109);
   U1466 : NAND3_X1 port map( A1 => n1111, A2 => n1110, A3 => n1109, ZN => 
                           curr_proc_regs(414));
   U1467 : NAND2_X1 port map( A1 => regs(927), A2 => n15, ZN => n1114);
   U1468 : AOI22_X1 port map( A1 => n30, A2 => regs(1439), B1 => n1596, B2 => 
                           regs(415), ZN => n1113);
   U1469 : AOI22_X1 port map( A1 => n43, A2 => regs(2463), B1 => n38, B2 => 
                           regs(1951), ZN => n1112);
   U1470 : NAND3_X1 port map( A1 => n1114, A2 => n1113, A3 => n1112, ZN => 
                           curr_proc_regs(415));
   U1471 : NAND2_X1 port map( A1 => regs(928), A2 => n12, ZN => n1117);
   U1472 : AOI22_X1 port map( A1 => n29, A2 => regs(1440), B1 => n23, B2 => 
                           regs(416), ZN => n1116);
   U1473 : AOI22_X1 port map( A1 => n43, A2 => regs(2464), B1 => n40, B2 => 
                           regs(1952), ZN => n1115);
   U1474 : NAND3_X1 port map( A1 => n1117, A2 => n1116, A3 => n1115, ZN => 
                           curr_proc_regs(416));
   U1475 : NAND2_X1 port map( A1 => regs(929), A2 => n14, ZN => n1120);
   U1476 : AOI22_X1 port map( A1 => n30, A2 => regs(1441), B1 => n23, B2 => 
                           regs(417), ZN => n1119);
   U1477 : AOI22_X1 port map( A1 => n43, A2 => regs(2465), B1 => n40, B2 => 
                           regs(1953), ZN => n1118);
   U1478 : NAND3_X1 port map( A1 => n1120, A2 => n1119, A3 => n1118, ZN => 
                           curr_proc_regs(417));
   U1479 : NAND2_X1 port map( A1 => regs(930), A2 => n14, ZN => n1123);
   U1480 : AOI22_X1 port map( A1 => n29, A2 => regs(1442), B1 => n1596, B2 => 
                           regs(418), ZN => n1122);
   U1481 : AOI22_X1 port map( A1 => n43, A2 => regs(2466), B1 => n36, B2 => 
                           regs(1954), ZN => n1121);
   U1482 : NAND3_X1 port map( A1 => n1123, A2 => n1122, A3 => n1121, ZN => 
                           curr_proc_regs(418));
   U1483 : NAND2_X1 port map( A1 => regs(931), A2 => n12, ZN => n1126);
   U1484 : AOI22_X1 port map( A1 => n30, A2 => regs(1443), B1 => n23, B2 => 
                           regs(419), ZN => n1125);
   U1485 : AOI22_X1 port map( A1 => n43, A2 => regs(2467), B1 => n40, B2 => 
                           regs(1955), ZN => n1124);
   U1486 : NAND3_X1 port map( A1 => n1126, A2 => n1125, A3 => n1124, ZN => 
                           curr_proc_regs(419));
   U1487 : NAND2_X1 port map( A1 => regs(553), A2 => n15, ZN => n1129);
   U1488 : AOI22_X1 port map( A1 => n29, A2 => regs(1065), B1 => n23, B2 => 
                           regs(41), ZN => n1128);
   U1489 : AOI22_X1 port map( A1 => n43, A2 => regs(2089), B1 => n40, B2 => 
                           regs(1577), ZN => n1127);
   U1490 : NAND3_X1 port map( A1 => n1129, A2 => n1128, A3 => n1127, ZN => 
                           curr_proc_regs(41));
   U1491 : NAND2_X1 port map( A1 => regs(932), A2 => n1, ZN => n1132);
   U1492 : AOI22_X1 port map( A1 => n29, A2 => regs(1444), B1 => n26, B2 => 
                           regs(420), ZN => n1131);
   U1493 : AOI22_X1 port map( A1 => n43, A2 => regs(2468), B1 => n35, B2 => 
                           regs(1956), ZN => n1130);
   U1494 : NAND3_X1 port map( A1 => n1132, A2 => n1131, A3 => n1130, ZN => 
                           curr_proc_regs(420));
   U1495 : NAND2_X1 port map( A1 => regs(933), A2 => n12, ZN => n1135);
   U1496 : AOI22_X1 port map( A1 => n29, A2 => regs(1445), B1 => n23, B2 => 
                           regs(421), ZN => n1134);
   U1497 : AOI22_X1 port map( A1 => n43, A2 => regs(2469), B1 => n40, B2 => 
                           regs(1957), ZN => n1133);
   U1498 : NAND3_X1 port map( A1 => n1135, A2 => n1134, A3 => n1133, ZN => 
                           curr_proc_regs(421));
   U1499 : NAND2_X1 port map( A1 => regs(934), A2 => n4, ZN => n1138);
   U1500 : AOI22_X1 port map( A1 => n31, A2 => regs(1446), B1 => n23, B2 => 
                           regs(422), ZN => n1137);
   U1501 : AOI22_X1 port map( A1 => n43, A2 => regs(2470), B1 => n40, B2 => 
                           regs(1958), ZN => n1136);
   U1502 : NAND3_X1 port map( A1 => n1138, A2 => n1137, A3 => n1136, ZN => 
                           curr_proc_regs(422));
   U1503 : NAND2_X1 port map( A1 => regs(935), A2 => n13, ZN => n1141);
   U1504 : AOI22_X1 port map( A1 => n31, A2 => regs(1447), B1 => n1596, B2 => 
                           regs(423), ZN => n1140);
   U1505 : AOI22_X1 port map( A1 => n43, A2 => regs(2471), B1 => n36, B2 => 
                           regs(1959), ZN => n1139);
   U1506 : NAND3_X1 port map( A1 => n1141, A2 => n1140, A3 => n1139, ZN => 
                           curr_proc_regs(423));
   U1507 : NAND2_X1 port map( A1 => regs(936), A2 => n12, ZN => n1144);
   U1508 : AOI22_X1 port map( A1 => n2, A2 => regs(1448), B1 => n23, B2 => 
                           regs(424), ZN => n1143);
   U1509 : AOI22_X1 port map( A1 => n49, A2 => regs(2472), B1 => n40, B2 => 
                           regs(1960), ZN => n1142);
   U1510 : NAND3_X1 port map( A1 => n1144, A2 => n1143, A3 => n1142, ZN => 
                           curr_proc_regs(424));
   U1511 : NAND2_X1 port map( A1 => regs(937), A2 => n12, ZN => n1147);
   U1512 : AOI22_X1 port map( A1 => n30, A2 => regs(1449), B1 => n23, B2 => 
                           regs(425), ZN => n1146);
   U1513 : AOI22_X1 port map( A1 => n51, A2 => regs(2473), B1 => n40, B2 => 
                           regs(1961), ZN => n1145);
   U1514 : NAND3_X1 port map( A1 => n1147, A2 => n1146, A3 => n1145, ZN => 
                           curr_proc_regs(425));
   U1515 : NAND2_X1 port map( A1 => regs(938), A2 => n12, ZN => n1150);
   U1516 : AOI22_X1 port map( A1 => n2, A2 => regs(1450), B1 => n23, B2 => 
                           regs(426), ZN => n1149);
   U1517 : AOI22_X1 port map( A1 => n50, A2 => regs(2474), B1 => n40, B2 => 
                           regs(1962), ZN => n1148);
   U1518 : NAND3_X1 port map( A1 => n1150, A2 => n1149, A3 => n1148, ZN => 
                           curr_proc_regs(426));
   U1519 : NAND2_X1 port map( A1 => regs(939), A2 => n12, ZN => n1153);
   U1520 : AOI22_X1 port map( A1 => n29, A2 => regs(1451), B1 => n23, B2 => 
                           regs(427), ZN => n1152);
   U1521 : AOI22_X1 port map( A1 => n46, A2 => regs(2475), B1 => n40, B2 => 
                           regs(1963), ZN => n1151);
   U1522 : NAND3_X1 port map( A1 => n1153, A2 => n1152, A3 => n1151, ZN => 
                           curr_proc_regs(427));
   U1523 : NAND2_X1 port map( A1 => regs(940), A2 => n12, ZN => n1156);
   U1524 : AOI22_X1 port map( A1 => n30, A2 => regs(1452), B1 => n23, B2 => 
                           regs(428), ZN => n1155);
   U1525 : AOI22_X1 port map( A1 => n54, A2 => regs(2476), B1 => n40, B2 => 
                           regs(1964), ZN => n1154);
   U1526 : NAND3_X1 port map( A1 => n1156, A2 => n1155, A3 => n1154, ZN => 
                           curr_proc_regs(428));
   U1527 : NAND2_X1 port map( A1 => regs(941), A2 => n12, ZN => n1159);
   U1528 : AOI22_X1 port map( A1 => n29, A2 => regs(1453), B1 => n23, B2 => 
                           regs(429), ZN => n1158);
   U1529 : AOI22_X1 port map( A1 => n47, A2 => regs(2477), B1 => n40, B2 => 
                           regs(1965), ZN => n1157);
   U1530 : NAND3_X1 port map( A1 => n1159, A2 => n1158, A3 => n1157, ZN => 
                           curr_proc_regs(429));
   U1531 : NAND2_X1 port map( A1 => regs(554), A2 => n12, ZN => n1162);
   U1532 : AOI22_X1 port map( A1 => n2, A2 => regs(1066), B1 => n23, B2 => 
                           regs(42), ZN => n1161);
   U1533 : AOI22_X1 port map( A1 => n48, A2 => regs(2090), B1 => n40, B2 => 
                           regs(1578), ZN => n1160);
   U1534 : NAND3_X1 port map( A1 => n1162, A2 => n1161, A3 => n1160, ZN => 
                           curr_proc_regs(42));
   U1535 : NAND2_X1 port map( A1 => regs(942), A2 => n12, ZN => n1165);
   U1536 : AOI22_X1 port map( A1 => n2, A2 => regs(1454), B1 => n23, B2 => 
                           regs(430), ZN => n1164);
   U1537 : AOI22_X1 port map( A1 => n44, A2 => regs(2478), B1 => n40, B2 => 
                           regs(1966), ZN => n1163);
   U1538 : NAND3_X1 port map( A1 => n1165, A2 => n1164, A3 => n1163, ZN => 
                           curr_proc_regs(430));
   U1539 : NAND2_X1 port map( A1 => regs(943), A2 => n12, ZN => n1168);
   U1540 : AOI22_X1 port map( A1 => n31, A2 => regs(1455), B1 => n23, B2 => 
                           regs(431), ZN => n1167);
   U1541 : AOI22_X1 port map( A1 => n50, A2 => regs(2479), B1 => n40, B2 => 
                           regs(1967), ZN => n1166);
   U1542 : NAND3_X1 port map( A1 => n1168, A2 => n1167, A3 => n1166, ZN => 
                           curr_proc_regs(431));
   U1543 : NAND2_X1 port map( A1 => regs(944), A2 => n12, ZN => n1171);
   U1544 : AOI22_X1 port map( A1 => n31, A2 => regs(1456), B1 => n23, B2 => 
                           regs(432), ZN => n1170);
   U1545 : AOI22_X1 port map( A1 => n46, A2 => regs(2480), B1 => n40, B2 => 
                           regs(1968), ZN => n1169);
   U1546 : NAND3_X1 port map( A1 => n1171, A2 => n1170, A3 => n1169, ZN => 
                           curr_proc_regs(432));
   U1547 : NAND2_X1 port map( A1 => regs(945), A2 => n12, ZN => n1174);
   U1548 : AOI22_X1 port map( A1 => n2, A2 => regs(1457), B1 => n23, B2 => 
                           regs(433), ZN => n1173);
   U1549 : AOI22_X1 port map( A1 => n47, A2 => regs(2481), B1 => n40, B2 => 
                           regs(1969), ZN => n1172);
   U1550 : NAND3_X1 port map( A1 => n1174, A2 => n1173, A3 => n1172, ZN => 
                           curr_proc_regs(433));
   U1551 : NAND2_X1 port map( A1 => regs(946), A2 => n12, ZN => n1177);
   U1552 : AOI22_X1 port map( A1 => n30, A2 => regs(1458), B1 => n23, B2 => 
                           regs(434), ZN => n1176);
   U1553 : AOI22_X1 port map( A1 => n44, A2 => regs(2482), B1 => n40, B2 => 
                           regs(1970), ZN => n1175);
   U1554 : NAND3_X1 port map( A1 => n1177, A2 => n1176, A3 => n1175, ZN => 
                           curr_proc_regs(434));
   U1555 : NAND2_X1 port map( A1 => regs(947), A2 => n1, ZN => n1180);
   U1556 : AOI22_X1 port map( A1 => n2, A2 => regs(1459), B1 => n23, B2 => 
                           regs(435), ZN => n1179);
   U1557 : AOI22_X1 port map( A1 => n54, A2 => regs(2483), B1 => n35, B2 => 
                           regs(1971), ZN => n1178);
   U1558 : NAND3_X1 port map( A1 => n1180, A2 => n1179, A3 => n1178, ZN => 
                           curr_proc_regs(435));
   U1559 : NAND2_X1 port map( A1 => regs(948), A2 => n12, ZN => n1183);
   U1560 : AOI22_X1 port map( A1 => n29, A2 => regs(1460), B1 => n23, B2 => 
                           regs(436), ZN => n1182);
   U1561 : AOI22_X1 port map( A1 => n47, A2 => regs(2484), B1 => n40, B2 => 
                           regs(1972), ZN => n1181);
   U1562 : NAND3_X1 port map( A1 => n1183, A2 => n1182, A3 => n1181, ZN => 
                           curr_proc_regs(436));
   U1563 : NAND2_X1 port map( A1 => regs(949), A2 => n13, ZN => n1186);
   U1564 : AOI22_X1 port map( A1 => n29, A2 => regs(1461), B1 => n23, B2 => 
                           regs(437), ZN => n1185);
   U1565 : AOI22_X1 port map( A1 => n48, A2 => regs(2485), B1 => n40, B2 => 
                           regs(1973), ZN => n1184);
   U1566 : NAND3_X1 port map( A1 => n1186, A2 => n1185, A3 => n1184, ZN => 
                           curr_proc_regs(437));
   U1567 : NAND2_X1 port map( A1 => regs(950), A2 => n12, ZN => n1189);
   U1568 : AOI22_X1 port map( A1 => n2, A2 => regs(1462), B1 => n23, B2 => 
                           regs(438), ZN => n1188);
   U1569 : AOI22_X1 port map( A1 => n44, A2 => regs(2486), B1 => n40, B2 => 
                           regs(1974), ZN => n1187);
   U1570 : NAND3_X1 port map( A1 => n1189, A2 => n1188, A3 => n1187, ZN => 
                           curr_proc_regs(438));
   U1571 : NAND2_X1 port map( A1 => regs(951), A2 => n13, ZN => n1192);
   U1572 : AOI22_X1 port map( A1 => n32, A2 => regs(1463), B1 => n21, B2 => 
                           regs(439), ZN => n1191);
   U1573 : AOI22_X1 port map( A1 => n52, A2 => regs(2487), B1 => n40, B2 => 
                           regs(1975), ZN => n1190);
   U1574 : NAND3_X1 port map( A1 => n1192, A2 => n1191, A3 => n1190, ZN => 
                           curr_proc_regs(439));
   U1575 : NAND2_X1 port map( A1 => regs(555), A2 => n12, ZN => n1195);
   U1576 : AOI22_X1 port map( A1 => n30, A2 => regs(1067), B1 => n23, B2 => 
                           regs(43), ZN => n1194);
   U1577 : AOI22_X1 port map( A1 => n53, A2 => regs(2091), B1 => n40, B2 => 
                           regs(1579), ZN => n1193);
   U1578 : NAND3_X1 port map( A1 => n1195, A2 => n1194, A3 => n1193, ZN => 
                           curr_proc_regs(43));
   U1579 : NAND2_X1 port map( A1 => regs(952), A2 => n1, ZN => n1198);
   U1580 : AOI22_X1 port map( A1 => n29, A2 => regs(1464), B1 => n23, B2 => 
                           regs(440), ZN => n1197);
   U1581 : AOI22_X1 port map( A1 => n55, A2 => regs(2488), B1 => n40, B2 => 
                           regs(1976), ZN => n1196);
   U1582 : NAND3_X1 port map( A1 => n1198, A2 => n1197, A3 => n1196, ZN => 
                           curr_proc_regs(440));
   U1583 : NAND2_X1 port map( A1 => regs(953), A2 => n14, ZN => n1201);
   U1584 : AOI22_X1 port map( A1 => n29, A2 => regs(1465), B1 => n23, B2 => 
                           regs(441), ZN => n1200);
   U1585 : AOI22_X1 port map( A1 => win(4), A2 => regs(2489), B1 => n40, B2 => 
                           regs(1977), ZN => n1199);
   U1586 : NAND3_X1 port map( A1 => n1201, A2 => n1200, A3 => n1199, ZN => 
                           curr_proc_regs(441));
   U1587 : NAND2_X1 port map( A1 => regs(954), A2 => n4, ZN => n1204);
   U1588 : AOI22_X1 port map( A1 => n2, A2 => regs(1466), B1 => n19, B2 => 
                           regs(442), ZN => n1203);
   U1589 : AOI22_X1 port map( A1 => n44, A2 => regs(2490), B1 => n39, B2 => 
                           regs(1978), ZN => n1202);
   U1590 : NAND3_X1 port map( A1 => n1204, A2 => n1203, A3 => n1202, ZN => 
                           curr_proc_regs(442));
   U1591 : NAND2_X1 port map( A1 => regs(955), A2 => n15, ZN => n1207);
   U1592 : AOI22_X1 port map( A1 => n31, A2 => regs(1467), B1 => n23, B2 => 
                           regs(443), ZN => n1206);
   U1593 : AOI22_X1 port map( A1 => n45, A2 => regs(2491), B1 => n40, B2 => 
                           regs(1979), ZN => n1205);
   U1594 : NAND3_X1 port map( A1 => n1207, A2 => n1206, A3 => n1205, ZN => 
                           curr_proc_regs(443));
   U1595 : NAND2_X1 port map( A1 => regs(956), A2 => n4, ZN => n1210);
   U1596 : AOI22_X1 port map( A1 => n30, A2 => regs(1468), B1 => n23, B2 => 
                           regs(444), ZN => n1209);
   U1597 : AOI22_X1 port map( A1 => n44, A2 => regs(2492), B1 => n40, B2 => 
                           regs(1980), ZN => n1208);
   U1598 : NAND3_X1 port map( A1 => n1210, A2 => n1209, A3 => n1208, ZN => 
                           curr_proc_regs(444));
   U1599 : NAND2_X1 port map( A1 => regs(957), A2 => n13, ZN => n1213);
   U1600 : AOI22_X1 port map( A1 => n2, A2 => regs(1469), B1 => n23, B2 => 
                           regs(445), ZN => n1212);
   U1601 : AOI22_X1 port map( A1 => n6, A2 => regs(2493), B1 => n40, B2 => 
                           regs(1981), ZN => n1211);
   U1602 : NAND3_X1 port map( A1 => n1213, A2 => n1212, A3 => n1211, ZN => 
                           curr_proc_regs(445));
   U1603 : NAND2_X1 port map( A1 => regs(958), A2 => n12, ZN => n1216);
   U1604 : AOI22_X1 port map( A1 => n29, A2 => regs(1470), B1 => n23, B2 => 
                           regs(446), ZN => n1215);
   U1605 : AOI22_X1 port map( A1 => n6, A2 => regs(2494), B1 => n40, B2 => 
                           regs(1982), ZN => n1214);
   U1606 : NAND3_X1 port map( A1 => n1216, A2 => n1215, A3 => n1214, ZN => 
                           curr_proc_regs(446));
   U1607 : NAND2_X1 port map( A1 => regs(959), A2 => n1, ZN => n1219);
   U1608 : AOI22_X1 port map( A1 => n32, A2 => regs(1471), B1 => n23, B2 => 
                           regs(447), ZN => n1218);
   U1609 : AOI22_X1 port map( A1 => n6, A2 => regs(2495), B1 => n40, B2 => 
                           regs(1983), ZN => n1217);
   U1610 : NAND3_X1 port map( A1 => n1219, A2 => n1218, A3 => n1217, ZN => 
                           curr_proc_regs(447));
   U1611 : NAND2_X1 port map( A1 => regs(960), A2 => n14, ZN => n1222);
   U1612 : AOI22_X1 port map( A1 => n2, A2 => regs(1472), B1 => n23, B2 => 
                           regs(448), ZN => n1221);
   U1613 : AOI22_X1 port map( A1 => n6, A2 => regs(2496), B1 => n40, B2 => 
                           regs(1984), ZN => n1220);
   U1614 : NAND3_X1 port map( A1 => n1222, A2 => n1221, A3 => n1220, ZN => 
                           curr_proc_regs(448));
   U1615 : NAND2_X1 port map( A1 => regs(961), A2 => n15, ZN => n1225);
   U1616 : AOI22_X1 port map( A1 => n30, A2 => regs(1473), B1 => n23, B2 => 
                           regs(449), ZN => n1224);
   U1617 : AOI22_X1 port map( A1 => n6, A2 => regs(2497), B1 => n40, B2 => 
                           regs(1985), ZN => n1223);
   U1618 : NAND3_X1 port map( A1 => n1225, A2 => n1224, A3 => n1223, ZN => 
                           curr_proc_regs(449));
   U1619 : NAND2_X1 port map( A1 => regs(556), A2 => n14, ZN => n1228);
   U1620 : AOI22_X1 port map( A1 => n29, A2 => regs(1068), B1 => n21, B2 => 
                           regs(44), ZN => n1227);
   U1621 : AOI22_X1 port map( A1 => n56, A2 => regs(2092), B1 => n36, B2 => 
                           regs(1580), ZN => n1226);
   U1622 : NAND3_X1 port map( A1 => n1228, A2 => n1227, A3 => n1226, ZN => 
                           curr_proc_regs(44));
   U1623 : NAND2_X1 port map( A1 => regs(962), A2 => n12, ZN => n1231);
   U1624 : AOI22_X1 port map( A1 => n29, A2 => regs(1474), B1 => n23, B2 => 
                           regs(450), ZN => n1230);
   U1625 : AOI22_X1 port map( A1 => n43, A2 => regs(2498), B1 => n40, B2 => 
                           regs(1986), ZN => n1229);
   U1626 : NAND3_X1 port map( A1 => n1231, A2 => n1230, A3 => n1229, ZN => 
                           curr_proc_regs(450));
   U1627 : NAND2_X1 port map( A1 => regs(963), A2 => n4, ZN => n1234);
   U1628 : AOI22_X1 port map( A1 => n2, A2 => regs(1475), B1 => n23, B2 => 
                           regs(451), ZN => n1233);
   U1629 : AOI22_X1 port map( A1 => n45, A2 => regs(2499), B1 => n40, B2 => 
                           regs(1987), ZN => n1232);
   U1630 : NAND3_X1 port map( A1 => n1234, A2 => n1233, A3 => n1232, ZN => 
                           curr_proc_regs(451));
   U1631 : NAND2_X1 port map( A1 => regs(964), A2 => n13, ZN => n1237);
   U1632 : AOI22_X1 port map( A1 => n29, A2 => regs(1476), B1 => n23, B2 => 
                           regs(452), ZN => n1236);
   U1633 : AOI22_X1 port map( A1 => n49, A2 => regs(2500), B1 => n40, B2 => 
                           regs(1988), ZN => n1235);
   U1634 : NAND3_X1 port map( A1 => n1237, A2 => n1236, A3 => n1235, ZN => 
                           curr_proc_regs(452));
   U1635 : NAND2_X1 port map( A1 => regs(965), A2 => n1, ZN => n1240);
   U1636 : AOI22_X1 port map( A1 => n28, A2 => regs(1477), B1 => n23, B2 => 
                           regs(453), ZN => n1239);
   U1637 : AOI22_X1 port map( A1 => n48, A2 => regs(2501), B1 => n40, B2 => 
                           regs(1989), ZN => n1238);
   U1638 : NAND3_X1 port map( A1 => n1240, A2 => n1239, A3 => n1238, ZN => 
                           curr_proc_regs(453));
   U1639 : NAND2_X1 port map( A1 => regs(966), A2 => n14, ZN => n1243);
   U1640 : AOI22_X1 port map( A1 => n28, A2 => regs(1478), B1 => n23, B2 => 
                           regs(454), ZN => n1242);
   U1641 : AOI22_X1 port map( A1 => n54, A2 => regs(2502), B1 => n40, B2 => 
                           regs(1990), ZN => n1241);
   U1642 : NAND3_X1 port map( A1 => n1243, A2 => n1242, A3 => n1241, ZN => 
                           curr_proc_regs(454));
   U1643 : NAND2_X1 port map( A1 => regs(967), A2 => n15, ZN => n1246);
   U1644 : AOI22_X1 port map( A1 => n28, A2 => regs(1479), B1 => n23, B2 => 
                           regs(455), ZN => n1245);
   U1645 : AOI22_X1 port map( A1 => n51, A2 => regs(2503), B1 => n40, B2 => 
                           regs(1991), ZN => n1244);
   U1646 : NAND3_X1 port map( A1 => n1246, A2 => n1245, A3 => n1244, ZN => 
                           curr_proc_regs(455));
   U1647 : NAND2_X1 port map( A1 => regs(968), A2 => n4, ZN => n1249);
   U1648 : AOI22_X1 port map( A1 => n28, A2 => regs(1480), B1 => n23, B2 => 
                           regs(456), ZN => n1248);
   U1649 : AOI22_X1 port map( A1 => n47, A2 => regs(2504), B1 => n40, B2 => 
                           regs(1992), ZN => n1247);
   U1650 : NAND3_X1 port map( A1 => n1249, A2 => n1248, A3 => n1247, ZN => 
                           curr_proc_regs(456));
   U1651 : NAND2_X1 port map( A1 => regs(969), A2 => n14, ZN => n1252);
   U1652 : AOI22_X1 port map( A1 => n28, A2 => regs(1481), B1 => n19, B2 => 
                           regs(457), ZN => n1251);
   U1653 : AOI22_X1 port map( A1 => n46, A2 => regs(2505), B1 => n40, B2 => 
                           regs(1993), ZN => n1250);
   U1654 : NAND3_X1 port map( A1 => n1252, A2 => n1251, A3 => n1250, ZN => 
                           curr_proc_regs(457));
   U1655 : NAND2_X1 port map( A1 => regs(970), A2 => n1595, ZN => n1255);
   U1656 : AOI22_X1 port map( A1 => n28, A2 => regs(1482), B1 => n20, B2 => 
                           regs(458), ZN => n1254);
   U1657 : AOI22_X1 port map( A1 => n50, A2 => regs(2506), B1 => n35, B2 => 
                           regs(1994), ZN => n1253);
   U1658 : NAND3_X1 port map( A1 => n1255, A2 => n1254, A3 => n1253, ZN => 
                           curr_proc_regs(458));
   U1659 : NAND2_X1 port map( A1 => regs(971), A2 => n14, ZN => n1258);
   U1660 : AOI22_X1 port map( A1 => n28, A2 => regs(1483), B1 => n19, B2 => 
                           regs(459), ZN => n1257);
   U1661 : AOI22_X1 port map( A1 => n53, A2 => regs(2507), B1 => n35, B2 => 
                           regs(1995), ZN => n1256);
   U1662 : NAND3_X1 port map( A1 => n1258, A2 => n1257, A3 => n1256, ZN => 
                           curr_proc_regs(459));
   U1663 : NAND2_X1 port map( A1 => regs(557), A2 => n14, ZN => n1261);
   U1664 : AOI22_X1 port map( A1 => n28, A2 => regs(1069), B1 => n1596, B2 => 
                           regs(45), ZN => n1260);
   U1665 : AOI22_X1 port map( A1 => n55, A2 => regs(2093), B1 => n36, B2 => 
                           regs(1581), ZN => n1259);
   U1666 : NAND3_X1 port map( A1 => n1261, A2 => n1260, A3 => n1259, ZN => 
                           curr_proc_regs(45));
   U1667 : NAND2_X1 port map( A1 => regs(972), A2 => n1595, ZN => n1264);
   U1668 : AOI22_X1 port map( A1 => n28, A2 => regs(1484), B1 => n19, B2 => 
                           regs(460), ZN => n1263);
   U1669 : AOI22_X1 port map( A1 => n43, A2 => regs(2508), B1 => n35, B2 => 
                           regs(1996), ZN => n1262);
   U1670 : NAND3_X1 port map( A1 => n1264, A2 => n1263, A3 => n1262, ZN => 
                           curr_proc_regs(460));
   U1671 : NAND2_X1 port map( A1 => regs(973), A2 => n14, ZN => n1267);
   U1672 : AOI22_X1 port map( A1 => n28, A2 => regs(1485), B1 => n18, B2 => 
                           regs(461), ZN => n1266);
   U1673 : AOI22_X1 port map( A1 => n45, A2 => regs(2509), B1 => n38, B2 => 
                           regs(1997), ZN => n1265);
   U1674 : NAND3_X1 port map( A1 => n1267, A2 => n1266, A3 => n1265, ZN => 
                           curr_proc_regs(461));
   U1675 : NAND2_X1 port map( A1 => regs(974), A2 => n14, ZN => n1270);
   U1676 : AOI22_X1 port map( A1 => n28, A2 => regs(1486), B1 => n19, B2 => 
                           regs(462), ZN => n1269);
   U1677 : AOI22_X1 port map( A1 => n49, A2 => regs(2510), B1 => n35, B2 => 
                           regs(1998), ZN => n1268);
   U1678 : NAND3_X1 port map( A1 => n1270, A2 => n1269, A3 => n1268, ZN => 
                           curr_proc_regs(462));
   U1679 : NAND2_X1 port map( A1 => regs(975), A2 => n1595, ZN => n1273);
   U1680 : AOI22_X1 port map( A1 => n28, A2 => regs(1487), B1 => n23, B2 => 
                           regs(463), ZN => n1272);
   U1681 : AOI22_X1 port map( A1 => n48, A2 => regs(2511), B1 => n39, B2 => 
                           regs(1999), ZN => n1271);
   U1682 : NAND3_X1 port map( A1 => n1273, A2 => n1272, A3 => n1271, ZN => 
                           curr_proc_regs(463));
   U1683 : NAND2_X1 port map( A1 => regs(976), A2 => n14, ZN => n1276);
   U1684 : AOI22_X1 port map( A1 => n2, A2 => regs(1488), B1 => n19, B2 => 
                           regs(464), ZN => n1275);
   U1685 : AOI22_X1 port map( A1 => n54, A2 => regs(2512), B1 => n35, B2 => 
                           regs(2000), ZN => n1274);
   U1686 : NAND3_X1 port map( A1 => n1276, A2 => n1275, A3 => n1274, ZN => 
                           curr_proc_regs(464));
   U1687 : NAND2_X1 port map( A1 => regs(977), A2 => n14, ZN => n1279);
   U1688 : AOI22_X1 port map( A1 => n29, A2 => regs(1489), B1 => n19, B2 => 
                           regs(465), ZN => n1278);
   U1689 : AOI22_X1 port map( A1 => n51, A2 => regs(2513), B1 => n35, B2 => 
                           regs(2001), ZN => n1277);
   U1690 : NAND3_X1 port map( A1 => n1279, A2 => n1278, A3 => n1277, ZN => 
                           curr_proc_regs(465));
   U1691 : NAND2_X1 port map( A1 => regs(978), A2 => n1595, ZN => n1282);
   U1692 : AOI22_X1 port map( A1 => n31, A2 => regs(1490), B1 => n19, B2 => 
                           regs(466), ZN => n1281);
   U1693 : AOI22_X1 port map( A1 => n47, A2 => regs(2514), B1 => n35, B2 => 
                           regs(2002), ZN => n1280);
   U1694 : NAND3_X1 port map( A1 => n1282, A2 => n1281, A3 => n1280, ZN => 
                           curr_proc_regs(466));
   U1695 : NAND2_X1 port map( A1 => regs(979), A2 => n14, ZN => n1285);
   U1696 : AOI22_X1 port map( A1 => n2, A2 => regs(1491), B1 => n19, B2 => 
                           regs(467), ZN => n1284);
   U1697 : AOI22_X1 port map( A1 => n46, A2 => regs(2515), B1 => n35, B2 => 
                           regs(2003), ZN => n1283);
   U1698 : NAND3_X1 port map( A1 => n1285, A2 => n1284, A3 => n1283, ZN => 
                           curr_proc_regs(467));
   U1699 : NAND2_X1 port map( A1 => regs(980), A2 => n1595, ZN => n1288);
   U1700 : AOI22_X1 port map( A1 => n29, A2 => regs(1492), B1 => n1596, B2 => 
                           regs(468), ZN => n1287);
   U1701 : AOI22_X1 port map( A1 => n50, A2 => regs(2516), B1 => n36, B2 => 
                           regs(2004), ZN => n1286);
   U1702 : NAND3_X1 port map( A1 => n1288, A2 => n1287, A3 => n1286, ZN => 
                           curr_proc_regs(468));
   U1703 : NAND2_X1 port map( A1 => regs(981), A2 => n14, ZN => n1291);
   U1704 : AOI22_X1 port map( A1 => n31, A2 => regs(1493), B1 => n19, B2 => 
                           regs(469), ZN => n1290);
   U1705 : AOI22_X1 port map( A1 => n53, A2 => regs(2517), B1 => n35, B2 => 
                           regs(2005), ZN => n1289);
   U1706 : NAND3_X1 port map( A1 => n1291, A2 => n1290, A3 => n1289, ZN => 
                           curr_proc_regs(469));
   U1707 : NAND2_X1 port map( A1 => regs(558), A2 => n14, ZN => n1294);
   U1708 : AOI22_X1 port map( A1 => n2, A2 => regs(1070), B1 => n17, B2 => 
                           regs(46), ZN => n1293);
   U1709 : AOI22_X1 port map( A1 => n55, A2 => regs(2094), B1 => n35, B2 => 
                           regs(1582), ZN => n1292);
   U1710 : NAND3_X1 port map( A1 => n1294, A2 => n1293, A3 => n1292, ZN => 
                           curr_proc_regs(46));
   U1711 : NAND2_X1 port map( A1 => regs(982), A2 => n1595, ZN => n1297);
   U1712 : AOI22_X1 port map( A1 => n29, A2 => regs(1494), B1 => n20, B2 => 
                           regs(470), ZN => n1296);
   U1713 : AOI22_X1 port map( A1 => n52, A2 => regs(2518), B1 => n36, B2 => 
                           regs(2006), ZN => n1295);
   U1714 : NAND3_X1 port map( A1 => n1297, A2 => n1296, A3 => n1295, ZN => 
                           curr_proc_regs(470));
   U1715 : NAND2_X1 port map( A1 => regs(983), A2 => n14, ZN => n1300);
   U1716 : AOI22_X1 port map( A1 => n31, A2 => regs(1495), B1 => n19, B2 => 
                           regs(471), ZN => n1299);
   U1717 : AOI22_X1 port map( A1 => n52, A2 => regs(2519), B1 => n35, B2 => 
                           regs(2007), ZN => n1298);
   U1718 : NAND3_X1 port map( A1 => n1300, A2 => n1299, A3 => n1298, ZN => 
                           curr_proc_regs(471));
   U1719 : NAND2_X1 port map( A1 => regs(984), A2 => n14, ZN => n1303);
   U1720 : AOI22_X1 port map( A1 => n2, A2 => regs(1496), B1 => n19, B2 => 
                           regs(472), ZN => n1302);
   U1721 : AOI22_X1 port map( A1 => n52, A2 => regs(2520), B1 => n39, B2 => 
                           regs(2008), ZN => n1301);
   U1722 : NAND3_X1 port map( A1 => n1303, A2 => n1302, A3 => n1301, ZN => 
                           curr_proc_regs(472));
   U1723 : NAND2_X1 port map( A1 => regs(985), A2 => n14, ZN => n1306);
   U1724 : AOI22_X1 port map( A1 => n29, A2 => regs(1497), B1 => n19, B2 => 
                           regs(473), ZN => n1305);
   U1725 : AOI22_X1 port map( A1 => n52, A2 => regs(2521), B1 => n38, B2 => 
                           regs(2009), ZN => n1304);
   U1726 : NAND3_X1 port map( A1 => n1306, A2 => n1305, A3 => n1304, ZN => 
                           curr_proc_regs(473));
   U1727 : NAND2_X1 port map( A1 => regs(986), A2 => n1595, ZN => n1309);
   U1728 : AOI22_X1 port map( A1 => n31, A2 => regs(1498), B1 => n19, B2 => 
                           regs(474), ZN => n1308);
   U1729 : AOI22_X1 port map( A1 => n52, A2 => regs(2522), B1 => n35, B2 => 
                           regs(2010), ZN => n1307);
   U1730 : NAND3_X1 port map( A1 => n1309, A2 => n1308, A3 => n1307, ZN => 
                           curr_proc_regs(474));
   U1731 : NAND2_X1 port map( A1 => regs(987), A2 => n14, ZN => n1312);
   U1732 : AOI22_X1 port map( A1 => n29, A2 => regs(1499), B1 => n21, B2 => 
                           regs(475), ZN => n1311);
   U1733 : AOI22_X1 port map( A1 => n52, A2 => regs(2523), B1 => n36, B2 => 
                           regs(2011), ZN => n1310);
   U1734 : NAND3_X1 port map( A1 => n1312, A2 => n1311, A3 => n1310, ZN => 
                           curr_proc_regs(475));
   U1735 : NAND2_X1 port map( A1 => regs(988), A2 => n14, ZN => n1315);
   U1736 : AOI22_X1 port map( A1 => n31, A2 => regs(1500), B1 => n26, B2 => 
                           regs(476), ZN => n1314);
   U1737 : AOI22_X1 port map( A1 => n52, A2 => regs(2524), B1 => n35, B2 => 
                           regs(2012), ZN => n1313);
   U1738 : NAND3_X1 port map( A1 => n1315, A2 => n1314, A3 => n1313, ZN => 
                           curr_proc_regs(476));
   U1739 : NAND2_X1 port map( A1 => regs(989), A2 => n14, ZN => n1318);
   U1740 : AOI22_X1 port map( A1 => n2, A2 => regs(1501), B1 => n19, B2 => 
                           regs(477), ZN => n1317);
   U1741 : AOI22_X1 port map( A1 => n52, A2 => regs(2525), B1 => n35, B2 => 
                           regs(2013), ZN => n1316);
   U1742 : NAND3_X1 port map( A1 => n1318, A2 => n1317, A3 => n1316, ZN => 
                           curr_proc_regs(477));
   U1743 : NAND2_X1 port map( A1 => regs(990), A2 => n14, ZN => n1321);
   U1744 : AOI22_X1 port map( A1 => n29, A2 => regs(1502), B1 => n18, B2 => 
                           regs(478), ZN => n1320);
   U1745 : AOI22_X1 port map( A1 => n52, A2 => regs(2526), B1 => n35, B2 => 
                           regs(2014), ZN => n1319);
   U1746 : NAND3_X1 port map( A1 => n1321, A2 => n1320, A3 => n1319, ZN => 
                           curr_proc_regs(478));
   U1747 : NAND2_X1 port map( A1 => regs(991), A2 => n14, ZN => n1324);
   U1748 : AOI22_X1 port map( A1 => n31, A2 => regs(1503), B1 => n26, B2 => 
                           regs(479), ZN => n1323);
   U1749 : AOI22_X1 port map( A1 => n52, A2 => regs(2527), B1 => n39, B2 => 
                           regs(2015), ZN => n1322);
   U1750 : NAND3_X1 port map( A1 => n1324, A2 => n1323, A3 => n1322, ZN => 
                           curr_proc_regs(479));
   U1751 : NAND2_X1 port map( A1 => regs(559), A2 => n14, ZN => n1327);
   U1752 : AOI22_X1 port map( A1 => n2, A2 => regs(1071), B1 => n19, B2 => 
                           regs(47), ZN => n1326);
   U1753 : AOI22_X1 port map( A1 => n52, A2 => regs(2095), B1 => n38, B2 => 
                           regs(1583), ZN => n1325);
   U1754 : NAND3_X1 port map( A1 => n1327, A2 => n1326, A3 => n1325, ZN => 
                           curr_proc_regs(47));
   U1755 : NAND2_X1 port map( A1 => regs(992), A2 => n14, ZN => n1330);
   U1756 : AOI22_X1 port map( A1 => n29, A2 => regs(1504), B1 => n1596, B2 => 
                           regs(480), ZN => n1329);
   U1757 : AOI22_X1 port map( A1 => n52, A2 => regs(2528), B1 => n36, B2 => 
                           regs(2016), ZN => n1328);
   U1758 : NAND3_X1 port map( A1 => n1330, A2 => n1329, A3 => n1328, ZN => 
                           curr_proc_regs(480));
   U1759 : NAND2_X1 port map( A1 => regs(993), A2 => n14, ZN => n1333);
   U1760 : AOI22_X1 port map( A1 => n31, A2 => regs(1505), B1 => n17, B2 => 
                           regs(481), ZN => n1332);
   U1761 : AOI22_X1 port map( A1 => n52, A2 => regs(2529), B1 => n35, B2 => 
                           regs(2017), ZN => n1331);
   U1762 : NAND3_X1 port map( A1 => n1333, A2 => n1332, A3 => n1331, ZN => 
                           curr_proc_regs(481));
   U1763 : NAND2_X1 port map( A1 => regs(994), A2 => n14, ZN => n1336);
   U1764 : AOI22_X1 port map( A1 => n2, A2 => regs(1506), B1 => n20, B2 => 
                           regs(482), ZN => n1335);
   U1765 : AOI22_X1 port map( A1 => n7, A2 => regs(2530), B1 => n36, B2 => 
                           regs(2018), ZN => n1334);
   U1766 : NAND3_X1 port map( A1 => n1336, A2 => n1335, A3 => n1334, ZN => 
                           curr_proc_regs(482));
   U1767 : NAND2_X1 port map( A1 => regs(995), A2 => n14, ZN => n1339);
   U1768 : AOI22_X1 port map( A1 => n29, A2 => regs(1507), B1 => n21, B2 => 
                           regs(483), ZN => n1338);
   U1769 : AOI22_X1 port map( A1 => n7, A2 => regs(2531), B1 => n39, B2 => 
                           regs(2019), ZN => n1337);
   U1770 : NAND3_X1 port map( A1 => n1339, A2 => n1338, A3 => n1337, ZN => 
                           curr_proc_regs(483));
   U1771 : NAND2_X1 port map( A1 => regs(996), A2 => n14, ZN => n1342);
   U1772 : AOI22_X1 port map( A1 => n31, A2 => regs(1508), B1 => n19, B2 => 
                           regs(484), ZN => n1341);
   U1773 : AOI22_X1 port map( A1 => n7, A2 => regs(2532), B1 => n38, B2 => 
                           regs(2020), ZN => n1340);
   U1774 : NAND3_X1 port map( A1 => n1342, A2 => n1341, A3 => n1340, ZN => 
                           curr_proc_regs(484));
   U1775 : NAND2_X1 port map( A1 => regs(997), A2 => n14, ZN => n1345);
   U1776 : AOI22_X1 port map( A1 => n2, A2 => regs(1509), B1 => n21, B2 => 
                           regs(485), ZN => n1344);
   U1777 : AOI22_X1 port map( A1 => n7, A2 => regs(2533), B1 => n36, B2 => 
                           regs(2021), ZN => n1343);
   U1778 : NAND3_X1 port map( A1 => n1345, A2 => n1344, A3 => n1343, ZN => 
                           curr_proc_regs(485));
   U1779 : NAND2_X1 port map( A1 => regs(998), A2 => n14, ZN => n1348);
   U1780 : AOI22_X1 port map( A1 => n30, A2 => regs(1510), B1 => n26, B2 => 
                           regs(486), ZN => n1347);
   U1781 : AOI22_X1 port map( A1 => n7, A2 => regs(2534), B1 => n35, B2 => 
                           regs(2022), ZN => n1346);
   U1782 : NAND3_X1 port map( A1 => n1348, A2 => n1347, A3 => n1346, ZN => 
                           curr_proc_regs(486));
   U1783 : NAND2_X1 port map( A1 => regs(999), A2 => n14, ZN => n1351);
   U1784 : AOI22_X1 port map( A1 => n27, A2 => regs(1511), B1 => n18, B2 => 
                           regs(487), ZN => n1350);
   U1785 : AOI22_X1 port map( A1 => n7, A2 => regs(2535), B1 => n35, B2 => 
                           regs(2023), ZN => n1349);
   U1786 : NAND3_X1 port map( A1 => n1351, A2 => n1350, A3 => n1349, ZN => 
                           curr_proc_regs(487));
   U1787 : NAND2_X1 port map( A1 => regs(1000), A2 => n14, ZN => n1354);
   U1788 : AOI22_X1 port map( A1 => n29, A2 => regs(1512), B1 => n23, B2 => 
                           regs(488), ZN => n1353);
   U1789 : AOI22_X1 port map( A1 => n7, A2 => regs(2536), B1 => n39, B2 => 
                           regs(2024), ZN => n1352);
   U1790 : NAND3_X1 port map( A1 => n1354, A2 => n1353, A3 => n1352, ZN => 
                           curr_proc_regs(488));
   U1791 : NAND2_X1 port map( A1 => regs(1001), A2 => n14, ZN => n1357);
   U1792 : AOI22_X1 port map( A1 => n30, A2 => regs(1513), B1 => n23, B2 => 
                           regs(489), ZN => n1356);
   U1793 : AOI22_X1 port map( A1 => n7, A2 => regs(2537), B1 => n38, B2 => 
                           regs(2025), ZN => n1355);
   U1794 : NAND3_X1 port map( A1 => n1357, A2 => n1356, A3 => n1355, ZN => 
                           curr_proc_regs(489));
   U1795 : NAND2_X1 port map( A1 => regs(560), A2 => n1595, ZN => n1360);
   U1796 : AOI22_X1 port map( A1 => n27, A2 => regs(1072), B1 => n26, B2 => 
                           regs(48), ZN => n1359);
   U1797 : AOI22_X1 port map( A1 => n7, A2 => regs(2096), B1 => n38, B2 => 
                           regs(1584), ZN => n1358);
   U1798 : NAND3_X1 port map( A1 => n1360, A2 => n1359, A3 => n1358, ZN => 
                           curr_proc_regs(48));
   U1799 : NAND2_X1 port map( A1 => regs(1002), A2 => n14, ZN => n1363);
   U1800 : AOI22_X1 port map( A1 => n29, A2 => regs(1514), B1 => n21, B2 => 
                           regs(490), ZN => n1362);
   U1801 : AOI22_X1 port map( A1 => n7, A2 => regs(2538), B1 => n36, B2 => 
                           regs(2026), ZN => n1361);
   U1802 : NAND3_X1 port map( A1 => n1363, A2 => n1362, A3 => n1361, ZN => 
                           curr_proc_regs(490));
   U1803 : NAND2_X1 port map( A1 => regs(1003), A2 => n14, ZN => n1366);
   U1804 : AOI22_X1 port map( A1 => n30, A2 => regs(1515), B1 => n19, B2 => 
                           regs(491), ZN => n1365);
   U1805 : AOI22_X1 port map( A1 => n7, A2 => regs(2539), B1 => n35, B2 => 
                           regs(2027), ZN => n1364);
   U1806 : NAND3_X1 port map( A1 => n1366, A2 => n1365, A3 => n1364, ZN => 
                           curr_proc_regs(491));
   U1807 : NAND2_X1 port map( A1 => regs(1004), A2 => n1595, ZN => n1369);
   U1808 : AOI22_X1 port map( A1 => n27, A2 => regs(1516), B1 => n1596, B2 => 
                           regs(492), ZN => n1368);
   U1809 : AOI22_X1 port map( A1 => n7, A2 => regs(2540), B1 => n35, B2 => 
                           regs(2028), ZN => n1367);
   U1810 : NAND3_X1 port map( A1 => n1369, A2 => n1368, A3 => n1367, ZN => 
                           curr_proc_regs(492));
   U1811 : NAND2_X1 port map( A1 => regs(1005), A2 => n14, ZN => n1372);
   U1812 : AOI22_X1 port map( A1 => n29, A2 => regs(1517), B1 => n21, B2 => 
                           regs(493), ZN => n1371);
   U1813 : AOI22_X1 port map( A1 => n7, A2 => regs(2541), B1 => n40, B2 => 
                           regs(2029), ZN => n1370);
   U1814 : NAND3_X1 port map( A1 => n1372, A2 => n1371, A3 => n1370, ZN => 
                           curr_proc_regs(493));
   U1815 : NAND2_X1 port map( A1 => regs(1006), A2 => n1595, ZN => n1375);
   U1816 : AOI22_X1 port map( A1 => n30, A2 => regs(1518), B1 => n20, B2 => 
                           regs(494), ZN => n1374);
   U1817 : AOI22_X1 port map( A1 => n7, A2 => regs(2542), B1 => n39, B2 => 
                           regs(2030), ZN => n1373);
   U1818 : NAND3_X1 port map( A1 => n1375, A2 => n1374, A3 => n1373, ZN => 
                           curr_proc_regs(494));
   U1819 : NAND2_X1 port map( A1 => regs(1007), A2 => n14, ZN => n1378);
   U1820 : AOI22_X1 port map( A1 => n27, A2 => regs(1519), B1 => n19, B2 => 
                           regs(495), ZN => n1377);
   U1821 : AOI22_X1 port map( A1 => n7, A2 => regs(2543), B1 => n35, B2 => 
                           regs(2031), ZN => n1376);
   U1822 : NAND3_X1 port map( A1 => n1378, A2 => n1377, A3 => n1376, ZN => 
                           curr_proc_regs(495));
   U1823 : NAND2_X1 port map( A1 => regs(1008), A2 => n14, ZN => n1381);
   U1824 : AOI22_X1 port map( A1 => n29, A2 => regs(1520), B1 => n19, B2 => 
                           regs(496), ZN => n1380);
   U1825 : AOI22_X1 port map( A1 => n7, A2 => regs(2544), B1 => n35, B2 => 
                           regs(2032), ZN => n1379);
   U1826 : NAND3_X1 port map( A1 => n1381, A2 => n1380, A3 => n1379, ZN => 
                           curr_proc_regs(496));
   U1827 : NAND2_X1 port map( A1 => regs(1009), A2 => n14, ZN => n1384);
   U1828 : AOI22_X1 port map( A1 => n29, A2 => regs(1521), B1 => n20, B2 => 
                           regs(497), ZN => n1383);
   U1829 : AOI22_X1 port map( A1 => n7, A2 => regs(2545), B1 => n38, B2 => 
                           regs(2033), ZN => n1382);
   U1830 : NAND3_X1 port map( A1 => n1384, A2 => n1383, A3 => n1382, ZN => 
                           curr_proc_regs(497));
   U1831 : NAND2_X1 port map( A1 => regs(1010), A2 => n14, ZN => n1387);
   U1832 : AOI22_X1 port map( A1 => n30, A2 => regs(1522), B1 => n19, B2 => 
                           regs(498), ZN => n1386);
   U1833 : AOI22_X1 port map( A1 => n7, A2 => regs(2546), B1 => n35, B2 => 
                           regs(2034), ZN => n1385);
   U1834 : NAND3_X1 port map( A1 => n1387, A2 => n1386, A3 => n1385, ZN => 
                           curr_proc_regs(498));
   U1835 : NAND2_X1 port map( A1 => regs(1011), A2 => n14, ZN => n1390);
   U1836 : AOI22_X1 port map( A1 => n27, A2 => regs(1523), B1 => n19, B2 => 
                           regs(499), ZN => n1389);
   U1837 : AOI22_X1 port map( A1 => n7, A2 => regs(2547), B1 => n35, B2 => 
                           regs(2035), ZN => n1388);
   U1838 : NAND3_X1 port map( A1 => n1390, A2 => n1389, A3 => n1388, ZN => 
                           curr_proc_regs(499));
   U1839 : NAND2_X1 port map( A1 => regs(561), A2 => n14, ZN => n1393);
   U1840 : AOI22_X1 port map( A1 => n30, A2 => regs(1073), B1 => n19, B2 => 
                           regs(49), ZN => n1392);
   U1841 : AOI22_X1 port map( A1 => n7, A2 => regs(2097), B1 => n35, B2 => 
                           regs(1585), ZN => n1391);
   U1842 : NAND3_X1 port map( A1 => n1393, A2 => n1392, A3 => n1391, ZN => 
                           curr_proc_regs(49));
   U1843 : NAND2_X1 port map( A1 => regs(516), A2 => n1595, ZN => n1396);
   U1844 : AOI22_X1 port map( A1 => n2, A2 => regs(1028), B1 => n26, B2 => 
                           regs(4), ZN => n1395);
   U1845 : AOI22_X1 port map( A1 => n7, A2 => regs(2052), B1 => n35, B2 => 
                           regs(1540), ZN => n1394);
   U1846 : NAND3_X1 port map( A1 => n1396, A2 => n1395, A3 => n1394, ZN => 
                           curr_proc_regs(4));
   U1847 : NAND2_X1 port map( A1 => regs(1012), A2 => n14, ZN => n1399);
   U1848 : AOI22_X1 port map( A1 => n29, A2 => regs(1524), B1 => n19, B2 => 
                           regs(500), ZN => n1398);
   U1849 : AOI22_X1 port map( A1 => n7, A2 => regs(2548), B1 => n35, B2 => 
                           regs(2036), ZN => n1397);
   U1850 : NAND3_X1 port map( A1 => n1399, A2 => n1398, A3 => n1397, ZN => 
                           curr_proc_regs(500));
   U1851 : NAND2_X1 port map( A1 => regs(1013), A2 => n1595, ZN => n1402);
   U1852 : AOI22_X1 port map( A1 => n27, A2 => regs(1525), B1 => n19, B2 => 
                           regs(501), ZN => n1401);
   U1853 : AOI22_X1 port map( A1 => n7, A2 => regs(2549), B1 => n35, B2 => 
                           regs(2037), ZN => n1400);
   U1854 : NAND3_X1 port map( A1 => n1402, A2 => n1401, A3 => n1400, ZN => 
                           curr_proc_regs(501));
   U1855 : NAND2_X1 port map( A1 => regs(1014), A2 => n14, ZN => n1405);
   U1856 : AOI22_X1 port map( A1 => n29, A2 => regs(1526), B1 => n19, B2 => 
                           regs(502), ZN => n1404);
   U1857 : AOI22_X1 port map( A1 => n51, A2 => regs(2550), B1 => n35, B2 => 
                           regs(2038), ZN => n1403);
   U1858 : NAND3_X1 port map( A1 => n1405, A2 => n1404, A3 => n1403, ZN => 
                           curr_proc_regs(502));
   U1859 : NAND2_X1 port map( A1 => regs(1015), A2 => n1595, ZN => n1408);
   U1860 : AOI22_X1 port map( A1 => n30, A2 => regs(1527), B1 => n18, B2 => 
                           regs(503), ZN => n1407);
   U1861 : AOI22_X1 port map( A1 => n51, A2 => regs(2551), B1 => n35, B2 => 
                           regs(2039), ZN => n1406);
   U1862 : NAND3_X1 port map( A1 => n1408, A2 => n1407, A3 => n1406, ZN => 
                           curr_proc_regs(503));
   U1863 : NAND2_X1 port map( A1 => regs(1016), A2 => n14, ZN => n1411);
   U1864 : AOI22_X1 port map( A1 => n29, A2 => regs(1528), B1 => n23, B2 => 
                           regs(504), ZN => n1410);
   U1865 : AOI22_X1 port map( A1 => n51, A2 => regs(2552), B1 => n39, B2 => 
                           regs(2040), ZN => n1409);
   U1866 : NAND3_X1 port map( A1 => n1411, A2 => n1410, A3 => n1409, ZN => 
                           curr_proc_regs(504));
   U1867 : NAND2_X1 port map( A1 => regs(1017), A2 => n1595, ZN => n1414);
   U1868 : AOI22_X1 port map( A1 => n27, A2 => regs(1529), B1 => n19, B2 => 
                           regs(505), ZN => n1413);
   U1869 : AOI22_X1 port map( A1 => n51, A2 => regs(2553), B1 => n35, B2 => 
                           regs(2041), ZN => n1412);
   U1870 : NAND3_X1 port map( A1 => n1414, A2 => n1413, A3 => n1412, ZN => 
                           curr_proc_regs(505));
   U1871 : NAND2_X1 port map( A1 => regs(1018), A2 => n14, ZN => n1417);
   U1872 : AOI22_X1 port map( A1 => n30, A2 => regs(1530), B1 => n19, B2 => 
                           regs(506), ZN => n1416);
   U1873 : AOI22_X1 port map( A1 => n51, A2 => regs(2554), B1 => n35, B2 => 
                           regs(2042), ZN => n1415);
   U1874 : NAND3_X1 port map( A1 => n1417, A2 => n1416, A3 => n1415, ZN => 
                           curr_proc_regs(506));
   U1875 : NAND2_X1 port map( A1 => regs(1019), A2 => n1595, ZN => n1420);
   U1876 : AOI22_X1 port map( A1 => n27, A2 => regs(1531), B1 => n19, B2 => 
                           regs(507), ZN => n1419);
   U1877 : AOI22_X1 port map( A1 => n51, A2 => regs(2555), B1 => n35, B2 => 
                           regs(2043), ZN => n1418);
   U1878 : NAND3_X1 port map( A1 => n1420, A2 => n1419, A3 => n1418, ZN => 
                           curr_proc_regs(507));
   U1879 : NAND2_X1 port map( A1 => regs(1020), A2 => n14, ZN => n1423);
   U1880 : AOI22_X1 port map( A1 => n27, A2 => regs(1532), B1 => n19, B2 => 
                           regs(508), ZN => n1422);
   U1881 : AOI22_X1 port map( A1 => n51, A2 => regs(2556), B1 => n35, B2 => 
                           regs(2044), ZN => n1421);
   U1882 : NAND3_X1 port map( A1 => n1423, A2 => n1422, A3 => n1421, ZN => 
                           curr_proc_regs(508));
   U1883 : NAND2_X1 port map( A1 => regs(1021), A2 => n1595, ZN => n1426);
   U1884 : AOI22_X1 port map( A1 => n27, A2 => regs(1533), B1 => n19, B2 => 
                           regs(509), ZN => n1425);
   U1885 : AOI22_X1 port map( A1 => n51, A2 => regs(2557), B1 => n35, B2 => 
                           regs(2045), ZN => n1424);
   U1886 : NAND3_X1 port map( A1 => n1426, A2 => n1425, A3 => n1424, ZN => 
                           curr_proc_regs(509));
   U1887 : NAND2_X1 port map( A1 => regs(562), A2 => n1595, ZN => n1429);
   U1888 : AOI22_X1 port map( A1 => n27, A2 => regs(1074), B1 => n19, B2 => 
                           regs(50), ZN => n1428);
   U1889 : AOI22_X1 port map( A1 => n51, A2 => regs(2098), B1 => n35, B2 => 
                           regs(1586), ZN => n1427);
   U1890 : NAND3_X1 port map( A1 => n1429, A2 => n1428, A3 => n1427, ZN => 
                           curr_proc_regs(50));
   U1891 : NAND2_X1 port map( A1 => regs(1022), A2 => n13, ZN => n1432);
   U1892 : AOI22_X1 port map( A1 => n27, A2 => regs(1534), B1 => n26, B2 => 
                           regs(510), ZN => n1431);
   U1893 : AOI22_X1 port map( A1 => n51, A2 => regs(2558), B1 => n35, B2 => 
                           regs(2046), ZN => n1430);
   U1894 : NAND3_X1 port map( A1 => n1432, A2 => n1431, A3 => n1430, ZN => 
                           curr_proc_regs(510));
   U1895 : NAND2_X1 port map( A1 => regs(1023), A2 => n3, ZN => n1435);
   U1896 : AOI22_X1 port map( A1 => n27, A2 => regs(1535), B1 => n22, B2 => 
                           regs(511), ZN => n1434);
   U1897 : AOI22_X1 port map( A1 => n51, A2 => regs(2559), B1 => n40, B2 => 
                           regs(2047), ZN => n1433);
   U1898 : NAND3_X1 port map( A1 => n1435, A2 => n1434, A3 => n1433, ZN => 
                           curr_proc_regs(511));
   U1899 : NAND2_X1 port map( A1 => regs(563), A2 => n13, ZN => n1438);
   U1900 : AOI22_X1 port map( A1 => n27, A2 => regs(1075), B1 => n18, B2 => 
                           regs(51), ZN => n1437);
   U1901 : AOI22_X1 port map( A1 => n51, A2 => regs(2099), B1 => n40, B2 => 
                           regs(1587), ZN => n1436);
   U1902 : NAND3_X1 port map( A1 => n1438, A2 => n1437, A3 => n1436, ZN => 
                           curr_proc_regs(51));
   U1903 : NAND2_X1 port map( A1 => regs(564), A2 => n13, ZN => n1441);
   U1904 : AOI22_X1 port map( A1 => n27, A2 => regs(1076), B1 => n22, B2 => 
                           regs(52), ZN => n1440);
   U1905 : AOI22_X1 port map( A1 => n50, A2 => regs(2100), B1 => n35, B2 => 
                           regs(1588), ZN => n1439);
   U1906 : NAND3_X1 port map( A1 => n1441, A2 => n1440, A3 => n1439, ZN => 
                           curr_proc_regs(52));
   U1907 : NAND2_X1 port map( A1 => regs(565), A2 => n3, ZN => n1444);
   U1908 : AOI22_X1 port map( A1 => n27, A2 => regs(1077), B1 => n22, B2 => 
                           regs(53), ZN => n1443);
   U1909 : AOI22_X1 port map( A1 => n50, A2 => regs(2101), B1 => n38, B2 => 
                           regs(1589), ZN => n1442);
   U1910 : NAND3_X1 port map( A1 => n1444, A2 => n1443, A3 => n1442, ZN => 
                           curr_proc_regs(53));
   U1911 : NAND2_X1 port map( A1 => regs(566), A2 => n13, ZN => n1447);
   U1912 : AOI22_X1 port map( A1 => n27, A2 => regs(1078), B1 => n23, B2 => 
                           regs(54), ZN => n1446);
   U1913 : AOI22_X1 port map( A1 => n50, A2 => regs(2102), B1 => n42, B2 => 
                           regs(1590), ZN => n1445);
   U1914 : NAND3_X1 port map( A1 => n1447, A2 => n1446, A3 => n1445, ZN => 
                           curr_proc_regs(54));
   U1915 : NAND2_X1 port map( A1 => regs(567), A2 => n13, ZN => n1450);
   U1916 : AOI22_X1 port map( A1 => n27, A2 => regs(1079), B1 => n26, B2 => 
                           regs(55), ZN => n1449);
   U1917 : AOI22_X1 port map( A1 => n50, A2 => regs(2103), B1 => n42, B2 => 
                           regs(1591), ZN => n1448);
   U1918 : NAND3_X1 port map( A1 => n1450, A2 => n1449, A3 => n1448, ZN => 
                           curr_proc_regs(55));
   U1919 : NAND2_X1 port map( A1 => regs(568), A2 => n3, ZN => n1453);
   U1920 : AOI22_X1 port map( A1 => n27, A2 => regs(1080), B1 => n22, B2 => 
                           regs(56), ZN => n1452);
   U1921 : AOI22_X1 port map( A1 => n50, A2 => regs(2104), B1 => n36, B2 => 
                           regs(1592), ZN => n1451);
   U1922 : NAND3_X1 port map( A1 => n1453, A2 => n1452, A3 => n1451, ZN => 
                           curr_proc_regs(56));
   U1923 : NAND2_X1 port map( A1 => regs(569), A2 => n13, ZN => n1456);
   U1924 : AOI22_X1 port map( A1 => n32, A2 => regs(1081), B1 => n1596, B2 => 
                           regs(57), ZN => n1455);
   U1925 : AOI22_X1 port map( A1 => n50, A2 => regs(2105), B1 => n42, B2 => 
                           regs(1593), ZN => n1454);
   U1926 : NAND3_X1 port map( A1 => n1456, A2 => n1455, A3 => n1454, ZN => 
                           curr_proc_regs(57));
   U1927 : NAND2_X1 port map( A1 => regs(570), A2 => n13, ZN => n1459);
   U1928 : AOI22_X1 port map( A1 => n2, A2 => regs(1082), B1 => n22, B2 => 
                           regs(58), ZN => n1458);
   U1929 : AOI22_X1 port map( A1 => n50, A2 => regs(2106), B1 => n40, B2 => 
                           regs(1594), ZN => n1457);
   U1930 : NAND3_X1 port map( A1 => n1459, A2 => n1458, A3 => n1457, ZN => 
                           curr_proc_regs(58));
   U1931 : NAND2_X1 port map( A1 => regs(571), A2 => n3, ZN => n1462);
   U1932 : AOI22_X1 port map( A1 => n29, A2 => regs(1083), B1 => n22, B2 => 
                           regs(59), ZN => n1461);
   U1933 : AOI22_X1 port map( A1 => n50, A2 => regs(2107), B1 => n35, B2 => 
                           regs(1595), ZN => n1460);
   U1934 : NAND3_X1 port map( A1 => n1462, A2 => n1461, A3 => n1460, ZN => 
                           curr_proc_regs(59));
   U1935 : NAND2_X1 port map( A1 => regs(517), A2 => n13, ZN => n1465);
   U1936 : AOI22_X1 port map( A1 => n2, A2 => regs(1029), B1 => n23, B2 => 
                           regs(5), ZN => n1464);
   U1937 : AOI22_X1 port map( A1 => n50, A2 => regs(2053), B1 => n39, B2 => 
                           regs(1541), ZN => n1463);
   U1938 : NAND3_X1 port map( A1 => n1465, A2 => n1464, A3 => n1463, ZN => 
                           curr_proc_regs(5));
   U1939 : NAND2_X1 port map( A1 => regs(572), A2 => n13, ZN => n1468);
   U1940 : AOI22_X1 port map( A1 => n29, A2 => regs(1084), B1 => n21, B2 => 
                           regs(60), ZN => n1467);
   U1941 : AOI22_X1 port map( A1 => n50, A2 => regs(2108), B1 => n36, B2 => 
                           regs(1596), ZN => n1466);
   U1942 : NAND3_X1 port map( A1 => n1468, A2 => n1467, A3 => n1466, ZN => 
                           curr_proc_regs(60));
   U1943 : NAND2_X1 port map( A1 => regs(573), A2 => n13, ZN => n1471);
   U1944 : AOI22_X1 port map( A1 => n29, A2 => regs(1085), B1 => n19, B2 => 
                           regs(61), ZN => n1470);
   U1945 : AOI22_X1 port map( A1 => n50, A2 => regs(2109), B1 => n38, B2 => 
                           regs(1597), ZN => n1469);
   U1946 : NAND3_X1 port map( A1 => n1471, A2 => n1470, A3 => n1469, ZN => 
                           curr_proc_regs(61));
   U1947 : NAND2_X1 port map( A1 => regs(574), A2 => n13, ZN => n1474);
   U1948 : AOI22_X1 port map( A1 => n32, A2 => regs(1086), B1 => n21, B2 => 
                           regs(62), ZN => n1473);
   U1949 : AOI22_X1 port map( A1 => n50, A2 => regs(2110), B1 => n39, B2 => 
                           regs(1598), ZN => n1472);
   U1950 : NAND3_X1 port map( A1 => n1474, A2 => n1473, A3 => n1472, ZN => 
                           curr_proc_regs(62));
   U1951 : NAND2_X1 port map( A1 => regs(575), A2 => n13, ZN => n1477);
   U1952 : AOI22_X1 port map( A1 => n30, A2 => regs(1087), B1 => n20, B2 => 
                           regs(63), ZN => n1476);
   U1953 : AOI22_X1 port map( A1 => n49, A2 => regs(2111), B1 => n42, B2 => 
                           regs(1599), ZN => n1475);
   U1954 : NAND3_X1 port map( A1 => n1477, A2 => n1476, A3 => n1475, ZN => 
                           curr_proc_regs(63));
   U1955 : NAND2_X1 port map( A1 => regs(576), A2 => n13, ZN => n1480);
   U1956 : AOI22_X1 port map( A1 => n31, A2 => regs(1088), B1 => n17, B2 => 
                           regs(64), ZN => n1479);
   U1957 : AOI22_X1 port map( A1 => n49, A2 => regs(2112), B1 => n42, B2 => 
                           regs(1600), ZN => n1478);
   U1958 : NAND3_X1 port map( A1 => n1480, A2 => n1479, A3 => n1478, ZN => 
                           curr_proc_regs(64));
   U1959 : NAND2_X1 port map( A1 => regs(577), A2 => n13, ZN => n1483);
   U1960 : AOI22_X1 port map( A1 => n31, A2 => regs(1089), B1 => n1596, B2 => 
                           regs(65), ZN => n1482);
   U1961 : AOI22_X1 port map( A1 => n49, A2 => regs(2113), B1 => n36, B2 => 
                           regs(1601), ZN => n1481);
   U1962 : NAND3_X1 port map( A1 => n1483, A2 => n1482, A3 => n1481, ZN => 
                           curr_proc_regs(65));
   U1963 : NAND2_X1 port map( A1 => regs(578), A2 => n13, ZN => n1486);
   U1964 : AOI22_X1 port map( A1 => n2, A2 => regs(1090), B1 => n20, B2 => 
                           regs(66), ZN => n1485);
   U1965 : AOI22_X1 port map( A1 => n49, A2 => regs(2114), B1 => n35, B2 => 
                           regs(1602), ZN => n1484);
   U1966 : NAND3_X1 port map( A1 => n1486, A2 => n1485, A3 => n1484, ZN => 
                           curr_proc_regs(66));
   U1967 : NAND2_X1 port map( A1 => regs(579), A2 => n13, ZN => n1489);
   U1968 : AOI22_X1 port map( A1 => n30, A2 => regs(1091), B1 => n22, B2 => 
                           regs(67), ZN => n1488);
   U1969 : AOI22_X1 port map( A1 => n49, A2 => regs(2115), B1 => n36, B2 => 
                           regs(1603), ZN => n1487);
   U1970 : NAND3_X1 port map( A1 => n1489, A2 => n1488, A3 => n1487, ZN => 
                           curr_proc_regs(67));
   U1971 : NAND2_X1 port map( A1 => regs(580), A2 => n13, ZN => n1492);
   U1972 : AOI22_X1 port map( A1 => n29, A2 => regs(1092), B1 => n21, B2 => 
                           regs(68), ZN => n1491);
   U1973 : AOI22_X1 port map( A1 => n49, A2 => regs(2116), B1 => n36, B2 => 
                           regs(1604), ZN => n1490);
   U1974 : NAND3_X1 port map( A1 => n1492, A2 => n1491, A3 => n1490, ZN => 
                           curr_proc_regs(68));
   U1975 : NAND2_X1 port map( A1 => regs(581), A2 => n13, ZN => n1495);
   U1976 : AOI22_X1 port map( A1 => n29, A2 => regs(1093), B1 => n22, B2 => 
                           regs(69), ZN => n1494);
   U1977 : AOI22_X1 port map( A1 => n49, A2 => regs(2117), B1 => n40, B2 => 
                           regs(1605), ZN => n1493);
   U1978 : NAND3_X1 port map( A1 => n1495, A2 => n1494, A3 => n1493, ZN => 
                           curr_proc_regs(69));
   U1979 : NAND2_X1 port map( A1 => regs(518), A2 => n13, ZN => n1498);
   U1980 : AOI22_X1 port map( A1 => n29, A2 => regs(1030), B1 => n19, B2 => 
                           regs(6), ZN => n1497);
   U1981 : AOI22_X1 port map( A1 => n49, A2 => regs(2054), B1 => n38, B2 => 
                           regs(1542), ZN => n1496);
   U1982 : NAND3_X1 port map( A1 => n1498, A2 => n1497, A3 => n1496, ZN => 
                           curr_proc_regs(6));
   U1983 : NAND2_X1 port map( A1 => regs(582), A2 => n13, ZN => n1501);
   U1984 : AOI22_X1 port map( A1 => n29, A2 => regs(1094), B1 => n22, B2 => 
                           regs(70), ZN => n1500);
   U1985 : AOI22_X1 port map( A1 => n49, A2 => regs(2118), B1 => n36, B2 => 
                           regs(1606), ZN => n1499);
   U1986 : NAND3_X1 port map( A1 => n1501, A2 => n1500, A3 => n1499, ZN => 
                           curr_proc_regs(70));
   U1987 : NAND2_X1 port map( A1 => regs(583), A2 => n13, ZN => n1504);
   U1988 : AOI22_X1 port map( A1 => n29, A2 => regs(1095), B1 => n22, B2 => 
                           regs(71), ZN => n1503);
   U1989 : AOI22_X1 port map( A1 => n49, A2 => regs(2119), B1 => n40, B2 => 
                           regs(1607), ZN => n1502);
   U1990 : NAND3_X1 port map( A1 => n1504, A2 => n1503, A3 => n1502, ZN => 
                           curr_proc_regs(71));
   U1991 : NAND2_X1 port map( A1 => regs(584), A2 => n13, ZN => n1507);
   U1992 : AOI22_X1 port map( A1 => n29, A2 => regs(1096), B1 => n20, B2 => 
                           regs(72), ZN => n1506);
   U1993 : AOI22_X1 port map( A1 => n49, A2 => regs(2120), B1 => n42, B2 => 
                           regs(1608), ZN => n1505);
   U1994 : NAND3_X1 port map( A1 => n1507, A2 => n1506, A3 => n1505, ZN => 
                           curr_proc_regs(72));
   U1995 : NAND2_X1 port map( A1 => regs(585), A2 => n3, ZN => n1510);
   U1996 : AOI22_X1 port map( A1 => n29, A2 => regs(1097), B1 => n22, B2 => 
                           regs(73), ZN => n1509);
   U1997 : AOI22_X1 port map( A1 => n49, A2 => regs(2121), B1 => n35, B2 => 
                           regs(1609), ZN => n1508);
   U1998 : NAND3_X1 port map( A1 => n1510, A2 => n1509, A3 => n1508, ZN => 
                           curr_proc_regs(73));
   U1999 : NAND2_X1 port map( A1 => regs(586), A2 => n13, ZN => n1513);
   U2000 : AOI22_X1 port map( A1 => n29, A2 => regs(1098), B1 => n26, B2 => 
                           regs(74), ZN => n1512);
   U2001 : AOI22_X1 port map( A1 => win(4), A2 => regs(2122), B1 => n39, B2 => 
                           regs(1610), ZN => n1511);
   U2002 : NAND3_X1 port map( A1 => n1513, A2 => n1512, A3 => n1511, ZN => 
                           curr_proc_regs(74));
   U2003 : NAND2_X1 port map( A1 => regs(587), A2 => n13, ZN => n1516);
   U2004 : AOI22_X1 port map( A1 => n29, A2 => regs(1099), B1 => n22, B2 => 
                           regs(75), ZN => n1515);
   U2005 : AOI22_X1 port map( A1 => win(4), A2 => regs(2123), B1 => n38, B2 => 
                           regs(1611), ZN => n1514);
   U2006 : NAND3_X1 port map( A1 => n1516, A2 => n1515, A3 => n1514, ZN => 
                           curr_proc_regs(75));
   U2007 : NAND2_X1 port map( A1 => regs(588), A2 => n13, ZN => n1519);
   U2008 : AOI22_X1 port map( A1 => n29, A2 => regs(1100), B1 => n22, B2 => 
                           regs(76), ZN => n1518);
   U2009 : AOI22_X1 port map( A1 => win(4), A2 => regs(2124), B1 => n36, B2 => 
                           regs(1612), ZN => n1517);
   U2010 : NAND3_X1 port map( A1 => n1519, A2 => n1518, A3 => n1517, ZN => 
                           curr_proc_regs(76));
   U2011 : NAND2_X1 port map( A1 => regs(589), A2 => n3, ZN => n1522);
   U2012 : AOI22_X1 port map( A1 => n29, A2 => regs(1101), B1 => n19, B2 => 
                           regs(77), ZN => n1521);
   U2013 : AOI22_X1 port map( A1 => win(4), A2 => regs(2125), B1 => n38, B2 => 
                           regs(1613), ZN => n1520);
   U2014 : NAND3_X1 port map( A1 => n1522, A2 => n1521, A3 => n1520, ZN => 
                           curr_proc_regs(77));
   U2015 : NAND2_X1 port map( A1 => regs(590), A2 => n13, ZN => n1525);
   U2016 : AOI22_X1 port map( A1 => n29, A2 => regs(1102), B1 => n21, B2 => 
                           regs(78), ZN => n1524);
   U2017 : AOI22_X1 port map( A1 => n53, A2 => regs(2126), B1 => n36, B2 => 
                           regs(1614), ZN => n1523);
   U2018 : NAND3_X1 port map( A1 => n1525, A2 => n1524, A3 => n1523, ZN => 
                           curr_proc_regs(78));
   U2019 : NAND2_X1 port map( A1 => regs(591), A2 => n3, ZN => n1528);
   U2020 : AOI22_X1 port map( A1 => n28, A2 => regs(1103), B1 => n22, B2 => 
                           regs(79), ZN => n1527);
   U2021 : AOI22_X1 port map( A1 => n55, A2 => regs(2127), B1 => n40, B2 => 
                           regs(1615), ZN => n1526);
   U2022 : NAND3_X1 port map( A1 => n1528, A2 => n1527, A3 => n1526, ZN => 
                           curr_proc_regs(79));
   U2023 : NAND2_X1 port map( A1 => regs(519), A2 => n13, ZN => n1531);
   U2024 : AOI22_X1 port map( A1 => n28, A2 => regs(1031), B1 => n22, B2 => 
                           regs(7), ZN => n1530);
   U2025 : AOI22_X1 port map( A1 => n52, A2 => regs(2055), B1 => n35, B2 => 
                           regs(1543), ZN => n1529);
   U2026 : NAND3_X1 port map( A1 => n1531, A2 => n1530, A3 => n1529, ZN => 
                           curr_proc_regs(7));
   U2027 : NAND2_X1 port map( A1 => regs(592), A2 => n13, ZN => n1534);
   U2028 : AOI22_X1 port map( A1 => n28, A2 => regs(1104), B1 => n22, B2 => 
                           regs(80), ZN => n1533);
   U2029 : AOI22_X1 port map( A1 => win(4), A2 => regs(2128), B1 => n38, B2 => 
                           regs(1616), ZN => n1532);
   U2030 : NAND3_X1 port map( A1 => n1534, A2 => n1533, A3 => n1532, ZN => 
                           curr_proc_regs(80));
   U2031 : NAND2_X1 port map( A1 => regs(593), A2 => n13, ZN => n1537);
   U2032 : AOI22_X1 port map( A1 => n28, A2 => regs(1105), B1 => n22, B2 => 
                           regs(81), ZN => n1536);
   U2033 : AOI22_X1 port map( A1 => n56, A2 => regs(2129), B1 => n36, B2 => 
                           regs(1617), ZN => n1535);
   U2034 : NAND3_X1 port map( A1 => n1537, A2 => n1536, A3 => n1535, ZN => 
                           curr_proc_regs(81));
   U2035 : NAND2_X1 port map( A1 => regs(594), A2 => n3, ZN => n1540);
   U2036 : AOI22_X1 port map( A1 => n28, A2 => regs(1106), B1 => n26, B2 => 
                           regs(82), ZN => n1539);
   U2037 : AOI22_X1 port map( A1 => n45, A2 => regs(2130), B1 => n36, B2 => 
                           regs(1618), ZN => n1538);
   U2038 : NAND3_X1 port map( A1 => n1540, A2 => n1539, A3 => n1538, ZN => 
                           curr_proc_regs(82));
   U2039 : NAND2_X1 port map( A1 => regs(595), A2 => n13, ZN => n1543);
   U2040 : AOI22_X1 port map( A1 => n28, A2 => regs(1107), B1 => n22, B2 => 
                           regs(83), ZN => n1542);
   U2041 : AOI22_X1 port map( A1 => n49, A2 => regs(2131), B1 => n42, B2 => 
                           regs(1619), ZN => n1541);
   U2042 : NAND3_X1 port map( A1 => n1543, A2 => n1542, A3 => n1541, ZN => 
                           curr_proc_regs(83));
   U2043 : NAND2_X1 port map( A1 => regs(596), A2 => n13, ZN => n1546);
   U2044 : AOI22_X1 port map( A1 => n28, A2 => regs(1108), B1 => n19, B2 => 
                           regs(84), ZN => n1545);
   U2045 : AOI22_X1 port map( A1 => n43, A2 => regs(2132), B1 => n35, B2 => 
                           regs(1620), ZN => n1544);
   U2046 : NAND3_X1 port map( A1 => n1546, A2 => n1545, A3 => n1544, ZN => 
                           curr_proc_regs(84));
   U2047 : NAND2_X1 port map( A1 => regs(597), A2 => n13, ZN => n1549);
   U2048 : AOI22_X1 port map( A1 => n28, A2 => regs(1109), B1 => n22, B2 => 
                           regs(85), ZN => n1548);
   U2049 : AOI22_X1 port map( A1 => n48, A2 => regs(2133), B1 => n38, B2 => 
                           regs(1621), ZN => n1547);
   U2050 : NAND3_X1 port map( A1 => n1549, A2 => n1548, A3 => n1547, ZN => 
                           curr_proc_regs(85));
   U2051 : NAND2_X1 port map( A1 => regs(598), A2 => n13, ZN => n1552);
   U2052 : AOI22_X1 port map( A1 => n28, A2 => regs(1110), B1 => n22, B2 => 
                           regs(86), ZN => n1551);
   U2053 : AOI22_X1 port map( A1 => n48, A2 => regs(2134), B1 => n36, B2 => 
                           regs(1622), ZN => n1550);
   U2054 : NAND3_X1 port map( A1 => n1552, A2 => n1551, A3 => n1550, ZN => 
                           curr_proc_regs(86));
   U2055 : NAND2_X1 port map( A1 => regs(599), A2 => n3, ZN => n1555);
   U2056 : AOI22_X1 port map( A1 => n28, A2 => regs(1111), B1 => n18, B2 => 
                           regs(87), ZN => n1554);
   U2057 : AOI22_X1 port map( A1 => n48, A2 => regs(2135), B1 => n35, B2 => 
                           regs(1623), ZN => n1553);
   U2058 : NAND3_X1 port map( A1 => n1555, A2 => n1554, A3 => n1553, ZN => 
                           curr_proc_regs(87));
   U2059 : NAND2_X1 port map( A1 => regs(600), A2 => n13, ZN => n1558);
   U2060 : AOI22_X1 port map( A1 => n28, A2 => regs(1112), B1 => n22, B2 => 
                           regs(88), ZN => n1557);
   U2061 : AOI22_X1 port map( A1 => n48, A2 => regs(2136), B1 => n40, B2 => 
                           regs(1624), ZN => n1556);
   U2062 : NAND3_X1 port map( A1 => n1558, A2 => n1557, A3 => n1556, ZN => 
                           curr_proc_regs(88));
   U2063 : NAND2_X1 port map( A1 => regs(601), A2 => n13, ZN => n1561);
   U2064 : AOI22_X1 port map( A1 => n28, A2 => regs(1113), B1 => n1596, B2 => 
                           regs(89), ZN => n1560);
   U2065 : AOI22_X1 port map( A1 => n48, A2 => regs(2137), B1 => n42, B2 => 
                           regs(1625), ZN => n1559);
   U2066 : NAND3_X1 port map( A1 => n1561, A2 => n1560, A3 => n1559, ZN => 
                           curr_proc_regs(89));
   U2067 : NAND2_X1 port map( A1 => regs(520), A2 => n3, ZN => n1564);
   U2068 : AOI22_X1 port map( A1 => n30, A2 => regs(1032), B1 => n22, B2 => 
                           regs(8), ZN => n1563);
   U2069 : AOI22_X1 port map( A1 => n48, A2 => regs(2056), B1 => n35, B2 => 
                           regs(1544), ZN => n1562);
   U2070 : NAND3_X1 port map( A1 => n1564, A2 => n1563, A3 => n1562, ZN => 
                           curr_proc_regs(8));
   U2071 : NAND2_X1 port map( A1 => regs(602), A2 => n13, ZN => n1567);
   U2072 : AOI22_X1 port map( A1 => n30, A2 => regs(1114), B1 => n17, B2 => 
                           regs(90), ZN => n1566);
   U2073 : AOI22_X1 port map( A1 => n48, A2 => regs(2138), B1 => n42, B2 => 
                           regs(1626), ZN => n1565);
   U2074 : NAND3_X1 port map( A1 => n1567, A2 => n1566, A3 => n1565, ZN => 
                           curr_proc_regs(90));
   U2075 : NAND2_X1 port map( A1 => regs(603), A2 => n3, ZN => n1570);
   U2076 : AOI22_X1 port map( A1 => n30, A2 => regs(1115), B1 => n22, B2 => 
                           regs(91), ZN => n1569);
   U2077 : AOI22_X1 port map( A1 => n48, A2 => regs(2139), B1 => n38, B2 => 
                           regs(1627), ZN => n1568);
   U2078 : NAND3_X1 port map( A1 => n1570, A2 => n1569, A3 => n1568, ZN => 
                           curr_proc_regs(91));
   U2079 : NAND2_X1 port map( A1 => regs(604), A2 => n13, ZN => n1573);
   U2080 : AOI22_X1 port map( A1 => n30, A2 => regs(1116), B1 => n22, B2 => 
                           regs(92), ZN => n1572);
   U2081 : AOI22_X1 port map( A1 => n48, A2 => regs(2140), B1 => n36, B2 => 
                           regs(1628), ZN => n1571);
   U2082 : NAND3_X1 port map( A1 => n1573, A2 => n1572, A3 => n1571, ZN => 
                           curr_proc_regs(92));
   U2083 : NAND2_X1 port map( A1 => regs(605), A2 => n13, ZN => n1576);
   U2084 : AOI22_X1 port map( A1 => n30, A2 => regs(1117), B1 => n26, B2 => 
                           regs(93), ZN => n1575);
   U2085 : AOI22_X1 port map( A1 => n48, A2 => regs(2141), B1 => n36, B2 => 
                           regs(1629), ZN => n1574);
   U2086 : NAND3_X1 port map( A1 => n1576, A2 => n1575, A3 => n1574, ZN => 
                           curr_proc_regs(93));
   U2087 : NAND2_X1 port map( A1 => regs(606), A2 => n3, ZN => n1579);
   U2088 : AOI22_X1 port map( A1 => n30, A2 => regs(1118), B1 => n22, B2 => 
                           regs(94), ZN => n1578);
   U2089 : AOI22_X1 port map( A1 => n48, A2 => regs(2142), B1 => n42, B2 => 
                           regs(1630), ZN => n1577);
   U2090 : NAND3_X1 port map( A1 => n1579, A2 => n1578, A3 => n1577, ZN => 
                           curr_proc_regs(94));
   U2091 : NAND2_X1 port map( A1 => regs(607), A2 => n3, ZN => n1582);
   U2092 : AOI22_X1 port map( A1 => n30, A2 => regs(1119), B1 => n18, B2 => 
                           regs(95), ZN => n1581);
   U2093 : AOI22_X1 port map( A1 => n48, A2 => regs(2143), B1 => n42, B2 => 
                           regs(1631), ZN => n1580);
   U2094 : NAND3_X1 port map( A1 => n1582, A2 => n1581, A3 => n1580, ZN => 
                           curr_proc_regs(95));
   U2095 : NAND2_X1 port map( A1 => regs(608), A2 => n13, ZN => n1585);
   U2096 : AOI22_X1 port map( A1 => n30, A2 => regs(1120), B1 => n22, B2 => 
                           regs(96), ZN => n1584);
   U2097 : AOI22_X1 port map( A1 => n5, A2 => regs(2144), B1 => n42, B2 => 
                           regs(1632), ZN => n1583);
   U2098 : NAND3_X1 port map( A1 => n1585, A2 => n1584, A3 => n1583, ZN => 
                           curr_proc_regs(96));
   U2099 : NAND2_X1 port map( A1 => regs(609), A2 => n3, ZN => n1588);
   U2100 : AOI22_X1 port map( A1 => n30, A2 => regs(1121), B1 => n23, B2 => 
                           regs(97), ZN => n1587);
   U2101 : AOI22_X1 port map( A1 => n5, A2 => regs(2145), B1 => n42, B2 => 
                           regs(1633), ZN => n1586);
   U2102 : NAND3_X1 port map( A1 => n1588, A2 => n1587, A3 => n1586, ZN => 
                           curr_proc_regs(97));
   U2103 : NAND2_X1 port map( A1 => regs(610), A2 => n13, ZN => n1591);
   U2104 : AOI22_X1 port map( A1 => n30, A2 => regs(1122), B1 => n17, B2 => 
                           regs(98), ZN => n1590);
   U2105 : AOI22_X1 port map( A1 => n7, A2 => regs(2146), B1 => n42, B2 => 
                           regs(1634), ZN => n1589);
   U2106 : NAND3_X1 port map( A1 => n1591, A2 => n1590, A3 => n1589, ZN => 
                           curr_proc_regs(98));
   U2107 : NAND2_X1 port map( A1 => regs(611), A2 => n3, ZN => n1594);
   U2108 : AOI22_X1 port map( A1 => n30, A2 => regs(1123), B1 => n26, B2 => 
                           regs(99), ZN => n1593);
   U2109 : AOI22_X1 port map( A1 => n56, A2 => regs(2147), B1 => n39, B2 => 
                           regs(1635), ZN => n1592);
   U2110 : NAND3_X1 port map( A1 => n1594, A2 => n1593, A3 => n1592, ZN => 
                           curr_proc_regs(99));
   U2111 : NAND2_X1 port map( A1 => regs(521), A2 => n13, ZN => n1601);
   U2112 : AOI22_X1 port map( A1 => n30, A2 => regs(1033), B1 => n26, B2 => 
                           regs(9), ZN => n1600);
   U2113 : AOI22_X1 port map( A1 => n6, A2 => regs(2057), B1 => n38, B2 => 
                           regs(1545), ZN => n1599);
   U2114 : NAND3_X1 port map( A1 => n1601, A2 => n1600, A3 => n1599, ZN => 
                           curr_proc_regs(9));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32.all;

entity hazard_table_N_REGS_LOG5 is

   port( CLK, RST, WR1, WR2 : in std_logic;  ADD_WR1, ADD_WR2, ADD_CHECK1, 
         ADD_CHECK2 : in std_logic_vector (4 downto 0);  BUSY, BUSY_WINDOW : 
         out std_logic);

end hazard_table_N_REGS_LOG5;

architecture SYN_behavioural of hazard_table_N_REGS_LOG5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Table_0_2_port, Table_0_1_port, Table_0_0_port, Table_1_2_port, 
      Table_1_1_port, Table_1_0_port, Table_2_2_port, Table_2_1_port, 
      Table_2_0_port, Table_3_2_port, Table_3_1_port, Table_3_0_port, 
      Table_4_2_port, Table_4_1_port, Table_4_0_port, Table_5_2_port, 
      Table_5_1_port, Table_5_0_port, Table_6_2_port, Table_6_1_port, 
      Table_6_0_port, Table_7_2_port, Table_7_1_port, Table_7_0_port, 
      Table_8_2_port, Table_8_1_port, Table_9_2_port, Table_9_1_port, 
      Table_9_0_port, Table_10_2_port, Table_10_1_port, Table_11_2_port, 
      Table_11_1_port, Table_11_0_port, Table_12_2_port, Table_13_2_port, 
      Table_13_1_port, Table_13_0_port, Table_14_2_port, Table_14_1_port, 
      Table_14_0_port, Table_15_2_port, Table_15_1_port, Table_15_0_port, 
      Table_16_2_port, Table_16_1_port, Table_16_0_port, Table_17_2_port, 
      Table_17_1_port, Table_18_2_port, Table_18_1_port, Table_18_0_port, 
      Table_19_2_port, Table_19_1_port, Table_19_0_port, Table_20_2_port, 
      Table_20_1_port, Table_21_2_port, Table_21_1_port, Table_22_2_port, 
      Table_22_1_port, Table_22_0_port, Table_23_2_port, Table_23_1_port, 
      Table_23_0_port, Table_24_2_port, Table_24_1_port, Table_24_0_port, 
      Table_25_2_port, Table_25_1_port, Table_25_0_port, Table_26_2_port, 
      Table_26_1_port, Table_26_0_port, Table_27_2_port, Table_27_1_port, 
      Table_27_0_port, Table_28_2_port, Table_28_1_port, Table_28_0_port, 
      Table_29_2_port, Table_29_1_port, Table_29_0_port, Table_30_2_port, 
      Table_30_1_port, Table_30_0_port, Table_31_2_port, Table_31_1_port, 
      Table_31_0_port, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
      n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, 
      n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, 
      n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, 
      n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, 
      n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, 
      n795, n796, n797, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, 
      n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, 
      n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, 
      n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, 
      n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, 
      n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, 
      n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, 
      n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, 
      n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, 
      n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, 
      n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, 
      n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, 
      n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, 
      n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, 
      n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, 
      n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, 
      n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, 
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, 
      n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, 
      n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, 
      n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, 
      n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, 
      n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, 
      n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, 
      n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, 
      n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, 
      n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, 
      n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, 
      n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, 
      n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, 
      n821, n822, n823, n824, n825, n826, n827, n828, n829, n830 : std_logic;

begin
   
   Table_reg_17_0_inst : DFF_X1 port map( D => n755, CK => CLK, Q => n11, QN =>
                           n60);
   Table_reg_21_0_inst : DFF_X1 port map( D => n767, CK => CLK, Q => n13, QN =>
                           n84);
   Table_reg_14_0_inst : DFF_X1 port map( D => n746, CK => CLK, Q => 
                           Table_14_0_port, QN => n606);
   Table_reg_14_1_inst : DFF_X1 port map( D => n745, CK => CLK, Q => 
                           Table_14_1_port, QN => n608);
   Table_reg_14_2_inst : DFF_X1 port map( D => n744, CK => CLK, Q => 
                           Table_14_2_port, QN => n613);
   Table_reg_8_2_inst : DFF_X1 port map( D => n726, CK => CLK, Q => 
                           Table_8_2_port, QN => n659);
   Table_reg_4_1_inst : DFF_X1 port map( D => n715, CK => CLK, Q => 
                           Table_4_1_port, QN => n45);
   Table_reg_2_1_inst : DFF_X1 port map( D => n709, CK => CLK, Q => 
                           Table_2_1_port, QN => n54);
   Table_reg_1_1_inst : DFF_X1 port map( D => n706, CK => CLK, Q => 
                           Table_1_1_port, QN => n57);
   Table_reg_6_1_inst : DFF_X1 port map( D => n721, CK => CLK, Q => 
                           Table_6_1_port, QN => n42);
   Table_reg_16_0_inst : DFF_X1 port map( D => n752, CK => CLK, Q => 
                           Table_16_0_port, QN => n31);
   Table_reg_30_0_inst : DFF_X1 port map( D => n794, CK => CLK, Q => 
                           Table_30_0_port, QN => n55);
   Table_reg_28_0_inst : DFF_X1 port map( D => n788, CK => CLK, Q => 
                           Table_28_0_port, QN => n248);
   Table_reg_27_0_inst : DFF_X1 port map( D => n785, CK => CLK, Q => 
                           Table_27_0_port, QN => n82);
   Table_reg_26_0_inst : DFF_X1 port map( D => n782, CK => CLK, Q => 
                           Table_26_0_port, QN => n108);
   Table_reg_25_0_inst : DFF_X1 port map( D => n779, CK => CLK, Q => 
                           Table_25_0_port, QN => n59);
   Table_reg_24_0_inst : DFF_X1 port map( D => n776, CK => CLK, Q => 
                           Table_24_0_port, QN => n85);
   Table_reg_19_0_inst : DFF_X1 port map( D => n761, CK => CLK, Q => 
                           Table_19_0_port, QN => n41);
   Table_reg_18_0_inst : DFF_X1 port map( D => n758, CK => CLK, Q => 
                           Table_18_0_port, QN => n572);
   Table_reg_15_0_inst : DFF_X1 port map( D => n749, CK => CLK, Q => 
                           Table_15_0_port, QN => n101);
   Table_reg_13_0_inst : DFF_X1 port map( D => n743, CK => CLK, Q => 
                           Table_13_0_port, QN => n83);
   Table_reg_12_0_inst : DFF_X1 port map( D => n740, CK => CLK, Q => n39, QN =>
                           n123);
   Table_reg_11_0_inst : DFF_X1 port map( D => n737, CK => CLK, Q => 
                           Table_11_0_port, QN => n19);
   Table_reg_10_0_inst : DFF_X1 port map( D => n734, CK => CLK, Q => n37, QN =>
                           n17);
   Table_reg_9_0_inst : DFF_X1 port map( D => n731, CK => CLK, Q => 
                           Table_9_0_port, QN => n80);
   Table_reg_8_0_inst : DFF_X1 port map( D => n728, CK => CLK, Q => n4, QN => 
                           n105);
   Table_reg_1_0_inst : DFF_X1 port map( D => n707, CK => CLK, Q => 
                           Table_1_0_port, QN => n62);
   Table_reg_29_0_inst : DFF_X1 port map( D => n791, CK => CLK, Q => 
                           Table_29_0_port, QN => n120);
   Table_reg_23_0_inst : DFF_X1 port map( D => n773, CK => CLK, Q => 
                           Table_23_0_port, QN => n116);
   Table_reg_22_0_inst : DFF_X1 port map( D => n770, CK => CLK, Q => 
                           Table_22_0_port, QN => n100);
   Table_reg_20_0_inst : DFF_X1 port map( D => n764, CK => CLK, Q => n38, QN =>
                           n122);
   Table_reg_7_0_inst : DFF_X1 port map( D => n725, CK => CLK, Q => 
                           Table_7_0_port, QN => n27);
   Table_reg_6_0_inst : DFF_X1 port map( D => n722, CK => CLK, Q => 
                           Table_6_0_port, QN => n43);
   Table_reg_5_0_inst : DFF_X1 port map( D => n719, CK => CLK, Q => 
                           Table_5_0_port, QN => n61);
   Table_reg_4_0_inst : DFF_X1 port map( D => n716, CK => CLK, Q => 
                           Table_4_0_port, QN => n47);
   Table_reg_3_0_inst : DFF_X1 port map( D => n713, CK => CLK, Q => 
                           Table_3_0_port, QN => n28);
   Table_reg_2_0_inst : DFF_X1 port map( D => n710, CK => CLK, Q => 
                           Table_2_0_port, QN => n52);
   Table_reg_0_0_inst : DFF_X1 port map( D => n704, CK => CLK, Q => 
                           Table_0_0_port, QN => n29);
   Table_reg_31_0_inst : DFF_X1 port map( D => n797, CK => CLK, Q => 
                           Table_31_0_port, QN => n360);
   Table_reg_29_2_inst : DFF_X1 port map( D => n789, CK => CLK, Q => 
                           Table_29_2_port, QN => n487);
   Table_reg_23_2_inst : DFF_X1 port map( D => n771, CK => CLK, Q => 
                           Table_23_2_port, QN => n539);
   Table_reg_21_2_inst : DFF_X1 port map( D => n765, CK => CLK, Q => 
                           Table_21_2_port, QN => n87);
   Table_reg_20_2_inst : DFF_X1 port map( D => n762, CK => CLK, Q => 
                           Table_20_2_port, QN => n111);
   Table_reg_7_2_inst : DFF_X1 port map( D => n723, CK => CLK, Q => 
                           Table_7_2_port, QN => n24);
   Table_reg_6_2_inst : DFF_X1 port map( D => n720, CK => CLK, Q => 
                           Table_6_2_port, QN => n44);
   Table_reg_5_2_inst : DFF_X1 port map( D => n717, CK => CLK, Q => 
                           Table_5_2_port, QN => n64);
   Table_reg_4_2_inst : DFF_X1 port map( D => n714, CK => CLK, Q => 
                           Table_4_2_port, QN => n48);
   Table_reg_3_2_inst : DFF_X1 port map( D => n711, CK => CLK, Q => 
                           Table_3_2_port, QN => n25);
   Table_reg_1_2_inst : DFF_X1 port map( D => n705, CK => CLK, Q => 
                           Table_1_2_port, QN => n65);
   Table_reg_0_2_inst : DFF_X1 port map( D => n702, CK => CLK, Q => 
                           Table_0_2_port, QN => n36);
   Table_reg_16_1_inst : DFF_X1 port map( D => n751, CK => CLK, Q => 
                           Table_16_1_port, QN => n51);
   Table_reg_31_1_inst : DFF_X1 port map( D => n796, CK => CLK, Q => 
                           Table_31_1_port, QN => n412);
   Table_reg_30_1_inst : DFF_X1 port map( D => n793, CK => CLK, Q => 
                           Table_30_1_port, QN => n58);
   Table_reg_29_1_inst : DFF_X1 port map( D => n790, CK => CLK, Q => 
                           Table_29_1_port, QN => n93);
   Table_reg_28_1_inst : DFF_X1 port map( D => n787, CK => CLK, Q => 
                           Table_28_1_port, QN => n94);
   Table_reg_27_1_inst : DFF_X1 port map( D => n784, CK => CLK, Q => 
                           Table_27_1_port, QN => n90);
   Table_reg_26_1_inst : DFF_X1 port map( D => n781, CK => CLK, Q => 
                           Table_26_1_port, QN => n114);
   Table_reg_25_1_inst : DFF_X1 port map( D => n778, CK => CLK, Q => 
                           Table_25_1_port, QN => n63);
   Table_reg_24_1_inst : DFF_X1 port map( D => n775, CK => CLK, Q => 
                           Table_24_1_port, QN => n30);
   Table_reg_23_1_inst : DFF_X1 port map( D => n772, CK => CLK, Q => 
                           Table_23_1_port, QN => n121);
   Table_reg_22_1_inst : DFF_X1 port map( D => n769, CK => CLK, Q => 
                           Table_22_1_port, QN => n10);
   Table_reg_21_1_inst : DFF_X1 port map( D => n766, CK => CLK, Q => 
                           Table_21_1_port, QN => n32);
   Table_reg_20_1_inst : DFF_X1 port map( D => n763, CK => CLK, Q => 
                           Table_20_1_port, QN => n124);
   Table_reg_19_1_inst : DFF_X1 port map( D => n760, CK => CLK, Q => 
                           Table_19_1_port, QN => n106);
   Table_reg_18_1_inst : DFF_X1 port map( D => n757, CK => CLK, Q => 
                           Table_18_1_port, QN => n574);
   Table_reg_17_1_inst : DFF_X1 port map( D => n754, CK => CLK, Q => 
                           Table_17_1_port, QN => n91);
   Table_reg_15_1_inst : DFF_X1 port map( D => n748, CK => CLK, Q => 
                           Table_15_1_port, QN => n3);
   Table_reg_13_1_inst : DFF_X1 port map( D => n742, CK => CLK, Q => 
                           Table_13_1_port, QN => n92);
   Table_reg_12_1_inst : DFF_X1 port map( D => n739, CK => CLK, Q => n7, QN => 
                           n126);
   Table_reg_11_1_inst : DFF_X1 port map( D => n736, CK => CLK, Q => 
                           Table_11_1_port, QN => n86);
   Table_reg_10_1_inst : DFF_X1 port map( D => n733, CK => CLK, Q => 
                           Table_10_1_port, QN => n125);
   Table_reg_9_1_inst : DFF_X1 port map( D => n730, CK => CLK, Q => 
                           Table_9_1_port, QN => n89);
   Table_reg_8_1_inst : DFF_X1 port map( D => n727, CK => CLK, Q => 
                           Table_8_1_port, QN => n109);
   Table_reg_3_1_inst : DFF_X1 port map( D => n712, CK => CLK, Q => 
                           Table_3_1_port, QN => n35);
   Table_reg_7_1_inst : DFF_X1 port map( D => n724, CK => CLK, Q => 
                           Table_7_1_port, QN => n34);
   Table_reg_5_1_inst : DFF_X1 port map( D => n718, CK => CLK, Q => 
                           Table_5_1_port, QN => n56);
   Table_reg_0_1_inst : DFF_X1 port map( D => n703, CK => CLK, Q => 
                           Table_0_1_port, QN => n26);
   Table_reg_31_2_inst : DFF_X1 port map( D => n795, CK => CLK, Q => 
                           Table_31_2_port, QN => n104);
   Table_reg_16_2_inst : DFF_X1 port map( D => n750, CK => CLK, Q => 
                           Table_16_2_port, QN => n40);
   Table_reg_28_2_inst : DFF_X1 port map( D => n786, CK => CLK, Q => 
                           Table_28_2_port, QN => n249);
   Table_reg_27_2_inst : DFF_X1 port map( D => n783, CK => CLK, Q => 
                           Table_27_2_port, QN => n504);
   Table_reg_25_2_inst : DFF_X1 port map( D => n777, CK => CLK, Q => 
                           Table_25_2_port, QN => n50);
   Table_reg_19_2_inst : DFF_X1 port map( D => n759, CK => CLK, Q => 
                           Table_19_2_port, QN => n569);
   Table_reg_17_2_inst : DFF_X1 port map( D => n753, CK => CLK, Q => 
                           Table_17_2_port, QN => n586);
   Table_reg_13_2_inst : DFF_X1 port map( D => n741, CK => CLK, Q => 
                           Table_13_2_port, QN => n621);
   Table_reg_11_2_inst : DFF_X1 port map( D => n735, CK => CLK, Q => 
                           Table_11_2_port, QN => n636);
   Table_reg_9_2_inst : DFF_X1 port map( D => n729, CK => CLK, Q => 
                           Table_9_2_port, QN => n49);
   Table_reg_15_2_inst : DFF_X1 port map( D => n747, CK => CLK, Q => 
                           Table_15_2_port, QN => n603);
   Table_reg_30_2_inst : DFF_X1 port map( D => n792, CK => CLK, Q => 
                           Table_30_2_port, QN => n478);
   Table_reg_26_2_inst : DFF_X1 port map( D => n780, CK => CLK, Q => 
                           Table_26_2_port, QN => n513);
   Table_reg_24_2_inst : DFF_X1 port map( D => n774, CK => CLK, Q => 
                           Table_24_2_port, QN => n88);
   Table_reg_22_2_inst : DFF_X1 port map( D => n768, CK => CLK, Q => 
                           Table_22_2_port, QN => n547);
   Table_reg_18_2_inst : DFF_X1 port map( D => n756, CK => CLK, Q => 
                           Table_18_2_port, QN => n53);
   Table_reg_12_2_inst : DFF_X1 port map( D => n738, CK => CLK, Q => 
                           Table_12_2_port, QN => n115);
   Table_reg_10_2_inst : DFF_X1 port map( D => n732, CK => CLK, Q => 
                           Table_10_2_port, QN => n113);
   Table_reg_2_2_inst : DFF_X1 port map( D => n708, CK => CLK, Q => 
                           Table_2_2_port, QN => n46);
   U3 : AND2_X2 port map( A1 => n460, A2 => n383, ZN => n819);
   U4 : AOI211_X4 port map( C1 => n439, C2 => n438, A => RST, B => n437, ZN => 
                           n827);
   U5 : NAND2_X1 port map( A1 => n22, A2 => n100, ZN => n212);
   U6 : BUF_X1 port map( A => n824, Z => n130);
   U7 : BUF_X2 port map( A => n822, Z => n1);
   U8 : BUF_X1 port map( A => n815, Z => n128);
   U9 : AOI21_X1 port map( B1 => n291, B2 => WR1, A => n290, ZN => n815);
   U10 : BUF_X2 port map( A => n821, Z => n2);
   U11 : INV_X1 port map( A => ADD_WR1(1), ZN => n333);
   U12 : AND2_X1 port map( A1 => n103, A2 => n120, ZN => n119);
   U13 : NOR2_X1 port map( A1 => n8, A2 => Table_17_1_port, ZN => n227);
   U14 : AND3_X1 port map( A1 => n49, A2 => n89, A3 => n80, ZN => n228);
   U15 : INV_X1 port map( A => ADD_WR1(2), ZN => n334);
   U16 : BUF_X1 port map( A => n818, Z => n129);
   U17 : NOR2_X2 port map( A1 => ADD_WR1(1), A2 => n331, ZN => n480);
   U18 : NOR3_X2 port map( A1 => n333, A2 => n334, A3 => n332, ZN => n427);
   U19 : INV_X1 port map( A => ADD_WR1(0), ZN => n332);
   U20 : AND4_X1 port map( A1 => n97, A2 => n227, A3 => n228, A4 => n139, ZN =>
                           n143);
   U21 : AND2_X1 port map( A1 => n85, A2 => n88, ZN => n76);
   U22 : NOR2_X1 port map( A1 => n5, A2 => n6, ZN => n69);
   U23 : NAND2_X1 port map( A1 => n41, A2 => n19, ZN => n5);
   U24 : NAND2_X1 port map( A1 => n90, A2 => n92, ZN => n6);
   U25 : NAND2_X1 port map( A1 => n60, A2 => n586, ZN => n8);
   U26 : AND2_X1 port map( A1 => n138, A2 => n50, ZN => n97);
   U27 : OR2_X1 port map( A1 => n16, A2 => n39, ZN => n9);
   U28 : AND2_X1 port map( A1 => n134, A2 => n412, ZN => n12);
   U29 : NOR2_X1 port map( A1 => n14, A2 => Table_21_2_port, ZN => n73);
   U30 : NAND2_X1 port map( A1 => n84, A2 => n32, ZN => n14);
   U31 : AND2_X1 port map( A1 => n95, A2 => n101, ZN => n15);
   U32 : NOR2_X1 port map( A1 => n16, A2 => n39, ZN => n198);
   U33 : NAND2_X1 port map( A1 => n115, A2 => n126, ZN => n16);
   U34 : AND2_X1 port map( A1 => n23, A2 => n113, ZN => n18);
   U35 : AND2_X1 port map( A1 => n106, A2 => n86, ZN => n72);
   U36 : AND2_X1 port map( A1 => n82, A2 => n83, ZN => n71);
   U37 : NOR2_X1 port map( A1 => n20, A2 => Table_8_2_port, ZN => n200);
   U38 : NAND2_X1 port map( A1 => n105, A2 => n109, ZN => n20);
   U39 : AND2_X1 port map( A1 => n478, A2 => n58, ZN => n21);
   U40 : AND2_X1 port map( A1 => n547, A2 => n10, ZN => n22);
   U41 : AND2_X1 port map( A1 => n17, A2 => n125, ZN => n23);
   U42 : NOR2_X1 port map( A1 => Table_10_2_port, A2 => Table_10_1_port, ZN => 
                           n118);
   U43 : INV_X1 port map( A => ADD_CHECK2(4), ZN => n250);
   U44 : NOR4_X1 port map( A1 => n209, A2 => n112, A3 => n210, A4 => n212, ZN 
                           => n142);
   U45 : AND2_X1 port map( A1 => n572, A2 => n574, ZN => n141);
   U46 : AOI21_X1 port map( B1 => n463, B2 => n462, A => n461, ZN => n824);
   U47 : NAND4_X1 port map( A1 => n144, A2 => n145, A3 => n143, A4 => n142, ZN 
                           => BUSY_WINDOW);
   U48 : NOR2_X1 port map( A1 => n136, A2 => n135, ZN => n144);
   U49 : AND2_X1 port map( A1 => n360, A2 => n104, ZN => n134);
   U50 : AND3_X1 port map( A1 => n539, A2 => n116, A3 => n121, ZN => n110);
   U51 : AND2_X1 port map( A1 => n3, A2 => n603, ZN => n95);
   U52 : NOR2_X1 port map( A1 => RST, A2 => n407, ZN => n818);
   U53 : AOI221_X1 port map( B1 => ADD_WR1(4), B2 => n313, C1 => n344, C2 => 
                           ADD_WR2(4), A => n288, ZN => n291);
   U54 : AND2_X1 port map( A1 => n248, A2 => n249, ZN => n137);
   U55 : NOR2_X1 port map( A1 => n77, A2 => n75, ZN => n145);
   U56 : AND2_X1 port map( A1 => n81, A2 => n30, ZN => n74);
   U57 : AND2_X1 port map( A1 => n487, A2 => n93, ZN => n103);
   U58 : AND2_X1 port map( A1 => n636, A2 => n569, ZN => n33);
   U59 : INV_X1 port map( A => n497, ZN => n695);
   U60 : INV_X1 port map( A => n515, ZN => n807);
   U61 : INV_X1 port map( A => n489, ZN => n687);
   U62 : INV_X1 port map( A => n469, ZN => n671);
   U63 : INV_X1 port map( A => n506, ZN => n799);
   U64 : INV_X1 port map( A => n523, ZN => n817);
   U65 : INV_X1 port map( A => n427, ZN => n663);
   U66 : INV_X1 port map( A => n480, ZN => n679);
   U67 : INV_X1 port map( A => RST, ZN => n131);
   U68 : INV_X1 port map( A => RST, ZN => n132);
   U69 : INV_X1 port map( A => ADD_WR2(2), ZN => n293);
   U70 : INV_X1 port map( A => ADD_WR2(4), ZN => n313);
   U71 : NOR3_X2 port map( A1 => ADD_WR1(0), A2 => n334, A3 => n333, ZN => n469
                           );
   U72 : NOR3_X2 port map( A1 => ADD_WR1(1), A2 => ADD_WR1(0), A3 => n334, ZN 
                           => n489);
   U73 : NOR3_X2 port map( A1 => ADD_WR1(2), A2 => n333, A3 => n332, ZN => n497
                           );
   U74 : NOR3_X2 port map( A1 => ADD_WR1(2), A2 => ADD_WR1(0), A3 => n333, ZN 
                           => n506);
   U75 : NOR3_X2 port map( A1 => ADD_WR1(1), A2 => ADD_WR1(2), A3 => n332, ZN 
                           => n515);
   U76 : NOR3_X2 port map( A1 => ADD_WR1(1), A2 => ADD_WR1(2), A3 => ADD_WR1(0)
                           , ZN => n523);
   U77 : AOI22_X1 port map( A1 => n590, A2 => n593, B1 => n595, B2 => n51, ZN 
                           => n751);
   U78 : AOI22_X1 port map( A1 => n589, A2 => n593, B1 => n595, B2 => n31, ZN 
                           => n752);
   U79 : AOI22_X1 port map( A1 => n594, A2 => n593, B1 => n595, B2 => n40, ZN 
                           => n750);
   U80 : OAI211_X1 port map( C1 => n247, C2 => n246, A => n245, B => n244, ZN 
                           => BUSY);
   U81 : AOI22_X1 port map( A1 => n243, A2 => n242, B1 => n241, B2 => n240, ZN 
                           => n244);
   U82 : OAI211_X1 port map( C1 => n278, C2 => n279, A => n239, B => n238, ZN 
                           => n241);
   U83 : AOI21_X1 port map( B1 => n237, B2 => n236, A => n235, ZN => n238);
   U84 : INV_X1 port map( A => n73, ZN => n236);
   U85 : NAND2_X1 port map( A1 => n284, A2 => n233, ZN => n239);
   U86 : OAI211_X1 port map( C1 => n280, C2 => n279, A => n232, B => n231, ZN 
                           => n242);
   U87 : AOI21_X1 port map( B1 => n237, B2 => n230, A => n229, ZN => n231);
   U88 : AOI211_X1 port map( C1 => n225, C2 => n224, A => n223, B => n222, ZN 
                           => n245);
   U89 : AOI211_X1 port map( C1 => ADD_CHECK2(3), C2 => n221, A => 
                           ADD_CHECK2(0), B => n220, ZN => n222);
   U90 : AOI21_X1 port map( B1 => n219, B2 => n218, A => ADD_CHECK2(3), ZN => 
                           n220);
   U91 : INV_X1 port map( A => n211, ZN => n213);
   U92 : OAI211_X1 port map( C1 => n254, C2 => n208, A => n207, B => n206, ZN 
                           => n219);
   U93 : NAND2_X1 port map( A1 => n243, A2 => n257, ZN => n206);
   U94 : AOI211_X1 port map( C1 => n240, C2 => n205, A => ADD_CHECK2(4), B => 
                           n204, ZN => n207);
   U95 : NOR2_X1 port map( A1 => n211, A2 => n255, ZN => n204);
   U96 : OAI21_X1 port map( B1 => n203, B2 => n202, A => n250, ZN => n221);
   U97 : INV_X1 port map( A => n240, ZN => n216);
   U98 : AND2_X1 port map( A1 => n197, A2 => ADD_CHECK2(2), ZN => n240);
   U99 : INV_X1 port map( A => ADD_CHECK2(1), ZN => n197);
   U100 : INV_X1 port map( A => n243, ZN => n199);
   U101 : NOR2_X1 port map( A1 => ADD_CHECK2(2), A2 => ADD_CHECK2(1), ZN => 
                           n243);
   U102 : OAI211_X1 port map( C1 => n196, C2 => n211, A => n195, B => n194, ZN 
                           => n223);
   U103 : OAI21_X1 port map( B1 => n193, B2 => n192, A => n265, ZN => n194);
   U104 : AOI21_X1 port map( B1 => n262, B2 => n188, A => n187, ZN => n195);
   U105 : OAI21_X1 port map( B1 => n186, B2 => n259, A => n185, ZN => n187);
   U106 : OAI21_X1 port map( B1 => n184, B2 => n183, A => n272, ZN => n185);
   U107 : OAI22_X1 port map( A1 => n15, A2 => n270, B1 => n268, B2 => n269, ZN 
                           => n183);
   U108 : OAI22_X1 port map( A1 => n110, A2 => n266, B1 => n12, B2 => n267, ZN 
                           => n184);
   U109 : AOI211_X1 port map( C1 => n182, C2 => n181, A => n180, B => n179, ZN 
                           => n186);
   U110 : NOR2_X1 port map( A1 => n278, A2 => n268, ZN => n179);
   U111 : OAI22_X1 port map( A1 => n266, A2 => n73, B1 => n270, B2 => n234, ZN 
                           => n180);
   U112 : INV_X1 port map( A => n119, ZN => n181);
   U113 : OAI21_X1 port map( B1 => n268, B2 => n280, A => n178, ZN => n188);
   U114 : AOI21_X1 port map( B1 => n182, B2 => n177, A => n176, ZN => n178);
   U115 : INV_X1 port map( A => n97, ZN => n177);
   U116 : INV_X1 port map( A => n267, ZN => n182);
   U117 : INV_X1 port map( A => ADD_CHECK1(4), ZN => n261);
   U118 : NAND2_X1 port map( A1 => ADD_CHECK2(1), A2 => ADD_CHECK2(2), ZN => 
                           n211);
   U119 : AOI21_X1 port map( B1 => n237, B2 => n175, A => n174, ZN => n196);
   U120 : NAND2_X1 port map( A1 => n276, A2 => n277, ZN => n171);
   U121 : INV_X1 port map( A => n282, ZN => n167);
   U122 : INV_X1 port map( A => n281, ZN => n170);
   U123 : INV_X1 port map( A => n110, ZN => n175);
   U124 : INV_X1 port map( A => n283, ZN => n237);
   U125 : AOI211_X1 port map( C1 => n274, C2 => n277, A => n165, B => n164, ZN 
                           => n166);
   U126 : NOR3_X1 port map( A1 => Table_27_2_port, A2 => Table_27_0_port, A3 =>
                           Table_27_1_port, ZN => n190);
   U127 : AND2_X1 port map( A1 => n66, A2 => n636, ZN => n189);
   U128 : NOR2_X1 port map( A1 => Table_11_0_port, A2 => Table_11_1_port, ZN =>
                           n66);
   U129 : AND2_X1 port map( A1 => n67, A2 => n569, ZN => n191);
   U130 : NOR2_X1 port map( A1 => Table_19_0_port, A2 => Table_19_1_port, ZN =>
                           n67);
   U131 : INV_X1 port map( A => n208, ZN => n225);
   U132 : NAND2_X1 port map( A1 => n163, A2 => ADD_CHECK2(1), ZN => n208);
   U133 : INV_X1 port map( A => ADD_CHECK2(2), ZN => n163);
   U134 : NAND2_X1 port map( A1 => n162, A2 => n161, ZN => n246);
   U135 : INV_X1 port map( A => ADD_CHECK1(0), ZN => n161);
   U136 : OAI21_X1 port map( B1 => n160, B2 => n159, A => ADD_CHECK1(4), ZN => 
                           n162);
   U137 : AOI211_X1 port map( C1 => n263, C2 => n233, A => n260, B => n156, ZN 
                           => n157);
   U138 : INV_X1 port map( A => n112, ZN => n173);
   U139 : NAND2_X1 port map( A1 => n76, A2 => n30, ZN => n226);
   U140 : NOR2_X1 port map( A1 => n107, A2 => n253, ZN => n153);
   U141 : AOI21_X1 port map( B1 => n152, B2 => n151, A => ADD_CHECK1(4), ZN => 
                           n247);
   U142 : AOI211_X1 port map( C1 => n96, C2 => n265, A => n149, B => n260, ZN 
                           => n150);
   U143 : NAND2_X1 port map( A1 => n9, A2 => n263, ZN => n148);
   U144 : OAI21_X1 port map( B1 => n259, B2 => n147, A => n258, ZN => n152);
   U145 : NOR2_X1 port map( A1 => n133, A2 => Table_2_2_port, ZN => n254);
   U146 : OR2_X1 port map( A1 => Table_2_0_port, A2 => Table_2_1_port, ZN => 
                           n133);
   U147 : NOR3_X1 port map( A1 => Table_6_2_port, A2 => Table_6_0_port, A3 => 
                           Table_6_1_port, ZN => n255);
   U148 : INV_X1 port map( A => n205, ZN => n147);
   U149 : NAND2_X1 port map( A1 => n146, A2 => n48, ZN => n205);
   U150 : NOR2_X1 port map( A1 => Table_4_0_port, A2 => Table_4_1_port, ZN => 
                           n146);
   U151 : INV_X1 port map( A => n233, ZN => n139);
   U152 : NAND2_X1 port map( A1 => n137, A2 => n94, ZN => n233);
   U153 : NOR3_X1 port map( A1 => Table_13_2_port, A2 => Table_13_0_port, A3 =>
                           Table_13_1_port, ZN => n234);
   U154 : NAND4_X1 port map( A1 => n70, A2 => n69, A3 => n68, A4 => n33, ZN => 
                           n135);
   U155 : NOR2_X1 port map( A1 => Table_13_2_port, A2 => Table_27_2_port, ZN =>
                           n68);
   U156 : AND2_X1 port map( A1 => n72, A2 => n71, ZN => n70);
   U157 : NAND4_X1 port map( A1 => n15, A2 => n73, A3 => n110, A4 => n12, ZN =>
                           n136);
   U158 : NAND4_X1 port map( A1 => n74, A2 => n200, A3 => n76, A4 => n198, ZN 
                           => n75);
   U159 : NAND4_X1 port map( A1 => n18, A2 => n119, A3 => n78, A4 => n98, ZN =>
                           n77);
   U160 : NOR2_X1 port map( A1 => n79, A2 => n99, ZN => n78);
   U161 : NAND2_X1 port map( A1 => n108, A2 => n122, ZN => n79);
   U162 : NAND2_X1 port map( A1 => n23, A2 => n113, ZN => n96);
   U163 : AND3_X1 port map( A1 => n613, A2 => n606, A3 => n608, ZN => n81);
   U164 : AOI22_X1 port map( A1 => n225, A2 => n210, B1 => n243, B2 => n209, ZN
                           => n215);
   U165 : AOI21_X1 port map( B1 => n262, B2 => n209, A => n155, ZN => n160);
   U166 : AOI21_X1 port map( B1 => n213, B2 => n212, A => n250, ZN => n214);
   U167 : AOI211_X1 port map( C1 => n272, C2 => n212, A => n153, B => 
                           ADD_CHECK1(3), ZN => n154);
   U168 : NAND2_X1 port map( A1 => n140, A2 => n31, ZN => n209);
   U169 : OAI22_X1 port map( A1 => n281, A2 => n228, B1 => n97, B2 => n282, ZN 
                           => n229);
   U170 : NOR2_X1 port map( A1 => Table_20_2_port, A2 => Table_20_1_port, ZN =>
                           n98);
   U171 : NAND2_X1 port map( A1 => n513, A2 => n114, ZN => n99);
   U172 : NAND2_X1 port map( A1 => n284, A2 => n226, ZN => n232);
   U173 : AOI21_X1 port map( B1 => n262, B2 => n226, A => n158, ZN => n159);
   U174 : NOR2_X1 port map( A1 => Table_16_1_port, A2 => Table_16_2_port, ZN =>
                           n140);
   U175 : AND2_X1 port map( A1 => n127, A2 => n513, ZN => n102);
   U176 : AND2_X1 port map( A1 => n141, A2 => n53, ZN => n107);
   U177 : NAND2_X1 port map( A1 => n21, A2 => n55, ZN => n112);
   U178 : OAI21_X1 port map( B1 => n283, B2 => n191, A => n166, ZN => n224);
   U179 : AOI22_X1 port map( A1 => n170, A2 => n169, B1 => n168, B2 => n167, ZN
                           => n172);
   U180 : INV_X1 port map( A => n227, ZN => n230);
   U181 : OAI22_X1 port map( A1 => n270, A2 => n228, B1 => n266, B2 => n227, ZN
                           => n176);
   U182 : OAI22_X1 port map( A1 => n189, A2 => n270, B1 => n268, B2 => n264, ZN
                           => n193);
   U183 : NAND2_X1 port map( A1 => n141, A2 => n53, ZN => n210);
   U184 : NOR2_X1 port map( A1 => Table_25_0_port, A2 => Table_25_1_port, ZN =>
                           n138);
   U185 : NAND2_X1 port map( A1 => n134, A2 => n412, ZN => n168);
   U186 : AND2_X1 port map( A1 => n122, A2 => n117, ZN => n217);
   U187 : NOR2_X1 port map( A1 => Table_20_1_port, A2 => Table_20_2_port, ZN =>
                           n117);
   U188 : AND2_X1 port map( A1 => n118, A2 => n17, ZN => n201);
   U189 : OAI22_X1 port map( A1 => n191, A2 => n266, B1 => n190, B2 => n267, ZN
                           => n192);
   U190 : OAI22_X1 port map( A1 => n189, A2 => n281, B1 => n190, B2 => n282, ZN
                           => n164);
   U191 : OAI21_X1 port map( B1 => n81, B2 => n271, A => n150, ZN => n151);
   U192 : NAND2_X1 port map( A1 => n95, A2 => n101, ZN => n169);
   U193 : OAI21_X1 port map( B1 => n271, B2 => n173, A => n157, ZN => n158);
   U194 : OAI211_X1 port map( C1 => n173, C2 => n275, A => n172, B => n171, ZN 
                           => n174);
   U195 : NOR2_X1 port map( A1 => Table_26_0_port, A2 => Table_26_1_port, ZN =>
                           n127);
   U196 : OAI21_X1 port map( B1 => n200, B2 => n252, A => n148, ZN => n149);
   U197 : OAI22_X1 port map( A1 => n282, A2 => n119, B1 => n234, B2 => n281, ZN
                           => n235);
   U198 : OAI22_X1 port map( A1 => n208, A2 => n201, B1 => n81, B2 => n211, ZN 
                           => n202);
   U199 : OAI22_X1 port map( A1 => n200, A2 => n199, B1 => n216, B2 => n198, ZN
                           => n203);
   U200 : OAI21_X1 port map( B1 => n259, B2 => n217, A => n154, ZN => n155);
   U201 : OAI211_X1 port map( C1 => n217, C2 => n216, A => n215, B => n214, ZN 
                           => n218);
   U202 : NOR2_X1 port map( A1 => n102, A2 => n253, ZN => n156);
   U203 : NOR2_X1 port map( A1 => n102, A2 => n275, ZN => n165);
   U204 : NAND3_X1 port map( A1 => n36, A2 => n29, A3 => n26, ZN => n257);
   U205 : NOR2_X1 port map( A1 => ADD_CHECK1(1), A2 => ADD_CHECK1(2), ZN => 
                           n262);
   U206 : INV_X1 port map( A => ADD_CHECK1(3), ZN => n260);
   U207 : NAND2_X1 port map( A1 => ADD_CHECK1(1), A2 => ADD_CHECK1(2), ZN => 
                           n271);
   U208 : INV_X1 port map( A => ADD_CHECK1(1), ZN => n251);
   U209 : NOR2_X1 port map( A1 => ADD_CHECK1(2), A2 => n251, ZN => n265);
   U210 : INV_X1 port map( A => n265, ZN => n253);
   U211 : NAND2_X1 port map( A1 => n251, A2 => ADD_CHECK1(2), ZN => n259);
   U212 : INV_X1 port map( A => n259, ZN => n263);
   U213 : INV_X1 port map( A => n262, ZN => n252);
   U214 : OAI22_X1 port map( A1 => n255, A2 => n271, B1 => n254, B2 => n253, ZN
                           => n256);
   U215 : AOI211_X1 port map( C1 => n262, C2 => n257, A => ADD_CHECK1(3), B => 
                           n256, ZN => n258);
   U216 : NAND3_X1 port map( A1 => ADD_CHECK1(4), A2 => ADD_CHECK1(0), A3 => 
                           n260, ZN => n266);
   U217 : NAND3_X1 port map( A1 => ADD_CHECK1(0), A2 => ADD_CHECK1(4), A3 => 
                           ADD_CHECK1(3), ZN => n267);
   U218 : NAND3_X1 port map( A1 => ADD_CHECK1(0), A2 => ADD_CHECK1(3), A3 => 
                           n261, ZN => n270);
   U219 : NOR3_X1 port map( A1 => Table_1_1_port, A2 => Table_1_0_port, A3 => 
                           Table_1_2_port, ZN => n280);
   U220 : NAND3_X1 port map( A1 => ADD_CHECK1(0), A2 => n261, A3 => n260, ZN =>
                           n268);
   U221 : NOR3_X1 port map( A1 => Table_5_1_port, A2 => Table_5_0_port, A3 => 
                           Table_5_2_port, ZN => n278);
   U222 : NAND3_X1 port map( A1 => n35, A2 => n28, A3 => n25, ZN => n274);
   U223 : INV_X1 port map( A => n274, ZN => n264);
   U224 : NAND3_X1 port map( A1 => n34, A2 => n27, A3 => n24, ZN => n276);
   U225 : INV_X1 port map( A => n276, ZN => n269);
   U226 : INV_X1 port map( A => n271, ZN => n272);
   U227 : INV_X1 port map( A => ADD_CHECK2(3), ZN => n273);
   U228 : NAND3_X1 port map( A1 => n273, A2 => n250, A3 => ADD_CHECK2(0), ZN =>
                           n279);
   U229 : INV_X1 port map( A => n279, ZN => n277);
   U230 : NAND3_X1 port map( A1 => ADD_CHECK2(0), A2 => ADD_CHECK2(3), A3 => 
                           ADD_CHECK2(4), ZN => n282);
   U231 : NAND3_X1 port map( A1 => ADD_CHECK2(3), A2 => ADD_CHECK2(0), A3 => 
                           n250, ZN => n281);
   U232 : NAND3_X1 port map( A1 => ADD_CHECK2(0), A2 => ADD_CHECK2(4), A3 => 
                           n273, ZN => n283);
   U233 : NOR3_X1 port map( A1 => n273, A2 => n250, A3 => ADD_CHECK2(0), ZN => 
                           n284);
   U234 : INV_X1 port map( A => n284, ZN => n275);
   U235 : NAND2_X1 port map( A1 => ADD_WR1(3), A2 => ADD_WR1(4), ZN => n470);
   U236 : NOR2_X1 port map( A1 => n663, A2 => n470, ZN => n421);
   U237 : INV_X1 port map( A => ADD_WR1(4), ZN => n344);
   U238 : INV_X1 port map( A => ADD_WR2(0), ZN => n296);
   U239 : INV_X1 port map( A => ADD_WR1(3), ZN => n349);
   U240 : AOI22_X1 port map( A1 => n333, A2 => ADD_WR2(1), B1 => ADD_WR2(3), B2
                           => n349, ZN => n285);
   U241 : OAI221_X1 port map( B1 => n333, B2 => ADD_WR2(1), C1 => n349, C2 => 
                           ADD_WR2(3), A => n285, ZN => n286);
   U242 : AOI221_X1 port map( B1 => ADD_WR1(0), B2 => n296, C1 => n332, C2 => 
                           ADD_WR2(0), A => n286, ZN => n287);
   U243 : OAI221_X1 port map( B1 => ADD_WR1(2), B2 => n293, C1 => n334, C2 => 
                           ADD_WR2(2), A => n287, ZN => n288);
   U244 : INV_X1 port map( A => WR1, ZN => n289);
   U245 : AOI21_X1 port map( B1 => n291, B2 => WR2, A => n289, ZN => n661);
   U246 : INV_X1 port map( A => WR2, ZN => n290);
   U247 : NAND2_X1 port map( A1 => ADD_WR2(4), A2 => ADD_WR2(3), ZN => n297);
   U248 : NAND3_X1 port map( A1 => ADD_WR2(2), A2 => ADD_WR2(0), A3 => 
                           ADD_WR2(1), ZN => n322);
   U249 : NOR2_X1 port map( A1 => n297, A2 => n322, ZN => n464);
   U250 : NAND2_X1 port map( A1 => n128, A2 => n464, ZN => n465);
   U251 : INV_X1 port map( A => n465, ZN => n292);
   U252 : AOI211_X1 port map( C1 => n421, C2 => n661, A => RST, B => n292, ZN 
                           => n468);
   U253 : NAND2_X1 port map( A1 => n132, A2 => n128, ZN => n381);
   U254 : INV_X1 port map( A => n381, ZN => n460);
   U255 : NOR2_X1 port map( A1 => ADD_WR2(0), A2 => ADD_WR2(1), ZN => n295);
   U256 : NAND2_X1 port map( A1 => n295, A2 => n293, ZN => n314);
   U257 : NOR2_X1 port map( A1 => n297, A2 => n314, ZN => n527);
   U258 : INV_X1 port map( A => ADD_WR2(1), ZN => n294);
   U259 : NAND3_X1 port map( A1 => ADD_WR2(0), A2 => n293, A3 => n294, ZN => 
                           n315);
   U260 : NOR2_X1 port map( A1 => n297, A2 => n315, ZN => n518);
   U261 : AOI22_X1 port map( A1 => Table_24_0_port, A2 => n527, B1 => 
                           Table_25_0_port, B2 => n518, ZN => n301);
   U262 : NAND3_X1 port map( A1 => ADD_WR2(1), A2 => n293, A3 => n296, ZN => 
                           n316);
   U263 : NOR2_X1 port map( A1 => n297, A2 => n316, ZN => n509);
   U264 : NAND3_X1 port map( A1 => ADD_WR2(0), A2 => ADD_WR2(1), A3 => n293, ZN
                           => n317);
   U265 : NOR2_X1 port map( A1 => n297, A2 => n317, ZN => n500);
   U266 : AOI22_X1 port map( A1 => Table_26_0_port, A2 => n509, B1 => 
                           Table_27_0_port, B2 => n500, ZN => n300);
   U267 : NAND3_X1 port map( A1 => ADD_WR2(0), A2 => ADD_WR2(2), A3 => n294, ZN
                           => n319);
   U268 : NOR2_X1 port map( A1 => n297, A2 => n319, ZN => n483);
   U269 : NAND2_X1 port map( A1 => ADD_WR2(2), A2 => n295, ZN => n318);
   U270 : NOR2_X1 port map( A1 => n297, A2 => n318, ZN => n492);
   U271 : AOI22_X1 port map( A1 => Table_29_0_port, A2 => n483, B1 => 
                           Table_28_0_port, B2 => n492, ZN => n299);
   U272 : NAND3_X1 port map( A1 => ADD_WR2(2), A2 => ADD_WR2(1), A3 => n296, ZN
                           => n320);
   U273 : NOR2_X1 port map( A1 => n297, A2 => n320, ZN => n474);
   U274 : AOI22_X1 port map( A1 => Table_30_0_port, A2 => n474, B1 => 
                           Table_31_0_port, B2 => n464, ZN => n298);
   U275 : NAND4_X1 port map( A1 => n301, A2 => n300, A3 => n299, A4 => n298, ZN
                           => n330);
   U276 : INV_X1 port map( A => ADD_WR2(3), ZN => n312);
   U277 : NAND2_X1 port map( A1 => ADD_WR2(4), A2 => n312, ZN => n302);
   U278 : NOR2_X1 port map( A1 => n314, A2 => n302, ZN => n591);
   U279 : NOR2_X1 port map( A1 => n315, A2 => n302, ZN => n582);
   U280 : AOI22_X1 port map( A1 => Table_16_0_port, A2 => n591, B1 => n11, B2 
                           => n582, ZN => n306);
   U281 : NOR2_X1 port map( A1 => n316, A2 => n302, ZN => n575);
   U282 : NOR2_X1 port map( A1 => n317, A2 => n302, ZN => n565);
   U283 : AOI22_X1 port map( A1 => Table_18_0_port, A2 => n575, B1 => 
                           Table_19_0_port, B2 => n565, ZN => n305);
   U284 : NOR2_X1 port map( A1 => n318, A2 => n302, ZN => n558);
   U285 : NOR2_X1 port map( A1 => n319, A2 => n302, ZN => n551);
   U286 : AOI22_X1 port map( A1 => n38, A2 => n558, B1 => n13, B2 => n551, ZN 
                           => n304);
   U287 : NOR2_X1 port map( A1 => n320, A2 => n302, ZN => n543);
   U288 : NOR2_X1 port map( A1 => n322, A2 => n302, ZN => n535);
   U289 : AOI22_X1 port map( A1 => Table_22_0_port, A2 => n543, B1 => 
                           Table_23_0_port, B2 => n535, ZN => n303);
   U290 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => n329);
   U291 : NAND2_X1 port map( A1 => ADD_WR2(3), A2 => n313, ZN => n307);
   U292 : NOR2_X1 port map( A1 => n314, A2 => n307, ZN => n655);
   U293 : NOR2_X1 port map( A1 => n315, A2 => n307, ZN => n647);
   U294 : AOI22_X1 port map( A1 => n4, A2 => n655, B1 => Table_9_0_port, B2 => 
                           n647, ZN => n311);
   U295 : NOR2_X1 port map( A1 => n316, A2 => n307, ZN => n640);
   U296 : NOR2_X1 port map( A1 => n317, A2 => n307, ZN => n632);
   U297 : AOI22_X1 port map( A1 => n37, A2 => n640, B1 => Table_11_0_port, B2 
                           => n632, ZN => n310);
   U298 : NOR2_X1 port map( A1 => n318, A2 => n307, ZN => n625);
   U299 : NOR2_X1 port map( A1 => n319, A2 => n307, ZN => n617);
   U300 : AOI22_X1 port map( A1 => n39, A2 => n625, B1 => Table_13_0_port, B2 
                           => n617, ZN => n309);
   U301 : NOR2_X1 port map( A1 => n320, A2 => n307, ZN => n609);
   U302 : NOR2_X1 port map( A1 => n322, A2 => n307, ZN => n599);
   U303 : AOI22_X1 port map( A1 => Table_14_0_port, A2 => n609, B1 => 
                           Table_15_0_port, B2 => n599, ZN => n308);
   U304 : NAND4_X1 port map( A1 => n311, A2 => n310, A3 => n309, A4 => n308, ZN
                           => n328);
   U305 : NAND2_X1 port map( A1 => n313, A2 => n312, ZN => n321);
   U306 : NOR2_X1 port map( A1 => n314, A2 => n321, ZN => n825);
   U307 : NOR2_X1 port map( A1 => n315, A2 => n321, ZN => n810);
   U308 : AOI22_X1 port map( A1 => Table_0_0_port, A2 => n825, B1 => 
                           Table_1_0_port, B2 => n810, ZN => n326);
   U309 : NOR2_X1 port map( A1 => n316, A2 => n321, ZN => n802);
   U310 : NOR2_X1 port map( A1 => n317, A2 => n321, ZN => n698);
   U311 : AOI22_X1 port map( A1 => Table_2_0_port, A2 => n802, B1 => 
                           Table_3_0_port, B2 => n698, ZN => n325);
   U312 : NOR2_X1 port map( A1 => n318, A2 => n321, ZN => n690);
   U313 : NOR2_X1 port map( A1 => n319, A2 => n321, ZN => n682);
   U314 : AOI22_X1 port map( A1 => Table_4_0_port, A2 => n690, B1 => 
                           Table_5_0_port, B2 => n682, ZN => n324);
   U315 : NOR2_X1 port map( A1 => n320, A2 => n321, ZN => n674);
   U316 : NOR2_X1 port map( A1 => n322, A2 => n321, ZN => n666);
   U317 : AOI22_X1 port map( A1 => Table_6_0_port, A2 => n674, B1 => 
                           Table_7_0_port, B2 => n666, ZN => n323);
   U318 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => n327);
   U319 : NOR4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN 
                           => n383);
   U320 : NAND2_X1 port map( A1 => ADD_WR1(2), A2 => ADD_WR1(0), ZN => n331);
   U321 : AOI22_X1 port map( A1 => n523, A2 => Table_24_0_port, B1 => n515, B2 
                           => Table_25_0_port, ZN => n337);
   U322 : AOI22_X1 port map( A1 => n506, A2 => Table_26_0_port, B1 => n497, B2 
                           => Table_27_0_port, ZN => n336);
   U323 : AOI22_X1 port map( A1 => n489, A2 => Table_28_0_port, B1 => n469, B2 
                           => Table_30_0_port, ZN => n335);
   U324 : NAND3_X1 port map( A1 => n337, A2 => n336, A3 => n335, ZN => n338);
   U325 : AOI21_X1 port map( B1 => n480, B2 => Table_29_0_port, A => n338, ZN 
                           => n358);
   U326 : NOR2_X1 port map( A1 => ADD_WR1(3), A2 => ADD_WR1(4), ZN => n662);
   U327 : AOI22_X1 port map( A1 => n523, A2 => Table_0_0_port, B1 => n515, B2 
                           => Table_1_0_port, ZN => n342);
   U328 : AOI22_X1 port map( A1 => n506, A2 => Table_2_0_port, B1 => n497, B2 
                           => Table_3_0_port, ZN => n341);
   U329 : AOI22_X1 port map( A1 => n489, A2 => Table_4_0_port, B1 => n480, B2 
                           => Table_5_0_port, ZN => n340);
   U330 : AOI22_X1 port map( A1 => n469, A2 => Table_6_0_port, B1 => n427, B2 
                           => Table_7_0_port, ZN => n339);
   U331 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => n343);
   U332 : AOI22_X1 port map( A1 => n662, A2 => n343, B1 => n421, B2 => 
                           Table_31_0_port, ZN => n357);
   U333 : NOR2_X1 port map( A1 => ADD_WR1(3), A2 => n344, ZN => n532);
   U334 : AOI22_X1 port map( A1 => n523, A2 => Table_16_0_port, B1 => n515, B2 
                           => n11, ZN => n348);
   U335 : AOI22_X1 port map( A1 => n506, A2 => Table_18_0_port, B1 => n497, B2 
                           => Table_19_0_port, ZN => n347);
   U336 : AOI22_X1 port map( A1 => n489, A2 => n38, B1 => n480, B2 => n13, ZN 
                           => n346);
   U337 : AOI22_X1 port map( A1 => n469, A2 => Table_22_0_port, B1 => n427, B2 
                           => Table_23_0_port, ZN => n345);
   U338 : NAND4_X1 port map( A1 => n348, A2 => n347, A3 => n346, A4 => n345, ZN
                           => n355);
   U339 : NOR2_X1 port map( A1 => ADD_WR1(4), A2 => n349, ZN => n596);
   U340 : AOI22_X1 port map( A1 => n523, A2 => n4, B1 => n515, B2 => 
                           Table_9_0_port, ZN => n353);
   U341 : AOI22_X1 port map( A1 => n506, A2 => n37, B1 => n497, B2 => 
                           Table_11_0_port, ZN => n352);
   U342 : AOI22_X1 port map( A1 => n489, A2 => n39, B1 => n480, B2 => 
                           Table_13_0_port, ZN => n351);
   U343 : AOI22_X1 port map( A1 => n469, A2 => Table_14_0_port, B1 => n427, B2 
                           => Table_15_0_port, ZN => n350);
   U344 : NAND4_X1 port map( A1 => n353, A2 => n352, A3 => n351, A4 => n350, ZN
                           => n354);
   U345 : AOI22_X1 port map( A1 => n532, A2 => n355, B1 => n596, B2 => n354, ZN
                           => n356);
   U346 : OAI211_X1 port map( C1 => n358, C2 => n470, A => n357, B => n356, ZN 
                           => n407);
   U347 : AOI22_X1 port map( A1 => n464, A2 => n819, B1 => n129, B2 => n465, ZN
                           => n359);
   U348 : INV_X1 port map( A => n468, ZN => n410);
   U349 : AOI22_X1 port map( A1 => n468, A2 => n360, B1 => n359, B2 => n410, ZN
                           => n797);
   U350 : AOI22_X1 port map( A1 => Table_24_1_port, A2 => n527, B1 => 
                           Table_25_1_port, B2 => n518, ZN => n364);
   U351 : AOI22_X1 port map( A1 => Table_26_1_port, A2 => n509, B1 => 
                           Table_27_1_port, B2 => n500, ZN => n363);
   U352 : AOI22_X1 port map( A1 => Table_29_1_port, A2 => n483, B1 => 
                           Table_28_1_port, B2 => n492, ZN => n362);
   U353 : AOI22_X1 port map( A1 => Table_30_1_port, A2 => n474, B1 => 
                           Table_31_1_port, B2 => n464, ZN => n361);
   U354 : NAND4_X1 port map( A1 => n364, A2 => n363, A3 => n362, A4 => n361, ZN
                           => n380);
   U355 : AOI22_X1 port map( A1 => Table_16_1_port, A2 => n591, B1 => 
                           Table_17_1_port, B2 => n582, ZN => n368);
   U356 : AOI22_X1 port map( A1 => Table_18_1_port, A2 => n575, B1 => 
                           Table_19_1_port, B2 => n565, ZN => n367);
   U357 : AOI22_X1 port map( A1 => Table_20_1_port, A2 => n558, B1 => 
                           Table_21_1_port, B2 => n551, ZN => n366);
   U358 : AOI22_X1 port map( A1 => Table_22_1_port, A2 => n543, B1 => 
                           Table_23_1_port, B2 => n535, ZN => n365);
   U359 : NAND4_X1 port map( A1 => n368, A2 => n367, A3 => n366, A4 => n365, ZN
                           => n379);
   U360 : AOI22_X1 port map( A1 => Table_8_1_port, A2 => n655, B1 => 
                           Table_9_1_port, B2 => n647, ZN => n372);
   U361 : AOI22_X1 port map( A1 => Table_10_1_port, A2 => n640, B1 => 
                           Table_11_1_port, B2 => n632, ZN => n371);
   U362 : AOI22_X1 port map( A1 => n7, A2 => n625, B1 => Table_13_1_port, B2 =>
                           n617, ZN => n370);
   U363 : AOI22_X1 port map( A1 => Table_14_1_port, A2 => n609, B1 => 
                           Table_15_1_port, B2 => n599, ZN => n369);
   U364 : NAND4_X1 port map( A1 => n372, A2 => n371, A3 => n370, A4 => n369, ZN
                           => n378);
   U365 : AOI22_X1 port map( A1 => Table_0_1_port, A2 => n825, B1 => 
                           Table_1_1_port, B2 => n810, ZN => n376);
   U366 : AOI22_X1 port map( A1 => Table_2_1_port, A2 => n802, B1 => 
                           Table_3_1_port, B2 => n698, ZN => n375);
   U367 : AOI22_X1 port map( A1 => Table_4_1_port, A2 => n690, B1 => 
                           Table_5_1_port, B2 => n682, ZN => n374);
   U368 : AOI22_X1 port map( A1 => Table_6_1_port, A2 => n674, B1 => 
                           Table_7_1_port, B2 => n666, ZN => n373);
   U369 : NAND4_X1 port map( A1 => n376, A2 => n375, A3 => n374, A4 => n373, ZN
                           => n377);
   U370 : NOR4_X1 port map( A1 => n380, A2 => n379, A3 => n378, A4 => n377, ZN 
                           => n382);
   U371 : NAND2_X1 port map( A1 => n382, A2 => n383, ZN => n462);
   U372 : AOI221_X1 port map( B1 => n383, B2 => n462, C1 => n382, C2 => n462, A
                           => n381, ZN => n822);
   U373 : AOI22_X1 port map( A1 => n523, A2 => Table_24_1_port, B1 => n515, B2 
                           => Table_25_1_port, ZN => n386);
   U374 : AOI22_X1 port map( A1 => n506, A2 => Table_26_1_port, B1 => n497, B2 
                           => Table_27_1_port, ZN => n385);
   U375 : AOI22_X1 port map( A1 => n489, A2 => Table_28_1_port, B1 => n469, B2 
                           => Table_30_1_port, ZN => n384);
   U376 : NAND3_X1 port map( A1 => n386, A2 => n385, A3 => n384, ZN => n387);
   U377 : AOI21_X1 port map( B1 => n480, B2 => Table_29_1_port, A => n387, ZN 
                           => n405);
   U378 : AOI22_X1 port map( A1 => n523, A2 => Table_0_1_port, B1 => n515, B2 
                           => Table_1_1_port, ZN => n391);
   U379 : AOI22_X1 port map( A1 => n506, A2 => Table_2_1_port, B1 => n497, B2 
                           => Table_3_1_port, ZN => n390);
   U380 : AOI22_X1 port map( A1 => n489, A2 => Table_4_1_port, B1 => n480, B2 
                           => Table_5_1_port, ZN => n389);
   U381 : AOI22_X1 port map( A1 => n469, A2 => Table_6_1_port, B1 => n427, B2 
                           => Table_7_1_port, ZN => n388);
   U382 : NAND4_X1 port map( A1 => n391, A2 => n390, A3 => n389, A4 => n388, ZN
                           => n392);
   U383 : AOI22_X1 port map( A1 => Table_31_1_port, A2 => n421, B1 => n662, B2 
                           => n392, ZN => n404);
   U384 : AOI22_X1 port map( A1 => n523, A2 => Table_8_1_port, B1 => n515, B2 
                           => Table_9_1_port, ZN => n396);
   U385 : AOI22_X1 port map( A1 => n506, A2 => Table_10_1_port, B1 => n497, B2 
                           => Table_11_1_port, ZN => n395);
   U386 : AOI22_X1 port map( A1 => n489, A2 => n7, B1 => n480, B2 => 
                           Table_13_1_port, ZN => n394);
   U387 : AOI22_X1 port map( A1 => n469, A2 => Table_14_1_port, B1 => n427, B2 
                           => Table_15_1_port, ZN => n393);
   U388 : NAND4_X1 port map( A1 => n396, A2 => n395, A3 => n394, A4 => n393, ZN
                           => n402);
   U389 : AOI22_X1 port map( A1 => n523, A2 => Table_16_1_port, B1 => n515, B2 
                           => Table_17_1_port, ZN => n400);
   U390 : AOI22_X1 port map( A1 => n506, A2 => Table_18_1_port, B1 => n497, B2 
                           => Table_19_1_port, ZN => n399);
   U391 : AOI22_X1 port map( A1 => n489, A2 => Table_20_1_port, B1 => n480, B2 
                           => Table_21_1_port, ZN => n398);
   U392 : AOI22_X1 port map( A1 => n469, A2 => Table_22_1_port, B1 => n427, B2 
                           => Table_23_1_port, ZN => n397);
   U393 : NAND4_X1 port map( A1 => n400, A2 => n399, A3 => n398, A4 => n397, ZN
                           => n401);
   U394 : AOI22_X1 port map( A1 => n596, A2 => n402, B1 => n532, B2 => n401, ZN
                           => n403);
   U395 : OAI211_X1 port map( C1 => n405, C2 => n470, A => n404, B => n403, ZN 
                           => n406);
   U396 : INV_X1 port map( A => n406, ZN => n409);
   U397 : INV_X1 port map( A => n407, ZN => n408);
   U398 : NOR2_X1 port map( A1 => n409, A2 => n408, ZN => n439);
   U399 : AOI211_X1 port map( C1 => n409, C2 => n408, A => RST, B => n439, ZN 
                           => n821);
   U400 : AOI22_X1 port map( A1 => n464, A2 => n1, B1 => n2, B2 => n465, ZN => 
                           n411);
   U401 : AOI22_X1 port map( A1 => n468, A2 => n412, B1 => n411, B2 => n410, ZN
                           => n796);
   U402 : AOI22_X1 port map( A1 => n523, A2 => Table_24_2_port, B1 => n515, B2 
                           => Table_25_2_port, ZN => n415);
   U403 : AOI22_X1 port map( A1 => n506, A2 => Table_26_2_port, B1 => n497, B2 
                           => Table_27_2_port, ZN => n414);
   U404 : AOI22_X1 port map( A1 => n489, A2 => Table_28_2_port, B1 => n469, B2 
                           => Table_30_2_port, ZN => n413);
   U405 : NAND3_X1 port map( A1 => n415, A2 => n414, A3 => n413, ZN => n416);
   U406 : AOI21_X1 port map( B1 => n480, B2 => Table_29_2_port, A => n416, ZN 
                           => n436);
   U407 : AOI22_X1 port map( A1 => n523, A2 => Table_0_2_port, B1 => n515, B2 
                           => Table_1_2_port, ZN => n420);
   U408 : AOI22_X1 port map( A1 => n506, A2 => Table_2_2_port, B1 => n497, B2 
                           => Table_3_2_port, ZN => n419);
   U409 : AOI22_X1 port map( A1 => n489, A2 => Table_4_2_port, B1 => n480, B2 
                           => Table_5_2_port, ZN => n418);
   U410 : AOI22_X1 port map( A1 => n469, A2 => Table_6_2_port, B1 => n427, B2 
                           => Table_7_2_port, ZN => n417);
   U411 : NAND4_X1 port map( A1 => n420, A2 => n419, A3 => n418, A4 => n417, ZN
                           => n422);
   U412 : AOI22_X1 port map( A1 => n662, A2 => n422, B1 => n421, B2 => 
                           Table_31_2_port, ZN => n435);
   U413 : AOI22_X1 port map( A1 => n523, A2 => Table_16_2_port, B1 => n515, B2 
                           => Table_17_2_port, ZN => n426);
   U414 : AOI22_X1 port map( A1 => n506, A2 => Table_18_2_port, B1 => n497, B2 
                           => Table_19_2_port, ZN => n425);
   U415 : AOI22_X1 port map( A1 => n489, A2 => Table_20_2_port, B1 => n480, B2 
                           => Table_21_2_port, ZN => n424);
   U416 : AOI22_X1 port map( A1 => n469, A2 => Table_22_2_port, B1 => n427, B2 
                           => Table_23_2_port, ZN => n423);
   U417 : NAND4_X1 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN
                           => n433);
   U418 : AOI22_X1 port map( A1 => n523, A2 => Table_8_2_port, B1 => n515, B2 
                           => Table_9_2_port, ZN => n431);
   U419 : AOI22_X1 port map( A1 => n506, A2 => Table_10_2_port, B1 => n497, B2 
                           => Table_11_2_port, ZN => n430);
   U420 : AOI22_X1 port map( A1 => n489, A2 => Table_12_2_port, B1 => n480, B2 
                           => Table_13_2_port, ZN => n429);
   U421 : AOI22_X1 port map( A1 => n469, A2 => Table_14_2_port, B1 => n427, B2 
                           => Table_15_2_port, ZN => n428);
   U422 : NAND4_X1 port map( A1 => n431, A2 => n430, A3 => n429, A4 => n428, ZN
                           => n432);
   U423 : AOI22_X1 port map( A1 => n532, A2 => n433, B1 => n596, B2 => n432, ZN
                           => n434);
   U424 : OAI211_X1 port map( C1 => n436, C2 => n470, A => n435, B => n434, ZN 
                           => n438);
   U425 : NOR2_X1 port map( A1 => n439, A2 => n438, ZN => n437);
   U426 : AOI22_X1 port map( A1 => Table_24_2_port, A2 => n527, B1 => 
                           Table_25_2_port, B2 => n518, ZN => n443);
   U427 : AOI22_X1 port map( A1 => Table_26_2_port, A2 => n509, B1 => 
                           Table_27_2_port, B2 => n500, ZN => n442);
   U428 : AOI22_X1 port map( A1 => Table_29_2_port, A2 => n483, B1 => 
                           Table_28_2_port, B2 => n492, ZN => n441);
   U429 : AOI22_X1 port map( A1 => Table_30_2_port, A2 => n474, B1 => 
                           Table_31_2_port, B2 => n464, ZN => n440);
   U430 : NAND4_X1 port map( A1 => n443, A2 => n442, A3 => n441, A4 => n440, ZN
                           => n459);
   U431 : AOI22_X1 port map( A1 => Table_16_2_port, A2 => n591, B1 => 
                           Table_17_2_port, B2 => n582, ZN => n447);
   U432 : AOI22_X1 port map( A1 => Table_18_2_port, A2 => n575, B1 => 
                           Table_19_2_port, B2 => n565, ZN => n446);
   U433 : AOI22_X1 port map( A1 => Table_20_2_port, A2 => n558, B1 => 
                           Table_21_2_port, B2 => n551, ZN => n445);
   U434 : AOI22_X1 port map( A1 => Table_22_2_port, A2 => n543, B1 => 
                           Table_23_2_port, B2 => n535, ZN => n444);
   U435 : NAND4_X1 port map( A1 => n447, A2 => n446, A3 => n445, A4 => n444, ZN
                           => n458);
   U436 : AOI22_X1 port map( A1 => Table_8_2_port, A2 => n655, B1 => 
                           Table_9_2_port, B2 => n647, ZN => n451);
   U437 : AOI22_X1 port map( A1 => Table_10_2_port, A2 => n640, B1 => 
                           Table_11_2_port, B2 => n632, ZN => n450);
   U438 : AOI22_X1 port map( A1 => Table_12_2_port, A2 => n625, B1 => 
                           Table_13_2_port, B2 => n617, ZN => n449);
   U439 : AOI22_X1 port map( A1 => Table_14_2_port, A2 => n609, B1 => 
                           Table_15_2_port, B2 => n599, ZN => n448);
   U440 : NAND4_X1 port map( A1 => n451, A2 => n450, A3 => n449, A4 => n448, ZN
                           => n457);
   U441 : AOI22_X1 port map( A1 => Table_0_2_port, A2 => n825, B1 => 
                           Table_1_2_port, B2 => n810, ZN => n455);
   U442 : AOI22_X1 port map( A1 => Table_2_2_port, A2 => n802, B1 => 
                           Table_3_2_port, B2 => n698, ZN => n454);
   U443 : AOI22_X1 port map( A1 => Table_4_2_port, A2 => n690, B1 => 
                           Table_5_2_port, B2 => n682, ZN => n453);
   U444 : AOI22_X1 port map( A1 => Table_6_2_port, A2 => n674, B1 => 
                           Table_7_2_port, B2 => n666, ZN => n452);
   U445 : NAND4_X1 port map( A1 => n455, A2 => n454, A3 => n453, A4 => n452, ZN
                           => n456);
   U446 : NOR4_X1 port map( A1 => n459, A2 => n458, A3 => n457, A4 => n456, ZN 
                           => n463);
   U447 : OAI21_X1 port map( B1 => n463, B2 => n462, A => n460, ZN => n461);
   U448 : AOI22_X1 port map( A1 => n827, A2 => n465, B1 => n464, B2 => n130, ZN
                           => n467);
   U449 : NAND2_X1 port map( A1 => n468, A2 => Table_31_2_port, ZN => n466);
   U450 : OAI21_X1 port map( B1 => n468, B2 => n467, A => n466, ZN => n795);
   U451 : INV_X1 port map( A => n470, ZN => n471);
   U452 : NAND2_X1 port map( A1 => n471, A2 => n661, ZN => n524);
   U453 : NAND2_X1 port map( A1 => n815, A2 => n474, ZN => n475);
   U454 : OAI211_X1 port map( C1 => n671, C2 => n524, A => n131, B => n475, ZN 
                           => n476);
   U455 : INV_X1 port map( A => n476, ZN => n479);
   U456 : AOI22_X1 port map( A1 => n474, A2 => n819, B1 => n129, B2 => n475, ZN
                           => n472);
   U457 : AOI22_X1 port map( A1 => n479, A2 => n55, B1 => n472, B2 => n476, ZN 
                           => n794);
   U458 : AOI22_X1 port map( A1 => n474, A2 => n1, B1 => n2, B2 => n475, ZN => 
                           n473);
   U459 : AOI22_X1 port map( A1 => n479, A2 => n58, B1 => n473, B2 => n476, ZN 
                           => n793);
   U460 : AOI22_X1 port map( A1 => n827, A2 => n475, B1 => n474, B2 => n130, ZN
                           => n477);
   U461 : AOI22_X1 port map( A1 => n479, A2 => n478, B1 => n477, B2 => n476, ZN
                           => n792);
   U462 : NAND2_X1 port map( A1 => n815, A2 => n483, ZN => n484);
   U463 : OAI211_X1 port map( C1 => n679, C2 => n524, A => n132, B => n484, ZN 
                           => n485);
   U464 : INV_X1 port map( A => n485, ZN => n488);
   U465 : AOI22_X1 port map( A1 => n483, A2 => n819, B1 => n818, B2 => n484, ZN
                           => n481);
   U466 : AOI22_X1 port map( A1 => n488, A2 => n120, B1 => n481, B2 => n485, ZN
                           => n791);
   U467 : AOI22_X1 port map( A1 => n483, A2 => n1, B1 => n2, B2 => n484, ZN => 
                           n482);
   U468 : AOI22_X1 port map( A1 => n488, A2 => n93, B1 => n482, B2 => n485, ZN 
                           => n790);
   U469 : AOI22_X1 port map( A1 => n827, A2 => n484, B1 => n483, B2 => n824, ZN
                           => n486);
   U470 : AOI22_X1 port map( A1 => n488, A2 => n487, B1 => n486, B2 => n485, ZN
                           => n789);
   U471 : NAND2_X1 port map( A1 => n815, A2 => n492, ZN => n493);
   U472 : OAI211_X1 port map( C1 => n687, C2 => n524, A => n131, B => n493, ZN 
                           => n494);
   U473 : INV_X1 port map( A => n494, ZN => n496);
   U474 : AOI22_X1 port map( A1 => n492, A2 => n819, B1 => n129, B2 => n493, ZN
                           => n490);
   U475 : AOI22_X1 port map( A1 => n496, A2 => n248, B1 => n490, B2 => n494, ZN
                           => n788);
   U476 : AOI22_X1 port map( A1 => n492, A2 => n1, B1 => n2, B2 => n493, ZN => 
                           n491);
   U477 : AOI22_X1 port map( A1 => n496, A2 => n94, B1 => n491, B2 => n494, ZN 
                           => n787);
   U478 : AOI22_X1 port map( A1 => n827, A2 => n493, B1 => n492, B2 => n130, ZN
                           => n495);
   U479 : AOI22_X1 port map( A1 => n496, A2 => n249, B1 => n495, B2 => n494, ZN
                           => n786);
   U480 : NAND2_X1 port map( A1 => n815, A2 => n500, ZN => n501);
   U481 : OAI211_X1 port map( C1 => n695, C2 => n524, A => n132, B => n501, ZN 
                           => n502);
   U482 : INV_X1 port map( A => n502, ZN => n505);
   U483 : AOI22_X1 port map( A1 => n500, A2 => n819, B1 => n129, B2 => n501, ZN
                           => n498);
   U484 : AOI22_X1 port map( A1 => n505, A2 => n82, B1 => n498, B2 => n502, ZN 
                           => n785);
   U485 : AOI22_X1 port map( A1 => n500, A2 => n1, B1 => n2, B2 => n501, ZN => 
                           n499);
   U486 : AOI22_X1 port map( A1 => n505, A2 => n90, B1 => n499, B2 => n502, ZN 
                           => n784);
   U487 : AOI22_X1 port map( A1 => n827, A2 => n501, B1 => n500, B2 => n130, ZN
                           => n503);
   U488 : AOI22_X1 port map( A1 => n505, A2 => n504, B1 => n503, B2 => n502, ZN
                           => n783);
   U489 : NAND2_X1 port map( A1 => n815, A2 => n509, ZN => n510);
   U490 : OAI211_X1 port map( C1 => n799, C2 => n524, A => n131, B => n510, ZN 
                           => n511);
   U491 : INV_X1 port map( A => n511, ZN => n514);
   U492 : AOI22_X1 port map( A1 => n509, A2 => n819, B1 => n129, B2 => n510, ZN
                           => n507);
   U493 : AOI22_X1 port map( A1 => n514, A2 => n108, B1 => n507, B2 => n511, ZN
                           => n782);
   U494 : AOI22_X1 port map( A1 => n509, A2 => n1, B1 => n2, B2 => n510, ZN => 
                           n508);
   U495 : AOI22_X1 port map( A1 => n514, A2 => n114, B1 => n508, B2 => n511, ZN
                           => n781);
   U496 : AOI22_X1 port map( A1 => n827, A2 => n510, B1 => n509, B2 => n130, ZN
                           => n512);
   U497 : AOI22_X1 port map( A1 => n514, A2 => n513, B1 => n512, B2 => n511, ZN
                           => n780);
   U498 : NAND2_X1 port map( A1 => n815, A2 => n518, ZN => n519);
   U499 : OAI211_X1 port map( C1 => n807, C2 => n524, A => n132, B => n519, ZN 
                           => n520);
   U500 : INV_X1 port map( A => n520, ZN => n522);
   U501 : AOI22_X1 port map( A1 => n518, A2 => n819, B1 => n129, B2 => n519, ZN
                           => n516);
   U502 : AOI22_X1 port map( A1 => n522, A2 => n59, B1 => n516, B2 => n520, ZN 
                           => n779);
   U503 : AOI22_X1 port map( A1 => n518, A2 => n1, B1 => n2, B2 => n519, ZN => 
                           n517);
   U504 : AOI22_X1 port map( A1 => n522, A2 => n63, B1 => n517, B2 => n520, ZN 
                           => n778);
   U505 : AOI22_X1 port map( A1 => n827, A2 => n519, B1 => n518, B2 => n130, ZN
                           => n521);
   U506 : AOI22_X1 port map( A1 => n522, A2 => n50, B1 => n521, B2 => n520, ZN 
                           => n777);
   U507 : NAND2_X1 port map( A1 => n815, A2 => n527, ZN => n528);
   U508 : OAI211_X1 port map( C1 => n817, C2 => n524, A => n131, B => n528, ZN 
                           => n529);
   U509 : INV_X1 port map( A => n529, ZN => n531);
   U510 : AOI22_X1 port map( A1 => n527, A2 => n819, B1 => n129, B2 => n528, ZN
                           => n525);
   U511 : AOI22_X1 port map( A1 => n531, A2 => n85, B1 => n525, B2 => n529, ZN 
                           => n776);
   U512 : AOI22_X1 port map( A1 => n527, A2 => n1, B1 => n2, B2 => n528, ZN => 
                           n526);
   U513 : AOI22_X1 port map( A1 => n531, A2 => n30, B1 => n526, B2 => n529, ZN 
                           => n775);
   U514 : AOI22_X1 port map( A1 => n827, A2 => n528, B1 => n527, B2 => n130, ZN
                           => n530);
   U515 : AOI22_X1 port map( A1 => n531, A2 => n88, B1 => n530, B2 => n529, ZN 
                           => n774);
   U516 : NAND2_X1 port map( A1 => n532, A2 => n661, ZN => n588);
   U517 : NAND2_X1 port map( A1 => n128, A2 => n535, ZN => n536);
   U518 : OAI211_X1 port map( C1 => n663, C2 => n588, A => n132, B => n536, ZN 
                           => n537);
   U519 : INV_X1 port map( A => n537, ZN => n540);
   U520 : AOI22_X1 port map( A1 => n535, A2 => n819, B1 => n818, B2 => n536, ZN
                           => n533);
   U521 : AOI22_X1 port map( A1 => n540, A2 => n116, B1 => n533, B2 => n537, ZN
                           => n773);
   U522 : AOI22_X1 port map( A1 => n535, A2 => n1, B1 => n2, B2 => n536, ZN => 
                           n534);
   U523 : AOI22_X1 port map( A1 => n540, A2 => n121, B1 => n534, B2 => n537, ZN
                           => n772);
   U524 : AOI22_X1 port map( A1 => n827, A2 => n536, B1 => n535, B2 => n824, ZN
                           => n538);
   U525 : AOI22_X1 port map( A1 => n540, A2 => n539, B1 => n538, B2 => n537, ZN
                           => n771);
   U526 : NAND2_X1 port map( A1 => n815, A2 => n543, ZN => n544);
   U527 : OAI211_X1 port map( C1 => n671, C2 => n588, A => n132, B => n544, ZN 
                           => n545);
   U528 : INV_X1 port map( A => n545, ZN => n548);
   U529 : AOI22_X1 port map( A1 => n543, A2 => n819, B1 => n818, B2 => n544, ZN
                           => n541);
   U530 : AOI22_X1 port map( A1 => n548, A2 => n100, B1 => n541, B2 => n545, ZN
                           => n770);
   U531 : AOI22_X1 port map( A1 => n543, A2 => n1, B1 => n2, B2 => n544, ZN => 
                           n542);
   U532 : AOI22_X1 port map( A1 => n548, A2 => n10, B1 => n542, B2 => n545, ZN 
                           => n769);
   U533 : AOI22_X1 port map( A1 => n827, A2 => n544, B1 => n543, B2 => n130, ZN
                           => n546);
   U534 : AOI22_X1 port map( A1 => n548, A2 => n547, B1 => n546, B2 => n545, ZN
                           => n768);
   U535 : NAND2_X1 port map( A1 => n128, A2 => n551, ZN => n552);
   U536 : OAI211_X1 port map( C1 => n679, C2 => n588, A => n132, B => n552, ZN 
                           => n553);
   U537 : INV_X1 port map( A => n553, ZN => n555);
   U538 : AOI22_X1 port map( A1 => n551, A2 => n819, B1 => n818, B2 => n552, ZN
                           => n549);
   U539 : AOI22_X1 port map( A1 => n555, A2 => n84, B1 => n549, B2 => n553, ZN 
                           => n767);
   U540 : AOI22_X1 port map( A1 => n551, A2 => n1, B1 => n2, B2 => n552, ZN => 
                           n550);
   U541 : AOI22_X1 port map( A1 => n555, A2 => n32, B1 => n550, B2 => n553, ZN 
                           => n766);
   U542 : AOI22_X1 port map( A1 => n827, A2 => n552, B1 => n551, B2 => n824, ZN
                           => n554);
   U543 : AOI22_X1 port map( A1 => n555, A2 => n87, B1 => n554, B2 => n553, ZN 
                           => n765);
   U544 : NAND2_X1 port map( A1 => n128, A2 => n558, ZN => n559);
   U545 : OAI211_X1 port map( C1 => n687, C2 => n588, A => n132, B => n559, ZN 
                           => n560);
   U546 : INV_X1 port map( A => n560, ZN => n562);
   U547 : AOI22_X1 port map( A1 => n558, A2 => n819, B1 => n818, B2 => n559, ZN
                           => n556);
   U548 : AOI22_X1 port map( A1 => n562, A2 => n122, B1 => n556, B2 => n560, ZN
                           => n764);
   U549 : AOI22_X1 port map( A1 => n558, A2 => n1, B1 => n2, B2 => n559, ZN => 
                           n557);
   U550 : AOI22_X1 port map( A1 => n562, A2 => n124, B1 => n557, B2 => n560, ZN
                           => n763);
   U551 : AOI22_X1 port map( A1 => n827, A2 => n559, B1 => n558, B2 => n824, ZN
                           => n561);
   U552 : AOI22_X1 port map( A1 => n562, A2 => n111, B1 => n561, B2 => n560, ZN
                           => n762);
   U553 : NAND2_X1 port map( A1 => n128, A2 => n565, ZN => n566);
   U554 : OAI211_X1 port map( C1 => n695, C2 => n588, A => n132, B => n566, ZN 
                           => n567);
   U555 : INV_X1 port map( A => n567, ZN => n570);
   U556 : AOI22_X1 port map( A1 => n565, A2 => n819, B1 => n129, B2 => n566, ZN
                           => n563);
   U557 : AOI22_X1 port map( A1 => n570, A2 => n41, B1 => n563, B2 => n567, ZN 
                           => n761);
   U558 : AOI22_X1 port map( A1 => n565, A2 => n1, B1 => n2, B2 => n566, ZN => 
                           n564);
   U559 : AOI22_X1 port map( A1 => n570, A2 => n106, B1 => n564, B2 => n567, ZN
                           => n760);
   U560 : AOI22_X1 port map( A1 => n827, A2 => n566, B1 => n565, B2 => n130, ZN
                           => n568);
   U561 : AOI22_X1 port map( A1 => n570, A2 => n569, B1 => n568, B2 => n567, ZN
                           => n759);
   U562 : NAND2_X1 port map( A1 => n128, A2 => n575, ZN => n576);
   U563 : OAI211_X1 port map( C1 => n799, C2 => n588, A => n132, B => n576, ZN 
                           => n577);
   U564 : INV_X1 port map( A => n577, ZN => n579);
   U565 : AOI22_X1 port map( A1 => n575, A2 => n819, B1 => n129, B2 => n576, ZN
                           => n571);
   U566 : AOI22_X1 port map( A1 => n579, A2 => n572, B1 => n571, B2 => n577, ZN
                           => n758);
   U567 : AOI22_X1 port map( A1 => n575, A2 => n1, B1 => n2, B2 => n576, ZN => 
                           n573);
   U568 : AOI22_X1 port map( A1 => n579, A2 => n574, B1 => n573, B2 => n577, ZN
                           => n757);
   U569 : AOI22_X1 port map( A1 => n827, A2 => n576, B1 => n575, B2 => n130, ZN
                           => n578);
   U570 : AOI22_X1 port map( A1 => n579, A2 => n53, B1 => n578, B2 => n577, ZN 
                           => n756);
   U571 : NAND2_X1 port map( A1 => n128, A2 => n582, ZN => n583);
   U572 : OAI211_X1 port map( C1 => n807, C2 => n588, A => n132, B => n583, ZN 
                           => n584);
   U573 : INV_X1 port map( A => n584, ZN => n587);
   U574 : AOI22_X1 port map( A1 => n582, A2 => n819, B1 => n129, B2 => n583, ZN
                           => n580);
   U575 : AOI22_X1 port map( A1 => n587, A2 => n60, B1 => n580, B2 => n584, ZN 
                           => n755);
   U576 : AOI22_X1 port map( A1 => n582, A2 => n1, B1 => n2, B2 => n583, ZN => 
                           n581);
   U577 : AOI22_X1 port map( A1 => n587, A2 => n91, B1 => n581, B2 => n584, ZN 
                           => n754);
   U578 : AOI22_X1 port map( A1 => n827, A2 => n583, B1 => n582, B2 => n130, ZN
                           => n585);
   U579 : AOI22_X1 port map( A1 => n587, A2 => n586, B1 => n585, B2 => n584, ZN
                           => n753);
   U580 : NAND2_X1 port map( A1 => n128, A2 => n591, ZN => n592);
   U581 : OAI211_X1 port map( C1 => n817, C2 => n588, A => n132, B => n592, ZN 
                           => n593);
   U582 : INV_X1 port map( A => n593, ZN => n595);
   U583 : AOI22_X1 port map( A1 => n591, A2 => n819, B1 => n129, B2 => n592, ZN
                           => n589);
   U584 : AOI22_X1 port map( A1 => n591, A2 => n1, B1 => n2, B2 => n592, ZN => 
                           n590);
   U585 : AOI22_X1 port map( A1 => n827, A2 => n592, B1 => n591, B2 => n130, ZN
                           => n594);
   U586 : NAND2_X1 port map( A1 => n596, A2 => n661, ZN => n652);
   U587 : NAND2_X1 port map( A1 => n815, A2 => n599, ZN => n600);
   U588 : OAI211_X1 port map( C1 => n663, C2 => n652, A => n132, B => n600, ZN 
                           => n601);
   U589 : INV_X1 port map( A => n601, ZN => n604);
   U590 : AOI22_X1 port map( A1 => n599, A2 => n819, B1 => n129, B2 => n600, ZN
                           => n597);
   U591 : AOI22_X1 port map( A1 => n604, A2 => n101, B1 => n597, B2 => n601, ZN
                           => n749);
   U592 : AOI22_X1 port map( A1 => n599, A2 => n1, B1 => n2, B2 => n600, ZN => 
                           n598);
   U593 : AOI22_X1 port map( A1 => n604, A2 => n3, B1 => n598, B2 => n601, ZN 
                           => n748);
   U594 : AOI22_X1 port map( A1 => n827, A2 => n600, B1 => n599, B2 => n130, ZN
                           => n602);
   U595 : AOI22_X1 port map( A1 => n604, A2 => n603, B1 => n602, B2 => n601, ZN
                           => n747);
   U596 : NAND2_X1 port map( A1 => n128, A2 => n609, ZN => n610);
   U597 : OAI211_X1 port map( C1 => n671, C2 => n652, A => n132, B => n610, ZN 
                           => n611);
   U598 : INV_X1 port map( A => n611, ZN => n614);
   U599 : AOI22_X1 port map( A1 => n609, A2 => n819, B1 => n129, B2 => n610, ZN
                           => n605);
   U600 : AOI22_X1 port map( A1 => n614, A2 => n606, B1 => n605, B2 => n611, ZN
                           => n746);
   U601 : AOI22_X1 port map( A1 => n609, A2 => n1, B1 => n2, B2 => n610, ZN => 
                           n607);
   U602 : AOI22_X1 port map( A1 => n614, A2 => n608, B1 => n607, B2 => n611, ZN
                           => n745);
   U603 : AOI22_X1 port map( A1 => n827, A2 => n610, B1 => n609, B2 => n130, ZN
                           => n612);
   U604 : AOI22_X1 port map( A1 => n614, A2 => n613, B1 => n612, B2 => n611, ZN
                           => n744);
   U605 : NAND2_X1 port map( A1 => n128, A2 => n617, ZN => n618);
   U606 : OAI211_X1 port map( C1 => n679, C2 => n652, A => n132, B => n618, ZN 
                           => n619);
   U607 : INV_X1 port map( A => n619, ZN => n622);
   U608 : AOI22_X1 port map( A1 => n617, A2 => n819, B1 => n129, B2 => n618, ZN
                           => n615);
   U609 : AOI22_X1 port map( A1 => n622, A2 => n83, B1 => n615, B2 => n619, ZN 
                           => n743);
   U610 : AOI22_X1 port map( A1 => n617, A2 => n1, B1 => n2, B2 => n618, ZN => 
                           n616);
   U611 : AOI22_X1 port map( A1 => n622, A2 => n92, B1 => n616, B2 => n619, ZN 
                           => n742);
   U612 : AOI22_X1 port map( A1 => n827, A2 => n618, B1 => n617, B2 => n130, ZN
                           => n620);
   U613 : AOI22_X1 port map( A1 => n622, A2 => n621, B1 => n620, B2 => n619, ZN
                           => n741);
   U614 : NAND2_X1 port map( A1 => n128, A2 => n625, ZN => n626);
   U615 : OAI211_X1 port map( C1 => n687, C2 => n652, A => n132, B => n626, ZN 
                           => n627);
   U616 : INV_X1 port map( A => n627, ZN => n629);
   U617 : AOI22_X1 port map( A1 => n625, A2 => n819, B1 => n129, B2 => n626, ZN
                           => n623);
   U618 : AOI22_X1 port map( A1 => n629, A2 => n123, B1 => n623, B2 => n627, ZN
                           => n740);
   U619 : AOI22_X1 port map( A1 => n625, A2 => n1, B1 => n2, B2 => n626, ZN => 
                           n624);
   U620 : AOI22_X1 port map( A1 => n629, A2 => n126, B1 => n624, B2 => n627, ZN
                           => n739);
   U621 : AOI22_X1 port map( A1 => n827, A2 => n626, B1 => n625, B2 => n130, ZN
                           => n628);
   U622 : AOI22_X1 port map( A1 => n629, A2 => n115, B1 => n628, B2 => n627, ZN
                           => n738);
   U623 : NAND2_X1 port map( A1 => n815, A2 => n632, ZN => n633);
   U624 : OAI211_X1 port map( C1 => n695, C2 => n652, A => n131, B => n633, ZN 
                           => n634);
   U625 : INV_X1 port map( A => n634, ZN => n637);
   U626 : AOI22_X1 port map( A1 => n632, A2 => n819, B1 => n129, B2 => n633, ZN
                           => n630);
   U627 : AOI22_X1 port map( A1 => n637, A2 => n19, B1 => n630, B2 => n634, ZN 
                           => n737);
   U628 : AOI22_X1 port map( A1 => n632, A2 => n1, B1 => n2, B2 => n633, ZN => 
                           n631);
   U629 : AOI22_X1 port map( A1 => n637, A2 => n86, B1 => n631, B2 => n634, ZN 
                           => n736);
   U630 : AOI22_X1 port map( A1 => n827, A2 => n633, B1 => n632, B2 => n130, ZN
                           => n635);
   U631 : AOI22_X1 port map( A1 => n637, A2 => n636, B1 => n635, B2 => n634, ZN
                           => n735);
   U632 : NAND2_X1 port map( A1 => n128, A2 => n640, ZN => n641);
   U633 : OAI211_X1 port map( C1 => n799, C2 => n652, A => n131, B => n641, ZN 
                           => n642);
   U634 : INV_X1 port map( A => n642, ZN => n644);
   U635 : AOI22_X1 port map( A1 => n640, A2 => n819, B1 => n129, B2 => n641, ZN
                           => n638);
   U636 : AOI22_X1 port map( A1 => n644, A2 => n17, B1 => n638, B2 => n642, ZN 
                           => n734);
   U637 : AOI22_X1 port map( A1 => n640, A2 => n1, B1 => n2, B2 => n641, ZN => 
                           n639);
   U638 : AOI22_X1 port map( A1 => n644, A2 => n125, B1 => n639, B2 => n642, ZN
                           => n733);
   U639 : AOI22_X1 port map( A1 => n827, A2 => n641, B1 => n640, B2 => n130, ZN
                           => n643);
   U640 : AOI22_X1 port map( A1 => n644, A2 => n113, B1 => n643, B2 => n642, ZN
                           => n732);
   U641 : NAND2_X1 port map( A1 => n128, A2 => n647, ZN => n648);
   U642 : OAI211_X1 port map( C1 => n807, C2 => n652, A => n131, B => n648, ZN 
                           => n649);
   U643 : INV_X1 port map( A => n649, ZN => n651);
   U644 : AOI22_X1 port map( A1 => n647, A2 => n819, B1 => n129, B2 => n648, ZN
                           => n645);
   U645 : AOI22_X1 port map( A1 => n651, A2 => n80, B1 => n645, B2 => n649, ZN 
                           => n731);
   U646 : AOI22_X1 port map( A1 => n647, A2 => n1, B1 => n2, B2 => n648, ZN => 
                           n646);
   U647 : AOI22_X1 port map( A1 => n651, A2 => n89, B1 => n646, B2 => n649, ZN 
                           => n730);
   U648 : AOI22_X1 port map( A1 => n827, A2 => n648, B1 => n647, B2 => n130, ZN
                           => n650);
   U649 : AOI22_X1 port map( A1 => n651, A2 => n49, B1 => n650, B2 => n649, ZN 
                           => n729);
   U650 : NAND2_X1 port map( A1 => n128, A2 => n655, ZN => n656);
   U651 : OAI211_X1 port map( C1 => n817, C2 => n652, A => n131, B => n656, ZN 
                           => n657);
   U652 : INV_X1 port map( A => n657, ZN => n660);
   U653 : AOI22_X1 port map( A1 => n655, A2 => n819, B1 => n129, B2 => n656, ZN
                           => n653);
   U654 : AOI22_X1 port map( A1 => n660, A2 => n105, B1 => n653, B2 => n657, ZN
                           => n728);
   U655 : AOI22_X1 port map( A1 => n655, A2 => n1, B1 => n2, B2 => n656, ZN => 
                           n654);
   U656 : AOI22_X1 port map( A1 => n660, A2 => n109, B1 => n654, B2 => n657, ZN
                           => n727);
   U657 : AOI22_X1 port map( A1 => n827, A2 => n656, B1 => n655, B2 => n130, ZN
                           => n658);
   U658 : AOI22_X1 port map( A1 => n660, A2 => n659, B1 => n658, B2 => n657, ZN
                           => n726);
   U659 : NAND2_X1 port map( A1 => n662, A2 => n661, ZN => n816);
   U660 : NAND2_X1 port map( A1 => n128, A2 => n666, ZN => n667);
   U661 : OAI211_X1 port map( C1 => n663, C2 => n816, A => n131, B => n667, ZN 
                           => n668);
   U662 : INV_X1 port map( A => n668, ZN => n670);
   U663 : AOI22_X1 port map( A1 => n666, A2 => n819, B1 => n818, B2 => n667, ZN
                           => n664);
   U664 : AOI22_X1 port map( A1 => n670, A2 => n27, B1 => n664, B2 => n668, ZN 
                           => n725);
   U665 : AOI22_X1 port map( A1 => n666, A2 => n1, B1 => n821, B2 => n667, ZN 
                           => n665);
   U666 : AOI22_X1 port map( A1 => n670, A2 => n34, B1 => n665, B2 => n668, ZN 
                           => n724);
   U667 : AOI22_X1 port map( A1 => n827, A2 => n667, B1 => n666, B2 => n824, ZN
                           => n669);
   U668 : AOI22_X1 port map( A1 => n670, A2 => n24, B1 => n669, B2 => n668, ZN 
                           => n723);
   U669 : NAND2_X1 port map( A1 => n128, A2 => n674, ZN => n675);
   U670 : OAI211_X1 port map( C1 => n671, C2 => n816, A => n131, B => n675, ZN 
                           => n676);
   U671 : INV_X1 port map( A => n676, ZN => n678);
   U672 : AOI22_X1 port map( A1 => n674, A2 => n819, B1 => n818, B2 => n675, ZN
                           => n672);
   U673 : AOI22_X1 port map( A1 => n678, A2 => n43, B1 => n672, B2 => n676, ZN 
                           => n722);
   U674 : AOI22_X1 port map( A1 => n674, A2 => n822, B1 => n821, B2 => n675, ZN
                           => n673);
   U675 : AOI22_X1 port map( A1 => n678, A2 => n42, B1 => n673, B2 => n676, ZN 
                           => n721);
   U676 : AOI22_X1 port map( A1 => n827, A2 => n675, B1 => n674, B2 => n824, ZN
                           => n677);
   U677 : AOI22_X1 port map( A1 => n678, A2 => n44, B1 => n677, B2 => n676, ZN 
                           => n720);
   U678 : NAND2_X1 port map( A1 => n128, A2 => n682, ZN => n683);
   U679 : OAI211_X1 port map( C1 => n679, C2 => n816, A => n131, B => n683, ZN 
                           => n684);
   U680 : INV_X1 port map( A => n684, ZN => n686);
   U681 : AOI22_X1 port map( A1 => n682, A2 => n819, B1 => n818, B2 => n683, ZN
                           => n680);
   U682 : AOI22_X1 port map( A1 => n686, A2 => n61, B1 => n680, B2 => n684, ZN 
                           => n719);
   U683 : AOI22_X1 port map( A1 => n682, A2 => n1, B1 => n821, B2 => n683, ZN 
                           => n681);
   U684 : AOI22_X1 port map( A1 => n686, A2 => n56, B1 => n681, B2 => n684, ZN 
                           => n718);
   U685 : AOI22_X1 port map( A1 => n827, A2 => n683, B1 => n682, B2 => n824, ZN
                           => n685);
   U686 : AOI22_X1 port map( A1 => n686, A2 => n64, B1 => n685, B2 => n684, ZN 
                           => n717);
   U687 : NAND2_X1 port map( A1 => n128, A2 => n690, ZN => n691);
   U688 : OAI211_X1 port map( C1 => n687, C2 => n816, A => n131, B => n691, ZN 
                           => n692);
   U689 : INV_X1 port map( A => n692, ZN => n694);
   U690 : AOI22_X1 port map( A1 => n690, A2 => n819, B1 => n818, B2 => n691, ZN
                           => n688);
   U691 : AOI22_X1 port map( A1 => n694, A2 => n47, B1 => n688, B2 => n692, ZN 
                           => n716);
   U692 : AOI22_X1 port map( A1 => n690, A2 => n822, B1 => n2, B2 => n691, ZN 
                           => n689);
   U693 : AOI22_X1 port map( A1 => n694, A2 => n45, B1 => n689, B2 => n692, ZN 
                           => n715);
   U694 : AOI22_X1 port map( A1 => n827, A2 => n691, B1 => n690, B2 => n824, ZN
                           => n693);
   U695 : AOI22_X1 port map( A1 => n694, A2 => n48, B1 => n693, B2 => n692, ZN 
                           => n714);
   U696 : NAND2_X1 port map( A1 => n128, A2 => n698, ZN => n699);
   U697 : OAI211_X1 port map( C1 => n695, C2 => n816, A => n131, B => n699, ZN 
                           => n700);
   U698 : INV_X1 port map( A => n700, ZN => n798);
   U699 : AOI22_X1 port map( A1 => n698, A2 => n819, B1 => n818, B2 => n699, ZN
                           => n696);
   U700 : AOI22_X1 port map( A1 => n798, A2 => n28, B1 => n696, B2 => n700, ZN 
                           => n713);
   U701 : AOI22_X1 port map( A1 => n698, A2 => n1, B1 => n2, B2 => n699, ZN => 
                           n697);
   U702 : AOI22_X1 port map( A1 => n798, A2 => n35, B1 => n697, B2 => n700, ZN 
                           => n712);
   U703 : AOI22_X1 port map( A1 => n827, A2 => n699, B1 => n698, B2 => n824, ZN
                           => n701);
   U704 : AOI22_X1 port map( A1 => n798, A2 => n25, B1 => n701, B2 => n700, ZN 
                           => n711);
   U705 : NAND2_X1 port map( A1 => n128, A2 => n802, ZN => n803);
   U706 : OAI211_X1 port map( C1 => n799, C2 => n816, A => n131, B => n803, ZN 
                           => n804);
   U707 : INV_X1 port map( A => n804, ZN => n806);
   U708 : AOI22_X1 port map( A1 => n802, A2 => n819, B1 => n818, B2 => n803, ZN
                           => n800);
   U709 : AOI22_X1 port map( A1 => n806, A2 => n52, B1 => n800, B2 => n804, ZN 
                           => n710);
   U710 : AOI22_X1 port map( A1 => n802, A2 => n822, B1 => n2, B2 => n803, ZN 
                           => n801);
   U711 : AOI22_X1 port map( A1 => n806, A2 => n54, B1 => n801, B2 => n804, ZN 
                           => n709);
   U712 : AOI22_X1 port map( A1 => n827, A2 => n803, B1 => n802, B2 => n130, ZN
                           => n805);
   U713 : AOI22_X1 port map( A1 => n806, A2 => n46, B1 => n805, B2 => n804, ZN 
                           => n708);
   U714 : NAND2_X1 port map( A1 => n128, A2 => n810, ZN => n811);
   U715 : OAI211_X1 port map( C1 => n807, C2 => n816, A => n131, B => n811, ZN 
                           => n812);
   U716 : INV_X1 port map( A => n812, ZN => n814);
   U717 : AOI22_X1 port map( A1 => n810, A2 => n819, B1 => n129, B2 => n811, ZN
                           => n808);
   U718 : AOI22_X1 port map( A1 => n814, A2 => n62, B1 => n808, B2 => n812, ZN 
                           => n707);
   U719 : AOI22_X1 port map( A1 => n810, A2 => n822, B1 => n2, B2 => n811, ZN 
                           => n809);
   U720 : AOI22_X1 port map( A1 => n814, A2 => n57, B1 => n809, B2 => n812, ZN 
                           => n706);
   U721 : AOI22_X1 port map( A1 => n827, A2 => n811, B1 => n810, B2 => n824, ZN
                           => n813);
   U722 : AOI22_X1 port map( A1 => n814, A2 => n65, B1 => n813, B2 => n812, ZN 
                           => n705);
   U723 : NAND2_X1 port map( A1 => n815, A2 => n825, ZN => n826);
   U724 : OAI211_X1 port map( C1 => n817, C2 => n816, A => n131, B => n826, ZN 
                           => n828);
   U725 : INV_X1 port map( A => n828, ZN => n830);
   U726 : AOI22_X1 port map( A1 => n825, A2 => n819, B1 => n818, B2 => n826, ZN
                           => n820);
   U727 : AOI22_X1 port map( A1 => n830, A2 => n29, B1 => n820, B2 => n828, ZN 
                           => n704);
   U728 : AOI22_X1 port map( A1 => n825, A2 => n1, B1 => n821, B2 => n826, ZN 
                           => n823);
   U729 : AOI22_X1 port map( A1 => n830, A2 => n26, B1 => n823, B2 => n828, ZN 
                           => n703);
   U730 : AOI22_X1 port map( A1 => n827, A2 => n826, B1 => n825, B2 => n824, ZN
                           => n829);
   U731 : AOI22_X1 port map( A1 => n830, A2 => n36, B1 => n829, B2 => n828, ZN 
                           => n702);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32.all;

entity DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ISSUE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ISSUE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA_IN : in 
         std_logic_vector (31 downto 0);  DRAM_DATA_OUT : out std_logic_vector 
         (31 downto 0);  DATA_SIZE : out std_logic_vector (1 downto 0);  
         DRAMRF_ADDRESS : out std_logic_vector (31 downto 0);  DRAMRF_ISSUE, 
         DRAMRF_READNOTWRITE : out std_logic;  DRAMRF_READY : in std_logic;  
         DRAMRF_DATA_IN : in std_logic_vector (31 downto 0);  DRAMRF_DATA_OUT :
         out std_logic_vector (31 downto 0);  DATA_SIZE_RF : out 
         std_logic_vector (1 downto 0));

end DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X4
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X2
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X2
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component select_block_NBIT_DATA32_N8_F5
      port( regs : in std_logic_vector (2559 downto 0);  win : in 
            std_logic_vector (4 downto 0);  curr_proc_regs : out 
            std_logic_vector (767 downto 0));
   end component;
   
   component mux_N32_M5_0
      port( S : in std_logic_vector (4 downto 0);  Q : in std_logic_vector 
            (1023 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component mux_N32_M5_1
      port( S : in std_logic_vector (4 downto 0);  Q : in std_logic_vector 
            (1023 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component in_loc_selblock_NBIT_DATA32_N8_F5
      port( regs : in std_logic_vector (2559 downto 0);  win : in 
            std_logic_vector (4 downto 0);  curr_proc_regs : out 
            std_logic_vector (511 downto 0));
   end component;
   
   component hazard_table_N_REGS_LOG5
      port( CLK, RST, WR1, WR2 : in std_logic;  ADD_WR1, ADD_WR2, ADD_CHECK1, 
            ADD_CHECK2 : in std_logic_vector (4 downto 0);  BUSY, BUSY_WINDOW :
            out std_logic);
   end component;
   
   signal IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, IRAM_ADDRESS_29_port, 
      IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, IRAM_ADDRESS_26_port, 
      IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, IRAM_ADDRESS_23_port, 
      IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_20_port, 
      IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, IRAM_ADDRESS_17_port, 
      IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, IRAM_ADDRESS_14_port, 
      IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, IRAM_ADDRESS_11_port, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, IRAM_ADDRESS_8_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port, DRAM_ADDRESS_31_port, 
      DRAM_ADDRESS_30_port, DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, 
      DRAM_ADDRESS_27_port, DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, 
      DRAM_ADDRESS_24_port, DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, 
      DRAM_ADDRESS_21_port, DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, 
      DRAM_ADDRESS_18_port, DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, 
      DRAM_ADDRESS_15_port, DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, 
      DRAM_ADDRESS_12_port, DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, 
      DRAM_ADDRESS_9_port, DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, 
      DRAM_ADDRESS_6_port, DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, 
      DRAM_ADDRESS_3_port, DRAM_ADDRESS_2_port, DRAM_ADDRESS_1_port, 
      DRAM_ADDRESS_0_port, DRAM_DATA_OUT_31_port, DRAM_DATA_OUT_30_port, 
      DRAM_DATA_OUT_29_port, DRAM_DATA_OUT_28_port, DRAM_DATA_OUT_27_port, 
      DRAM_DATA_OUT_26_port, DRAM_DATA_OUT_25_port, DRAM_DATA_OUT_24_port, 
      DRAM_DATA_OUT_23_port, DRAM_DATA_OUT_22_port, DRAM_DATA_OUT_21_port, 
      DRAM_DATA_OUT_20_port, DRAM_DATA_OUT_19_port, DRAM_DATA_OUT_18_port, 
      DRAM_DATA_OUT_17_port, DRAM_DATA_OUT_16_port, DRAM_DATA_OUT_15_port, 
      DRAM_DATA_OUT_14_port, DRAM_DATA_OUT_13_port, DRAM_DATA_OUT_12_port, 
      DRAM_DATA_OUT_11_port, DRAM_DATA_OUT_10_port, DRAM_DATA_OUT_9_port, 
      DRAM_DATA_OUT_8_port, DRAM_DATA_OUT_7_port, DRAM_DATA_OUT_6_port, 
      DRAM_DATA_OUT_5_port, DRAM_DATA_OUT_4_port, DRAM_DATA_OUT_3_port, 
      DRAM_DATA_OUT_2_port, DRAM_DATA_OUT_1_port, DRAM_DATA_OUT_0_port, 
      DATA_SIZE_1_port, DATA_SIZE_0_port, DRAMRF_ADDRESS_31_port, 
      DRAMRF_ADDRESS_30_port, DRAMRF_ADDRESS_29_port, DRAMRF_ADDRESS_28_port, 
      DRAMRF_ADDRESS_27_port, DRAMRF_ADDRESS_26_port, DRAMRF_ADDRESS_25_port, 
      DRAMRF_ADDRESS_24_port, DRAMRF_ADDRESS_23_port, DRAMRF_ADDRESS_22_port, 
      DRAMRF_ADDRESS_21_port, DRAMRF_ADDRESS_20_port, DRAMRF_ADDRESS_19_port, 
      DRAMRF_ADDRESS_18_port, DRAMRF_ADDRESS_17_port, DRAMRF_ADDRESS_16_port, 
      DRAMRF_ADDRESS_15_port, DRAMRF_ADDRESS_14_port, DRAMRF_ADDRESS_13_port, 
      DRAMRF_ADDRESS_12_port, DRAMRF_ADDRESS_11_port, DRAMRF_ADDRESS_10_port, 
      DRAMRF_ADDRESS_9_port, DRAMRF_ADDRESS_8_port, DRAMRF_ADDRESS_7_port, 
      DRAMRF_ADDRESS_6_port, DRAMRF_ADDRESS_5_port, DRAMRF_ADDRESS_4_port, 
      DRAMRF_ADDRESS_3_port, DRAMRF_ADDRESS_2_port, DRAMRF_ADDRESS_1_port, 
      DRAMRF_ADDRESS_0_port, DRAMRF_READNOTWRITE_port, i_DATAMEM_WM, IR_30_port
      , IR_26_port, IR_13_port, IR_10_port, IR_9_port, IR_8_port, IR_7_port, 
      IR_6_port, IR_5_port, IR_4_port, IR_3_port, IR_2_port, IR_1_port, 
      i_HAZARD_SIG_CU, i_BUSY_WINDOW, i_SEL_CMPB, i_NPC_SEL, i_S2, 
      i_ALU_OP_3_port, i_ALU_OP_2_port, i_ALU_OP_1_port, i_ALU_OP_0_port, 
      i_SEL_LGET_1_port, i_SEL_LGET_0_port, i_DATAMEM_RM, i_UNSIG_SIGN_N, i_WF,
      i_RF1, i_RF2, i_ADD_WB_4_port, i_ADD_WB_3_port, i_ADD_WB_2_port, 
      i_ADD_WB_1_port, i_ADD_WB_0_port, i_RD1_31_port, i_RD1_30_port, 
      i_RD1_29_port, i_RD1_28_port, i_RD1_27_port, i_RD1_26_port, i_RD1_25_port
      , i_RD1_24_port, i_RD1_23_port, i_RD1_22_port, i_RD1_21_port, 
      i_RD1_20_port, i_RD1_19_port, i_RD1_18_port, i_RD1_17_port, i_RD1_16_port
      , i_RD1_15_port, i_RD1_14_port, i_RD1_13_port, i_RD1_12_port, 
      i_RD1_11_port, i_RD1_10_port, i_RD1_9_port, i_RD1_8_port, i_RD1_7_port, 
      i_RD1_6_port, i_RD1_5_port, i_RD1_4_port, i_RD1_3_port, i_RD1_2_port, 
      i_RD1_1_port, i_RD1_0_port, i_RD2_31_port, i_RD2_30_port, i_RD2_29_port, 
      i_RD2_28_port, i_RD2_27_port, i_RD2_26_port, i_RD2_25_port, i_RD2_24_port
      , i_RD2_23_port, i_RD2_22_port, i_RD2_21_port, i_RD2_20_port, 
      i_RD2_19_port, i_RD2_18_port, i_RD2_17_port, i_RD2_16_port, i_RD2_15_port
      , i_RD2_14_port, i_RD2_13_port, i_RD2_12_port, i_RD2_11_port, 
      i_RD2_10_port, i_RD2_9_port, i_RD2_8_port, i_RD2_7_port, i_RD2_6_port, 
      i_RD2_5_port, i_RD2_4_port, i_RD2_3_port, i_RD2_2_port, i_RD2_1_port, 
      i_RD2_0_port, i_ADD_WS1_4_port, i_ADD_WS1_3_port, i_ADD_WS1_2_port, 
      i_ADD_WS1_1_port, i_ADD_WS1_0_port, CU_I_N184, CU_I_N171, CU_I_N170, 
      CU_I_i_SPILL_delay, CU_I_unsigned_1, CU_I_i_FILL_delay, 
      CU_I_CW_MEM_0_port, CU_I_CW_MEM_1_port, CU_I_CW_MEM_2_port, 
      CU_I_CW_EX_0_port, CU_I_CW_EX_1_port, CU_I_CW_EX_2_port, 
      CU_I_CW_EX_3_port, CU_I_CW_EX_4_port, CU_I_CW_EX_5_port, 
      CU_I_CW_EX_6_port, CU_I_CW_EX_18, CU_I_CW_ID_0_port, CU_I_CW_ID_1_port, 
      CU_I_CW_ID_2_port, CU_I_CW_ID_3_port, CU_I_CW_ID_4_port, 
      CU_I_CW_ID_5_port, CU_I_CW_ID_6_port, CU_I_CW_ID_16, CU_I_CW_ID_17, 
      CU_I_CW_ID_18, CU_I_CW_ID_19, CU_I_CW_ID_22, CU_I_CW_IF_0, CU_I_CW_3_port
      , CU_I_CW_4_port, CU_I_CW_5_port, CU_I_CW_6_port, CU_I_CW_16_port, 
      CU_I_CW_21_port, CU_I_CW_22_port, CU_I_CW_23_port, CU_I_CW_24_port, 
      CU_I_CW_25_port, DECODEhw_i_tickcounter_2_port, 
      DECODEhw_i_tickcounter_4_port, DECODEhw_i_tickcounter_6_port, 
      DECODEhw_i_tickcounter_8_port, DECODEhw_i_tickcounter_10_port, 
      DECODEhw_i_tickcounter_12_port, DECODEhw_i_tickcounter_14_port, 
      DECODEhw_i_tickcounter_16_port, DECODEhw_i_tickcounter_18_port, 
      DECODEhw_i_tickcounter_20_port, DECODEhw_i_tickcounter_22_port, 
      DECODEhw_i_tickcounter_24_port, DECODEhw_i_tickcounter_26_port, 
      DECODEhw_i_tickcounter_29_port, DECODEhw_i_tickcounter_31_port, 
      DECODEhw_i_WR1, DataPath_i_PIPLIN_WRB2_0_port, 
      DataPath_i_PIPLIN_WRB2_1_port, DataPath_i_PIPLIN_WRB2_2_port, 
      DataPath_i_PIPLIN_WRB2_3_port, DataPath_i_PIPLIN_WRB2_4_port, 
      DataPath_i_PIPLIN_WRB1_0_port, DataPath_i_PIPLIN_WRB1_1_port, 
      DataPath_i_PIPLIN_WRB1_2_port, DataPath_i_PIPLIN_WRB1_3_port, 
      DataPath_i_PIPLIN_WRB1_4_port, DataPath_i_REG_MEM_ALUOUT_0_port, 
      DataPath_i_REG_MEM_ALUOUT_1_port, DataPath_i_REG_MEM_ALUOUT_2_port, 
      DataPath_i_REG_MEM_ALUOUT_3_port, DataPath_i_REG_MEM_ALUOUT_4_port, 
      DataPath_i_REG_MEM_ALUOUT_5_port, DataPath_i_REG_MEM_ALUOUT_6_port, 
      DataPath_i_REG_MEM_ALUOUT_7_port, DataPath_i_REG_MEM_ALUOUT_8_port, 
      DataPath_i_REG_MEM_ALUOUT_9_port, DataPath_i_REG_MEM_ALUOUT_10_port, 
      DataPath_i_REG_MEM_ALUOUT_11_port, DataPath_i_REG_MEM_ALUOUT_12_port, 
      DataPath_i_REG_MEM_ALUOUT_13_port, DataPath_i_REG_MEM_ALUOUT_14_port, 
      DataPath_i_REG_MEM_ALUOUT_15_port, DataPath_i_REG_MEM_ALUOUT_16_port, 
      DataPath_i_REG_MEM_ALUOUT_17_port, DataPath_i_REG_MEM_ALUOUT_18_port, 
      DataPath_i_REG_MEM_ALUOUT_19_port, DataPath_i_REG_MEM_ALUOUT_20_port, 
      DataPath_i_REG_MEM_ALUOUT_21_port, DataPath_i_REG_MEM_ALUOUT_22_port, 
      DataPath_i_REG_MEM_ALUOUT_23_port, DataPath_i_REG_MEM_ALUOUT_24_port, 
      DataPath_i_REG_MEM_ALUOUT_25_port, DataPath_i_REG_MEM_ALUOUT_26_port, 
      DataPath_i_REG_MEM_ALUOUT_27_port, DataPath_i_REG_MEM_ALUOUT_28_port, 
      DataPath_i_REG_MEM_ALUOUT_29_port, DataPath_i_REG_MEM_ALUOUT_30_port, 
      DataPath_i_REG_MEM_ALUOUT_31_port, DataPath_i_REG_LDSTR_OUT_0_port, 
      DataPath_i_REG_LDSTR_OUT_1_port, DataPath_i_REG_LDSTR_OUT_2_port, 
      DataPath_i_REG_LDSTR_OUT_3_port, DataPath_i_REG_LDSTR_OUT_4_port, 
      DataPath_i_REG_LDSTR_OUT_5_port, DataPath_i_REG_LDSTR_OUT_6_port, 
      DataPath_i_REG_LDSTR_OUT_7_port, DataPath_i_REG_LDSTR_OUT_8_port, 
      DataPath_i_REG_LDSTR_OUT_9_port, DataPath_i_REG_LDSTR_OUT_10_port, 
      DataPath_i_REG_LDSTR_OUT_11_port, DataPath_i_REG_LDSTR_OUT_12_port, 
      DataPath_i_REG_LDSTR_OUT_13_port, DataPath_i_REG_LDSTR_OUT_14_port, 
      DataPath_i_REG_LDSTR_OUT_15_port, DataPath_i_REG_LDSTR_OUT_16_port, 
      DataPath_i_REG_LDSTR_OUT_17_port, DataPath_i_REG_LDSTR_OUT_18_port, 
      DataPath_i_REG_LDSTR_OUT_19_port, DataPath_i_REG_LDSTR_OUT_20_port, 
      DataPath_i_REG_LDSTR_OUT_21_port, DataPath_i_REG_LDSTR_OUT_22_port, 
      DataPath_i_REG_LDSTR_OUT_23_port, DataPath_i_REG_LDSTR_OUT_24_port, 
      DataPath_i_REG_LDSTR_OUT_25_port, DataPath_i_REG_LDSTR_OUT_26_port, 
      DataPath_i_REG_LDSTR_OUT_27_port, DataPath_i_REG_LDSTR_OUT_28_port, 
      DataPath_i_REG_LDSTR_OUT_29_port, DataPath_i_REG_LDSTR_OUT_30_port, 
      DataPath_i_REG_LDSTR_OUT_31_port, DataPath_i_REG_ME_DATA_DATAMEM_0_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_1_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_2_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_3_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_4_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_5_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_6_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_7_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_8_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_9_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_10_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_11_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_12_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_13_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_14_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_15_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_16_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_17_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_18_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_19_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_20_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_21_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_22_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_23_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_24_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_25_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_26_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_27_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_28_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_29_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_30_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_31_port, DataPath_i_LGET_0_port, 
      DataPath_i_PIPLIN_IN2_0_port, DataPath_i_PIPLIN_IN2_1_port, 
      DataPath_i_PIPLIN_IN2_2_port, DataPath_i_PIPLIN_IN2_3_port, 
      DataPath_i_PIPLIN_IN2_4_port, DataPath_i_PIPLIN_IN2_5_port, 
      DataPath_i_PIPLIN_IN2_6_port, DataPath_i_PIPLIN_IN2_7_port, 
      DataPath_i_PIPLIN_IN2_8_port, DataPath_i_PIPLIN_IN2_9_port, 
      DataPath_i_PIPLIN_IN2_10_port, DataPath_i_PIPLIN_IN2_11_port, 
      DataPath_i_PIPLIN_IN2_12_port, DataPath_i_PIPLIN_IN2_13_port, 
      DataPath_i_PIPLIN_IN2_14_port, DataPath_i_PIPLIN_IN2_15_port, 
      DataPath_i_PIPLIN_IN2_16_port, DataPath_i_PIPLIN_IN2_17_port, 
      DataPath_i_PIPLIN_IN2_18_port, DataPath_i_PIPLIN_IN2_19_port, 
      DataPath_i_PIPLIN_IN2_20_port, DataPath_i_PIPLIN_IN2_21_port, 
      DataPath_i_PIPLIN_IN2_22_port, DataPath_i_PIPLIN_IN2_23_port, 
      DataPath_i_PIPLIN_IN2_24_port, DataPath_i_PIPLIN_IN2_25_port, 
      DataPath_i_PIPLIN_IN2_26_port, DataPath_i_PIPLIN_IN2_27_port, 
      DataPath_i_PIPLIN_IN2_28_port, DataPath_i_PIPLIN_IN2_29_port, 
      DataPath_i_PIPLIN_IN2_30_port, DataPath_i_PIPLIN_IN2_31_port, 
      DataPath_i_PIPLIN_IN1_0_port, DataPath_i_PIPLIN_IN1_1_port, 
      DataPath_i_PIPLIN_IN1_2_port, DataPath_i_PIPLIN_IN1_3_port, 
      DataPath_i_PIPLIN_IN1_4_port, DataPath_i_PIPLIN_IN1_5_port, 
      DataPath_i_PIPLIN_IN1_6_port, DataPath_i_PIPLIN_IN1_7_port, 
      DataPath_i_PIPLIN_IN1_8_port, DataPath_i_PIPLIN_IN1_9_port, 
      DataPath_i_PIPLIN_IN1_10_port, DataPath_i_PIPLIN_IN1_11_port, 
      DataPath_i_PIPLIN_IN1_12_port, DataPath_i_PIPLIN_IN1_13_port, 
      DataPath_i_PIPLIN_IN1_14_port, DataPath_i_PIPLIN_IN1_15_port, 
      DataPath_i_PIPLIN_B_0_port, DataPath_i_PIPLIN_B_1_port, 
      DataPath_i_PIPLIN_B_2_port, DataPath_i_PIPLIN_B_3_port, 
      DataPath_i_PIPLIN_B_4_port, DataPath_i_PIPLIN_B_5_port, 
      DataPath_i_PIPLIN_B_6_port, DataPath_i_PIPLIN_B_7_port, 
      DataPath_i_PIPLIN_B_8_port, DataPath_i_PIPLIN_B_9_port, 
      DataPath_i_PIPLIN_B_10_port, DataPath_i_PIPLIN_B_11_port, 
      DataPath_i_PIPLIN_B_12_port, DataPath_i_PIPLIN_B_13_port, 
      DataPath_i_PIPLIN_B_14_port, DataPath_i_PIPLIN_B_15_port, 
      DataPath_i_PIPLIN_B_16_port, DataPath_i_PIPLIN_B_17_port, 
      DataPath_i_PIPLIN_B_18_port, DataPath_i_PIPLIN_B_19_port, 
      DataPath_i_PIPLIN_B_20_port, DataPath_i_PIPLIN_B_21_port, 
      DataPath_i_PIPLIN_B_22_port, DataPath_i_PIPLIN_B_23_port, 
      DataPath_i_PIPLIN_B_24_port, DataPath_i_PIPLIN_B_25_port, 
      DataPath_i_PIPLIN_B_26_port, DataPath_i_PIPLIN_B_27_port, 
      DataPath_i_PIPLIN_B_28_port, DataPath_i_PIPLIN_B_29_port, 
      DataPath_i_PIPLIN_B_30_port, DataPath_i_PIPLIN_B_31_port, 
      DataPath_i_PIPLIN_A_0_port, DataPath_i_PIPLIN_A_1_port, 
      DataPath_i_PIPLIN_A_2_port, DataPath_i_PIPLIN_A_3_port, 
      DataPath_i_PIPLIN_A_4_port, DataPath_i_PIPLIN_A_5_port, 
      DataPath_i_PIPLIN_A_6_port, DataPath_i_PIPLIN_A_7_port, 
      DataPath_i_PIPLIN_A_8_port, DataPath_i_PIPLIN_A_9_port, 
      DataPath_i_PIPLIN_A_10_port, DataPath_i_PIPLIN_A_11_port, 
      DataPath_i_PIPLIN_A_12_port, DataPath_i_PIPLIN_A_13_port, 
      DataPath_i_PIPLIN_A_14_port, DataPath_i_PIPLIN_A_15_port, 
      DataPath_i_PIPLIN_A_16_port, DataPath_i_PIPLIN_A_17_port, 
      DataPath_i_PIPLIN_A_18_port, DataPath_i_PIPLIN_A_19_port, 
      DataPath_i_PIPLIN_A_20_port, DataPath_i_PIPLIN_A_21_port, 
      DataPath_i_PIPLIN_A_22_port, DataPath_i_PIPLIN_A_23_port, 
      DataPath_i_PIPLIN_A_24_port, DataPath_i_PIPLIN_A_25_port, 
      DataPath_i_PIPLIN_A_26_port, DataPath_i_PIPLIN_A_27_port, 
      DataPath_i_PIPLIN_A_28_port, DataPath_i_PIPLIN_A_29_port, 
      DataPath_i_PIPLIN_A_30_port, DataPath_i_PIPLIN_A_31_port, 
      DataPath_RF_bus_sel_savedwin_data_0_port, 
      DataPath_RF_bus_sel_savedwin_data_1_port, 
      DataPath_RF_bus_sel_savedwin_data_2_port, 
      DataPath_RF_bus_sel_savedwin_data_3_port, 
      DataPath_RF_bus_sel_savedwin_data_4_port, 
      DataPath_RF_bus_sel_savedwin_data_5_port, 
      DataPath_RF_bus_sel_savedwin_data_6_port, 
      DataPath_RF_bus_sel_savedwin_data_7_port, 
      DataPath_RF_bus_sel_savedwin_data_8_port, 
      DataPath_RF_bus_sel_savedwin_data_9_port, 
      DataPath_RF_bus_sel_savedwin_data_10_port, 
      DataPath_RF_bus_sel_savedwin_data_11_port, 
      DataPath_RF_bus_sel_savedwin_data_12_port, 
      DataPath_RF_bus_sel_savedwin_data_13_port, 
      DataPath_RF_bus_sel_savedwin_data_14_port, 
      DataPath_RF_bus_sel_savedwin_data_15_port, 
      DataPath_RF_bus_sel_savedwin_data_16_port, 
      DataPath_RF_bus_sel_savedwin_data_17_port, 
      DataPath_RF_bus_sel_savedwin_data_18_port, 
      DataPath_RF_bus_sel_savedwin_data_19_port, 
      DataPath_RF_bus_sel_savedwin_data_20_port, 
      DataPath_RF_bus_sel_savedwin_data_21_port, 
      DataPath_RF_bus_sel_savedwin_data_22_port, 
      DataPath_RF_bus_sel_savedwin_data_23_port, 
      DataPath_RF_bus_sel_savedwin_data_24_port, 
      DataPath_RF_bus_sel_savedwin_data_25_port, 
      DataPath_RF_bus_sel_savedwin_data_26_port, 
      DataPath_RF_bus_sel_savedwin_data_27_port, 
      DataPath_RF_bus_sel_savedwin_data_28_port, 
      DataPath_RF_bus_sel_savedwin_data_29_port, 
      DataPath_RF_bus_sel_savedwin_data_30_port, 
      DataPath_RF_bus_sel_savedwin_data_31_port, 
      DataPath_RF_bus_sel_savedwin_data_32_port, 
      DataPath_RF_bus_sel_savedwin_data_33_port, 
      DataPath_RF_bus_sel_savedwin_data_34_port, 
      DataPath_RF_bus_sel_savedwin_data_35_port, 
      DataPath_RF_bus_sel_savedwin_data_36_port, 
      DataPath_RF_bus_sel_savedwin_data_37_port, 
      DataPath_RF_bus_sel_savedwin_data_38_port, 
      DataPath_RF_bus_sel_savedwin_data_39_port, 
      DataPath_RF_bus_sel_savedwin_data_40_port, 
      DataPath_RF_bus_sel_savedwin_data_41_port, 
      DataPath_RF_bus_sel_savedwin_data_42_port, 
      DataPath_RF_bus_sel_savedwin_data_43_port, 
      DataPath_RF_bus_sel_savedwin_data_44_port, 
      DataPath_RF_bus_sel_savedwin_data_45_port, 
      DataPath_RF_bus_sel_savedwin_data_46_port, 
      DataPath_RF_bus_sel_savedwin_data_47_port, 
      DataPath_RF_bus_sel_savedwin_data_48_port, 
      DataPath_RF_bus_sel_savedwin_data_49_port, 
      DataPath_RF_bus_sel_savedwin_data_50_port, 
      DataPath_RF_bus_sel_savedwin_data_51_port, 
      DataPath_RF_bus_sel_savedwin_data_52_port, 
      DataPath_RF_bus_sel_savedwin_data_53_port, 
      DataPath_RF_bus_sel_savedwin_data_54_port, 
      DataPath_RF_bus_sel_savedwin_data_55_port, 
      DataPath_RF_bus_sel_savedwin_data_56_port, 
      DataPath_RF_bus_sel_savedwin_data_57_port, 
      DataPath_RF_bus_sel_savedwin_data_58_port, 
      DataPath_RF_bus_sel_savedwin_data_59_port, 
      DataPath_RF_bus_sel_savedwin_data_60_port, 
      DataPath_RF_bus_sel_savedwin_data_61_port, 
      DataPath_RF_bus_sel_savedwin_data_62_port, 
      DataPath_RF_bus_sel_savedwin_data_63_port, 
      DataPath_RF_bus_sel_savedwin_data_64_port, 
      DataPath_RF_bus_sel_savedwin_data_65_port, 
      DataPath_RF_bus_sel_savedwin_data_66_port, 
      DataPath_RF_bus_sel_savedwin_data_67_port, 
      DataPath_RF_bus_sel_savedwin_data_68_port, 
      DataPath_RF_bus_sel_savedwin_data_69_port, 
      DataPath_RF_bus_sel_savedwin_data_70_port, 
      DataPath_RF_bus_sel_savedwin_data_71_port, 
      DataPath_RF_bus_sel_savedwin_data_72_port, 
      DataPath_RF_bus_sel_savedwin_data_73_port, 
      DataPath_RF_bus_sel_savedwin_data_74_port, 
      DataPath_RF_bus_sel_savedwin_data_75_port, 
      DataPath_RF_bus_sel_savedwin_data_76_port, 
      DataPath_RF_bus_sel_savedwin_data_77_port, 
      DataPath_RF_bus_sel_savedwin_data_78_port, 
      DataPath_RF_bus_sel_savedwin_data_79_port, 
      DataPath_RF_bus_sel_savedwin_data_80_port, 
      DataPath_RF_bus_sel_savedwin_data_81_port, 
      DataPath_RF_bus_sel_savedwin_data_82_port, 
      DataPath_RF_bus_sel_savedwin_data_83_port, 
      DataPath_RF_bus_sel_savedwin_data_84_port, 
      DataPath_RF_bus_sel_savedwin_data_85_port, 
      DataPath_RF_bus_sel_savedwin_data_86_port, 
      DataPath_RF_bus_sel_savedwin_data_87_port, 
      DataPath_RF_bus_sel_savedwin_data_88_port, 
      DataPath_RF_bus_sel_savedwin_data_89_port, 
      DataPath_RF_bus_sel_savedwin_data_90_port, 
      DataPath_RF_bus_sel_savedwin_data_91_port, 
      DataPath_RF_bus_sel_savedwin_data_92_port, 
      DataPath_RF_bus_sel_savedwin_data_93_port, 
      DataPath_RF_bus_sel_savedwin_data_94_port, 
      DataPath_RF_bus_sel_savedwin_data_95_port, 
      DataPath_RF_bus_sel_savedwin_data_96_port, 
      DataPath_RF_bus_sel_savedwin_data_97_port, 
      DataPath_RF_bus_sel_savedwin_data_98_port, 
      DataPath_RF_bus_sel_savedwin_data_99_port, 
      DataPath_RF_bus_sel_savedwin_data_100_port, 
      DataPath_RF_bus_sel_savedwin_data_101_port, 
      DataPath_RF_bus_sel_savedwin_data_102_port, 
      DataPath_RF_bus_sel_savedwin_data_103_port, 
      DataPath_RF_bus_sel_savedwin_data_104_port, 
      DataPath_RF_bus_sel_savedwin_data_105_port, 
      DataPath_RF_bus_sel_savedwin_data_106_port, 
      DataPath_RF_bus_sel_savedwin_data_107_port, 
      DataPath_RF_bus_sel_savedwin_data_108_port, 
      DataPath_RF_bus_sel_savedwin_data_109_port, 
      DataPath_RF_bus_sel_savedwin_data_110_port, 
      DataPath_RF_bus_sel_savedwin_data_111_port, 
      DataPath_RF_bus_sel_savedwin_data_112_port, 
      DataPath_RF_bus_sel_savedwin_data_113_port, 
      DataPath_RF_bus_sel_savedwin_data_114_port, 
      DataPath_RF_bus_sel_savedwin_data_115_port, 
      DataPath_RF_bus_sel_savedwin_data_116_port, 
      DataPath_RF_bus_sel_savedwin_data_117_port, 
      DataPath_RF_bus_sel_savedwin_data_118_port, 
      DataPath_RF_bus_sel_savedwin_data_119_port, 
      DataPath_RF_bus_sel_savedwin_data_120_port, 
      DataPath_RF_bus_sel_savedwin_data_121_port, 
      DataPath_RF_bus_sel_savedwin_data_122_port, 
      DataPath_RF_bus_sel_savedwin_data_123_port, 
      DataPath_RF_bus_sel_savedwin_data_124_port, 
      DataPath_RF_bus_sel_savedwin_data_125_port, 
      DataPath_RF_bus_sel_savedwin_data_126_port, 
      DataPath_RF_bus_sel_savedwin_data_127_port, 
      DataPath_RF_bus_sel_savedwin_data_128_port, 
      DataPath_RF_bus_sel_savedwin_data_129_port, 
      DataPath_RF_bus_sel_savedwin_data_130_port, 
      DataPath_RF_bus_sel_savedwin_data_131_port, 
      DataPath_RF_bus_sel_savedwin_data_132_port, 
      DataPath_RF_bus_sel_savedwin_data_133_port, 
      DataPath_RF_bus_sel_savedwin_data_134_port, 
      DataPath_RF_bus_sel_savedwin_data_135_port, 
      DataPath_RF_bus_sel_savedwin_data_136_port, 
      DataPath_RF_bus_sel_savedwin_data_137_port, 
      DataPath_RF_bus_sel_savedwin_data_138_port, 
      DataPath_RF_bus_sel_savedwin_data_139_port, 
      DataPath_RF_bus_sel_savedwin_data_140_port, 
      DataPath_RF_bus_sel_savedwin_data_141_port, 
      DataPath_RF_bus_sel_savedwin_data_142_port, 
      DataPath_RF_bus_sel_savedwin_data_143_port, 
      DataPath_RF_bus_sel_savedwin_data_144_port, 
      DataPath_RF_bus_sel_savedwin_data_145_port, 
      DataPath_RF_bus_sel_savedwin_data_146_port, 
      DataPath_RF_bus_sel_savedwin_data_147_port, 
      DataPath_RF_bus_sel_savedwin_data_148_port, 
      DataPath_RF_bus_sel_savedwin_data_149_port, 
      DataPath_RF_bus_sel_savedwin_data_150_port, 
      DataPath_RF_bus_sel_savedwin_data_151_port, 
      DataPath_RF_bus_sel_savedwin_data_152_port, 
      DataPath_RF_bus_sel_savedwin_data_153_port, 
      DataPath_RF_bus_sel_savedwin_data_154_port, 
      DataPath_RF_bus_sel_savedwin_data_155_port, 
      DataPath_RF_bus_sel_savedwin_data_156_port, 
      DataPath_RF_bus_sel_savedwin_data_157_port, 
      DataPath_RF_bus_sel_savedwin_data_158_port, 
      DataPath_RF_bus_sel_savedwin_data_159_port, 
      DataPath_RF_bus_sel_savedwin_data_160_port, 
      DataPath_RF_bus_sel_savedwin_data_161_port, 
      DataPath_RF_bus_sel_savedwin_data_162_port, 
      DataPath_RF_bus_sel_savedwin_data_163_port, 
      DataPath_RF_bus_sel_savedwin_data_164_port, 
      DataPath_RF_bus_sel_savedwin_data_165_port, 
      DataPath_RF_bus_sel_savedwin_data_166_port, 
      DataPath_RF_bus_sel_savedwin_data_167_port, 
      DataPath_RF_bus_sel_savedwin_data_168_port, 
      DataPath_RF_bus_sel_savedwin_data_169_port, 
      DataPath_RF_bus_sel_savedwin_data_170_port, 
      DataPath_RF_bus_sel_savedwin_data_171_port, 
      DataPath_RF_bus_sel_savedwin_data_172_port, 
      DataPath_RF_bus_sel_savedwin_data_173_port, 
      DataPath_RF_bus_sel_savedwin_data_174_port, 
      DataPath_RF_bus_sel_savedwin_data_175_port, 
      DataPath_RF_bus_sel_savedwin_data_176_port, 
      DataPath_RF_bus_sel_savedwin_data_177_port, 
      DataPath_RF_bus_sel_savedwin_data_178_port, 
      DataPath_RF_bus_sel_savedwin_data_179_port, 
      DataPath_RF_bus_sel_savedwin_data_180_port, 
      DataPath_RF_bus_sel_savedwin_data_181_port, 
      DataPath_RF_bus_sel_savedwin_data_182_port, 
      DataPath_RF_bus_sel_savedwin_data_183_port, 
      DataPath_RF_bus_sel_savedwin_data_184_port, 
      DataPath_RF_bus_sel_savedwin_data_185_port, 
      DataPath_RF_bus_sel_savedwin_data_186_port, 
      DataPath_RF_bus_sel_savedwin_data_187_port, 
      DataPath_RF_bus_sel_savedwin_data_188_port, 
      DataPath_RF_bus_sel_savedwin_data_189_port, 
      DataPath_RF_bus_sel_savedwin_data_190_port, 
      DataPath_RF_bus_sel_savedwin_data_191_port, 
      DataPath_RF_bus_sel_savedwin_data_192_port, 
      DataPath_RF_bus_sel_savedwin_data_193_port, 
      DataPath_RF_bus_sel_savedwin_data_194_port, 
      DataPath_RF_bus_sel_savedwin_data_195_port, 
      DataPath_RF_bus_sel_savedwin_data_196_port, 
      DataPath_RF_bus_sel_savedwin_data_197_port, 
      DataPath_RF_bus_sel_savedwin_data_198_port, 
      DataPath_RF_bus_sel_savedwin_data_199_port, 
      DataPath_RF_bus_sel_savedwin_data_200_port, 
      DataPath_RF_bus_sel_savedwin_data_201_port, 
      DataPath_RF_bus_sel_savedwin_data_202_port, 
      DataPath_RF_bus_sel_savedwin_data_203_port, 
      DataPath_RF_bus_sel_savedwin_data_204_port, 
      DataPath_RF_bus_sel_savedwin_data_205_port, 
      DataPath_RF_bus_sel_savedwin_data_206_port, 
      DataPath_RF_bus_sel_savedwin_data_207_port, 
      DataPath_RF_bus_sel_savedwin_data_208_port, 
      DataPath_RF_bus_sel_savedwin_data_209_port, 
      DataPath_RF_bus_sel_savedwin_data_210_port, 
      DataPath_RF_bus_sel_savedwin_data_211_port, 
      DataPath_RF_bus_sel_savedwin_data_212_port, 
      DataPath_RF_bus_sel_savedwin_data_213_port, 
      DataPath_RF_bus_sel_savedwin_data_214_port, 
      DataPath_RF_bus_sel_savedwin_data_215_port, 
      DataPath_RF_bus_sel_savedwin_data_216_port, 
      DataPath_RF_bus_sel_savedwin_data_217_port, 
      DataPath_RF_bus_sel_savedwin_data_218_port, 
      DataPath_RF_bus_sel_savedwin_data_219_port, 
      DataPath_RF_bus_sel_savedwin_data_220_port, 
      DataPath_RF_bus_sel_savedwin_data_221_port, 
      DataPath_RF_bus_sel_savedwin_data_222_port, 
      DataPath_RF_bus_sel_savedwin_data_223_port, 
      DataPath_RF_bus_sel_savedwin_data_224_port, 
      DataPath_RF_bus_sel_savedwin_data_225_port, 
      DataPath_RF_bus_sel_savedwin_data_226_port, 
      DataPath_RF_bus_sel_savedwin_data_227_port, 
      DataPath_RF_bus_sel_savedwin_data_228_port, 
      DataPath_RF_bus_sel_savedwin_data_229_port, 
      DataPath_RF_bus_sel_savedwin_data_230_port, 
      DataPath_RF_bus_sel_savedwin_data_231_port, 
      DataPath_RF_bus_sel_savedwin_data_232_port, 
      DataPath_RF_bus_sel_savedwin_data_233_port, 
      DataPath_RF_bus_sel_savedwin_data_234_port, 
      DataPath_RF_bus_sel_savedwin_data_235_port, 
      DataPath_RF_bus_sel_savedwin_data_236_port, 
      DataPath_RF_bus_sel_savedwin_data_237_port, 
      DataPath_RF_bus_sel_savedwin_data_238_port, 
      DataPath_RF_bus_sel_savedwin_data_239_port, 
      DataPath_RF_bus_sel_savedwin_data_240_port, 
      DataPath_RF_bus_sel_savedwin_data_241_port, 
      DataPath_RF_bus_sel_savedwin_data_242_port, 
      DataPath_RF_bus_sel_savedwin_data_243_port, 
      DataPath_RF_bus_sel_savedwin_data_244_port, 
      DataPath_RF_bus_sel_savedwin_data_245_port, 
      DataPath_RF_bus_sel_savedwin_data_246_port, 
      DataPath_RF_bus_sel_savedwin_data_247_port, 
      DataPath_RF_bus_sel_savedwin_data_248_port, 
      DataPath_RF_bus_sel_savedwin_data_249_port, 
      DataPath_RF_bus_sel_savedwin_data_250_port, 
      DataPath_RF_bus_sel_savedwin_data_251_port, 
      DataPath_RF_bus_sel_savedwin_data_252_port, 
      DataPath_RF_bus_sel_savedwin_data_253_port, 
      DataPath_RF_bus_sel_savedwin_data_254_port, 
      DataPath_RF_bus_sel_savedwin_data_255_port, 
      DataPath_RF_bus_sel_savedwin_data_256_port, 
      DataPath_RF_bus_sel_savedwin_data_257_port, 
      DataPath_RF_bus_sel_savedwin_data_258_port, 
      DataPath_RF_bus_sel_savedwin_data_259_port, 
      DataPath_RF_bus_sel_savedwin_data_260_port, 
      DataPath_RF_bus_sel_savedwin_data_261_port, 
      DataPath_RF_bus_sel_savedwin_data_262_port, 
      DataPath_RF_bus_sel_savedwin_data_263_port, 
      DataPath_RF_bus_sel_savedwin_data_264_port, 
      DataPath_RF_bus_sel_savedwin_data_265_port, 
      DataPath_RF_bus_sel_savedwin_data_266_port, 
      DataPath_RF_bus_sel_savedwin_data_267_port, 
      DataPath_RF_bus_sel_savedwin_data_268_port, 
      DataPath_RF_bus_sel_savedwin_data_269_port, 
      DataPath_RF_bus_sel_savedwin_data_270_port, 
      DataPath_RF_bus_sel_savedwin_data_271_port, 
      DataPath_RF_bus_sel_savedwin_data_272_port, 
      DataPath_RF_bus_sel_savedwin_data_273_port, 
      DataPath_RF_bus_sel_savedwin_data_274_port, 
      DataPath_RF_bus_sel_savedwin_data_275_port, 
      DataPath_RF_bus_sel_savedwin_data_276_port, 
      DataPath_RF_bus_sel_savedwin_data_277_port, 
      DataPath_RF_bus_sel_savedwin_data_278_port, 
      DataPath_RF_bus_sel_savedwin_data_279_port, 
      DataPath_RF_bus_sel_savedwin_data_280_port, 
      DataPath_RF_bus_sel_savedwin_data_281_port, 
      DataPath_RF_bus_sel_savedwin_data_282_port, 
      DataPath_RF_bus_sel_savedwin_data_283_port, 
      DataPath_RF_bus_sel_savedwin_data_284_port, 
      DataPath_RF_bus_sel_savedwin_data_285_port, 
      DataPath_RF_bus_sel_savedwin_data_286_port, 
      DataPath_RF_bus_sel_savedwin_data_287_port, 
      DataPath_RF_bus_sel_savedwin_data_288_port, 
      DataPath_RF_bus_sel_savedwin_data_289_port, 
      DataPath_RF_bus_sel_savedwin_data_290_port, 
      DataPath_RF_bus_sel_savedwin_data_291_port, 
      DataPath_RF_bus_sel_savedwin_data_292_port, 
      DataPath_RF_bus_sel_savedwin_data_293_port, 
      DataPath_RF_bus_sel_savedwin_data_294_port, 
      DataPath_RF_bus_sel_savedwin_data_295_port, 
      DataPath_RF_bus_sel_savedwin_data_296_port, 
      DataPath_RF_bus_sel_savedwin_data_297_port, 
      DataPath_RF_bus_sel_savedwin_data_298_port, 
      DataPath_RF_bus_sel_savedwin_data_299_port, 
      DataPath_RF_bus_sel_savedwin_data_300_port, 
      DataPath_RF_bus_sel_savedwin_data_301_port, 
      DataPath_RF_bus_sel_savedwin_data_302_port, 
      DataPath_RF_bus_sel_savedwin_data_303_port, 
      DataPath_RF_bus_sel_savedwin_data_304_port, 
      DataPath_RF_bus_sel_savedwin_data_305_port, 
      DataPath_RF_bus_sel_savedwin_data_306_port, 
      DataPath_RF_bus_sel_savedwin_data_307_port, 
      DataPath_RF_bus_sel_savedwin_data_308_port, 
      DataPath_RF_bus_sel_savedwin_data_309_port, 
      DataPath_RF_bus_sel_savedwin_data_310_port, 
      DataPath_RF_bus_sel_savedwin_data_311_port, 
      DataPath_RF_bus_sel_savedwin_data_312_port, 
      DataPath_RF_bus_sel_savedwin_data_313_port, 
      DataPath_RF_bus_sel_savedwin_data_314_port, 
      DataPath_RF_bus_sel_savedwin_data_315_port, 
      DataPath_RF_bus_sel_savedwin_data_316_port, 
      DataPath_RF_bus_sel_savedwin_data_317_port, 
      DataPath_RF_bus_sel_savedwin_data_318_port, 
      DataPath_RF_bus_sel_savedwin_data_319_port, 
      DataPath_RF_bus_sel_savedwin_data_320_port, 
      DataPath_RF_bus_sel_savedwin_data_321_port, 
      DataPath_RF_bus_sel_savedwin_data_322_port, 
      DataPath_RF_bus_sel_savedwin_data_323_port, 
      DataPath_RF_bus_sel_savedwin_data_324_port, 
      DataPath_RF_bus_sel_savedwin_data_325_port, 
      DataPath_RF_bus_sel_savedwin_data_326_port, 
      DataPath_RF_bus_sel_savedwin_data_327_port, 
      DataPath_RF_bus_sel_savedwin_data_328_port, 
      DataPath_RF_bus_sel_savedwin_data_329_port, 
      DataPath_RF_bus_sel_savedwin_data_330_port, 
      DataPath_RF_bus_sel_savedwin_data_331_port, 
      DataPath_RF_bus_sel_savedwin_data_332_port, 
      DataPath_RF_bus_sel_savedwin_data_333_port, 
      DataPath_RF_bus_sel_savedwin_data_334_port, 
      DataPath_RF_bus_sel_savedwin_data_335_port, 
      DataPath_RF_bus_sel_savedwin_data_336_port, 
      DataPath_RF_bus_sel_savedwin_data_337_port, 
      DataPath_RF_bus_sel_savedwin_data_338_port, 
      DataPath_RF_bus_sel_savedwin_data_339_port, 
      DataPath_RF_bus_sel_savedwin_data_340_port, 
      DataPath_RF_bus_sel_savedwin_data_341_port, 
      DataPath_RF_bus_sel_savedwin_data_342_port, 
      DataPath_RF_bus_sel_savedwin_data_343_port, 
      DataPath_RF_bus_sel_savedwin_data_344_port, 
      DataPath_RF_bus_sel_savedwin_data_345_port, 
      DataPath_RF_bus_sel_savedwin_data_346_port, 
      DataPath_RF_bus_sel_savedwin_data_347_port, 
      DataPath_RF_bus_sel_savedwin_data_348_port, 
      DataPath_RF_bus_sel_savedwin_data_349_port, 
      DataPath_RF_bus_sel_savedwin_data_350_port, 
      DataPath_RF_bus_sel_savedwin_data_351_port, 
      DataPath_RF_bus_sel_savedwin_data_352_port, 
      DataPath_RF_bus_sel_savedwin_data_353_port, 
      DataPath_RF_bus_sel_savedwin_data_354_port, 
      DataPath_RF_bus_sel_savedwin_data_355_port, 
      DataPath_RF_bus_sel_savedwin_data_356_port, 
      DataPath_RF_bus_sel_savedwin_data_357_port, 
      DataPath_RF_bus_sel_savedwin_data_358_port, 
      DataPath_RF_bus_sel_savedwin_data_359_port, 
      DataPath_RF_bus_sel_savedwin_data_360_port, 
      DataPath_RF_bus_sel_savedwin_data_361_port, 
      DataPath_RF_bus_sel_savedwin_data_362_port, 
      DataPath_RF_bus_sel_savedwin_data_363_port, 
      DataPath_RF_bus_sel_savedwin_data_364_port, 
      DataPath_RF_bus_sel_savedwin_data_365_port, 
      DataPath_RF_bus_sel_savedwin_data_366_port, 
      DataPath_RF_bus_sel_savedwin_data_367_port, 
      DataPath_RF_bus_sel_savedwin_data_368_port, 
      DataPath_RF_bus_sel_savedwin_data_369_port, 
      DataPath_RF_bus_sel_savedwin_data_370_port, 
      DataPath_RF_bus_sel_savedwin_data_371_port, 
      DataPath_RF_bus_sel_savedwin_data_372_port, 
      DataPath_RF_bus_sel_savedwin_data_373_port, 
      DataPath_RF_bus_sel_savedwin_data_374_port, 
      DataPath_RF_bus_sel_savedwin_data_375_port, 
      DataPath_RF_bus_sel_savedwin_data_376_port, 
      DataPath_RF_bus_sel_savedwin_data_377_port, 
      DataPath_RF_bus_sel_savedwin_data_378_port, 
      DataPath_RF_bus_sel_savedwin_data_379_port, 
      DataPath_RF_bus_sel_savedwin_data_380_port, 
      DataPath_RF_bus_sel_savedwin_data_381_port, 
      DataPath_RF_bus_sel_savedwin_data_382_port, 
      DataPath_RF_bus_sel_savedwin_data_383_port, 
      DataPath_RF_bus_sel_savedwin_data_384_port, 
      DataPath_RF_bus_sel_savedwin_data_385_port, 
      DataPath_RF_bus_sel_savedwin_data_386_port, 
      DataPath_RF_bus_sel_savedwin_data_387_port, 
      DataPath_RF_bus_sel_savedwin_data_388_port, 
      DataPath_RF_bus_sel_savedwin_data_389_port, 
      DataPath_RF_bus_sel_savedwin_data_390_port, 
      DataPath_RF_bus_sel_savedwin_data_391_port, 
      DataPath_RF_bus_sel_savedwin_data_392_port, 
      DataPath_RF_bus_sel_savedwin_data_393_port, 
      DataPath_RF_bus_sel_savedwin_data_394_port, 
      DataPath_RF_bus_sel_savedwin_data_395_port, 
      DataPath_RF_bus_sel_savedwin_data_396_port, 
      DataPath_RF_bus_sel_savedwin_data_397_port, 
      DataPath_RF_bus_sel_savedwin_data_398_port, 
      DataPath_RF_bus_sel_savedwin_data_399_port, 
      DataPath_RF_bus_sel_savedwin_data_400_port, 
      DataPath_RF_bus_sel_savedwin_data_401_port, 
      DataPath_RF_bus_sel_savedwin_data_402_port, 
      DataPath_RF_bus_sel_savedwin_data_403_port, 
      DataPath_RF_bus_sel_savedwin_data_404_port, 
      DataPath_RF_bus_sel_savedwin_data_405_port, 
      DataPath_RF_bus_sel_savedwin_data_406_port, 
      DataPath_RF_bus_sel_savedwin_data_407_port, 
      DataPath_RF_bus_sel_savedwin_data_408_port, 
      DataPath_RF_bus_sel_savedwin_data_409_port, 
      DataPath_RF_bus_sel_savedwin_data_410_port, 
      DataPath_RF_bus_sel_savedwin_data_411_port, 
      DataPath_RF_bus_sel_savedwin_data_412_port, 
      DataPath_RF_bus_sel_savedwin_data_413_port, 
      DataPath_RF_bus_sel_savedwin_data_414_port, 
      DataPath_RF_bus_sel_savedwin_data_415_port, 
      DataPath_RF_bus_sel_savedwin_data_416_port, 
      DataPath_RF_bus_sel_savedwin_data_417_port, 
      DataPath_RF_bus_sel_savedwin_data_418_port, 
      DataPath_RF_bus_sel_savedwin_data_419_port, 
      DataPath_RF_bus_sel_savedwin_data_420_port, 
      DataPath_RF_bus_sel_savedwin_data_421_port, 
      DataPath_RF_bus_sel_savedwin_data_422_port, 
      DataPath_RF_bus_sel_savedwin_data_423_port, 
      DataPath_RF_bus_sel_savedwin_data_424_port, 
      DataPath_RF_bus_sel_savedwin_data_425_port, 
      DataPath_RF_bus_sel_savedwin_data_426_port, 
      DataPath_RF_bus_sel_savedwin_data_427_port, 
      DataPath_RF_bus_sel_savedwin_data_428_port, 
      DataPath_RF_bus_sel_savedwin_data_429_port, 
      DataPath_RF_bus_sel_savedwin_data_430_port, 
      DataPath_RF_bus_sel_savedwin_data_431_port, 
      DataPath_RF_bus_sel_savedwin_data_432_port, 
      DataPath_RF_bus_sel_savedwin_data_433_port, 
      DataPath_RF_bus_sel_savedwin_data_434_port, 
      DataPath_RF_bus_sel_savedwin_data_435_port, 
      DataPath_RF_bus_sel_savedwin_data_436_port, 
      DataPath_RF_bus_sel_savedwin_data_437_port, 
      DataPath_RF_bus_sel_savedwin_data_438_port, 
      DataPath_RF_bus_sel_savedwin_data_439_port, 
      DataPath_RF_bus_sel_savedwin_data_440_port, 
      DataPath_RF_bus_sel_savedwin_data_441_port, 
      DataPath_RF_bus_sel_savedwin_data_442_port, 
      DataPath_RF_bus_sel_savedwin_data_443_port, 
      DataPath_RF_bus_sel_savedwin_data_444_port, 
      DataPath_RF_bus_sel_savedwin_data_445_port, 
      DataPath_RF_bus_sel_savedwin_data_446_port, 
      DataPath_RF_bus_sel_savedwin_data_447_port, 
      DataPath_RF_bus_sel_savedwin_data_448_port, 
      DataPath_RF_bus_sel_savedwin_data_449_port, 
      DataPath_RF_bus_sel_savedwin_data_450_port, 
      DataPath_RF_bus_sel_savedwin_data_451_port, 
      DataPath_RF_bus_sel_savedwin_data_452_port, 
      DataPath_RF_bus_sel_savedwin_data_453_port, 
      DataPath_RF_bus_sel_savedwin_data_454_port, 
      DataPath_RF_bus_sel_savedwin_data_455_port, 
      DataPath_RF_bus_sel_savedwin_data_456_port, 
      DataPath_RF_bus_sel_savedwin_data_457_port, 
      DataPath_RF_bus_sel_savedwin_data_458_port, 
      DataPath_RF_bus_sel_savedwin_data_459_port, 
      DataPath_RF_bus_sel_savedwin_data_460_port, 
      DataPath_RF_bus_sel_savedwin_data_461_port, 
      DataPath_RF_bus_sel_savedwin_data_462_port, 
      DataPath_RF_bus_sel_savedwin_data_463_port, 
      DataPath_RF_bus_sel_savedwin_data_464_port, 
      DataPath_RF_bus_sel_savedwin_data_465_port, 
      DataPath_RF_bus_sel_savedwin_data_466_port, 
      DataPath_RF_bus_sel_savedwin_data_467_port, 
      DataPath_RF_bus_sel_savedwin_data_468_port, 
      DataPath_RF_bus_sel_savedwin_data_469_port, 
      DataPath_RF_bus_sel_savedwin_data_470_port, 
      DataPath_RF_bus_sel_savedwin_data_471_port, 
      DataPath_RF_bus_sel_savedwin_data_472_port, 
      DataPath_RF_bus_sel_savedwin_data_473_port, 
      DataPath_RF_bus_sel_savedwin_data_474_port, 
      DataPath_RF_bus_sel_savedwin_data_475_port, 
      DataPath_RF_bus_sel_savedwin_data_476_port, 
      DataPath_RF_bus_sel_savedwin_data_477_port, 
      DataPath_RF_bus_sel_savedwin_data_478_port, 
      DataPath_RF_bus_sel_savedwin_data_479_port, 
      DataPath_RF_bus_sel_savedwin_data_480_port, 
      DataPath_RF_bus_sel_savedwin_data_481_port, 
      DataPath_RF_bus_sel_savedwin_data_482_port, 
      DataPath_RF_bus_sel_savedwin_data_483_port, 
      DataPath_RF_bus_sel_savedwin_data_484_port, 
      DataPath_RF_bus_sel_savedwin_data_485_port, 
      DataPath_RF_bus_sel_savedwin_data_486_port, 
      DataPath_RF_bus_sel_savedwin_data_487_port, 
      DataPath_RF_bus_sel_savedwin_data_488_port, 
      DataPath_RF_bus_sel_savedwin_data_489_port, 
      DataPath_RF_bus_sel_savedwin_data_490_port, 
      DataPath_RF_bus_sel_savedwin_data_491_port, 
      DataPath_RF_bus_sel_savedwin_data_492_port, 
      DataPath_RF_bus_sel_savedwin_data_493_port, 
      DataPath_RF_bus_sel_savedwin_data_494_port, 
      DataPath_RF_bus_sel_savedwin_data_495_port, 
      DataPath_RF_bus_sel_savedwin_data_496_port, 
      DataPath_RF_bus_sel_savedwin_data_497_port, 
      DataPath_RF_bus_sel_savedwin_data_498_port, 
      DataPath_RF_bus_sel_savedwin_data_499_port, 
      DataPath_RF_bus_sel_savedwin_data_500_port, 
      DataPath_RF_bus_sel_savedwin_data_501_port, 
      DataPath_RF_bus_sel_savedwin_data_502_port, 
      DataPath_RF_bus_sel_savedwin_data_503_port, 
      DataPath_RF_bus_sel_savedwin_data_504_port, 
      DataPath_RF_bus_sel_savedwin_data_505_port, 
      DataPath_RF_bus_sel_savedwin_data_506_port, 
      DataPath_RF_bus_sel_savedwin_data_507_port, 
      DataPath_RF_bus_sel_savedwin_data_508_port, 
      DataPath_RF_bus_sel_savedwin_data_509_port, 
      DataPath_RF_bus_sel_savedwin_data_510_port, 
      DataPath_RF_bus_sel_savedwin_data_511_port, DataPath_RF_c_swin_0_port, 
      DataPath_RF_c_swin_1_port, DataPath_RF_c_swin_2_port, 
      DataPath_RF_c_swin_3_port, DataPath_RF_c_swin_4_port, 
      DataPath_RF_internal_out2_0_port, DataPath_RF_internal_out2_1_port, 
      DataPath_RF_internal_out2_2_port, DataPath_RF_internal_out2_3_port, 
      DataPath_RF_internal_out2_4_port, DataPath_RF_internal_out2_5_port, 
      DataPath_RF_internal_out2_6_port, DataPath_RF_internal_out2_7_port, 
      DataPath_RF_internal_out2_8_port, DataPath_RF_internal_out2_9_port, 
      DataPath_RF_internal_out2_10_port, DataPath_RF_internal_out2_11_port, 
      DataPath_RF_internal_out2_12_port, DataPath_RF_internal_out2_13_port, 
      DataPath_RF_internal_out2_14_port, DataPath_RF_internal_out2_15_port, 
      DataPath_RF_internal_out2_16_port, DataPath_RF_internal_out2_17_port, 
      DataPath_RF_internal_out2_18_port, DataPath_RF_internal_out2_19_port, 
      DataPath_RF_internal_out2_20_port, DataPath_RF_internal_out2_21_port, 
      DataPath_RF_internal_out2_22_port, DataPath_RF_internal_out2_23_port, 
      DataPath_RF_internal_out2_24_port, DataPath_RF_internal_out2_25_port, 
      DataPath_RF_internal_out2_26_port, DataPath_RF_internal_out2_27_port, 
      DataPath_RF_internal_out2_28_port, DataPath_RF_internal_out2_29_port, 
      DataPath_RF_internal_out2_30_port, DataPath_RF_internal_out2_31_port, 
      DataPath_RF_internal_out1_0_port, DataPath_RF_internal_out1_1_port, 
      DataPath_RF_internal_out1_2_port, DataPath_RF_internal_out1_3_port, 
      DataPath_RF_internal_out1_4_port, DataPath_RF_internal_out1_5_port, 
      DataPath_RF_internal_out1_6_port, DataPath_RF_internal_out1_7_port, 
      DataPath_RF_internal_out1_8_port, DataPath_RF_internal_out1_9_port, 
      DataPath_RF_internal_out1_10_port, DataPath_RF_internal_out1_11_port, 
      DataPath_RF_internal_out1_12_port, DataPath_RF_internal_out1_13_port, 
      DataPath_RF_internal_out1_14_port, DataPath_RF_internal_out1_15_port, 
      DataPath_RF_internal_out1_16_port, DataPath_RF_internal_out1_17_port, 
      DataPath_RF_internal_out1_18_port, DataPath_RF_internal_out1_19_port, 
      DataPath_RF_internal_out1_20_port, DataPath_RF_internal_out1_21_port, 
      DataPath_RF_internal_out1_22_port, DataPath_RF_internal_out1_23_port, 
      DataPath_RF_internal_out1_24_port, DataPath_RF_internal_out1_25_port, 
      DataPath_RF_internal_out1_26_port, DataPath_RF_internal_out1_27_port, 
      DataPath_RF_internal_out1_28_port, DataPath_RF_internal_out1_29_port, 
      DataPath_RF_internal_out1_30_port, DataPath_RF_internal_out1_31_port, 
      DataPath_RF_bus_complete_win_data_0_port, 
      DataPath_RF_bus_complete_win_data_32_port, 
      DataPath_RF_bus_complete_win_data_33_port, 
      DataPath_RF_bus_complete_win_data_34_port, 
      DataPath_RF_bus_complete_win_data_35_port, 
      DataPath_RF_bus_complete_win_data_36_port, 
      DataPath_RF_bus_complete_win_data_37_port, 
      DataPath_RF_bus_complete_win_data_38_port, 
      DataPath_RF_bus_complete_win_data_39_port, 
      DataPath_RF_bus_complete_win_data_40_port, 
      DataPath_RF_bus_complete_win_data_41_port, 
      DataPath_RF_bus_complete_win_data_42_port, 
      DataPath_RF_bus_complete_win_data_43_port, 
      DataPath_RF_bus_complete_win_data_44_port, 
      DataPath_RF_bus_complete_win_data_45_port, 
      DataPath_RF_bus_complete_win_data_46_port, 
      DataPath_RF_bus_complete_win_data_47_port, 
      DataPath_RF_bus_complete_win_data_48_port, 
      DataPath_RF_bus_complete_win_data_49_port, 
      DataPath_RF_bus_complete_win_data_50_port, 
      DataPath_RF_bus_complete_win_data_51_port, 
      DataPath_RF_bus_complete_win_data_52_port, 
      DataPath_RF_bus_complete_win_data_53_port, 
      DataPath_RF_bus_complete_win_data_54_port, 
      DataPath_RF_bus_complete_win_data_55_port, 
      DataPath_RF_bus_complete_win_data_56_port, 
      DataPath_RF_bus_complete_win_data_57_port, 
      DataPath_RF_bus_complete_win_data_58_port, 
      DataPath_RF_bus_complete_win_data_59_port, 
      DataPath_RF_bus_complete_win_data_60_port, 
      DataPath_RF_bus_complete_win_data_61_port, 
      DataPath_RF_bus_complete_win_data_62_port, 
      DataPath_RF_bus_complete_win_data_63_port, 
      DataPath_RF_bus_complete_win_data_64_port, 
      DataPath_RF_bus_complete_win_data_65_port, 
      DataPath_RF_bus_complete_win_data_66_port, 
      DataPath_RF_bus_complete_win_data_67_port, 
      DataPath_RF_bus_complete_win_data_68_port, 
      DataPath_RF_bus_complete_win_data_69_port, 
      DataPath_RF_bus_complete_win_data_70_port, 
      DataPath_RF_bus_complete_win_data_71_port, 
      DataPath_RF_bus_complete_win_data_72_port, 
      DataPath_RF_bus_complete_win_data_73_port, 
      DataPath_RF_bus_complete_win_data_74_port, 
      DataPath_RF_bus_complete_win_data_75_port, 
      DataPath_RF_bus_complete_win_data_76_port, 
      DataPath_RF_bus_complete_win_data_77_port, 
      DataPath_RF_bus_complete_win_data_78_port, 
      DataPath_RF_bus_complete_win_data_79_port, 
      DataPath_RF_bus_complete_win_data_80_port, 
      DataPath_RF_bus_complete_win_data_81_port, 
      DataPath_RF_bus_complete_win_data_82_port, 
      DataPath_RF_bus_complete_win_data_83_port, 
      DataPath_RF_bus_complete_win_data_84_port, 
      DataPath_RF_bus_complete_win_data_85_port, 
      DataPath_RF_bus_complete_win_data_86_port, 
      DataPath_RF_bus_complete_win_data_87_port, 
      DataPath_RF_bus_complete_win_data_88_port, 
      DataPath_RF_bus_complete_win_data_89_port, 
      DataPath_RF_bus_complete_win_data_90_port, 
      DataPath_RF_bus_complete_win_data_91_port, 
      DataPath_RF_bus_complete_win_data_92_port, 
      DataPath_RF_bus_complete_win_data_93_port, 
      DataPath_RF_bus_complete_win_data_94_port, 
      DataPath_RF_bus_complete_win_data_95_port, 
      DataPath_RF_bus_complete_win_data_96_port, 
      DataPath_RF_bus_complete_win_data_97_port, 
      DataPath_RF_bus_complete_win_data_98_port, 
      DataPath_RF_bus_complete_win_data_99_port, 
      DataPath_RF_bus_complete_win_data_100_port, 
      DataPath_RF_bus_complete_win_data_101_port, 
      DataPath_RF_bus_complete_win_data_102_port, 
      DataPath_RF_bus_complete_win_data_103_port, 
      DataPath_RF_bus_complete_win_data_104_port, 
      DataPath_RF_bus_complete_win_data_105_port, 
      DataPath_RF_bus_complete_win_data_106_port, 
      DataPath_RF_bus_complete_win_data_107_port, 
      DataPath_RF_bus_complete_win_data_108_port, 
      DataPath_RF_bus_complete_win_data_109_port, 
      DataPath_RF_bus_complete_win_data_110_port, 
      DataPath_RF_bus_complete_win_data_111_port, 
      DataPath_RF_bus_complete_win_data_112_port, 
      DataPath_RF_bus_complete_win_data_113_port, 
      DataPath_RF_bus_complete_win_data_114_port, 
      DataPath_RF_bus_complete_win_data_115_port, 
      DataPath_RF_bus_complete_win_data_116_port, 
      DataPath_RF_bus_complete_win_data_117_port, 
      DataPath_RF_bus_complete_win_data_118_port, 
      DataPath_RF_bus_complete_win_data_119_port, 
      DataPath_RF_bus_complete_win_data_120_port, 
      DataPath_RF_bus_complete_win_data_121_port, 
      DataPath_RF_bus_complete_win_data_122_port, 
      DataPath_RF_bus_complete_win_data_123_port, 
      DataPath_RF_bus_complete_win_data_124_port, 
      DataPath_RF_bus_complete_win_data_125_port, 
      DataPath_RF_bus_complete_win_data_126_port, 
      DataPath_RF_bus_complete_win_data_127_port, 
      DataPath_RF_bus_complete_win_data_128_port, 
      DataPath_RF_bus_complete_win_data_129_port, 
      DataPath_RF_bus_complete_win_data_130_port, 
      DataPath_RF_bus_complete_win_data_131_port, 
      DataPath_RF_bus_complete_win_data_132_port, 
      DataPath_RF_bus_complete_win_data_133_port, 
      DataPath_RF_bus_complete_win_data_134_port, 
      DataPath_RF_bus_complete_win_data_135_port, 
      DataPath_RF_bus_complete_win_data_136_port, 
      DataPath_RF_bus_complete_win_data_137_port, 
      DataPath_RF_bus_complete_win_data_138_port, 
      DataPath_RF_bus_complete_win_data_139_port, 
      DataPath_RF_bus_complete_win_data_140_port, 
      DataPath_RF_bus_complete_win_data_141_port, 
      DataPath_RF_bus_complete_win_data_142_port, 
      DataPath_RF_bus_complete_win_data_143_port, 
      DataPath_RF_bus_complete_win_data_144_port, 
      DataPath_RF_bus_complete_win_data_145_port, 
      DataPath_RF_bus_complete_win_data_146_port, 
      DataPath_RF_bus_complete_win_data_147_port, 
      DataPath_RF_bus_complete_win_data_148_port, 
      DataPath_RF_bus_complete_win_data_149_port, 
      DataPath_RF_bus_complete_win_data_150_port, 
      DataPath_RF_bus_complete_win_data_151_port, 
      DataPath_RF_bus_complete_win_data_152_port, 
      DataPath_RF_bus_complete_win_data_153_port, 
      DataPath_RF_bus_complete_win_data_154_port, 
      DataPath_RF_bus_complete_win_data_155_port, 
      DataPath_RF_bus_complete_win_data_156_port, 
      DataPath_RF_bus_complete_win_data_157_port, 
      DataPath_RF_bus_complete_win_data_158_port, 
      DataPath_RF_bus_complete_win_data_159_port, 
      DataPath_RF_bus_complete_win_data_160_port, 
      DataPath_RF_bus_complete_win_data_161_port, 
      DataPath_RF_bus_complete_win_data_162_port, 
      DataPath_RF_bus_complete_win_data_163_port, 
      DataPath_RF_bus_complete_win_data_164_port, 
      DataPath_RF_bus_complete_win_data_165_port, 
      DataPath_RF_bus_complete_win_data_166_port, 
      DataPath_RF_bus_complete_win_data_167_port, 
      DataPath_RF_bus_complete_win_data_168_port, 
      DataPath_RF_bus_complete_win_data_169_port, 
      DataPath_RF_bus_complete_win_data_170_port, 
      DataPath_RF_bus_complete_win_data_171_port, 
      DataPath_RF_bus_complete_win_data_172_port, 
      DataPath_RF_bus_complete_win_data_173_port, 
      DataPath_RF_bus_complete_win_data_174_port, 
      DataPath_RF_bus_complete_win_data_175_port, 
      DataPath_RF_bus_complete_win_data_176_port, 
      DataPath_RF_bus_complete_win_data_177_port, 
      DataPath_RF_bus_complete_win_data_178_port, 
      DataPath_RF_bus_complete_win_data_179_port, 
      DataPath_RF_bus_complete_win_data_180_port, 
      DataPath_RF_bus_complete_win_data_181_port, 
      DataPath_RF_bus_complete_win_data_182_port, 
      DataPath_RF_bus_complete_win_data_183_port, 
      DataPath_RF_bus_complete_win_data_184_port, 
      DataPath_RF_bus_complete_win_data_185_port, 
      DataPath_RF_bus_complete_win_data_186_port, 
      DataPath_RF_bus_complete_win_data_187_port, 
      DataPath_RF_bus_complete_win_data_188_port, 
      DataPath_RF_bus_complete_win_data_189_port, 
      DataPath_RF_bus_complete_win_data_190_port, 
      DataPath_RF_bus_complete_win_data_191_port, 
      DataPath_RF_bus_complete_win_data_192_port, 
      DataPath_RF_bus_complete_win_data_193_port, 
      DataPath_RF_bus_complete_win_data_194_port, 
      DataPath_RF_bus_complete_win_data_195_port, 
      DataPath_RF_bus_complete_win_data_196_port, 
      DataPath_RF_bus_complete_win_data_197_port, 
      DataPath_RF_bus_complete_win_data_198_port, 
      DataPath_RF_bus_complete_win_data_199_port, 
      DataPath_RF_bus_complete_win_data_200_port, 
      DataPath_RF_bus_complete_win_data_201_port, 
      DataPath_RF_bus_complete_win_data_202_port, 
      DataPath_RF_bus_complete_win_data_203_port, 
      DataPath_RF_bus_complete_win_data_204_port, 
      DataPath_RF_bus_complete_win_data_205_port, 
      DataPath_RF_bus_complete_win_data_206_port, 
      DataPath_RF_bus_complete_win_data_207_port, 
      DataPath_RF_bus_complete_win_data_208_port, 
      DataPath_RF_bus_complete_win_data_209_port, 
      DataPath_RF_bus_complete_win_data_210_port, 
      DataPath_RF_bus_complete_win_data_211_port, 
      DataPath_RF_bus_complete_win_data_212_port, 
      DataPath_RF_bus_complete_win_data_213_port, 
      DataPath_RF_bus_complete_win_data_214_port, 
      DataPath_RF_bus_complete_win_data_215_port, 
      DataPath_RF_bus_complete_win_data_216_port, 
      DataPath_RF_bus_complete_win_data_217_port, 
      DataPath_RF_bus_complete_win_data_218_port, 
      DataPath_RF_bus_complete_win_data_219_port, 
      DataPath_RF_bus_complete_win_data_220_port, 
      DataPath_RF_bus_complete_win_data_221_port, 
      DataPath_RF_bus_complete_win_data_222_port, 
      DataPath_RF_bus_complete_win_data_223_port, 
      DataPath_RF_bus_complete_win_data_224_port, 
      DataPath_RF_bus_complete_win_data_225_port, 
      DataPath_RF_bus_complete_win_data_226_port, 
      DataPath_RF_bus_complete_win_data_227_port, 
      DataPath_RF_bus_complete_win_data_228_port, 
      DataPath_RF_bus_complete_win_data_229_port, 
      DataPath_RF_bus_complete_win_data_230_port, 
      DataPath_RF_bus_complete_win_data_231_port, 
      DataPath_RF_bus_complete_win_data_232_port, 
      DataPath_RF_bus_complete_win_data_233_port, 
      DataPath_RF_bus_complete_win_data_234_port, 
      DataPath_RF_bus_complete_win_data_235_port, 
      DataPath_RF_bus_complete_win_data_236_port, 
      DataPath_RF_bus_complete_win_data_237_port, 
      DataPath_RF_bus_complete_win_data_238_port, 
      DataPath_RF_bus_complete_win_data_239_port, 
      DataPath_RF_bus_complete_win_data_240_port, 
      DataPath_RF_bus_complete_win_data_241_port, 
      DataPath_RF_bus_complete_win_data_242_port, 
      DataPath_RF_bus_complete_win_data_243_port, 
      DataPath_RF_bus_complete_win_data_244_port, 
      DataPath_RF_bus_complete_win_data_245_port, 
      DataPath_RF_bus_complete_win_data_246_port, 
      DataPath_RF_bus_complete_win_data_247_port, 
      DataPath_RF_bus_complete_win_data_248_port, 
      DataPath_RF_bus_complete_win_data_249_port, 
      DataPath_RF_bus_complete_win_data_250_port, 
      DataPath_RF_bus_complete_win_data_251_port, 
      DataPath_RF_bus_complete_win_data_252_port, 
      DataPath_RF_bus_complete_win_data_253_port, 
      DataPath_RF_bus_complete_win_data_254_port, 
      DataPath_RF_bus_complete_win_data_255_port, 
      DataPath_RF_bus_selected_win_data_0_port, 
      DataPath_RF_bus_selected_win_data_1_port, 
      DataPath_RF_bus_selected_win_data_2_port, 
      DataPath_RF_bus_selected_win_data_3_port, 
      DataPath_RF_bus_selected_win_data_4_port, 
      DataPath_RF_bus_selected_win_data_5_port, 
      DataPath_RF_bus_selected_win_data_6_port, 
      DataPath_RF_bus_selected_win_data_7_port, 
      DataPath_RF_bus_selected_win_data_8_port, 
      DataPath_RF_bus_selected_win_data_9_port, 
      DataPath_RF_bus_selected_win_data_10_port, 
      DataPath_RF_bus_selected_win_data_11_port, 
      DataPath_RF_bus_selected_win_data_12_port, 
      DataPath_RF_bus_selected_win_data_13_port, 
      DataPath_RF_bus_selected_win_data_14_port, 
      DataPath_RF_bus_selected_win_data_15_port, 
      DataPath_RF_bus_selected_win_data_16_port, 
      DataPath_RF_bus_selected_win_data_17_port, 
      DataPath_RF_bus_selected_win_data_18_port, 
      DataPath_RF_bus_selected_win_data_19_port, 
      DataPath_RF_bus_selected_win_data_20_port, 
      DataPath_RF_bus_selected_win_data_21_port, 
      DataPath_RF_bus_selected_win_data_22_port, 
      DataPath_RF_bus_selected_win_data_23_port, 
      DataPath_RF_bus_selected_win_data_24_port, 
      DataPath_RF_bus_selected_win_data_25_port, 
      DataPath_RF_bus_selected_win_data_26_port, 
      DataPath_RF_bus_selected_win_data_27_port, 
      DataPath_RF_bus_selected_win_data_28_port, 
      DataPath_RF_bus_selected_win_data_29_port, 
      DataPath_RF_bus_selected_win_data_30_port, 
      DataPath_RF_bus_selected_win_data_31_port, 
      DataPath_RF_bus_selected_win_data_32_port, 
      DataPath_RF_bus_selected_win_data_33_port, 
      DataPath_RF_bus_selected_win_data_34_port, 
      DataPath_RF_bus_selected_win_data_35_port, 
      DataPath_RF_bus_selected_win_data_36_port, 
      DataPath_RF_bus_selected_win_data_37_port, 
      DataPath_RF_bus_selected_win_data_38_port, 
      DataPath_RF_bus_selected_win_data_39_port, 
      DataPath_RF_bus_selected_win_data_40_port, 
      DataPath_RF_bus_selected_win_data_41_port, 
      DataPath_RF_bus_selected_win_data_42_port, 
      DataPath_RF_bus_selected_win_data_43_port, 
      DataPath_RF_bus_selected_win_data_44_port, 
      DataPath_RF_bus_selected_win_data_45_port, 
      DataPath_RF_bus_selected_win_data_46_port, 
      DataPath_RF_bus_selected_win_data_47_port, 
      DataPath_RF_bus_selected_win_data_48_port, 
      DataPath_RF_bus_selected_win_data_49_port, 
      DataPath_RF_bus_selected_win_data_50_port, 
      DataPath_RF_bus_selected_win_data_51_port, 
      DataPath_RF_bus_selected_win_data_52_port, 
      DataPath_RF_bus_selected_win_data_53_port, 
      DataPath_RF_bus_selected_win_data_54_port, 
      DataPath_RF_bus_selected_win_data_55_port, 
      DataPath_RF_bus_selected_win_data_56_port, 
      DataPath_RF_bus_selected_win_data_57_port, 
      DataPath_RF_bus_selected_win_data_58_port, 
      DataPath_RF_bus_selected_win_data_59_port, 
      DataPath_RF_bus_selected_win_data_60_port, 
      DataPath_RF_bus_selected_win_data_61_port, 
      DataPath_RF_bus_selected_win_data_62_port, 
      DataPath_RF_bus_selected_win_data_63_port, 
      DataPath_RF_bus_selected_win_data_64_port, 
      DataPath_RF_bus_selected_win_data_65_port, 
      DataPath_RF_bus_selected_win_data_66_port, 
      DataPath_RF_bus_selected_win_data_67_port, 
      DataPath_RF_bus_selected_win_data_68_port, 
      DataPath_RF_bus_selected_win_data_69_port, 
      DataPath_RF_bus_selected_win_data_70_port, 
      DataPath_RF_bus_selected_win_data_71_port, 
      DataPath_RF_bus_selected_win_data_72_port, 
      DataPath_RF_bus_selected_win_data_73_port, 
      DataPath_RF_bus_selected_win_data_74_port, 
      DataPath_RF_bus_selected_win_data_75_port, 
      DataPath_RF_bus_selected_win_data_76_port, 
      DataPath_RF_bus_selected_win_data_77_port, 
      DataPath_RF_bus_selected_win_data_78_port, 
      DataPath_RF_bus_selected_win_data_79_port, 
      DataPath_RF_bus_selected_win_data_80_port, 
      DataPath_RF_bus_selected_win_data_81_port, 
      DataPath_RF_bus_selected_win_data_82_port, 
      DataPath_RF_bus_selected_win_data_83_port, 
      DataPath_RF_bus_selected_win_data_84_port, 
      DataPath_RF_bus_selected_win_data_85_port, 
      DataPath_RF_bus_selected_win_data_86_port, 
      DataPath_RF_bus_selected_win_data_87_port, 
      DataPath_RF_bus_selected_win_data_88_port, 
      DataPath_RF_bus_selected_win_data_89_port, 
      DataPath_RF_bus_selected_win_data_90_port, 
      DataPath_RF_bus_selected_win_data_91_port, 
      DataPath_RF_bus_selected_win_data_92_port, 
      DataPath_RF_bus_selected_win_data_93_port, 
      DataPath_RF_bus_selected_win_data_94_port, 
      DataPath_RF_bus_selected_win_data_95_port, 
      DataPath_RF_bus_selected_win_data_96_port, 
      DataPath_RF_bus_selected_win_data_97_port, 
      DataPath_RF_bus_selected_win_data_98_port, 
      DataPath_RF_bus_selected_win_data_99_port, 
      DataPath_RF_bus_selected_win_data_100_port, 
      DataPath_RF_bus_selected_win_data_101_port, 
      DataPath_RF_bus_selected_win_data_102_port, 
      DataPath_RF_bus_selected_win_data_103_port, 
      DataPath_RF_bus_selected_win_data_104_port, 
      DataPath_RF_bus_selected_win_data_105_port, 
      DataPath_RF_bus_selected_win_data_106_port, 
      DataPath_RF_bus_selected_win_data_107_port, 
      DataPath_RF_bus_selected_win_data_108_port, 
      DataPath_RF_bus_selected_win_data_109_port, 
      DataPath_RF_bus_selected_win_data_110_port, 
      DataPath_RF_bus_selected_win_data_111_port, 
      DataPath_RF_bus_selected_win_data_112_port, 
      DataPath_RF_bus_selected_win_data_113_port, 
      DataPath_RF_bus_selected_win_data_114_port, 
      DataPath_RF_bus_selected_win_data_115_port, 
      DataPath_RF_bus_selected_win_data_116_port, 
      DataPath_RF_bus_selected_win_data_117_port, 
      DataPath_RF_bus_selected_win_data_118_port, 
      DataPath_RF_bus_selected_win_data_119_port, 
      DataPath_RF_bus_selected_win_data_120_port, 
      DataPath_RF_bus_selected_win_data_121_port, 
      DataPath_RF_bus_selected_win_data_122_port, 
      DataPath_RF_bus_selected_win_data_123_port, 
      DataPath_RF_bus_selected_win_data_124_port, 
      DataPath_RF_bus_selected_win_data_125_port, 
      DataPath_RF_bus_selected_win_data_126_port, 
      DataPath_RF_bus_selected_win_data_127_port, 
      DataPath_RF_bus_selected_win_data_128_port, 
      DataPath_RF_bus_selected_win_data_129_port, 
      DataPath_RF_bus_selected_win_data_130_port, 
      DataPath_RF_bus_selected_win_data_131_port, 
      DataPath_RF_bus_selected_win_data_132_port, 
      DataPath_RF_bus_selected_win_data_133_port, 
      DataPath_RF_bus_selected_win_data_134_port, 
      DataPath_RF_bus_selected_win_data_135_port, 
      DataPath_RF_bus_selected_win_data_136_port, 
      DataPath_RF_bus_selected_win_data_137_port, 
      DataPath_RF_bus_selected_win_data_138_port, 
      DataPath_RF_bus_selected_win_data_139_port, 
      DataPath_RF_bus_selected_win_data_140_port, 
      DataPath_RF_bus_selected_win_data_141_port, 
      DataPath_RF_bus_selected_win_data_142_port, 
      DataPath_RF_bus_selected_win_data_143_port, 
      DataPath_RF_bus_selected_win_data_144_port, 
      DataPath_RF_bus_selected_win_data_145_port, 
      DataPath_RF_bus_selected_win_data_146_port, 
      DataPath_RF_bus_selected_win_data_147_port, 
      DataPath_RF_bus_selected_win_data_148_port, 
      DataPath_RF_bus_selected_win_data_149_port, 
      DataPath_RF_bus_selected_win_data_150_port, 
      DataPath_RF_bus_selected_win_data_151_port, 
      DataPath_RF_bus_selected_win_data_152_port, 
      DataPath_RF_bus_selected_win_data_153_port, 
      DataPath_RF_bus_selected_win_data_154_port, 
      DataPath_RF_bus_selected_win_data_155_port, 
      DataPath_RF_bus_selected_win_data_156_port, 
      DataPath_RF_bus_selected_win_data_157_port, 
      DataPath_RF_bus_selected_win_data_158_port, 
      DataPath_RF_bus_selected_win_data_159_port, 
      DataPath_RF_bus_selected_win_data_160_port, 
      DataPath_RF_bus_selected_win_data_161_port, 
      DataPath_RF_bus_selected_win_data_162_port, 
      DataPath_RF_bus_selected_win_data_163_port, 
      DataPath_RF_bus_selected_win_data_164_port, 
      DataPath_RF_bus_selected_win_data_165_port, 
      DataPath_RF_bus_selected_win_data_166_port, 
      DataPath_RF_bus_selected_win_data_167_port, 
      DataPath_RF_bus_selected_win_data_168_port, 
      DataPath_RF_bus_selected_win_data_169_port, 
      DataPath_RF_bus_selected_win_data_170_port, 
      DataPath_RF_bus_selected_win_data_171_port, 
      DataPath_RF_bus_selected_win_data_172_port, 
      DataPath_RF_bus_selected_win_data_173_port, 
      DataPath_RF_bus_selected_win_data_174_port, 
      DataPath_RF_bus_selected_win_data_175_port, 
      DataPath_RF_bus_selected_win_data_176_port, 
      DataPath_RF_bus_selected_win_data_177_port, 
      DataPath_RF_bus_selected_win_data_178_port, 
      DataPath_RF_bus_selected_win_data_179_port, 
      DataPath_RF_bus_selected_win_data_180_port, 
      DataPath_RF_bus_selected_win_data_181_port, 
      DataPath_RF_bus_selected_win_data_182_port, 
      DataPath_RF_bus_selected_win_data_183_port, 
      DataPath_RF_bus_selected_win_data_184_port, 
      DataPath_RF_bus_selected_win_data_185_port, 
      DataPath_RF_bus_selected_win_data_186_port, 
      DataPath_RF_bus_selected_win_data_187_port, 
      DataPath_RF_bus_selected_win_data_188_port, 
      DataPath_RF_bus_selected_win_data_189_port, 
      DataPath_RF_bus_selected_win_data_190_port, 
      DataPath_RF_bus_selected_win_data_191_port, 
      DataPath_RF_bus_selected_win_data_192_port, 
      DataPath_RF_bus_selected_win_data_193_port, 
      DataPath_RF_bus_selected_win_data_194_port, 
      DataPath_RF_bus_selected_win_data_195_port, 
      DataPath_RF_bus_selected_win_data_196_port, 
      DataPath_RF_bus_selected_win_data_197_port, 
      DataPath_RF_bus_selected_win_data_198_port, 
      DataPath_RF_bus_selected_win_data_199_port, 
      DataPath_RF_bus_selected_win_data_200_port, 
      DataPath_RF_bus_selected_win_data_201_port, 
      DataPath_RF_bus_selected_win_data_202_port, 
      DataPath_RF_bus_selected_win_data_203_port, 
      DataPath_RF_bus_selected_win_data_204_port, 
      DataPath_RF_bus_selected_win_data_205_port, 
      DataPath_RF_bus_selected_win_data_206_port, 
      DataPath_RF_bus_selected_win_data_207_port, 
      DataPath_RF_bus_selected_win_data_208_port, 
      DataPath_RF_bus_selected_win_data_209_port, 
      DataPath_RF_bus_selected_win_data_210_port, 
      DataPath_RF_bus_selected_win_data_211_port, 
      DataPath_RF_bus_selected_win_data_212_port, 
      DataPath_RF_bus_selected_win_data_213_port, 
      DataPath_RF_bus_selected_win_data_214_port, 
      DataPath_RF_bus_selected_win_data_215_port, 
      DataPath_RF_bus_selected_win_data_216_port, 
      DataPath_RF_bus_selected_win_data_217_port, 
      DataPath_RF_bus_selected_win_data_218_port, 
      DataPath_RF_bus_selected_win_data_219_port, 
      DataPath_RF_bus_selected_win_data_220_port, 
      DataPath_RF_bus_selected_win_data_221_port, 
      DataPath_RF_bus_selected_win_data_222_port, 
      DataPath_RF_bus_selected_win_data_223_port, 
      DataPath_RF_bus_selected_win_data_224_port, 
      DataPath_RF_bus_selected_win_data_225_port, 
      DataPath_RF_bus_selected_win_data_226_port, 
      DataPath_RF_bus_selected_win_data_227_port, 
      DataPath_RF_bus_selected_win_data_228_port, 
      DataPath_RF_bus_selected_win_data_229_port, 
      DataPath_RF_bus_selected_win_data_230_port, 
      DataPath_RF_bus_selected_win_data_231_port, 
      DataPath_RF_bus_selected_win_data_232_port, 
      DataPath_RF_bus_selected_win_data_233_port, 
      DataPath_RF_bus_selected_win_data_234_port, 
      DataPath_RF_bus_selected_win_data_235_port, 
      DataPath_RF_bus_selected_win_data_236_port, 
      DataPath_RF_bus_selected_win_data_237_port, 
      DataPath_RF_bus_selected_win_data_238_port, 
      DataPath_RF_bus_selected_win_data_239_port, 
      DataPath_RF_bus_selected_win_data_240_port, 
      DataPath_RF_bus_selected_win_data_241_port, 
      DataPath_RF_bus_selected_win_data_242_port, 
      DataPath_RF_bus_selected_win_data_243_port, 
      DataPath_RF_bus_selected_win_data_244_port, 
      DataPath_RF_bus_selected_win_data_245_port, 
      DataPath_RF_bus_selected_win_data_246_port, 
      DataPath_RF_bus_selected_win_data_247_port, 
      DataPath_RF_bus_selected_win_data_248_port, 
      DataPath_RF_bus_selected_win_data_249_port, 
      DataPath_RF_bus_selected_win_data_250_port, 
      DataPath_RF_bus_selected_win_data_251_port, 
      DataPath_RF_bus_selected_win_data_252_port, 
      DataPath_RF_bus_selected_win_data_253_port, 
      DataPath_RF_bus_selected_win_data_254_port, 
      DataPath_RF_bus_selected_win_data_255_port, 
      DataPath_RF_bus_selected_win_data_256_port, 
      DataPath_RF_bus_selected_win_data_257_port, 
      DataPath_RF_bus_selected_win_data_258_port, 
      DataPath_RF_bus_selected_win_data_259_port, 
      DataPath_RF_bus_selected_win_data_260_port, 
      DataPath_RF_bus_selected_win_data_261_port, 
      DataPath_RF_bus_selected_win_data_262_port, 
      DataPath_RF_bus_selected_win_data_263_port, 
      DataPath_RF_bus_selected_win_data_264_port, 
      DataPath_RF_bus_selected_win_data_265_port, 
      DataPath_RF_bus_selected_win_data_266_port, 
      DataPath_RF_bus_selected_win_data_267_port, 
      DataPath_RF_bus_selected_win_data_268_port, 
      DataPath_RF_bus_selected_win_data_269_port, 
      DataPath_RF_bus_selected_win_data_270_port, 
      DataPath_RF_bus_selected_win_data_271_port, 
      DataPath_RF_bus_selected_win_data_272_port, 
      DataPath_RF_bus_selected_win_data_273_port, 
      DataPath_RF_bus_selected_win_data_274_port, 
      DataPath_RF_bus_selected_win_data_275_port, 
      DataPath_RF_bus_selected_win_data_276_port, 
      DataPath_RF_bus_selected_win_data_277_port, 
      DataPath_RF_bus_selected_win_data_278_port, 
      DataPath_RF_bus_selected_win_data_279_port, 
      DataPath_RF_bus_selected_win_data_280_port, 
      DataPath_RF_bus_selected_win_data_281_port, 
      DataPath_RF_bus_selected_win_data_282_port, 
      DataPath_RF_bus_selected_win_data_283_port, 
      DataPath_RF_bus_selected_win_data_284_port, 
      DataPath_RF_bus_selected_win_data_285_port, 
      DataPath_RF_bus_selected_win_data_286_port, 
      DataPath_RF_bus_selected_win_data_287_port, 
      DataPath_RF_bus_selected_win_data_288_port, 
      DataPath_RF_bus_selected_win_data_289_port, 
      DataPath_RF_bus_selected_win_data_290_port, 
      DataPath_RF_bus_selected_win_data_291_port, 
      DataPath_RF_bus_selected_win_data_292_port, 
      DataPath_RF_bus_selected_win_data_293_port, 
      DataPath_RF_bus_selected_win_data_294_port, 
      DataPath_RF_bus_selected_win_data_295_port, 
      DataPath_RF_bus_selected_win_data_296_port, 
      DataPath_RF_bus_selected_win_data_297_port, 
      DataPath_RF_bus_selected_win_data_298_port, 
      DataPath_RF_bus_selected_win_data_299_port, 
      DataPath_RF_bus_selected_win_data_300_port, 
      DataPath_RF_bus_selected_win_data_301_port, 
      DataPath_RF_bus_selected_win_data_302_port, 
      DataPath_RF_bus_selected_win_data_303_port, 
      DataPath_RF_bus_selected_win_data_304_port, 
      DataPath_RF_bus_selected_win_data_305_port, 
      DataPath_RF_bus_selected_win_data_306_port, 
      DataPath_RF_bus_selected_win_data_307_port, 
      DataPath_RF_bus_selected_win_data_308_port, 
      DataPath_RF_bus_selected_win_data_309_port, 
      DataPath_RF_bus_selected_win_data_310_port, 
      DataPath_RF_bus_selected_win_data_311_port, 
      DataPath_RF_bus_selected_win_data_312_port, 
      DataPath_RF_bus_selected_win_data_313_port, 
      DataPath_RF_bus_selected_win_data_314_port, 
      DataPath_RF_bus_selected_win_data_315_port, 
      DataPath_RF_bus_selected_win_data_316_port, 
      DataPath_RF_bus_selected_win_data_317_port, 
      DataPath_RF_bus_selected_win_data_318_port, 
      DataPath_RF_bus_selected_win_data_319_port, 
      DataPath_RF_bus_selected_win_data_320_port, 
      DataPath_RF_bus_selected_win_data_321_port, 
      DataPath_RF_bus_selected_win_data_322_port, 
      DataPath_RF_bus_selected_win_data_323_port, 
      DataPath_RF_bus_selected_win_data_324_port, 
      DataPath_RF_bus_selected_win_data_325_port, 
      DataPath_RF_bus_selected_win_data_326_port, 
      DataPath_RF_bus_selected_win_data_327_port, 
      DataPath_RF_bus_selected_win_data_328_port, 
      DataPath_RF_bus_selected_win_data_329_port, 
      DataPath_RF_bus_selected_win_data_330_port, 
      DataPath_RF_bus_selected_win_data_331_port, 
      DataPath_RF_bus_selected_win_data_332_port, 
      DataPath_RF_bus_selected_win_data_333_port, 
      DataPath_RF_bus_selected_win_data_334_port, 
      DataPath_RF_bus_selected_win_data_335_port, 
      DataPath_RF_bus_selected_win_data_336_port, 
      DataPath_RF_bus_selected_win_data_337_port, 
      DataPath_RF_bus_selected_win_data_338_port, 
      DataPath_RF_bus_selected_win_data_339_port, 
      DataPath_RF_bus_selected_win_data_340_port, 
      DataPath_RF_bus_selected_win_data_341_port, 
      DataPath_RF_bus_selected_win_data_342_port, 
      DataPath_RF_bus_selected_win_data_343_port, 
      DataPath_RF_bus_selected_win_data_344_port, 
      DataPath_RF_bus_selected_win_data_345_port, 
      DataPath_RF_bus_selected_win_data_346_port, 
      DataPath_RF_bus_selected_win_data_347_port, 
      DataPath_RF_bus_selected_win_data_348_port, 
      DataPath_RF_bus_selected_win_data_349_port, 
      DataPath_RF_bus_selected_win_data_350_port, 
      DataPath_RF_bus_selected_win_data_351_port, 
      DataPath_RF_bus_selected_win_data_352_port, 
      DataPath_RF_bus_selected_win_data_353_port, 
      DataPath_RF_bus_selected_win_data_354_port, 
      DataPath_RF_bus_selected_win_data_355_port, 
      DataPath_RF_bus_selected_win_data_356_port, 
      DataPath_RF_bus_selected_win_data_357_port, 
      DataPath_RF_bus_selected_win_data_358_port, 
      DataPath_RF_bus_selected_win_data_359_port, 
      DataPath_RF_bus_selected_win_data_360_port, 
      DataPath_RF_bus_selected_win_data_361_port, 
      DataPath_RF_bus_selected_win_data_362_port, 
      DataPath_RF_bus_selected_win_data_363_port, 
      DataPath_RF_bus_selected_win_data_364_port, 
      DataPath_RF_bus_selected_win_data_365_port, 
      DataPath_RF_bus_selected_win_data_366_port, 
      DataPath_RF_bus_selected_win_data_367_port, 
      DataPath_RF_bus_selected_win_data_368_port, 
      DataPath_RF_bus_selected_win_data_369_port, 
      DataPath_RF_bus_selected_win_data_370_port, 
      DataPath_RF_bus_selected_win_data_371_port, 
      DataPath_RF_bus_selected_win_data_372_port, 
      DataPath_RF_bus_selected_win_data_373_port, 
      DataPath_RF_bus_selected_win_data_374_port, 
      DataPath_RF_bus_selected_win_data_375_port, 
      DataPath_RF_bus_selected_win_data_376_port, 
      DataPath_RF_bus_selected_win_data_377_port, 
      DataPath_RF_bus_selected_win_data_378_port, 
      DataPath_RF_bus_selected_win_data_379_port, 
      DataPath_RF_bus_selected_win_data_380_port, 
      DataPath_RF_bus_selected_win_data_381_port, 
      DataPath_RF_bus_selected_win_data_382_port, 
      DataPath_RF_bus_selected_win_data_383_port, 
      DataPath_RF_bus_selected_win_data_384_port, 
      DataPath_RF_bus_selected_win_data_385_port, 
      DataPath_RF_bus_selected_win_data_386_port, 
      DataPath_RF_bus_selected_win_data_387_port, 
      DataPath_RF_bus_selected_win_data_388_port, 
      DataPath_RF_bus_selected_win_data_389_port, 
      DataPath_RF_bus_selected_win_data_390_port, 
      DataPath_RF_bus_selected_win_data_391_port, 
      DataPath_RF_bus_selected_win_data_392_port, 
      DataPath_RF_bus_selected_win_data_393_port, 
      DataPath_RF_bus_selected_win_data_394_port, 
      DataPath_RF_bus_selected_win_data_395_port, 
      DataPath_RF_bus_selected_win_data_396_port, 
      DataPath_RF_bus_selected_win_data_397_port, 
      DataPath_RF_bus_selected_win_data_398_port, 
      DataPath_RF_bus_selected_win_data_399_port, 
      DataPath_RF_bus_selected_win_data_400_port, 
      DataPath_RF_bus_selected_win_data_401_port, 
      DataPath_RF_bus_selected_win_data_402_port, 
      DataPath_RF_bus_selected_win_data_403_port, 
      DataPath_RF_bus_selected_win_data_404_port, 
      DataPath_RF_bus_selected_win_data_405_port, 
      DataPath_RF_bus_selected_win_data_406_port, 
      DataPath_RF_bus_selected_win_data_407_port, 
      DataPath_RF_bus_selected_win_data_408_port, 
      DataPath_RF_bus_selected_win_data_409_port, 
      DataPath_RF_bus_selected_win_data_410_port, 
      DataPath_RF_bus_selected_win_data_411_port, 
      DataPath_RF_bus_selected_win_data_412_port, 
      DataPath_RF_bus_selected_win_data_413_port, 
      DataPath_RF_bus_selected_win_data_414_port, 
      DataPath_RF_bus_selected_win_data_415_port, 
      DataPath_RF_bus_selected_win_data_416_port, 
      DataPath_RF_bus_selected_win_data_417_port, 
      DataPath_RF_bus_selected_win_data_418_port, 
      DataPath_RF_bus_selected_win_data_419_port, 
      DataPath_RF_bus_selected_win_data_420_port, 
      DataPath_RF_bus_selected_win_data_421_port, 
      DataPath_RF_bus_selected_win_data_422_port, 
      DataPath_RF_bus_selected_win_data_423_port, 
      DataPath_RF_bus_selected_win_data_424_port, 
      DataPath_RF_bus_selected_win_data_425_port, 
      DataPath_RF_bus_selected_win_data_426_port, 
      DataPath_RF_bus_selected_win_data_427_port, 
      DataPath_RF_bus_selected_win_data_428_port, 
      DataPath_RF_bus_selected_win_data_429_port, 
      DataPath_RF_bus_selected_win_data_430_port, 
      DataPath_RF_bus_selected_win_data_431_port, 
      DataPath_RF_bus_selected_win_data_432_port, 
      DataPath_RF_bus_selected_win_data_433_port, 
      DataPath_RF_bus_selected_win_data_434_port, 
      DataPath_RF_bus_selected_win_data_435_port, 
      DataPath_RF_bus_selected_win_data_436_port, 
      DataPath_RF_bus_selected_win_data_437_port, 
      DataPath_RF_bus_selected_win_data_438_port, 
      DataPath_RF_bus_selected_win_data_439_port, 
      DataPath_RF_bus_selected_win_data_440_port, 
      DataPath_RF_bus_selected_win_data_441_port, 
      DataPath_RF_bus_selected_win_data_442_port, 
      DataPath_RF_bus_selected_win_data_443_port, 
      DataPath_RF_bus_selected_win_data_444_port, 
      DataPath_RF_bus_selected_win_data_445_port, 
      DataPath_RF_bus_selected_win_data_446_port, 
      DataPath_RF_bus_selected_win_data_447_port, 
      DataPath_RF_bus_selected_win_data_448_port, 
      DataPath_RF_bus_selected_win_data_449_port, 
      DataPath_RF_bus_selected_win_data_450_port, 
      DataPath_RF_bus_selected_win_data_451_port, 
      DataPath_RF_bus_selected_win_data_452_port, 
      DataPath_RF_bus_selected_win_data_453_port, 
      DataPath_RF_bus_selected_win_data_454_port, 
      DataPath_RF_bus_selected_win_data_455_port, 
      DataPath_RF_bus_selected_win_data_456_port, 
      DataPath_RF_bus_selected_win_data_457_port, 
      DataPath_RF_bus_selected_win_data_458_port, 
      DataPath_RF_bus_selected_win_data_459_port, 
      DataPath_RF_bus_selected_win_data_460_port, 
      DataPath_RF_bus_selected_win_data_461_port, 
      DataPath_RF_bus_selected_win_data_462_port, 
      DataPath_RF_bus_selected_win_data_463_port, 
      DataPath_RF_bus_selected_win_data_464_port, 
      DataPath_RF_bus_selected_win_data_465_port, 
      DataPath_RF_bus_selected_win_data_466_port, 
      DataPath_RF_bus_selected_win_data_467_port, 
      DataPath_RF_bus_selected_win_data_468_port, 
      DataPath_RF_bus_selected_win_data_469_port, 
      DataPath_RF_bus_selected_win_data_470_port, 
      DataPath_RF_bus_selected_win_data_471_port, 
      DataPath_RF_bus_selected_win_data_472_port, 
      DataPath_RF_bus_selected_win_data_473_port, 
      DataPath_RF_bus_selected_win_data_474_port, 
      DataPath_RF_bus_selected_win_data_475_port, 
      DataPath_RF_bus_selected_win_data_476_port, 
      DataPath_RF_bus_selected_win_data_477_port, 
      DataPath_RF_bus_selected_win_data_478_port, 
      DataPath_RF_bus_selected_win_data_479_port, 
      DataPath_RF_bus_selected_win_data_480_port, 
      DataPath_RF_bus_selected_win_data_481_port, 
      DataPath_RF_bus_selected_win_data_482_port, 
      DataPath_RF_bus_selected_win_data_483_port, 
      DataPath_RF_bus_selected_win_data_484_port, 
      DataPath_RF_bus_selected_win_data_485_port, 
      DataPath_RF_bus_selected_win_data_486_port, 
      DataPath_RF_bus_selected_win_data_487_port, 
      DataPath_RF_bus_selected_win_data_488_port, 
      DataPath_RF_bus_selected_win_data_489_port, 
      DataPath_RF_bus_selected_win_data_490_port, 
      DataPath_RF_bus_selected_win_data_491_port, 
      DataPath_RF_bus_selected_win_data_492_port, 
      DataPath_RF_bus_selected_win_data_493_port, 
      DataPath_RF_bus_selected_win_data_494_port, 
      DataPath_RF_bus_selected_win_data_495_port, 
      DataPath_RF_bus_selected_win_data_496_port, 
      DataPath_RF_bus_selected_win_data_497_port, 
      DataPath_RF_bus_selected_win_data_498_port, 
      DataPath_RF_bus_selected_win_data_499_port, 
      DataPath_RF_bus_selected_win_data_500_port, 
      DataPath_RF_bus_selected_win_data_501_port, 
      DataPath_RF_bus_selected_win_data_502_port, 
      DataPath_RF_bus_selected_win_data_503_port, 
      DataPath_RF_bus_selected_win_data_504_port, 
      DataPath_RF_bus_selected_win_data_505_port, 
      DataPath_RF_bus_selected_win_data_506_port, 
      DataPath_RF_bus_selected_win_data_507_port, 
      DataPath_RF_bus_selected_win_data_508_port, 
      DataPath_RF_bus_selected_win_data_509_port, 
      DataPath_RF_bus_selected_win_data_510_port, 
      DataPath_RF_bus_selected_win_data_511_port, 
      DataPath_RF_bus_selected_win_data_512_port, 
      DataPath_RF_bus_selected_win_data_513_port, 
      DataPath_RF_bus_selected_win_data_514_port, 
      DataPath_RF_bus_selected_win_data_515_port, 
      DataPath_RF_bus_selected_win_data_516_port, 
      DataPath_RF_bus_selected_win_data_517_port, 
      DataPath_RF_bus_selected_win_data_518_port, 
      DataPath_RF_bus_selected_win_data_519_port, 
      DataPath_RF_bus_selected_win_data_520_port, 
      DataPath_RF_bus_selected_win_data_521_port, 
      DataPath_RF_bus_selected_win_data_522_port, 
      DataPath_RF_bus_selected_win_data_523_port, 
      DataPath_RF_bus_selected_win_data_524_port, 
      DataPath_RF_bus_selected_win_data_525_port, 
      DataPath_RF_bus_selected_win_data_526_port, 
      DataPath_RF_bus_selected_win_data_527_port, 
      DataPath_RF_bus_selected_win_data_528_port, 
      DataPath_RF_bus_selected_win_data_529_port, 
      DataPath_RF_bus_selected_win_data_530_port, 
      DataPath_RF_bus_selected_win_data_531_port, 
      DataPath_RF_bus_selected_win_data_532_port, 
      DataPath_RF_bus_selected_win_data_533_port, 
      DataPath_RF_bus_selected_win_data_534_port, 
      DataPath_RF_bus_selected_win_data_535_port, 
      DataPath_RF_bus_selected_win_data_536_port, 
      DataPath_RF_bus_selected_win_data_537_port, 
      DataPath_RF_bus_selected_win_data_538_port, 
      DataPath_RF_bus_selected_win_data_539_port, 
      DataPath_RF_bus_selected_win_data_540_port, 
      DataPath_RF_bus_selected_win_data_541_port, 
      DataPath_RF_bus_selected_win_data_542_port, 
      DataPath_RF_bus_selected_win_data_543_port, 
      DataPath_RF_bus_selected_win_data_544_port, 
      DataPath_RF_bus_selected_win_data_545_port, 
      DataPath_RF_bus_selected_win_data_546_port, 
      DataPath_RF_bus_selected_win_data_547_port, 
      DataPath_RF_bus_selected_win_data_548_port, 
      DataPath_RF_bus_selected_win_data_549_port, 
      DataPath_RF_bus_selected_win_data_550_port, 
      DataPath_RF_bus_selected_win_data_551_port, 
      DataPath_RF_bus_selected_win_data_552_port, 
      DataPath_RF_bus_selected_win_data_553_port, 
      DataPath_RF_bus_selected_win_data_554_port, 
      DataPath_RF_bus_selected_win_data_555_port, 
      DataPath_RF_bus_selected_win_data_556_port, 
      DataPath_RF_bus_selected_win_data_557_port, 
      DataPath_RF_bus_selected_win_data_558_port, 
      DataPath_RF_bus_selected_win_data_559_port, 
      DataPath_RF_bus_selected_win_data_560_port, 
      DataPath_RF_bus_selected_win_data_561_port, 
      DataPath_RF_bus_selected_win_data_562_port, 
      DataPath_RF_bus_selected_win_data_563_port, 
      DataPath_RF_bus_selected_win_data_564_port, 
      DataPath_RF_bus_selected_win_data_565_port, 
      DataPath_RF_bus_selected_win_data_566_port, 
      DataPath_RF_bus_selected_win_data_567_port, 
      DataPath_RF_bus_selected_win_data_568_port, 
      DataPath_RF_bus_selected_win_data_569_port, 
      DataPath_RF_bus_selected_win_data_570_port, 
      DataPath_RF_bus_selected_win_data_571_port, 
      DataPath_RF_bus_selected_win_data_572_port, 
      DataPath_RF_bus_selected_win_data_573_port, 
      DataPath_RF_bus_selected_win_data_574_port, 
      DataPath_RF_bus_selected_win_data_575_port, 
      DataPath_RF_bus_selected_win_data_576_port, 
      DataPath_RF_bus_selected_win_data_577_port, 
      DataPath_RF_bus_selected_win_data_578_port, 
      DataPath_RF_bus_selected_win_data_579_port, 
      DataPath_RF_bus_selected_win_data_580_port, 
      DataPath_RF_bus_selected_win_data_581_port, 
      DataPath_RF_bus_selected_win_data_582_port, 
      DataPath_RF_bus_selected_win_data_583_port, 
      DataPath_RF_bus_selected_win_data_584_port, 
      DataPath_RF_bus_selected_win_data_585_port, 
      DataPath_RF_bus_selected_win_data_586_port, 
      DataPath_RF_bus_selected_win_data_587_port, 
      DataPath_RF_bus_selected_win_data_588_port, 
      DataPath_RF_bus_selected_win_data_589_port, 
      DataPath_RF_bus_selected_win_data_590_port, 
      DataPath_RF_bus_selected_win_data_591_port, 
      DataPath_RF_bus_selected_win_data_592_port, 
      DataPath_RF_bus_selected_win_data_593_port, 
      DataPath_RF_bus_selected_win_data_594_port, 
      DataPath_RF_bus_selected_win_data_595_port, 
      DataPath_RF_bus_selected_win_data_596_port, 
      DataPath_RF_bus_selected_win_data_597_port, 
      DataPath_RF_bus_selected_win_data_598_port, 
      DataPath_RF_bus_selected_win_data_599_port, 
      DataPath_RF_bus_selected_win_data_600_port, 
      DataPath_RF_bus_selected_win_data_601_port, 
      DataPath_RF_bus_selected_win_data_602_port, 
      DataPath_RF_bus_selected_win_data_603_port, 
      DataPath_RF_bus_selected_win_data_604_port, 
      DataPath_RF_bus_selected_win_data_605_port, 
      DataPath_RF_bus_selected_win_data_606_port, 
      DataPath_RF_bus_selected_win_data_607_port, 
      DataPath_RF_bus_selected_win_data_608_port, 
      DataPath_RF_bus_selected_win_data_609_port, 
      DataPath_RF_bus_selected_win_data_610_port, 
      DataPath_RF_bus_selected_win_data_611_port, 
      DataPath_RF_bus_selected_win_data_612_port, 
      DataPath_RF_bus_selected_win_data_613_port, 
      DataPath_RF_bus_selected_win_data_614_port, 
      DataPath_RF_bus_selected_win_data_615_port, 
      DataPath_RF_bus_selected_win_data_616_port, 
      DataPath_RF_bus_selected_win_data_617_port, 
      DataPath_RF_bus_selected_win_data_618_port, 
      DataPath_RF_bus_selected_win_data_619_port, 
      DataPath_RF_bus_selected_win_data_620_port, 
      DataPath_RF_bus_selected_win_data_621_port, 
      DataPath_RF_bus_selected_win_data_622_port, 
      DataPath_RF_bus_selected_win_data_623_port, 
      DataPath_RF_bus_selected_win_data_624_port, 
      DataPath_RF_bus_selected_win_data_625_port, 
      DataPath_RF_bus_selected_win_data_626_port, 
      DataPath_RF_bus_selected_win_data_627_port, 
      DataPath_RF_bus_selected_win_data_628_port, 
      DataPath_RF_bus_selected_win_data_629_port, 
      DataPath_RF_bus_selected_win_data_630_port, 
      DataPath_RF_bus_selected_win_data_631_port, 
      DataPath_RF_bus_selected_win_data_632_port, 
      DataPath_RF_bus_selected_win_data_633_port, 
      DataPath_RF_bus_selected_win_data_634_port, 
      DataPath_RF_bus_selected_win_data_635_port, 
      DataPath_RF_bus_selected_win_data_636_port, 
      DataPath_RF_bus_selected_win_data_637_port, 
      DataPath_RF_bus_selected_win_data_638_port, 
      DataPath_RF_bus_selected_win_data_639_port, 
      DataPath_RF_bus_selected_win_data_640_port, 
      DataPath_RF_bus_selected_win_data_641_port, 
      DataPath_RF_bus_selected_win_data_642_port, 
      DataPath_RF_bus_selected_win_data_643_port, 
      DataPath_RF_bus_selected_win_data_644_port, 
      DataPath_RF_bus_selected_win_data_645_port, 
      DataPath_RF_bus_selected_win_data_646_port, 
      DataPath_RF_bus_selected_win_data_647_port, 
      DataPath_RF_bus_selected_win_data_648_port, 
      DataPath_RF_bus_selected_win_data_649_port, 
      DataPath_RF_bus_selected_win_data_650_port, 
      DataPath_RF_bus_selected_win_data_651_port, 
      DataPath_RF_bus_selected_win_data_652_port, 
      DataPath_RF_bus_selected_win_data_653_port, 
      DataPath_RF_bus_selected_win_data_654_port, 
      DataPath_RF_bus_selected_win_data_655_port, 
      DataPath_RF_bus_selected_win_data_656_port, 
      DataPath_RF_bus_selected_win_data_657_port, 
      DataPath_RF_bus_selected_win_data_658_port, 
      DataPath_RF_bus_selected_win_data_659_port, 
      DataPath_RF_bus_selected_win_data_660_port, 
      DataPath_RF_bus_selected_win_data_661_port, 
      DataPath_RF_bus_selected_win_data_662_port, 
      DataPath_RF_bus_selected_win_data_663_port, 
      DataPath_RF_bus_selected_win_data_664_port, 
      DataPath_RF_bus_selected_win_data_665_port, 
      DataPath_RF_bus_selected_win_data_666_port, 
      DataPath_RF_bus_selected_win_data_667_port, 
      DataPath_RF_bus_selected_win_data_668_port, 
      DataPath_RF_bus_selected_win_data_669_port, 
      DataPath_RF_bus_selected_win_data_670_port, 
      DataPath_RF_bus_selected_win_data_671_port, 
      DataPath_RF_bus_selected_win_data_672_port, 
      DataPath_RF_bus_selected_win_data_673_port, 
      DataPath_RF_bus_selected_win_data_674_port, 
      DataPath_RF_bus_selected_win_data_675_port, 
      DataPath_RF_bus_selected_win_data_676_port, 
      DataPath_RF_bus_selected_win_data_677_port, 
      DataPath_RF_bus_selected_win_data_678_port, 
      DataPath_RF_bus_selected_win_data_679_port, 
      DataPath_RF_bus_selected_win_data_680_port, 
      DataPath_RF_bus_selected_win_data_681_port, 
      DataPath_RF_bus_selected_win_data_682_port, 
      DataPath_RF_bus_selected_win_data_683_port, 
      DataPath_RF_bus_selected_win_data_684_port, 
      DataPath_RF_bus_selected_win_data_685_port, 
      DataPath_RF_bus_selected_win_data_686_port, 
      DataPath_RF_bus_selected_win_data_687_port, 
      DataPath_RF_bus_selected_win_data_688_port, 
      DataPath_RF_bus_selected_win_data_689_port, 
      DataPath_RF_bus_selected_win_data_690_port, 
      DataPath_RF_bus_selected_win_data_691_port, 
      DataPath_RF_bus_selected_win_data_692_port, 
      DataPath_RF_bus_selected_win_data_693_port, 
      DataPath_RF_bus_selected_win_data_694_port, 
      DataPath_RF_bus_selected_win_data_695_port, 
      DataPath_RF_bus_selected_win_data_696_port, 
      DataPath_RF_bus_selected_win_data_697_port, 
      DataPath_RF_bus_selected_win_data_698_port, 
      DataPath_RF_bus_selected_win_data_699_port, 
      DataPath_RF_bus_selected_win_data_700_port, 
      DataPath_RF_bus_selected_win_data_701_port, 
      DataPath_RF_bus_selected_win_data_702_port, 
      DataPath_RF_bus_selected_win_data_703_port, 
      DataPath_RF_bus_selected_win_data_704_port, 
      DataPath_RF_bus_selected_win_data_705_port, 
      DataPath_RF_bus_selected_win_data_706_port, 
      DataPath_RF_bus_selected_win_data_707_port, 
      DataPath_RF_bus_selected_win_data_708_port, 
      DataPath_RF_bus_selected_win_data_709_port, 
      DataPath_RF_bus_selected_win_data_710_port, 
      DataPath_RF_bus_selected_win_data_711_port, 
      DataPath_RF_bus_selected_win_data_712_port, 
      DataPath_RF_bus_selected_win_data_713_port, 
      DataPath_RF_bus_selected_win_data_714_port, 
      DataPath_RF_bus_selected_win_data_715_port, 
      DataPath_RF_bus_selected_win_data_716_port, 
      DataPath_RF_bus_selected_win_data_717_port, 
      DataPath_RF_bus_selected_win_data_718_port, 
      DataPath_RF_bus_selected_win_data_719_port, 
      DataPath_RF_bus_selected_win_data_720_port, 
      DataPath_RF_bus_selected_win_data_721_port, 
      DataPath_RF_bus_selected_win_data_722_port, 
      DataPath_RF_bus_selected_win_data_723_port, 
      DataPath_RF_bus_selected_win_data_724_port, 
      DataPath_RF_bus_selected_win_data_725_port, 
      DataPath_RF_bus_selected_win_data_726_port, 
      DataPath_RF_bus_selected_win_data_727_port, 
      DataPath_RF_bus_selected_win_data_728_port, 
      DataPath_RF_bus_selected_win_data_729_port, 
      DataPath_RF_bus_selected_win_data_730_port, 
      DataPath_RF_bus_selected_win_data_731_port, 
      DataPath_RF_bus_selected_win_data_732_port, 
      DataPath_RF_bus_selected_win_data_733_port, 
      DataPath_RF_bus_selected_win_data_734_port, 
      DataPath_RF_bus_selected_win_data_735_port, 
      DataPath_RF_bus_selected_win_data_736_port, 
      DataPath_RF_bus_selected_win_data_737_port, 
      DataPath_RF_bus_selected_win_data_738_port, 
      DataPath_RF_bus_selected_win_data_739_port, 
      DataPath_RF_bus_selected_win_data_740_port, 
      DataPath_RF_bus_selected_win_data_741_port, 
      DataPath_RF_bus_selected_win_data_742_port, 
      DataPath_RF_bus_selected_win_data_743_port, 
      DataPath_RF_bus_selected_win_data_744_port, 
      DataPath_RF_bus_selected_win_data_745_port, 
      DataPath_RF_bus_selected_win_data_746_port, 
      DataPath_RF_bus_selected_win_data_747_port, 
      DataPath_RF_bus_selected_win_data_748_port, 
      DataPath_RF_bus_selected_win_data_749_port, 
      DataPath_RF_bus_selected_win_data_750_port, 
      DataPath_RF_bus_selected_win_data_751_port, 
      DataPath_RF_bus_selected_win_data_752_port, 
      DataPath_RF_bus_selected_win_data_753_port, 
      DataPath_RF_bus_selected_win_data_754_port, 
      DataPath_RF_bus_selected_win_data_755_port, 
      DataPath_RF_bus_selected_win_data_756_port, 
      DataPath_RF_bus_selected_win_data_757_port, 
      DataPath_RF_bus_selected_win_data_758_port, 
      DataPath_RF_bus_selected_win_data_759_port, 
      DataPath_RF_bus_selected_win_data_760_port, 
      DataPath_RF_bus_selected_win_data_761_port, 
      DataPath_RF_bus_selected_win_data_762_port, 
      DataPath_RF_bus_selected_win_data_763_port, 
      DataPath_RF_bus_selected_win_data_764_port, 
      DataPath_RF_bus_selected_win_data_765_port, 
      DataPath_RF_bus_selected_win_data_766_port, 
      DataPath_RF_bus_selected_win_data_767_port, 
      DataPath_RF_bus_reg_dataout_0_port, DataPath_RF_bus_reg_dataout_1_port, 
      DataPath_RF_bus_reg_dataout_2_port, DataPath_RF_bus_reg_dataout_3_port, 
      DataPath_RF_bus_reg_dataout_4_port, DataPath_RF_bus_reg_dataout_5_port, 
      DataPath_RF_bus_reg_dataout_6_port, DataPath_RF_bus_reg_dataout_7_port, 
      DataPath_RF_bus_reg_dataout_8_port, DataPath_RF_bus_reg_dataout_9_port, 
      DataPath_RF_bus_reg_dataout_10_port, DataPath_RF_bus_reg_dataout_11_port,
      DataPath_RF_bus_reg_dataout_12_port, DataPath_RF_bus_reg_dataout_13_port,
      DataPath_RF_bus_reg_dataout_14_port, DataPath_RF_bus_reg_dataout_15_port,
      DataPath_RF_bus_reg_dataout_16_port, DataPath_RF_bus_reg_dataout_17_port,
      DataPath_RF_bus_reg_dataout_18_port, DataPath_RF_bus_reg_dataout_19_port,
      DataPath_RF_bus_reg_dataout_20_port, DataPath_RF_bus_reg_dataout_21_port,
      DataPath_RF_bus_reg_dataout_22_port, DataPath_RF_bus_reg_dataout_23_port,
      DataPath_RF_bus_reg_dataout_24_port, DataPath_RF_bus_reg_dataout_25_port,
      DataPath_RF_bus_reg_dataout_26_port, DataPath_RF_bus_reg_dataout_27_port,
      DataPath_RF_bus_reg_dataout_28_port, DataPath_RF_bus_reg_dataout_29_port,
      DataPath_RF_bus_reg_dataout_30_port, DataPath_RF_bus_reg_dataout_31_port,
      DataPath_RF_bus_reg_dataout_32_port, DataPath_RF_bus_reg_dataout_33_port,
      DataPath_RF_bus_reg_dataout_34_port, DataPath_RF_bus_reg_dataout_35_port,
      DataPath_RF_bus_reg_dataout_36_port, DataPath_RF_bus_reg_dataout_37_port,
      DataPath_RF_bus_reg_dataout_38_port, DataPath_RF_bus_reg_dataout_39_port,
      DataPath_RF_bus_reg_dataout_40_port, DataPath_RF_bus_reg_dataout_41_port,
      DataPath_RF_bus_reg_dataout_42_port, DataPath_RF_bus_reg_dataout_43_port,
      DataPath_RF_bus_reg_dataout_44_port, DataPath_RF_bus_reg_dataout_45_port,
      DataPath_RF_bus_reg_dataout_46_port, DataPath_RF_bus_reg_dataout_47_port,
      DataPath_RF_bus_reg_dataout_48_port, DataPath_RF_bus_reg_dataout_49_port,
      DataPath_RF_bus_reg_dataout_50_port, DataPath_RF_bus_reg_dataout_51_port,
      DataPath_RF_bus_reg_dataout_52_port, DataPath_RF_bus_reg_dataout_53_port,
      DataPath_RF_bus_reg_dataout_54_port, DataPath_RF_bus_reg_dataout_55_port,
      DataPath_RF_bus_reg_dataout_56_port, DataPath_RF_bus_reg_dataout_57_port,
      DataPath_RF_bus_reg_dataout_58_port, DataPath_RF_bus_reg_dataout_59_port,
      DataPath_RF_bus_reg_dataout_60_port, DataPath_RF_bus_reg_dataout_61_port,
      DataPath_RF_bus_reg_dataout_62_port, DataPath_RF_bus_reg_dataout_63_port,
      DataPath_RF_bus_reg_dataout_64_port, DataPath_RF_bus_reg_dataout_65_port,
      DataPath_RF_bus_reg_dataout_66_port, DataPath_RF_bus_reg_dataout_67_port,
      DataPath_RF_bus_reg_dataout_68_port, DataPath_RF_bus_reg_dataout_69_port,
      DataPath_RF_bus_reg_dataout_70_port, DataPath_RF_bus_reg_dataout_71_port,
      DataPath_RF_bus_reg_dataout_72_port, DataPath_RF_bus_reg_dataout_73_port,
      DataPath_RF_bus_reg_dataout_74_port, DataPath_RF_bus_reg_dataout_75_port,
      DataPath_RF_bus_reg_dataout_76_port, DataPath_RF_bus_reg_dataout_77_port,
      DataPath_RF_bus_reg_dataout_78_port, DataPath_RF_bus_reg_dataout_79_port,
      DataPath_RF_bus_reg_dataout_80_port, DataPath_RF_bus_reg_dataout_81_port,
      DataPath_RF_bus_reg_dataout_82_port, DataPath_RF_bus_reg_dataout_83_port,
      DataPath_RF_bus_reg_dataout_84_port, DataPath_RF_bus_reg_dataout_85_port,
      DataPath_RF_bus_reg_dataout_86_port, DataPath_RF_bus_reg_dataout_87_port,
      DataPath_RF_bus_reg_dataout_88_port, DataPath_RF_bus_reg_dataout_89_port,
      DataPath_RF_bus_reg_dataout_90_port, DataPath_RF_bus_reg_dataout_91_port,
      DataPath_RF_bus_reg_dataout_92_port, DataPath_RF_bus_reg_dataout_93_port,
      DataPath_RF_bus_reg_dataout_94_port, DataPath_RF_bus_reg_dataout_95_port,
      DataPath_RF_bus_reg_dataout_96_port, DataPath_RF_bus_reg_dataout_97_port,
      DataPath_RF_bus_reg_dataout_98_port, DataPath_RF_bus_reg_dataout_99_port,
      DataPath_RF_bus_reg_dataout_100_port, 
      DataPath_RF_bus_reg_dataout_101_port, 
      DataPath_RF_bus_reg_dataout_102_port, 
      DataPath_RF_bus_reg_dataout_103_port, 
      DataPath_RF_bus_reg_dataout_104_port, 
      DataPath_RF_bus_reg_dataout_105_port, 
      DataPath_RF_bus_reg_dataout_106_port, 
      DataPath_RF_bus_reg_dataout_107_port, 
      DataPath_RF_bus_reg_dataout_108_port, 
      DataPath_RF_bus_reg_dataout_109_port, 
      DataPath_RF_bus_reg_dataout_110_port, 
      DataPath_RF_bus_reg_dataout_111_port, 
      DataPath_RF_bus_reg_dataout_112_port, 
      DataPath_RF_bus_reg_dataout_113_port, 
      DataPath_RF_bus_reg_dataout_114_port, 
      DataPath_RF_bus_reg_dataout_115_port, 
      DataPath_RF_bus_reg_dataout_116_port, 
      DataPath_RF_bus_reg_dataout_117_port, 
      DataPath_RF_bus_reg_dataout_118_port, 
      DataPath_RF_bus_reg_dataout_119_port, 
      DataPath_RF_bus_reg_dataout_120_port, 
      DataPath_RF_bus_reg_dataout_121_port, 
      DataPath_RF_bus_reg_dataout_122_port, 
      DataPath_RF_bus_reg_dataout_123_port, 
      DataPath_RF_bus_reg_dataout_124_port, 
      DataPath_RF_bus_reg_dataout_125_port, 
      DataPath_RF_bus_reg_dataout_126_port, 
      DataPath_RF_bus_reg_dataout_127_port, 
      DataPath_RF_bus_reg_dataout_128_port, 
      DataPath_RF_bus_reg_dataout_129_port, 
      DataPath_RF_bus_reg_dataout_130_port, 
      DataPath_RF_bus_reg_dataout_131_port, 
      DataPath_RF_bus_reg_dataout_132_port, 
      DataPath_RF_bus_reg_dataout_133_port, 
      DataPath_RF_bus_reg_dataout_134_port, 
      DataPath_RF_bus_reg_dataout_135_port, 
      DataPath_RF_bus_reg_dataout_136_port, 
      DataPath_RF_bus_reg_dataout_137_port, 
      DataPath_RF_bus_reg_dataout_138_port, 
      DataPath_RF_bus_reg_dataout_139_port, 
      DataPath_RF_bus_reg_dataout_140_port, 
      DataPath_RF_bus_reg_dataout_141_port, 
      DataPath_RF_bus_reg_dataout_142_port, 
      DataPath_RF_bus_reg_dataout_143_port, 
      DataPath_RF_bus_reg_dataout_144_port, 
      DataPath_RF_bus_reg_dataout_145_port, 
      DataPath_RF_bus_reg_dataout_146_port, 
      DataPath_RF_bus_reg_dataout_147_port, 
      DataPath_RF_bus_reg_dataout_148_port, 
      DataPath_RF_bus_reg_dataout_149_port, 
      DataPath_RF_bus_reg_dataout_150_port, 
      DataPath_RF_bus_reg_dataout_151_port, 
      DataPath_RF_bus_reg_dataout_152_port, 
      DataPath_RF_bus_reg_dataout_153_port, 
      DataPath_RF_bus_reg_dataout_154_port, 
      DataPath_RF_bus_reg_dataout_155_port, 
      DataPath_RF_bus_reg_dataout_156_port, 
      DataPath_RF_bus_reg_dataout_157_port, 
      DataPath_RF_bus_reg_dataout_158_port, 
      DataPath_RF_bus_reg_dataout_159_port, 
      DataPath_RF_bus_reg_dataout_160_port, 
      DataPath_RF_bus_reg_dataout_161_port, 
      DataPath_RF_bus_reg_dataout_162_port, 
      DataPath_RF_bus_reg_dataout_163_port, 
      DataPath_RF_bus_reg_dataout_164_port, 
      DataPath_RF_bus_reg_dataout_165_port, 
      DataPath_RF_bus_reg_dataout_166_port, 
      DataPath_RF_bus_reg_dataout_167_port, 
      DataPath_RF_bus_reg_dataout_168_port, 
      DataPath_RF_bus_reg_dataout_169_port, 
      DataPath_RF_bus_reg_dataout_170_port, 
      DataPath_RF_bus_reg_dataout_171_port, 
      DataPath_RF_bus_reg_dataout_172_port, 
      DataPath_RF_bus_reg_dataout_173_port, 
      DataPath_RF_bus_reg_dataout_174_port, 
      DataPath_RF_bus_reg_dataout_175_port, 
      DataPath_RF_bus_reg_dataout_176_port, 
      DataPath_RF_bus_reg_dataout_177_port, 
      DataPath_RF_bus_reg_dataout_178_port, 
      DataPath_RF_bus_reg_dataout_179_port, 
      DataPath_RF_bus_reg_dataout_180_port, 
      DataPath_RF_bus_reg_dataout_181_port, 
      DataPath_RF_bus_reg_dataout_182_port, 
      DataPath_RF_bus_reg_dataout_183_port, 
      DataPath_RF_bus_reg_dataout_184_port, 
      DataPath_RF_bus_reg_dataout_185_port, 
      DataPath_RF_bus_reg_dataout_186_port, 
      DataPath_RF_bus_reg_dataout_187_port, 
      DataPath_RF_bus_reg_dataout_188_port, 
      DataPath_RF_bus_reg_dataout_189_port, 
      DataPath_RF_bus_reg_dataout_190_port, 
      DataPath_RF_bus_reg_dataout_191_port, 
      DataPath_RF_bus_reg_dataout_192_port, 
      DataPath_RF_bus_reg_dataout_193_port, 
      DataPath_RF_bus_reg_dataout_194_port, 
      DataPath_RF_bus_reg_dataout_195_port, 
      DataPath_RF_bus_reg_dataout_196_port, 
      DataPath_RF_bus_reg_dataout_197_port, 
      DataPath_RF_bus_reg_dataout_198_port, 
      DataPath_RF_bus_reg_dataout_199_port, 
      DataPath_RF_bus_reg_dataout_200_port, 
      DataPath_RF_bus_reg_dataout_201_port, 
      DataPath_RF_bus_reg_dataout_202_port, 
      DataPath_RF_bus_reg_dataout_203_port, 
      DataPath_RF_bus_reg_dataout_204_port, 
      DataPath_RF_bus_reg_dataout_205_port, 
      DataPath_RF_bus_reg_dataout_206_port, 
      DataPath_RF_bus_reg_dataout_207_port, 
      DataPath_RF_bus_reg_dataout_208_port, 
      DataPath_RF_bus_reg_dataout_209_port, 
      DataPath_RF_bus_reg_dataout_210_port, 
      DataPath_RF_bus_reg_dataout_211_port, 
      DataPath_RF_bus_reg_dataout_212_port, 
      DataPath_RF_bus_reg_dataout_213_port, 
      DataPath_RF_bus_reg_dataout_214_port, 
      DataPath_RF_bus_reg_dataout_215_port, 
      DataPath_RF_bus_reg_dataout_216_port, 
      DataPath_RF_bus_reg_dataout_217_port, 
      DataPath_RF_bus_reg_dataout_218_port, 
      DataPath_RF_bus_reg_dataout_219_port, 
      DataPath_RF_bus_reg_dataout_220_port, 
      DataPath_RF_bus_reg_dataout_221_port, 
      DataPath_RF_bus_reg_dataout_222_port, 
      DataPath_RF_bus_reg_dataout_223_port, 
      DataPath_RF_bus_reg_dataout_224_port, 
      DataPath_RF_bus_reg_dataout_225_port, 
      DataPath_RF_bus_reg_dataout_226_port, 
      DataPath_RF_bus_reg_dataout_227_port, 
      DataPath_RF_bus_reg_dataout_228_port, 
      DataPath_RF_bus_reg_dataout_229_port, 
      DataPath_RF_bus_reg_dataout_230_port, 
      DataPath_RF_bus_reg_dataout_231_port, 
      DataPath_RF_bus_reg_dataout_232_port, 
      DataPath_RF_bus_reg_dataout_233_port, 
      DataPath_RF_bus_reg_dataout_234_port, 
      DataPath_RF_bus_reg_dataout_235_port, 
      DataPath_RF_bus_reg_dataout_236_port, 
      DataPath_RF_bus_reg_dataout_237_port, 
      DataPath_RF_bus_reg_dataout_238_port, 
      DataPath_RF_bus_reg_dataout_239_port, 
      DataPath_RF_bus_reg_dataout_240_port, 
      DataPath_RF_bus_reg_dataout_241_port, 
      DataPath_RF_bus_reg_dataout_242_port, 
      DataPath_RF_bus_reg_dataout_243_port, 
      DataPath_RF_bus_reg_dataout_244_port, 
      DataPath_RF_bus_reg_dataout_245_port, 
      DataPath_RF_bus_reg_dataout_246_port, 
      DataPath_RF_bus_reg_dataout_247_port, 
      DataPath_RF_bus_reg_dataout_248_port, 
      DataPath_RF_bus_reg_dataout_249_port, 
      DataPath_RF_bus_reg_dataout_250_port, 
      DataPath_RF_bus_reg_dataout_251_port, 
      DataPath_RF_bus_reg_dataout_252_port, 
      DataPath_RF_bus_reg_dataout_253_port, 
      DataPath_RF_bus_reg_dataout_254_port, 
      DataPath_RF_bus_reg_dataout_255_port, 
      DataPath_RF_bus_reg_dataout_256_port, 
      DataPath_RF_bus_reg_dataout_257_port, 
      DataPath_RF_bus_reg_dataout_258_port, 
      DataPath_RF_bus_reg_dataout_259_port, 
      DataPath_RF_bus_reg_dataout_260_port, 
      DataPath_RF_bus_reg_dataout_261_port, 
      DataPath_RF_bus_reg_dataout_262_port, 
      DataPath_RF_bus_reg_dataout_263_port, 
      DataPath_RF_bus_reg_dataout_264_port, 
      DataPath_RF_bus_reg_dataout_265_port, 
      DataPath_RF_bus_reg_dataout_266_port, 
      DataPath_RF_bus_reg_dataout_267_port, 
      DataPath_RF_bus_reg_dataout_268_port, 
      DataPath_RF_bus_reg_dataout_269_port, 
      DataPath_RF_bus_reg_dataout_270_port, 
      DataPath_RF_bus_reg_dataout_271_port, 
      DataPath_RF_bus_reg_dataout_272_port, 
      DataPath_RF_bus_reg_dataout_273_port, 
      DataPath_RF_bus_reg_dataout_274_port, 
      DataPath_RF_bus_reg_dataout_275_port, 
      DataPath_RF_bus_reg_dataout_276_port, 
      DataPath_RF_bus_reg_dataout_277_port, 
      DataPath_RF_bus_reg_dataout_278_port, 
      DataPath_RF_bus_reg_dataout_279_port, 
      DataPath_RF_bus_reg_dataout_280_port, 
      DataPath_RF_bus_reg_dataout_281_port, 
      DataPath_RF_bus_reg_dataout_282_port, 
      DataPath_RF_bus_reg_dataout_283_port, 
      DataPath_RF_bus_reg_dataout_284_port, 
      DataPath_RF_bus_reg_dataout_285_port, 
      DataPath_RF_bus_reg_dataout_286_port, 
      DataPath_RF_bus_reg_dataout_287_port, 
      DataPath_RF_bus_reg_dataout_288_port, 
      DataPath_RF_bus_reg_dataout_289_port, 
      DataPath_RF_bus_reg_dataout_290_port, 
      DataPath_RF_bus_reg_dataout_291_port, 
      DataPath_RF_bus_reg_dataout_292_port, 
      DataPath_RF_bus_reg_dataout_293_port, 
      DataPath_RF_bus_reg_dataout_294_port, 
      DataPath_RF_bus_reg_dataout_295_port, 
      DataPath_RF_bus_reg_dataout_296_port, 
      DataPath_RF_bus_reg_dataout_297_port, 
      DataPath_RF_bus_reg_dataout_298_port, 
      DataPath_RF_bus_reg_dataout_299_port, 
      DataPath_RF_bus_reg_dataout_300_port, 
      DataPath_RF_bus_reg_dataout_301_port, 
      DataPath_RF_bus_reg_dataout_302_port, 
      DataPath_RF_bus_reg_dataout_303_port, 
      DataPath_RF_bus_reg_dataout_304_port, 
      DataPath_RF_bus_reg_dataout_305_port, 
      DataPath_RF_bus_reg_dataout_306_port, 
      DataPath_RF_bus_reg_dataout_307_port, 
      DataPath_RF_bus_reg_dataout_308_port, 
      DataPath_RF_bus_reg_dataout_309_port, 
      DataPath_RF_bus_reg_dataout_310_port, 
      DataPath_RF_bus_reg_dataout_311_port, 
      DataPath_RF_bus_reg_dataout_312_port, 
      DataPath_RF_bus_reg_dataout_313_port, 
      DataPath_RF_bus_reg_dataout_314_port, 
      DataPath_RF_bus_reg_dataout_315_port, 
      DataPath_RF_bus_reg_dataout_316_port, 
      DataPath_RF_bus_reg_dataout_317_port, 
      DataPath_RF_bus_reg_dataout_318_port, 
      DataPath_RF_bus_reg_dataout_319_port, 
      DataPath_RF_bus_reg_dataout_320_port, 
      DataPath_RF_bus_reg_dataout_321_port, 
      DataPath_RF_bus_reg_dataout_322_port, 
      DataPath_RF_bus_reg_dataout_323_port, 
      DataPath_RF_bus_reg_dataout_324_port, 
      DataPath_RF_bus_reg_dataout_325_port, 
      DataPath_RF_bus_reg_dataout_326_port, 
      DataPath_RF_bus_reg_dataout_327_port, 
      DataPath_RF_bus_reg_dataout_328_port, 
      DataPath_RF_bus_reg_dataout_329_port, 
      DataPath_RF_bus_reg_dataout_330_port, 
      DataPath_RF_bus_reg_dataout_331_port, 
      DataPath_RF_bus_reg_dataout_332_port, 
      DataPath_RF_bus_reg_dataout_333_port, 
      DataPath_RF_bus_reg_dataout_334_port, 
      DataPath_RF_bus_reg_dataout_335_port, 
      DataPath_RF_bus_reg_dataout_336_port, 
      DataPath_RF_bus_reg_dataout_337_port, 
      DataPath_RF_bus_reg_dataout_338_port, 
      DataPath_RF_bus_reg_dataout_339_port, 
      DataPath_RF_bus_reg_dataout_340_port, 
      DataPath_RF_bus_reg_dataout_341_port, 
      DataPath_RF_bus_reg_dataout_342_port, 
      DataPath_RF_bus_reg_dataout_343_port, 
      DataPath_RF_bus_reg_dataout_344_port, 
      DataPath_RF_bus_reg_dataout_345_port, 
      DataPath_RF_bus_reg_dataout_346_port, 
      DataPath_RF_bus_reg_dataout_347_port, 
      DataPath_RF_bus_reg_dataout_348_port, 
      DataPath_RF_bus_reg_dataout_349_port, 
      DataPath_RF_bus_reg_dataout_350_port, 
      DataPath_RF_bus_reg_dataout_351_port, 
      DataPath_RF_bus_reg_dataout_352_port, 
      DataPath_RF_bus_reg_dataout_353_port, 
      DataPath_RF_bus_reg_dataout_354_port, 
      DataPath_RF_bus_reg_dataout_355_port, 
      DataPath_RF_bus_reg_dataout_356_port, 
      DataPath_RF_bus_reg_dataout_357_port, 
      DataPath_RF_bus_reg_dataout_358_port, 
      DataPath_RF_bus_reg_dataout_359_port, 
      DataPath_RF_bus_reg_dataout_360_port, 
      DataPath_RF_bus_reg_dataout_361_port, 
      DataPath_RF_bus_reg_dataout_362_port, 
      DataPath_RF_bus_reg_dataout_363_port, 
      DataPath_RF_bus_reg_dataout_364_port, 
      DataPath_RF_bus_reg_dataout_365_port, 
      DataPath_RF_bus_reg_dataout_366_port, 
      DataPath_RF_bus_reg_dataout_367_port, 
      DataPath_RF_bus_reg_dataout_368_port, 
      DataPath_RF_bus_reg_dataout_369_port, 
      DataPath_RF_bus_reg_dataout_370_port, 
      DataPath_RF_bus_reg_dataout_371_port, 
      DataPath_RF_bus_reg_dataout_372_port, 
      DataPath_RF_bus_reg_dataout_373_port, 
      DataPath_RF_bus_reg_dataout_374_port, 
      DataPath_RF_bus_reg_dataout_375_port, 
      DataPath_RF_bus_reg_dataout_376_port, 
      DataPath_RF_bus_reg_dataout_377_port, 
      DataPath_RF_bus_reg_dataout_378_port, 
      DataPath_RF_bus_reg_dataout_379_port, 
      DataPath_RF_bus_reg_dataout_380_port, 
      DataPath_RF_bus_reg_dataout_381_port, 
      DataPath_RF_bus_reg_dataout_382_port, 
      DataPath_RF_bus_reg_dataout_383_port, 
      DataPath_RF_bus_reg_dataout_384_port, 
      DataPath_RF_bus_reg_dataout_385_port, 
      DataPath_RF_bus_reg_dataout_386_port, 
      DataPath_RF_bus_reg_dataout_387_port, 
      DataPath_RF_bus_reg_dataout_388_port, 
      DataPath_RF_bus_reg_dataout_389_port, 
      DataPath_RF_bus_reg_dataout_390_port, 
      DataPath_RF_bus_reg_dataout_391_port, 
      DataPath_RF_bus_reg_dataout_392_port, 
      DataPath_RF_bus_reg_dataout_393_port, 
      DataPath_RF_bus_reg_dataout_394_port, 
      DataPath_RF_bus_reg_dataout_395_port, 
      DataPath_RF_bus_reg_dataout_396_port, 
      DataPath_RF_bus_reg_dataout_397_port, 
      DataPath_RF_bus_reg_dataout_398_port, 
      DataPath_RF_bus_reg_dataout_399_port, 
      DataPath_RF_bus_reg_dataout_400_port, 
      DataPath_RF_bus_reg_dataout_401_port, 
      DataPath_RF_bus_reg_dataout_402_port, 
      DataPath_RF_bus_reg_dataout_403_port, 
      DataPath_RF_bus_reg_dataout_404_port, 
      DataPath_RF_bus_reg_dataout_405_port, 
      DataPath_RF_bus_reg_dataout_406_port, 
      DataPath_RF_bus_reg_dataout_407_port, 
      DataPath_RF_bus_reg_dataout_408_port, 
      DataPath_RF_bus_reg_dataout_409_port, 
      DataPath_RF_bus_reg_dataout_410_port, 
      DataPath_RF_bus_reg_dataout_411_port, 
      DataPath_RF_bus_reg_dataout_412_port, 
      DataPath_RF_bus_reg_dataout_413_port, 
      DataPath_RF_bus_reg_dataout_414_port, 
      DataPath_RF_bus_reg_dataout_415_port, 
      DataPath_RF_bus_reg_dataout_416_port, 
      DataPath_RF_bus_reg_dataout_417_port, 
      DataPath_RF_bus_reg_dataout_418_port, 
      DataPath_RF_bus_reg_dataout_419_port, 
      DataPath_RF_bus_reg_dataout_420_port, 
      DataPath_RF_bus_reg_dataout_421_port, 
      DataPath_RF_bus_reg_dataout_422_port, 
      DataPath_RF_bus_reg_dataout_423_port, 
      DataPath_RF_bus_reg_dataout_424_port, 
      DataPath_RF_bus_reg_dataout_425_port, 
      DataPath_RF_bus_reg_dataout_426_port, 
      DataPath_RF_bus_reg_dataout_427_port, 
      DataPath_RF_bus_reg_dataout_428_port, 
      DataPath_RF_bus_reg_dataout_429_port, 
      DataPath_RF_bus_reg_dataout_430_port, 
      DataPath_RF_bus_reg_dataout_431_port, 
      DataPath_RF_bus_reg_dataout_432_port, 
      DataPath_RF_bus_reg_dataout_433_port, 
      DataPath_RF_bus_reg_dataout_434_port, 
      DataPath_RF_bus_reg_dataout_435_port, 
      DataPath_RF_bus_reg_dataout_436_port, 
      DataPath_RF_bus_reg_dataout_437_port, 
      DataPath_RF_bus_reg_dataout_438_port, 
      DataPath_RF_bus_reg_dataout_439_port, 
      DataPath_RF_bus_reg_dataout_440_port, 
      DataPath_RF_bus_reg_dataout_441_port, 
      DataPath_RF_bus_reg_dataout_442_port, 
      DataPath_RF_bus_reg_dataout_443_port, 
      DataPath_RF_bus_reg_dataout_444_port, 
      DataPath_RF_bus_reg_dataout_445_port, 
      DataPath_RF_bus_reg_dataout_446_port, 
      DataPath_RF_bus_reg_dataout_447_port, 
      DataPath_RF_bus_reg_dataout_448_port, 
      DataPath_RF_bus_reg_dataout_449_port, 
      DataPath_RF_bus_reg_dataout_450_port, 
      DataPath_RF_bus_reg_dataout_451_port, 
      DataPath_RF_bus_reg_dataout_452_port, 
      DataPath_RF_bus_reg_dataout_453_port, 
      DataPath_RF_bus_reg_dataout_454_port, 
      DataPath_RF_bus_reg_dataout_455_port, 
      DataPath_RF_bus_reg_dataout_456_port, 
      DataPath_RF_bus_reg_dataout_457_port, 
      DataPath_RF_bus_reg_dataout_458_port, 
      DataPath_RF_bus_reg_dataout_459_port, 
      DataPath_RF_bus_reg_dataout_460_port, 
      DataPath_RF_bus_reg_dataout_461_port, 
      DataPath_RF_bus_reg_dataout_462_port, 
      DataPath_RF_bus_reg_dataout_463_port, 
      DataPath_RF_bus_reg_dataout_464_port, 
      DataPath_RF_bus_reg_dataout_465_port, 
      DataPath_RF_bus_reg_dataout_466_port, 
      DataPath_RF_bus_reg_dataout_467_port, 
      DataPath_RF_bus_reg_dataout_468_port, 
      DataPath_RF_bus_reg_dataout_469_port, 
      DataPath_RF_bus_reg_dataout_470_port, 
      DataPath_RF_bus_reg_dataout_471_port, 
      DataPath_RF_bus_reg_dataout_472_port, 
      DataPath_RF_bus_reg_dataout_473_port, 
      DataPath_RF_bus_reg_dataout_474_port, 
      DataPath_RF_bus_reg_dataout_475_port, 
      DataPath_RF_bus_reg_dataout_476_port, 
      DataPath_RF_bus_reg_dataout_477_port, 
      DataPath_RF_bus_reg_dataout_478_port, 
      DataPath_RF_bus_reg_dataout_479_port, 
      DataPath_RF_bus_reg_dataout_480_port, 
      DataPath_RF_bus_reg_dataout_481_port, 
      DataPath_RF_bus_reg_dataout_482_port, 
      DataPath_RF_bus_reg_dataout_483_port, 
      DataPath_RF_bus_reg_dataout_484_port, 
      DataPath_RF_bus_reg_dataout_485_port, 
      DataPath_RF_bus_reg_dataout_486_port, 
      DataPath_RF_bus_reg_dataout_487_port, 
      DataPath_RF_bus_reg_dataout_488_port, 
      DataPath_RF_bus_reg_dataout_489_port, 
      DataPath_RF_bus_reg_dataout_490_port, 
      DataPath_RF_bus_reg_dataout_491_port, 
      DataPath_RF_bus_reg_dataout_492_port, 
      DataPath_RF_bus_reg_dataout_493_port, 
      DataPath_RF_bus_reg_dataout_494_port, 
      DataPath_RF_bus_reg_dataout_495_port, 
      DataPath_RF_bus_reg_dataout_496_port, 
      DataPath_RF_bus_reg_dataout_497_port, 
      DataPath_RF_bus_reg_dataout_498_port, 
      DataPath_RF_bus_reg_dataout_499_port, 
      DataPath_RF_bus_reg_dataout_500_port, 
      DataPath_RF_bus_reg_dataout_501_port, 
      DataPath_RF_bus_reg_dataout_502_port, 
      DataPath_RF_bus_reg_dataout_503_port, 
      DataPath_RF_bus_reg_dataout_504_port, 
      DataPath_RF_bus_reg_dataout_505_port, 
      DataPath_RF_bus_reg_dataout_506_port, 
      DataPath_RF_bus_reg_dataout_507_port, 
      DataPath_RF_bus_reg_dataout_508_port, 
      DataPath_RF_bus_reg_dataout_509_port, 
      DataPath_RF_bus_reg_dataout_510_port, 
      DataPath_RF_bus_reg_dataout_511_port, 
      DataPath_RF_bus_reg_dataout_512_port, 
      DataPath_RF_bus_reg_dataout_513_port, 
      DataPath_RF_bus_reg_dataout_514_port, 
      DataPath_RF_bus_reg_dataout_515_port, 
      DataPath_RF_bus_reg_dataout_516_port, 
      DataPath_RF_bus_reg_dataout_517_port, 
      DataPath_RF_bus_reg_dataout_518_port, 
      DataPath_RF_bus_reg_dataout_519_port, 
      DataPath_RF_bus_reg_dataout_520_port, 
      DataPath_RF_bus_reg_dataout_521_port, 
      DataPath_RF_bus_reg_dataout_522_port, 
      DataPath_RF_bus_reg_dataout_523_port, 
      DataPath_RF_bus_reg_dataout_524_port, 
      DataPath_RF_bus_reg_dataout_525_port, 
      DataPath_RF_bus_reg_dataout_526_port, 
      DataPath_RF_bus_reg_dataout_527_port, 
      DataPath_RF_bus_reg_dataout_528_port, 
      DataPath_RF_bus_reg_dataout_529_port, 
      DataPath_RF_bus_reg_dataout_530_port, 
      DataPath_RF_bus_reg_dataout_531_port, 
      DataPath_RF_bus_reg_dataout_532_port, 
      DataPath_RF_bus_reg_dataout_533_port, 
      DataPath_RF_bus_reg_dataout_534_port, 
      DataPath_RF_bus_reg_dataout_535_port, 
      DataPath_RF_bus_reg_dataout_536_port, 
      DataPath_RF_bus_reg_dataout_537_port, 
      DataPath_RF_bus_reg_dataout_538_port, 
      DataPath_RF_bus_reg_dataout_539_port, 
      DataPath_RF_bus_reg_dataout_540_port, 
      DataPath_RF_bus_reg_dataout_541_port, 
      DataPath_RF_bus_reg_dataout_542_port, 
      DataPath_RF_bus_reg_dataout_543_port, 
      DataPath_RF_bus_reg_dataout_544_port, 
      DataPath_RF_bus_reg_dataout_545_port, 
      DataPath_RF_bus_reg_dataout_546_port, 
      DataPath_RF_bus_reg_dataout_547_port, 
      DataPath_RF_bus_reg_dataout_548_port, 
      DataPath_RF_bus_reg_dataout_549_port, 
      DataPath_RF_bus_reg_dataout_550_port, 
      DataPath_RF_bus_reg_dataout_551_port, 
      DataPath_RF_bus_reg_dataout_552_port, 
      DataPath_RF_bus_reg_dataout_553_port, 
      DataPath_RF_bus_reg_dataout_554_port, 
      DataPath_RF_bus_reg_dataout_555_port, 
      DataPath_RF_bus_reg_dataout_556_port, 
      DataPath_RF_bus_reg_dataout_557_port, 
      DataPath_RF_bus_reg_dataout_558_port, 
      DataPath_RF_bus_reg_dataout_559_port, 
      DataPath_RF_bus_reg_dataout_560_port, 
      DataPath_RF_bus_reg_dataout_561_port, 
      DataPath_RF_bus_reg_dataout_562_port, 
      DataPath_RF_bus_reg_dataout_563_port, 
      DataPath_RF_bus_reg_dataout_564_port, 
      DataPath_RF_bus_reg_dataout_565_port, 
      DataPath_RF_bus_reg_dataout_566_port, 
      DataPath_RF_bus_reg_dataout_567_port, 
      DataPath_RF_bus_reg_dataout_568_port, 
      DataPath_RF_bus_reg_dataout_569_port, 
      DataPath_RF_bus_reg_dataout_570_port, 
      DataPath_RF_bus_reg_dataout_571_port, 
      DataPath_RF_bus_reg_dataout_572_port, 
      DataPath_RF_bus_reg_dataout_573_port, 
      DataPath_RF_bus_reg_dataout_574_port, 
      DataPath_RF_bus_reg_dataout_575_port, 
      DataPath_RF_bus_reg_dataout_576_port, 
      DataPath_RF_bus_reg_dataout_577_port, 
      DataPath_RF_bus_reg_dataout_578_port, 
      DataPath_RF_bus_reg_dataout_579_port, 
      DataPath_RF_bus_reg_dataout_580_port, 
      DataPath_RF_bus_reg_dataout_581_port, 
      DataPath_RF_bus_reg_dataout_582_port, 
      DataPath_RF_bus_reg_dataout_583_port, 
      DataPath_RF_bus_reg_dataout_584_port, 
      DataPath_RF_bus_reg_dataout_585_port, 
      DataPath_RF_bus_reg_dataout_586_port, 
      DataPath_RF_bus_reg_dataout_587_port, 
      DataPath_RF_bus_reg_dataout_588_port, 
      DataPath_RF_bus_reg_dataout_589_port, 
      DataPath_RF_bus_reg_dataout_590_port, 
      DataPath_RF_bus_reg_dataout_591_port, 
      DataPath_RF_bus_reg_dataout_592_port, 
      DataPath_RF_bus_reg_dataout_593_port, 
      DataPath_RF_bus_reg_dataout_594_port, 
      DataPath_RF_bus_reg_dataout_595_port, 
      DataPath_RF_bus_reg_dataout_596_port, 
      DataPath_RF_bus_reg_dataout_597_port, 
      DataPath_RF_bus_reg_dataout_598_port, 
      DataPath_RF_bus_reg_dataout_599_port, 
      DataPath_RF_bus_reg_dataout_600_port, 
      DataPath_RF_bus_reg_dataout_601_port, 
      DataPath_RF_bus_reg_dataout_602_port, 
      DataPath_RF_bus_reg_dataout_603_port, 
      DataPath_RF_bus_reg_dataout_604_port, 
      DataPath_RF_bus_reg_dataout_605_port, 
      DataPath_RF_bus_reg_dataout_606_port, 
      DataPath_RF_bus_reg_dataout_607_port, 
      DataPath_RF_bus_reg_dataout_608_port, 
      DataPath_RF_bus_reg_dataout_609_port, 
      DataPath_RF_bus_reg_dataout_610_port, 
      DataPath_RF_bus_reg_dataout_611_port, 
      DataPath_RF_bus_reg_dataout_612_port, 
      DataPath_RF_bus_reg_dataout_613_port, 
      DataPath_RF_bus_reg_dataout_614_port, 
      DataPath_RF_bus_reg_dataout_615_port, 
      DataPath_RF_bus_reg_dataout_616_port, 
      DataPath_RF_bus_reg_dataout_617_port, 
      DataPath_RF_bus_reg_dataout_618_port, 
      DataPath_RF_bus_reg_dataout_619_port, 
      DataPath_RF_bus_reg_dataout_620_port, 
      DataPath_RF_bus_reg_dataout_621_port, 
      DataPath_RF_bus_reg_dataout_622_port, 
      DataPath_RF_bus_reg_dataout_623_port, 
      DataPath_RF_bus_reg_dataout_624_port, 
      DataPath_RF_bus_reg_dataout_625_port, 
      DataPath_RF_bus_reg_dataout_626_port, 
      DataPath_RF_bus_reg_dataout_627_port, 
      DataPath_RF_bus_reg_dataout_628_port, 
      DataPath_RF_bus_reg_dataout_629_port, 
      DataPath_RF_bus_reg_dataout_630_port, 
      DataPath_RF_bus_reg_dataout_631_port, 
      DataPath_RF_bus_reg_dataout_632_port, 
      DataPath_RF_bus_reg_dataout_633_port, 
      DataPath_RF_bus_reg_dataout_634_port, 
      DataPath_RF_bus_reg_dataout_635_port, 
      DataPath_RF_bus_reg_dataout_636_port, 
      DataPath_RF_bus_reg_dataout_637_port, 
      DataPath_RF_bus_reg_dataout_638_port, 
      DataPath_RF_bus_reg_dataout_639_port, 
      DataPath_RF_bus_reg_dataout_640_port, 
      DataPath_RF_bus_reg_dataout_641_port, 
      DataPath_RF_bus_reg_dataout_642_port, 
      DataPath_RF_bus_reg_dataout_643_port, 
      DataPath_RF_bus_reg_dataout_644_port, 
      DataPath_RF_bus_reg_dataout_645_port, 
      DataPath_RF_bus_reg_dataout_646_port, 
      DataPath_RF_bus_reg_dataout_647_port, 
      DataPath_RF_bus_reg_dataout_648_port, 
      DataPath_RF_bus_reg_dataout_649_port, 
      DataPath_RF_bus_reg_dataout_650_port, 
      DataPath_RF_bus_reg_dataout_651_port, 
      DataPath_RF_bus_reg_dataout_652_port, 
      DataPath_RF_bus_reg_dataout_653_port, 
      DataPath_RF_bus_reg_dataout_654_port, 
      DataPath_RF_bus_reg_dataout_655_port, 
      DataPath_RF_bus_reg_dataout_656_port, 
      DataPath_RF_bus_reg_dataout_657_port, 
      DataPath_RF_bus_reg_dataout_658_port, 
      DataPath_RF_bus_reg_dataout_659_port, 
      DataPath_RF_bus_reg_dataout_660_port, 
      DataPath_RF_bus_reg_dataout_661_port, 
      DataPath_RF_bus_reg_dataout_662_port, 
      DataPath_RF_bus_reg_dataout_663_port, 
      DataPath_RF_bus_reg_dataout_664_port, 
      DataPath_RF_bus_reg_dataout_665_port, 
      DataPath_RF_bus_reg_dataout_666_port, 
      DataPath_RF_bus_reg_dataout_667_port, 
      DataPath_RF_bus_reg_dataout_668_port, 
      DataPath_RF_bus_reg_dataout_669_port, 
      DataPath_RF_bus_reg_dataout_670_port, 
      DataPath_RF_bus_reg_dataout_671_port, 
      DataPath_RF_bus_reg_dataout_672_port, 
      DataPath_RF_bus_reg_dataout_673_port, 
      DataPath_RF_bus_reg_dataout_674_port, 
      DataPath_RF_bus_reg_dataout_675_port, 
      DataPath_RF_bus_reg_dataout_676_port, 
      DataPath_RF_bus_reg_dataout_677_port, 
      DataPath_RF_bus_reg_dataout_678_port, 
      DataPath_RF_bus_reg_dataout_679_port, 
      DataPath_RF_bus_reg_dataout_680_port, 
      DataPath_RF_bus_reg_dataout_681_port, 
      DataPath_RF_bus_reg_dataout_682_port, 
      DataPath_RF_bus_reg_dataout_683_port, 
      DataPath_RF_bus_reg_dataout_684_port, 
      DataPath_RF_bus_reg_dataout_685_port, 
      DataPath_RF_bus_reg_dataout_686_port, 
      DataPath_RF_bus_reg_dataout_687_port, 
      DataPath_RF_bus_reg_dataout_688_port, 
      DataPath_RF_bus_reg_dataout_689_port, 
      DataPath_RF_bus_reg_dataout_690_port, 
      DataPath_RF_bus_reg_dataout_691_port, 
      DataPath_RF_bus_reg_dataout_692_port, 
      DataPath_RF_bus_reg_dataout_693_port, 
      DataPath_RF_bus_reg_dataout_694_port, 
      DataPath_RF_bus_reg_dataout_695_port, 
      DataPath_RF_bus_reg_dataout_696_port, 
      DataPath_RF_bus_reg_dataout_697_port, 
      DataPath_RF_bus_reg_dataout_698_port, 
      DataPath_RF_bus_reg_dataout_699_port, 
      DataPath_RF_bus_reg_dataout_700_port, 
      DataPath_RF_bus_reg_dataout_701_port, 
      DataPath_RF_bus_reg_dataout_702_port, 
      DataPath_RF_bus_reg_dataout_703_port, 
      DataPath_RF_bus_reg_dataout_704_port, 
      DataPath_RF_bus_reg_dataout_705_port, 
      DataPath_RF_bus_reg_dataout_706_port, 
      DataPath_RF_bus_reg_dataout_707_port, 
      DataPath_RF_bus_reg_dataout_708_port, 
      DataPath_RF_bus_reg_dataout_709_port, 
      DataPath_RF_bus_reg_dataout_710_port, 
      DataPath_RF_bus_reg_dataout_711_port, 
      DataPath_RF_bus_reg_dataout_712_port, 
      DataPath_RF_bus_reg_dataout_713_port, 
      DataPath_RF_bus_reg_dataout_714_port, 
      DataPath_RF_bus_reg_dataout_715_port, 
      DataPath_RF_bus_reg_dataout_716_port, 
      DataPath_RF_bus_reg_dataout_717_port, 
      DataPath_RF_bus_reg_dataout_718_port, 
      DataPath_RF_bus_reg_dataout_719_port, 
      DataPath_RF_bus_reg_dataout_720_port, 
      DataPath_RF_bus_reg_dataout_721_port, 
      DataPath_RF_bus_reg_dataout_722_port, 
      DataPath_RF_bus_reg_dataout_723_port, 
      DataPath_RF_bus_reg_dataout_724_port, 
      DataPath_RF_bus_reg_dataout_725_port, 
      DataPath_RF_bus_reg_dataout_726_port, 
      DataPath_RF_bus_reg_dataout_727_port, 
      DataPath_RF_bus_reg_dataout_728_port, 
      DataPath_RF_bus_reg_dataout_729_port, 
      DataPath_RF_bus_reg_dataout_730_port, 
      DataPath_RF_bus_reg_dataout_731_port, 
      DataPath_RF_bus_reg_dataout_732_port, 
      DataPath_RF_bus_reg_dataout_733_port, 
      DataPath_RF_bus_reg_dataout_734_port, 
      DataPath_RF_bus_reg_dataout_735_port, 
      DataPath_RF_bus_reg_dataout_736_port, 
      DataPath_RF_bus_reg_dataout_737_port, 
      DataPath_RF_bus_reg_dataout_738_port, 
      DataPath_RF_bus_reg_dataout_739_port, 
      DataPath_RF_bus_reg_dataout_740_port, 
      DataPath_RF_bus_reg_dataout_741_port, 
      DataPath_RF_bus_reg_dataout_742_port, 
      DataPath_RF_bus_reg_dataout_743_port, 
      DataPath_RF_bus_reg_dataout_744_port, 
      DataPath_RF_bus_reg_dataout_745_port, 
      DataPath_RF_bus_reg_dataout_746_port, 
      DataPath_RF_bus_reg_dataout_747_port, 
      DataPath_RF_bus_reg_dataout_748_port, 
      DataPath_RF_bus_reg_dataout_749_port, 
      DataPath_RF_bus_reg_dataout_750_port, 
      DataPath_RF_bus_reg_dataout_751_port, 
      DataPath_RF_bus_reg_dataout_752_port, 
      DataPath_RF_bus_reg_dataout_753_port, 
      DataPath_RF_bus_reg_dataout_754_port, 
      DataPath_RF_bus_reg_dataout_755_port, 
      DataPath_RF_bus_reg_dataout_756_port, 
      DataPath_RF_bus_reg_dataout_757_port, 
      DataPath_RF_bus_reg_dataout_758_port, 
      DataPath_RF_bus_reg_dataout_759_port, 
      DataPath_RF_bus_reg_dataout_760_port, 
      DataPath_RF_bus_reg_dataout_761_port, 
      DataPath_RF_bus_reg_dataout_762_port, 
      DataPath_RF_bus_reg_dataout_763_port, 
      DataPath_RF_bus_reg_dataout_764_port, 
      DataPath_RF_bus_reg_dataout_765_port, 
      DataPath_RF_bus_reg_dataout_766_port, 
      DataPath_RF_bus_reg_dataout_767_port, 
      DataPath_RF_bus_reg_dataout_768_port, 
      DataPath_RF_bus_reg_dataout_769_port, 
      DataPath_RF_bus_reg_dataout_770_port, 
      DataPath_RF_bus_reg_dataout_771_port, 
      DataPath_RF_bus_reg_dataout_772_port, 
      DataPath_RF_bus_reg_dataout_773_port, 
      DataPath_RF_bus_reg_dataout_774_port, 
      DataPath_RF_bus_reg_dataout_775_port, 
      DataPath_RF_bus_reg_dataout_776_port, 
      DataPath_RF_bus_reg_dataout_777_port, 
      DataPath_RF_bus_reg_dataout_778_port, 
      DataPath_RF_bus_reg_dataout_779_port, 
      DataPath_RF_bus_reg_dataout_780_port, 
      DataPath_RF_bus_reg_dataout_781_port, 
      DataPath_RF_bus_reg_dataout_782_port, 
      DataPath_RF_bus_reg_dataout_783_port, 
      DataPath_RF_bus_reg_dataout_784_port, 
      DataPath_RF_bus_reg_dataout_785_port, 
      DataPath_RF_bus_reg_dataout_786_port, 
      DataPath_RF_bus_reg_dataout_787_port, 
      DataPath_RF_bus_reg_dataout_788_port, 
      DataPath_RF_bus_reg_dataout_789_port, 
      DataPath_RF_bus_reg_dataout_790_port, 
      DataPath_RF_bus_reg_dataout_791_port, 
      DataPath_RF_bus_reg_dataout_792_port, 
      DataPath_RF_bus_reg_dataout_793_port, 
      DataPath_RF_bus_reg_dataout_794_port, 
      DataPath_RF_bus_reg_dataout_795_port, 
      DataPath_RF_bus_reg_dataout_796_port, 
      DataPath_RF_bus_reg_dataout_797_port, 
      DataPath_RF_bus_reg_dataout_798_port, 
      DataPath_RF_bus_reg_dataout_799_port, 
      DataPath_RF_bus_reg_dataout_800_port, 
      DataPath_RF_bus_reg_dataout_801_port, 
      DataPath_RF_bus_reg_dataout_802_port, 
      DataPath_RF_bus_reg_dataout_803_port, 
      DataPath_RF_bus_reg_dataout_804_port, 
      DataPath_RF_bus_reg_dataout_805_port, 
      DataPath_RF_bus_reg_dataout_806_port, 
      DataPath_RF_bus_reg_dataout_807_port, 
      DataPath_RF_bus_reg_dataout_808_port, 
      DataPath_RF_bus_reg_dataout_809_port, 
      DataPath_RF_bus_reg_dataout_810_port, 
      DataPath_RF_bus_reg_dataout_811_port, 
      DataPath_RF_bus_reg_dataout_812_port, 
      DataPath_RF_bus_reg_dataout_813_port, 
      DataPath_RF_bus_reg_dataout_814_port, 
      DataPath_RF_bus_reg_dataout_815_port, 
      DataPath_RF_bus_reg_dataout_816_port, 
      DataPath_RF_bus_reg_dataout_817_port, 
      DataPath_RF_bus_reg_dataout_818_port, 
      DataPath_RF_bus_reg_dataout_819_port, 
      DataPath_RF_bus_reg_dataout_820_port, 
      DataPath_RF_bus_reg_dataout_821_port, 
      DataPath_RF_bus_reg_dataout_822_port, 
      DataPath_RF_bus_reg_dataout_823_port, 
      DataPath_RF_bus_reg_dataout_824_port, 
      DataPath_RF_bus_reg_dataout_825_port, 
      DataPath_RF_bus_reg_dataout_826_port, 
      DataPath_RF_bus_reg_dataout_827_port, 
      DataPath_RF_bus_reg_dataout_828_port, 
      DataPath_RF_bus_reg_dataout_829_port, 
      DataPath_RF_bus_reg_dataout_830_port, 
      DataPath_RF_bus_reg_dataout_831_port, 
      DataPath_RF_bus_reg_dataout_832_port, 
      DataPath_RF_bus_reg_dataout_833_port, 
      DataPath_RF_bus_reg_dataout_834_port, 
      DataPath_RF_bus_reg_dataout_835_port, 
      DataPath_RF_bus_reg_dataout_836_port, 
      DataPath_RF_bus_reg_dataout_837_port, 
      DataPath_RF_bus_reg_dataout_838_port, 
      DataPath_RF_bus_reg_dataout_839_port, 
      DataPath_RF_bus_reg_dataout_840_port, 
      DataPath_RF_bus_reg_dataout_841_port, 
      DataPath_RF_bus_reg_dataout_842_port, 
      DataPath_RF_bus_reg_dataout_843_port, 
      DataPath_RF_bus_reg_dataout_844_port, 
      DataPath_RF_bus_reg_dataout_845_port, 
      DataPath_RF_bus_reg_dataout_846_port, 
      DataPath_RF_bus_reg_dataout_847_port, 
      DataPath_RF_bus_reg_dataout_848_port, 
      DataPath_RF_bus_reg_dataout_849_port, 
      DataPath_RF_bus_reg_dataout_850_port, 
      DataPath_RF_bus_reg_dataout_851_port, 
      DataPath_RF_bus_reg_dataout_852_port, 
      DataPath_RF_bus_reg_dataout_853_port, 
      DataPath_RF_bus_reg_dataout_854_port, 
      DataPath_RF_bus_reg_dataout_855_port, 
      DataPath_RF_bus_reg_dataout_856_port, 
      DataPath_RF_bus_reg_dataout_857_port, 
      DataPath_RF_bus_reg_dataout_858_port, 
      DataPath_RF_bus_reg_dataout_859_port, 
      DataPath_RF_bus_reg_dataout_860_port, 
      DataPath_RF_bus_reg_dataout_861_port, 
      DataPath_RF_bus_reg_dataout_862_port, 
      DataPath_RF_bus_reg_dataout_863_port, 
      DataPath_RF_bus_reg_dataout_864_port, 
      DataPath_RF_bus_reg_dataout_865_port, 
      DataPath_RF_bus_reg_dataout_866_port, 
      DataPath_RF_bus_reg_dataout_867_port, 
      DataPath_RF_bus_reg_dataout_868_port, 
      DataPath_RF_bus_reg_dataout_869_port, 
      DataPath_RF_bus_reg_dataout_870_port, 
      DataPath_RF_bus_reg_dataout_871_port, 
      DataPath_RF_bus_reg_dataout_872_port, 
      DataPath_RF_bus_reg_dataout_873_port, 
      DataPath_RF_bus_reg_dataout_874_port, 
      DataPath_RF_bus_reg_dataout_875_port, 
      DataPath_RF_bus_reg_dataout_876_port, 
      DataPath_RF_bus_reg_dataout_877_port, 
      DataPath_RF_bus_reg_dataout_878_port, 
      DataPath_RF_bus_reg_dataout_879_port, 
      DataPath_RF_bus_reg_dataout_880_port, 
      DataPath_RF_bus_reg_dataout_881_port, 
      DataPath_RF_bus_reg_dataout_882_port, 
      DataPath_RF_bus_reg_dataout_883_port, 
      DataPath_RF_bus_reg_dataout_884_port, 
      DataPath_RF_bus_reg_dataout_885_port, 
      DataPath_RF_bus_reg_dataout_886_port, 
      DataPath_RF_bus_reg_dataout_887_port, 
      DataPath_RF_bus_reg_dataout_888_port, 
      DataPath_RF_bus_reg_dataout_889_port, 
      DataPath_RF_bus_reg_dataout_890_port, 
      DataPath_RF_bus_reg_dataout_891_port, 
      DataPath_RF_bus_reg_dataout_892_port, 
      DataPath_RF_bus_reg_dataout_893_port, 
      DataPath_RF_bus_reg_dataout_894_port, 
      DataPath_RF_bus_reg_dataout_895_port, 
      DataPath_RF_bus_reg_dataout_896_port, 
      DataPath_RF_bus_reg_dataout_897_port, 
      DataPath_RF_bus_reg_dataout_898_port, 
      DataPath_RF_bus_reg_dataout_899_port, 
      DataPath_RF_bus_reg_dataout_900_port, 
      DataPath_RF_bus_reg_dataout_901_port, 
      DataPath_RF_bus_reg_dataout_902_port, 
      DataPath_RF_bus_reg_dataout_903_port, 
      DataPath_RF_bus_reg_dataout_904_port, 
      DataPath_RF_bus_reg_dataout_905_port, 
      DataPath_RF_bus_reg_dataout_906_port, 
      DataPath_RF_bus_reg_dataout_907_port, 
      DataPath_RF_bus_reg_dataout_908_port, 
      DataPath_RF_bus_reg_dataout_909_port, 
      DataPath_RF_bus_reg_dataout_910_port, 
      DataPath_RF_bus_reg_dataout_911_port, 
      DataPath_RF_bus_reg_dataout_912_port, 
      DataPath_RF_bus_reg_dataout_913_port, 
      DataPath_RF_bus_reg_dataout_914_port, 
      DataPath_RF_bus_reg_dataout_915_port, 
      DataPath_RF_bus_reg_dataout_916_port, 
      DataPath_RF_bus_reg_dataout_917_port, 
      DataPath_RF_bus_reg_dataout_918_port, 
      DataPath_RF_bus_reg_dataout_919_port, 
      DataPath_RF_bus_reg_dataout_920_port, 
      DataPath_RF_bus_reg_dataout_921_port, 
      DataPath_RF_bus_reg_dataout_922_port, 
      DataPath_RF_bus_reg_dataout_923_port, 
      DataPath_RF_bus_reg_dataout_924_port, 
      DataPath_RF_bus_reg_dataout_925_port, 
      DataPath_RF_bus_reg_dataout_926_port, 
      DataPath_RF_bus_reg_dataout_927_port, 
      DataPath_RF_bus_reg_dataout_928_port, 
      DataPath_RF_bus_reg_dataout_929_port, 
      DataPath_RF_bus_reg_dataout_930_port, 
      DataPath_RF_bus_reg_dataout_931_port, 
      DataPath_RF_bus_reg_dataout_932_port, 
      DataPath_RF_bus_reg_dataout_933_port, 
      DataPath_RF_bus_reg_dataout_934_port, 
      DataPath_RF_bus_reg_dataout_935_port, 
      DataPath_RF_bus_reg_dataout_936_port, 
      DataPath_RF_bus_reg_dataout_937_port, 
      DataPath_RF_bus_reg_dataout_938_port, 
      DataPath_RF_bus_reg_dataout_939_port, 
      DataPath_RF_bus_reg_dataout_940_port, 
      DataPath_RF_bus_reg_dataout_941_port, 
      DataPath_RF_bus_reg_dataout_942_port, 
      DataPath_RF_bus_reg_dataout_943_port, 
      DataPath_RF_bus_reg_dataout_944_port, 
      DataPath_RF_bus_reg_dataout_945_port, 
      DataPath_RF_bus_reg_dataout_946_port, 
      DataPath_RF_bus_reg_dataout_947_port, 
      DataPath_RF_bus_reg_dataout_948_port, 
      DataPath_RF_bus_reg_dataout_949_port, 
      DataPath_RF_bus_reg_dataout_950_port, 
      DataPath_RF_bus_reg_dataout_951_port, 
      DataPath_RF_bus_reg_dataout_952_port, 
      DataPath_RF_bus_reg_dataout_953_port, 
      DataPath_RF_bus_reg_dataout_954_port, 
      DataPath_RF_bus_reg_dataout_955_port, 
      DataPath_RF_bus_reg_dataout_956_port, 
      DataPath_RF_bus_reg_dataout_957_port, 
      DataPath_RF_bus_reg_dataout_958_port, 
      DataPath_RF_bus_reg_dataout_959_port, 
      DataPath_RF_bus_reg_dataout_960_port, 
      DataPath_RF_bus_reg_dataout_961_port, 
      DataPath_RF_bus_reg_dataout_962_port, 
      DataPath_RF_bus_reg_dataout_963_port, 
      DataPath_RF_bus_reg_dataout_964_port, 
      DataPath_RF_bus_reg_dataout_965_port, 
      DataPath_RF_bus_reg_dataout_966_port, 
      DataPath_RF_bus_reg_dataout_967_port, 
      DataPath_RF_bus_reg_dataout_968_port, 
      DataPath_RF_bus_reg_dataout_969_port, 
      DataPath_RF_bus_reg_dataout_970_port, 
      DataPath_RF_bus_reg_dataout_971_port, 
      DataPath_RF_bus_reg_dataout_972_port, 
      DataPath_RF_bus_reg_dataout_973_port, 
      DataPath_RF_bus_reg_dataout_974_port, 
      DataPath_RF_bus_reg_dataout_975_port, 
      DataPath_RF_bus_reg_dataout_976_port, 
      DataPath_RF_bus_reg_dataout_977_port, 
      DataPath_RF_bus_reg_dataout_978_port, 
      DataPath_RF_bus_reg_dataout_979_port, 
      DataPath_RF_bus_reg_dataout_980_port, 
      DataPath_RF_bus_reg_dataout_981_port, 
      DataPath_RF_bus_reg_dataout_982_port, 
      DataPath_RF_bus_reg_dataout_983_port, 
      DataPath_RF_bus_reg_dataout_984_port, 
      DataPath_RF_bus_reg_dataout_985_port, 
      DataPath_RF_bus_reg_dataout_986_port, 
      DataPath_RF_bus_reg_dataout_987_port, 
      DataPath_RF_bus_reg_dataout_988_port, 
      DataPath_RF_bus_reg_dataout_989_port, 
      DataPath_RF_bus_reg_dataout_990_port, 
      DataPath_RF_bus_reg_dataout_991_port, 
      DataPath_RF_bus_reg_dataout_992_port, 
      DataPath_RF_bus_reg_dataout_993_port, 
      DataPath_RF_bus_reg_dataout_994_port, 
      DataPath_RF_bus_reg_dataout_995_port, 
      DataPath_RF_bus_reg_dataout_996_port, 
      DataPath_RF_bus_reg_dataout_997_port, 
      DataPath_RF_bus_reg_dataout_998_port, 
      DataPath_RF_bus_reg_dataout_999_port, 
      DataPath_RF_bus_reg_dataout_1000_port, 
      DataPath_RF_bus_reg_dataout_1001_port, 
      DataPath_RF_bus_reg_dataout_1002_port, 
      DataPath_RF_bus_reg_dataout_1003_port, 
      DataPath_RF_bus_reg_dataout_1004_port, 
      DataPath_RF_bus_reg_dataout_1005_port, 
      DataPath_RF_bus_reg_dataout_1006_port, 
      DataPath_RF_bus_reg_dataout_1007_port, 
      DataPath_RF_bus_reg_dataout_1008_port, 
      DataPath_RF_bus_reg_dataout_1009_port, 
      DataPath_RF_bus_reg_dataout_1010_port, 
      DataPath_RF_bus_reg_dataout_1011_port, 
      DataPath_RF_bus_reg_dataout_1012_port, 
      DataPath_RF_bus_reg_dataout_1013_port, 
      DataPath_RF_bus_reg_dataout_1014_port, 
      DataPath_RF_bus_reg_dataout_1015_port, 
      DataPath_RF_bus_reg_dataout_1016_port, 
      DataPath_RF_bus_reg_dataout_1017_port, 
      DataPath_RF_bus_reg_dataout_1018_port, 
      DataPath_RF_bus_reg_dataout_1019_port, 
      DataPath_RF_bus_reg_dataout_1020_port, 
      DataPath_RF_bus_reg_dataout_1021_port, 
      DataPath_RF_bus_reg_dataout_1022_port, 
      DataPath_RF_bus_reg_dataout_1023_port, 
      DataPath_RF_bus_reg_dataout_1024_port, 
      DataPath_RF_bus_reg_dataout_1025_port, 
      DataPath_RF_bus_reg_dataout_1026_port, 
      DataPath_RF_bus_reg_dataout_1027_port, 
      DataPath_RF_bus_reg_dataout_1028_port, 
      DataPath_RF_bus_reg_dataout_1029_port, 
      DataPath_RF_bus_reg_dataout_1030_port, 
      DataPath_RF_bus_reg_dataout_1031_port, 
      DataPath_RF_bus_reg_dataout_1032_port, 
      DataPath_RF_bus_reg_dataout_1033_port, 
      DataPath_RF_bus_reg_dataout_1034_port, 
      DataPath_RF_bus_reg_dataout_1035_port, 
      DataPath_RF_bus_reg_dataout_1036_port, 
      DataPath_RF_bus_reg_dataout_1037_port, 
      DataPath_RF_bus_reg_dataout_1038_port, 
      DataPath_RF_bus_reg_dataout_1039_port, 
      DataPath_RF_bus_reg_dataout_1040_port, 
      DataPath_RF_bus_reg_dataout_1041_port, 
      DataPath_RF_bus_reg_dataout_1042_port, 
      DataPath_RF_bus_reg_dataout_1043_port, 
      DataPath_RF_bus_reg_dataout_1044_port, 
      DataPath_RF_bus_reg_dataout_1045_port, 
      DataPath_RF_bus_reg_dataout_1046_port, 
      DataPath_RF_bus_reg_dataout_1047_port, 
      DataPath_RF_bus_reg_dataout_1048_port, 
      DataPath_RF_bus_reg_dataout_1049_port, 
      DataPath_RF_bus_reg_dataout_1050_port, 
      DataPath_RF_bus_reg_dataout_1051_port, 
      DataPath_RF_bus_reg_dataout_1052_port, 
      DataPath_RF_bus_reg_dataout_1053_port, 
      DataPath_RF_bus_reg_dataout_1054_port, 
      DataPath_RF_bus_reg_dataout_1055_port, 
      DataPath_RF_bus_reg_dataout_1056_port, 
      DataPath_RF_bus_reg_dataout_1057_port, 
      DataPath_RF_bus_reg_dataout_1058_port, 
      DataPath_RF_bus_reg_dataout_1059_port, 
      DataPath_RF_bus_reg_dataout_1060_port, 
      DataPath_RF_bus_reg_dataout_1061_port, 
      DataPath_RF_bus_reg_dataout_1062_port, 
      DataPath_RF_bus_reg_dataout_1063_port, 
      DataPath_RF_bus_reg_dataout_1064_port, 
      DataPath_RF_bus_reg_dataout_1065_port, 
      DataPath_RF_bus_reg_dataout_1066_port, 
      DataPath_RF_bus_reg_dataout_1067_port, 
      DataPath_RF_bus_reg_dataout_1068_port, 
      DataPath_RF_bus_reg_dataout_1069_port, 
      DataPath_RF_bus_reg_dataout_1070_port, 
      DataPath_RF_bus_reg_dataout_1071_port, 
      DataPath_RF_bus_reg_dataout_1072_port, 
      DataPath_RF_bus_reg_dataout_1073_port, 
      DataPath_RF_bus_reg_dataout_1074_port, 
      DataPath_RF_bus_reg_dataout_1075_port, 
      DataPath_RF_bus_reg_dataout_1076_port, 
      DataPath_RF_bus_reg_dataout_1077_port, 
      DataPath_RF_bus_reg_dataout_1078_port, 
      DataPath_RF_bus_reg_dataout_1079_port, 
      DataPath_RF_bus_reg_dataout_1080_port, 
      DataPath_RF_bus_reg_dataout_1081_port, 
      DataPath_RF_bus_reg_dataout_1082_port, 
      DataPath_RF_bus_reg_dataout_1083_port, 
      DataPath_RF_bus_reg_dataout_1084_port, 
      DataPath_RF_bus_reg_dataout_1085_port, 
      DataPath_RF_bus_reg_dataout_1086_port, 
      DataPath_RF_bus_reg_dataout_1087_port, 
      DataPath_RF_bus_reg_dataout_1088_port, 
      DataPath_RF_bus_reg_dataout_1089_port, 
      DataPath_RF_bus_reg_dataout_1090_port, 
      DataPath_RF_bus_reg_dataout_1091_port, 
      DataPath_RF_bus_reg_dataout_1092_port, 
      DataPath_RF_bus_reg_dataout_1093_port, 
      DataPath_RF_bus_reg_dataout_1094_port, 
      DataPath_RF_bus_reg_dataout_1095_port, 
      DataPath_RF_bus_reg_dataout_1096_port, 
      DataPath_RF_bus_reg_dataout_1097_port, 
      DataPath_RF_bus_reg_dataout_1098_port, 
      DataPath_RF_bus_reg_dataout_1099_port, 
      DataPath_RF_bus_reg_dataout_1100_port, 
      DataPath_RF_bus_reg_dataout_1101_port, 
      DataPath_RF_bus_reg_dataout_1102_port, 
      DataPath_RF_bus_reg_dataout_1103_port, 
      DataPath_RF_bus_reg_dataout_1104_port, 
      DataPath_RF_bus_reg_dataout_1105_port, 
      DataPath_RF_bus_reg_dataout_1106_port, 
      DataPath_RF_bus_reg_dataout_1107_port, 
      DataPath_RF_bus_reg_dataout_1108_port, 
      DataPath_RF_bus_reg_dataout_1109_port, 
      DataPath_RF_bus_reg_dataout_1110_port, 
      DataPath_RF_bus_reg_dataout_1111_port, 
      DataPath_RF_bus_reg_dataout_1112_port, 
      DataPath_RF_bus_reg_dataout_1113_port, 
      DataPath_RF_bus_reg_dataout_1114_port, 
      DataPath_RF_bus_reg_dataout_1115_port, 
      DataPath_RF_bus_reg_dataout_1116_port, 
      DataPath_RF_bus_reg_dataout_1117_port, 
      DataPath_RF_bus_reg_dataout_1118_port, 
      DataPath_RF_bus_reg_dataout_1119_port, 
      DataPath_RF_bus_reg_dataout_1120_port, 
      DataPath_RF_bus_reg_dataout_1121_port, 
      DataPath_RF_bus_reg_dataout_1122_port, 
      DataPath_RF_bus_reg_dataout_1123_port, 
      DataPath_RF_bus_reg_dataout_1124_port, 
      DataPath_RF_bus_reg_dataout_1125_port, 
      DataPath_RF_bus_reg_dataout_1126_port, 
      DataPath_RF_bus_reg_dataout_1127_port, 
      DataPath_RF_bus_reg_dataout_1128_port, 
      DataPath_RF_bus_reg_dataout_1129_port, 
      DataPath_RF_bus_reg_dataout_1130_port, 
      DataPath_RF_bus_reg_dataout_1131_port, 
      DataPath_RF_bus_reg_dataout_1132_port, 
      DataPath_RF_bus_reg_dataout_1133_port, 
      DataPath_RF_bus_reg_dataout_1134_port, 
      DataPath_RF_bus_reg_dataout_1135_port, 
      DataPath_RF_bus_reg_dataout_1136_port, 
      DataPath_RF_bus_reg_dataout_1137_port, 
      DataPath_RF_bus_reg_dataout_1138_port, 
      DataPath_RF_bus_reg_dataout_1139_port, 
      DataPath_RF_bus_reg_dataout_1140_port, 
      DataPath_RF_bus_reg_dataout_1141_port, 
      DataPath_RF_bus_reg_dataout_1142_port, 
      DataPath_RF_bus_reg_dataout_1143_port, 
      DataPath_RF_bus_reg_dataout_1144_port, 
      DataPath_RF_bus_reg_dataout_1145_port, 
      DataPath_RF_bus_reg_dataout_1146_port, 
      DataPath_RF_bus_reg_dataout_1147_port, 
      DataPath_RF_bus_reg_dataout_1148_port, 
      DataPath_RF_bus_reg_dataout_1149_port, 
      DataPath_RF_bus_reg_dataout_1150_port, 
      DataPath_RF_bus_reg_dataout_1151_port, 
      DataPath_RF_bus_reg_dataout_1152_port, 
      DataPath_RF_bus_reg_dataout_1153_port, 
      DataPath_RF_bus_reg_dataout_1154_port, 
      DataPath_RF_bus_reg_dataout_1155_port, 
      DataPath_RF_bus_reg_dataout_1156_port, 
      DataPath_RF_bus_reg_dataout_1157_port, 
      DataPath_RF_bus_reg_dataout_1158_port, 
      DataPath_RF_bus_reg_dataout_1159_port, 
      DataPath_RF_bus_reg_dataout_1160_port, 
      DataPath_RF_bus_reg_dataout_1161_port, 
      DataPath_RF_bus_reg_dataout_1162_port, 
      DataPath_RF_bus_reg_dataout_1163_port, 
      DataPath_RF_bus_reg_dataout_1164_port, 
      DataPath_RF_bus_reg_dataout_1165_port, 
      DataPath_RF_bus_reg_dataout_1166_port, 
      DataPath_RF_bus_reg_dataout_1167_port, 
      DataPath_RF_bus_reg_dataout_1168_port, 
      DataPath_RF_bus_reg_dataout_1169_port, 
      DataPath_RF_bus_reg_dataout_1170_port, 
      DataPath_RF_bus_reg_dataout_1171_port, 
      DataPath_RF_bus_reg_dataout_1172_port, 
      DataPath_RF_bus_reg_dataout_1173_port, 
      DataPath_RF_bus_reg_dataout_1174_port, 
      DataPath_RF_bus_reg_dataout_1175_port, 
      DataPath_RF_bus_reg_dataout_1176_port, 
      DataPath_RF_bus_reg_dataout_1177_port, 
      DataPath_RF_bus_reg_dataout_1178_port, 
      DataPath_RF_bus_reg_dataout_1179_port, 
      DataPath_RF_bus_reg_dataout_1180_port, 
      DataPath_RF_bus_reg_dataout_1181_port, 
      DataPath_RF_bus_reg_dataout_1182_port, 
      DataPath_RF_bus_reg_dataout_1183_port, 
      DataPath_RF_bus_reg_dataout_1184_port, 
      DataPath_RF_bus_reg_dataout_1185_port, 
      DataPath_RF_bus_reg_dataout_1186_port, 
      DataPath_RF_bus_reg_dataout_1187_port, 
      DataPath_RF_bus_reg_dataout_1188_port, 
      DataPath_RF_bus_reg_dataout_1189_port, 
      DataPath_RF_bus_reg_dataout_1190_port, 
      DataPath_RF_bus_reg_dataout_1191_port, 
      DataPath_RF_bus_reg_dataout_1192_port, 
      DataPath_RF_bus_reg_dataout_1193_port, 
      DataPath_RF_bus_reg_dataout_1194_port, 
      DataPath_RF_bus_reg_dataout_1195_port, 
      DataPath_RF_bus_reg_dataout_1196_port, 
      DataPath_RF_bus_reg_dataout_1197_port, 
      DataPath_RF_bus_reg_dataout_1198_port, 
      DataPath_RF_bus_reg_dataout_1199_port, 
      DataPath_RF_bus_reg_dataout_1200_port, 
      DataPath_RF_bus_reg_dataout_1201_port, 
      DataPath_RF_bus_reg_dataout_1202_port, 
      DataPath_RF_bus_reg_dataout_1203_port, 
      DataPath_RF_bus_reg_dataout_1204_port, 
      DataPath_RF_bus_reg_dataout_1205_port, 
      DataPath_RF_bus_reg_dataout_1206_port, 
      DataPath_RF_bus_reg_dataout_1207_port, 
      DataPath_RF_bus_reg_dataout_1208_port, 
      DataPath_RF_bus_reg_dataout_1209_port, 
      DataPath_RF_bus_reg_dataout_1210_port, 
      DataPath_RF_bus_reg_dataout_1211_port, 
      DataPath_RF_bus_reg_dataout_1212_port, 
      DataPath_RF_bus_reg_dataout_1213_port, 
      DataPath_RF_bus_reg_dataout_1214_port, 
      DataPath_RF_bus_reg_dataout_1215_port, 
      DataPath_RF_bus_reg_dataout_1216_port, 
      DataPath_RF_bus_reg_dataout_1217_port, 
      DataPath_RF_bus_reg_dataout_1218_port, 
      DataPath_RF_bus_reg_dataout_1219_port, 
      DataPath_RF_bus_reg_dataout_1220_port, 
      DataPath_RF_bus_reg_dataout_1221_port, 
      DataPath_RF_bus_reg_dataout_1222_port, 
      DataPath_RF_bus_reg_dataout_1223_port, 
      DataPath_RF_bus_reg_dataout_1224_port, 
      DataPath_RF_bus_reg_dataout_1225_port, 
      DataPath_RF_bus_reg_dataout_1226_port, 
      DataPath_RF_bus_reg_dataout_1227_port, 
      DataPath_RF_bus_reg_dataout_1228_port, 
      DataPath_RF_bus_reg_dataout_1229_port, 
      DataPath_RF_bus_reg_dataout_1230_port, 
      DataPath_RF_bus_reg_dataout_1231_port, 
      DataPath_RF_bus_reg_dataout_1232_port, 
      DataPath_RF_bus_reg_dataout_1233_port, 
      DataPath_RF_bus_reg_dataout_1234_port, 
      DataPath_RF_bus_reg_dataout_1235_port, 
      DataPath_RF_bus_reg_dataout_1236_port, 
      DataPath_RF_bus_reg_dataout_1237_port, 
      DataPath_RF_bus_reg_dataout_1238_port, 
      DataPath_RF_bus_reg_dataout_1239_port, 
      DataPath_RF_bus_reg_dataout_1240_port, 
      DataPath_RF_bus_reg_dataout_1241_port, 
      DataPath_RF_bus_reg_dataout_1242_port, 
      DataPath_RF_bus_reg_dataout_1243_port, 
      DataPath_RF_bus_reg_dataout_1244_port, 
      DataPath_RF_bus_reg_dataout_1245_port, 
      DataPath_RF_bus_reg_dataout_1246_port, 
      DataPath_RF_bus_reg_dataout_1247_port, 
      DataPath_RF_bus_reg_dataout_1248_port, 
      DataPath_RF_bus_reg_dataout_1249_port, 
      DataPath_RF_bus_reg_dataout_1250_port, 
      DataPath_RF_bus_reg_dataout_1251_port, 
      DataPath_RF_bus_reg_dataout_1252_port, 
      DataPath_RF_bus_reg_dataout_1253_port, 
      DataPath_RF_bus_reg_dataout_1254_port, 
      DataPath_RF_bus_reg_dataout_1255_port, 
      DataPath_RF_bus_reg_dataout_1256_port, 
      DataPath_RF_bus_reg_dataout_1257_port, 
      DataPath_RF_bus_reg_dataout_1258_port, 
      DataPath_RF_bus_reg_dataout_1259_port, 
      DataPath_RF_bus_reg_dataout_1260_port, 
      DataPath_RF_bus_reg_dataout_1261_port, 
      DataPath_RF_bus_reg_dataout_1262_port, 
      DataPath_RF_bus_reg_dataout_1263_port, 
      DataPath_RF_bus_reg_dataout_1264_port, 
      DataPath_RF_bus_reg_dataout_1265_port, 
      DataPath_RF_bus_reg_dataout_1266_port, 
      DataPath_RF_bus_reg_dataout_1267_port, 
      DataPath_RF_bus_reg_dataout_1268_port, 
      DataPath_RF_bus_reg_dataout_1269_port, 
      DataPath_RF_bus_reg_dataout_1270_port, 
      DataPath_RF_bus_reg_dataout_1271_port, 
      DataPath_RF_bus_reg_dataout_1272_port, 
      DataPath_RF_bus_reg_dataout_1273_port, 
      DataPath_RF_bus_reg_dataout_1274_port, 
      DataPath_RF_bus_reg_dataout_1275_port, 
      DataPath_RF_bus_reg_dataout_1276_port, 
      DataPath_RF_bus_reg_dataout_1277_port, 
      DataPath_RF_bus_reg_dataout_1278_port, 
      DataPath_RF_bus_reg_dataout_1279_port, 
      DataPath_RF_bus_reg_dataout_1280_port, 
      DataPath_RF_bus_reg_dataout_1281_port, 
      DataPath_RF_bus_reg_dataout_1282_port, 
      DataPath_RF_bus_reg_dataout_1283_port, 
      DataPath_RF_bus_reg_dataout_1284_port, 
      DataPath_RF_bus_reg_dataout_1285_port, 
      DataPath_RF_bus_reg_dataout_1286_port, 
      DataPath_RF_bus_reg_dataout_1287_port, 
      DataPath_RF_bus_reg_dataout_1288_port, 
      DataPath_RF_bus_reg_dataout_1289_port, 
      DataPath_RF_bus_reg_dataout_1290_port, 
      DataPath_RF_bus_reg_dataout_1291_port, 
      DataPath_RF_bus_reg_dataout_1292_port, 
      DataPath_RF_bus_reg_dataout_1293_port, 
      DataPath_RF_bus_reg_dataout_1294_port, 
      DataPath_RF_bus_reg_dataout_1295_port, 
      DataPath_RF_bus_reg_dataout_1296_port, 
      DataPath_RF_bus_reg_dataout_1297_port, 
      DataPath_RF_bus_reg_dataout_1298_port, 
      DataPath_RF_bus_reg_dataout_1299_port, 
      DataPath_RF_bus_reg_dataout_1300_port, 
      DataPath_RF_bus_reg_dataout_1301_port, 
      DataPath_RF_bus_reg_dataout_1302_port, 
      DataPath_RF_bus_reg_dataout_1303_port, 
      DataPath_RF_bus_reg_dataout_1304_port, 
      DataPath_RF_bus_reg_dataout_1305_port, 
      DataPath_RF_bus_reg_dataout_1306_port, 
      DataPath_RF_bus_reg_dataout_1307_port, 
      DataPath_RF_bus_reg_dataout_1308_port, 
      DataPath_RF_bus_reg_dataout_1309_port, 
      DataPath_RF_bus_reg_dataout_1310_port, 
      DataPath_RF_bus_reg_dataout_1311_port, 
      DataPath_RF_bus_reg_dataout_1312_port, 
      DataPath_RF_bus_reg_dataout_1313_port, 
      DataPath_RF_bus_reg_dataout_1314_port, 
      DataPath_RF_bus_reg_dataout_1315_port, 
      DataPath_RF_bus_reg_dataout_1316_port, 
      DataPath_RF_bus_reg_dataout_1317_port, 
      DataPath_RF_bus_reg_dataout_1318_port, 
      DataPath_RF_bus_reg_dataout_1319_port, 
      DataPath_RF_bus_reg_dataout_1320_port, 
      DataPath_RF_bus_reg_dataout_1321_port, 
      DataPath_RF_bus_reg_dataout_1322_port, 
      DataPath_RF_bus_reg_dataout_1323_port, 
      DataPath_RF_bus_reg_dataout_1324_port, 
      DataPath_RF_bus_reg_dataout_1325_port, 
      DataPath_RF_bus_reg_dataout_1326_port, 
      DataPath_RF_bus_reg_dataout_1327_port, 
      DataPath_RF_bus_reg_dataout_1328_port, 
      DataPath_RF_bus_reg_dataout_1329_port, 
      DataPath_RF_bus_reg_dataout_1330_port, 
      DataPath_RF_bus_reg_dataout_1331_port, 
      DataPath_RF_bus_reg_dataout_1332_port, 
      DataPath_RF_bus_reg_dataout_1333_port, 
      DataPath_RF_bus_reg_dataout_1334_port, 
      DataPath_RF_bus_reg_dataout_1335_port, 
      DataPath_RF_bus_reg_dataout_1336_port, 
      DataPath_RF_bus_reg_dataout_1337_port, 
      DataPath_RF_bus_reg_dataout_1338_port, 
      DataPath_RF_bus_reg_dataout_1339_port, 
      DataPath_RF_bus_reg_dataout_1340_port, 
      DataPath_RF_bus_reg_dataout_1341_port, 
      DataPath_RF_bus_reg_dataout_1342_port, 
      DataPath_RF_bus_reg_dataout_1343_port, 
      DataPath_RF_bus_reg_dataout_1344_port, 
      DataPath_RF_bus_reg_dataout_1345_port, 
      DataPath_RF_bus_reg_dataout_1346_port, 
      DataPath_RF_bus_reg_dataout_1347_port, 
      DataPath_RF_bus_reg_dataout_1348_port, 
      DataPath_RF_bus_reg_dataout_1349_port, 
      DataPath_RF_bus_reg_dataout_1350_port, 
      DataPath_RF_bus_reg_dataout_1351_port, 
      DataPath_RF_bus_reg_dataout_1352_port, 
      DataPath_RF_bus_reg_dataout_1353_port, 
      DataPath_RF_bus_reg_dataout_1354_port, 
      DataPath_RF_bus_reg_dataout_1355_port, 
      DataPath_RF_bus_reg_dataout_1356_port, 
      DataPath_RF_bus_reg_dataout_1357_port, 
      DataPath_RF_bus_reg_dataout_1358_port, 
      DataPath_RF_bus_reg_dataout_1359_port, 
      DataPath_RF_bus_reg_dataout_1360_port, 
      DataPath_RF_bus_reg_dataout_1361_port, 
      DataPath_RF_bus_reg_dataout_1362_port, 
      DataPath_RF_bus_reg_dataout_1363_port, 
      DataPath_RF_bus_reg_dataout_1364_port, 
      DataPath_RF_bus_reg_dataout_1365_port, 
      DataPath_RF_bus_reg_dataout_1366_port, 
      DataPath_RF_bus_reg_dataout_1367_port, 
      DataPath_RF_bus_reg_dataout_1368_port, 
      DataPath_RF_bus_reg_dataout_1369_port, 
      DataPath_RF_bus_reg_dataout_1370_port, 
      DataPath_RF_bus_reg_dataout_1371_port, 
      DataPath_RF_bus_reg_dataout_1372_port, 
      DataPath_RF_bus_reg_dataout_1373_port, 
      DataPath_RF_bus_reg_dataout_1374_port, 
      DataPath_RF_bus_reg_dataout_1375_port, 
      DataPath_RF_bus_reg_dataout_1376_port, 
      DataPath_RF_bus_reg_dataout_1377_port, 
      DataPath_RF_bus_reg_dataout_1378_port, 
      DataPath_RF_bus_reg_dataout_1379_port, 
      DataPath_RF_bus_reg_dataout_1380_port, 
      DataPath_RF_bus_reg_dataout_1381_port, 
      DataPath_RF_bus_reg_dataout_1382_port, 
      DataPath_RF_bus_reg_dataout_1383_port, 
      DataPath_RF_bus_reg_dataout_1384_port, 
      DataPath_RF_bus_reg_dataout_1385_port, 
      DataPath_RF_bus_reg_dataout_1386_port, 
      DataPath_RF_bus_reg_dataout_1387_port, 
      DataPath_RF_bus_reg_dataout_1388_port, 
      DataPath_RF_bus_reg_dataout_1389_port, 
      DataPath_RF_bus_reg_dataout_1390_port, 
      DataPath_RF_bus_reg_dataout_1391_port, 
      DataPath_RF_bus_reg_dataout_1392_port, 
      DataPath_RF_bus_reg_dataout_1393_port, 
      DataPath_RF_bus_reg_dataout_1394_port, 
      DataPath_RF_bus_reg_dataout_1395_port, 
      DataPath_RF_bus_reg_dataout_1396_port, 
      DataPath_RF_bus_reg_dataout_1397_port, 
      DataPath_RF_bus_reg_dataout_1398_port, 
      DataPath_RF_bus_reg_dataout_1399_port, 
      DataPath_RF_bus_reg_dataout_1400_port, 
      DataPath_RF_bus_reg_dataout_1401_port, 
      DataPath_RF_bus_reg_dataout_1402_port, 
      DataPath_RF_bus_reg_dataout_1403_port, 
      DataPath_RF_bus_reg_dataout_1404_port, 
      DataPath_RF_bus_reg_dataout_1405_port, 
      DataPath_RF_bus_reg_dataout_1406_port, 
      DataPath_RF_bus_reg_dataout_1407_port, 
      DataPath_RF_bus_reg_dataout_1408_port, 
      DataPath_RF_bus_reg_dataout_1409_port, 
      DataPath_RF_bus_reg_dataout_1410_port, 
      DataPath_RF_bus_reg_dataout_1411_port, 
      DataPath_RF_bus_reg_dataout_1412_port, 
      DataPath_RF_bus_reg_dataout_1413_port, 
      DataPath_RF_bus_reg_dataout_1414_port, 
      DataPath_RF_bus_reg_dataout_1415_port, 
      DataPath_RF_bus_reg_dataout_1416_port, 
      DataPath_RF_bus_reg_dataout_1417_port, 
      DataPath_RF_bus_reg_dataout_1418_port, 
      DataPath_RF_bus_reg_dataout_1419_port, 
      DataPath_RF_bus_reg_dataout_1420_port, 
      DataPath_RF_bus_reg_dataout_1421_port, 
      DataPath_RF_bus_reg_dataout_1422_port, 
      DataPath_RF_bus_reg_dataout_1423_port, 
      DataPath_RF_bus_reg_dataout_1424_port, 
      DataPath_RF_bus_reg_dataout_1425_port, 
      DataPath_RF_bus_reg_dataout_1426_port, 
      DataPath_RF_bus_reg_dataout_1427_port, 
      DataPath_RF_bus_reg_dataout_1428_port, 
      DataPath_RF_bus_reg_dataout_1429_port, 
      DataPath_RF_bus_reg_dataout_1430_port, 
      DataPath_RF_bus_reg_dataout_1431_port, 
      DataPath_RF_bus_reg_dataout_1432_port, 
      DataPath_RF_bus_reg_dataout_1433_port, 
      DataPath_RF_bus_reg_dataout_1434_port, 
      DataPath_RF_bus_reg_dataout_1435_port, 
      DataPath_RF_bus_reg_dataout_1436_port, 
      DataPath_RF_bus_reg_dataout_1437_port, 
      DataPath_RF_bus_reg_dataout_1438_port, 
      DataPath_RF_bus_reg_dataout_1439_port, 
      DataPath_RF_bus_reg_dataout_1440_port, 
      DataPath_RF_bus_reg_dataout_1441_port, 
      DataPath_RF_bus_reg_dataout_1442_port, 
      DataPath_RF_bus_reg_dataout_1443_port, 
      DataPath_RF_bus_reg_dataout_1444_port, 
      DataPath_RF_bus_reg_dataout_1445_port, 
      DataPath_RF_bus_reg_dataout_1446_port, 
      DataPath_RF_bus_reg_dataout_1447_port, 
      DataPath_RF_bus_reg_dataout_1448_port, 
      DataPath_RF_bus_reg_dataout_1449_port, 
      DataPath_RF_bus_reg_dataout_1450_port, 
      DataPath_RF_bus_reg_dataout_1451_port, 
      DataPath_RF_bus_reg_dataout_1452_port, 
      DataPath_RF_bus_reg_dataout_1453_port, 
      DataPath_RF_bus_reg_dataout_1454_port, 
      DataPath_RF_bus_reg_dataout_1455_port, 
      DataPath_RF_bus_reg_dataout_1456_port, 
      DataPath_RF_bus_reg_dataout_1457_port, 
      DataPath_RF_bus_reg_dataout_1458_port, 
      DataPath_RF_bus_reg_dataout_1459_port, 
      DataPath_RF_bus_reg_dataout_1460_port, 
      DataPath_RF_bus_reg_dataout_1461_port, 
      DataPath_RF_bus_reg_dataout_1462_port, 
      DataPath_RF_bus_reg_dataout_1463_port, 
      DataPath_RF_bus_reg_dataout_1464_port, 
      DataPath_RF_bus_reg_dataout_1465_port, 
      DataPath_RF_bus_reg_dataout_1466_port, 
      DataPath_RF_bus_reg_dataout_1467_port, 
      DataPath_RF_bus_reg_dataout_1468_port, 
      DataPath_RF_bus_reg_dataout_1469_port, 
      DataPath_RF_bus_reg_dataout_1470_port, 
      DataPath_RF_bus_reg_dataout_1471_port, 
      DataPath_RF_bus_reg_dataout_1472_port, 
      DataPath_RF_bus_reg_dataout_1473_port, 
      DataPath_RF_bus_reg_dataout_1474_port, 
      DataPath_RF_bus_reg_dataout_1475_port, 
      DataPath_RF_bus_reg_dataout_1476_port, 
      DataPath_RF_bus_reg_dataout_1477_port, 
      DataPath_RF_bus_reg_dataout_1478_port, 
      DataPath_RF_bus_reg_dataout_1479_port, 
      DataPath_RF_bus_reg_dataout_1480_port, 
      DataPath_RF_bus_reg_dataout_1481_port, 
      DataPath_RF_bus_reg_dataout_1482_port, 
      DataPath_RF_bus_reg_dataout_1483_port, 
      DataPath_RF_bus_reg_dataout_1484_port, 
      DataPath_RF_bus_reg_dataout_1485_port, 
      DataPath_RF_bus_reg_dataout_1486_port, 
      DataPath_RF_bus_reg_dataout_1487_port, 
      DataPath_RF_bus_reg_dataout_1488_port, 
      DataPath_RF_bus_reg_dataout_1489_port, 
      DataPath_RF_bus_reg_dataout_1490_port, 
      DataPath_RF_bus_reg_dataout_1491_port, 
      DataPath_RF_bus_reg_dataout_1492_port, 
      DataPath_RF_bus_reg_dataout_1493_port, 
      DataPath_RF_bus_reg_dataout_1494_port, 
      DataPath_RF_bus_reg_dataout_1495_port, 
      DataPath_RF_bus_reg_dataout_1496_port, 
      DataPath_RF_bus_reg_dataout_1497_port, 
      DataPath_RF_bus_reg_dataout_1498_port, 
      DataPath_RF_bus_reg_dataout_1499_port, 
      DataPath_RF_bus_reg_dataout_1500_port, 
      DataPath_RF_bus_reg_dataout_1501_port, 
      DataPath_RF_bus_reg_dataout_1502_port, 
      DataPath_RF_bus_reg_dataout_1503_port, 
      DataPath_RF_bus_reg_dataout_1504_port, 
      DataPath_RF_bus_reg_dataout_1505_port, 
      DataPath_RF_bus_reg_dataout_1506_port, 
      DataPath_RF_bus_reg_dataout_1507_port, 
      DataPath_RF_bus_reg_dataout_1508_port, 
      DataPath_RF_bus_reg_dataout_1509_port, 
      DataPath_RF_bus_reg_dataout_1510_port, 
      DataPath_RF_bus_reg_dataout_1511_port, 
      DataPath_RF_bus_reg_dataout_1512_port, 
      DataPath_RF_bus_reg_dataout_1513_port, 
      DataPath_RF_bus_reg_dataout_1514_port, 
      DataPath_RF_bus_reg_dataout_1515_port, 
      DataPath_RF_bus_reg_dataout_1516_port, 
      DataPath_RF_bus_reg_dataout_1517_port, 
      DataPath_RF_bus_reg_dataout_1518_port, 
      DataPath_RF_bus_reg_dataout_1519_port, 
      DataPath_RF_bus_reg_dataout_1520_port, 
      DataPath_RF_bus_reg_dataout_1521_port, 
      DataPath_RF_bus_reg_dataout_1522_port, 
      DataPath_RF_bus_reg_dataout_1523_port, 
      DataPath_RF_bus_reg_dataout_1524_port, 
      DataPath_RF_bus_reg_dataout_1525_port, 
      DataPath_RF_bus_reg_dataout_1526_port, 
      DataPath_RF_bus_reg_dataout_1527_port, 
      DataPath_RF_bus_reg_dataout_1528_port, 
      DataPath_RF_bus_reg_dataout_1529_port, 
      DataPath_RF_bus_reg_dataout_1530_port, 
      DataPath_RF_bus_reg_dataout_1531_port, 
      DataPath_RF_bus_reg_dataout_1532_port, 
      DataPath_RF_bus_reg_dataout_1533_port, 
      DataPath_RF_bus_reg_dataout_1534_port, 
      DataPath_RF_bus_reg_dataout_1535_port, 
      DataPath_RF_bus_reg_dataout_1536_port, 
      DataPath_RF_bus_reg_dataout_1537_port, 
      DataPath_RF_bus_reg_dataout_1538_port, 
      DataPath_RF_bus_reg_dataout_1539_port, 
      DataPath_RF_bus_reg_dataout_1540_port, 
      DataPath_RF_bus_reg_dataout_1541_port, 
      DataPath_RF_bus_reg_dataout_1542_port, 
      DataPath_RF_bus_reg_dataout_1543_port, 
      DataPath_RF_bus_reg_dataout_1544_port, 
      DataPath_RF_bus_reg_dataout_1545_port, 
      DataPath_RF_bus_reg_dataout_1546_port, 
      DataPath_RF_bus_reg_dataout_1547_port, 
      DataPath_RF_bus_reg_dataout_1548_port, 
      DataPath_RF_bus_reg_dataout_1549_port, 
      DataPath_RF_bus_reg_dataout_1550_port, 
      DataPath_RF_bus_reg_dataout_1551_port, 
      DataPath_RF_bus_reg_dataout_1552_port, 
      DataPath_RF_bus_reg_dataout_1553_port, 
      DataPath_RF_bus_reg_dataout_1554_port, 
      DataPath_RF_bus_reg_dataout_1555_port, 
      DataPath_RF_bus_reg_dataout_1556_port, 
      DataPath_RF_bus_reg_dataout_1557_port, 
      DataPath_RF_bus_reg_dataout_1558_port, 
      DataPath_RF_bus_reg_dataout_1559_port, 
      DataPath_RF_bus_reg_dataout_1560_port, 
      DataPath_RF_bus_reg_dataout_1561_port, 
      DataPath_RF_bus_reg_dataout_1562_port, 
      DataPath_RF_bus_reg_dataout_1563_port, 
      DataPath_RF_bus_reg_dataout_1564_port, 
      DataPath_RF_bus_reg_dataout_1565_port, 
      DataPath_RF_bus_reg_dataout_1566_port, 
      DataPath_RF_bus_reg_dataout_1567_port, 
      DataPath_RF_bus_reg_dataout_1568_port, 
      DataPath_RF_bus_reg_dataout_1569_port, 
      DataPath_RF_bus_reg_dataout_1570_port, 
      DataPath_RF_bus_reg_dataout_1571_port, 
      DataPath_RF_bus_reg_dataout_1572_port, 
      DataPath_RF_bus_reg_dataout_1573_port, 
      DataPath_RF_bus_reg_dataout_1574_port, 
      DataPath_RF_bus_reg_dataout_1575_port, 
      DataPath_RF_bus_reg_dataout_1576_port, 
      DataPath_RF_bus_reg_dataout_1577_port, 
      DataPath_RF_bus_reg_dataout_1578_port, 
      DataPath_RF_bus_reg_dataout_1579_port, 
      DataPath_RF_bus_reg_dataout_1580_port, 
      DataPath_RF_bus_reg_dataout_1581_port, 
      DataPath_RF_bus_reg_dataout_1582_port, 
      DataPath_RF_bus_reg_dataout_1583_port, 
      DataPath_RF_bus_reg_dataout_1584_port, 
      DataPath_RF_bus_reg_dataout_1585_port, 
      DataPath_RF_bus_reg_dataout_1586_port, 
      DataPath_RF_bus_reg_dataout_1587_port, 
      DataPath_RF_bus_reg_dataout_1588_port, 
      DataPath_RF_bus_reg_dataout_1589_port, 
      DataPath_RF_bus_reg_dataout_1590_port, 
      DataPath_RF_bus_reg_dataout_1591_port, 
      DataPath_RF_bus_reg_dataout_1592_port, 
      DataPath_RF_bus_reg_dataout_1593_port, 
      DataPath_RF_bus_reg_dataout_1594_port, 
      DataPath_RF_bus_reg_dataout_1595_port, 
      DataPath_RF_bus_reg_dataout_1596_port, 
      DataPath_RF_bus_reg_dataout_1597_port, 
      DataPath_RF_bus_reg_dataout_1598_port, 
      DataPath_RF_bus_reg_dataout_1599_port, 
      DataPath_RF_bus_reg_dataout_1600_port, 
      DataPath_RF_bus_reg_dataout_1601_port, 
      DataPath_RF_bus_reg_dataout_1602_port, 
      DataPath_RF_bus_reg_dataout_1603_port, 
      DataPath_RF_bus_reg_dataout_1604_port, 
      DataPath_RF_bus_reg_dataout_1605_port, 
      DataPath_RF_bus_reg_dataout_1606_port, 
      DataPath_RF_bus_reg_dataout_1607_port, 
      DataPath_RF_bus_reg_dataout_1608_port, 
      DataPath_RF_bus_reg_dataout_1609_port, 
      DataPath_RF_bus_reg_dataout_1610_port, 
      DataPath_RF_bus_reg_dataout_1611_port, 
      DataPath_RF_bus_reg_dataout_1612_port, 
      DataPath_RF_bus_reg_dataout_1613_port, 
      DataPath_RF_bus_reg_dataout_1614_port, 
      DataPath_RF_bus_reg_dataout_1615_port, 
      DataPath_RF_bus_reg_dataout_1616_port, 
      DataPath_RF_bus_reg_dataout_1617_port, 
      DataPath_RF_bus_reg_dataout_1618_port, 
      DataPath_RF_bus_reg_dataout_1619_port, 
      DataPath_RF_bus_reg_dataout_1620_port, 
      DataPath_RF_bus_reg_dataout_1621_port, 
      DataPath_RF_bus_reg_dataout_1622_port, 
      DataPath_RF_bus_reg_dataout_1623_port, 
      DataPath_RF_bus_reg_dataout_1624_port, 
      DataPath_RF_bus_reg_dataout_1625_port, 
      DataPath_RF_bus_reg_dataout_1626_port, 
      DataPath_RF_bus_reg_dataout_1627_port, 
      DataPath_RF_bus_reg_dataout_1628_port, 
      DataPath_RF_bus_reg_dataout_1629_port, 
      DataPath_RF_bus_reg_dataout_1630_port, 
      DataPath_RF_bus_reg_dataout_1631_port, 
      DataPath_RF_bus_reg_dataout_1632_port, 
      DataPath_RF_bus_reg_dataout_1633_port, 
      DataPath_RF_bus_reg_dataout_1634_port, 
      DataPath_RF_bus_reg_dataout_1635_port, 
      DataPath_RF_bus_reg_dataout_1636_port, 
      DataPath_RF_bus_reg_dataout_1637_port, 
      DataPath_RF_bus_reg_dataout_1638_port, 
      DataPath_RF_bus_reg_dataout_1639_port, 
      DataPath_RF_bus_reg_dataout_1640_port, 
      DataPath_RF_bus_reg_dataout_1641_port, 
      DataPath_RF_bus_reg_dataout_1642_port, 
      DataPath_RF_bus_reg_dataout_1643_port, 
      DataPath_RF_bus_reg_dataout_1644_port, 
      DataPath_RF_bus_reg_dataout_1645_port, 
      DataPath_RF_bus_reg_dataout_1646_port, 
      DataPath_RF_bus_reg_dataout_1647_port, 
      DataPath_RF_bus_reg_dataout_1648_port, 
      DataPath_RF_bus_reg_dataout_1649_port, 
      DataPath_RF_bus_reg_dataout_1650_port, 
      DataPath_RF_bus_reg_dataout_1651_port, 
      DataPath_RF_bus_reg_dataout_1652_port, 
      DataPath_RF_bus_reg_dataout_1653_port, 
      DataPath_RF_bus_reg_dataout_1654_port, 
      DataPath_RF_bus_reg_dataout_1655_port, 
      DataPath_RF_bus_reg_dataout_1656_port, 
      DataPath_RF_bus_reg_dataout_1657_port, 
      DataPath_RF_bus_reg_dataout_1658_port, 
      DataPath_RF_bus_reg_dataout_1659_port, 
      DataPath_RF_bus_reg_dataout_1660_port, 
      DataPath_RF_bus_reg_dataout_1661_port, 
      DataPath_RF_bus_reg_dataout_1662_port, 
      DataPath_RF_bus_reg_dataout_1663_port, 
      DataPath_RF_bus_reg_dataout_1664_port, 
      DataPath_RF_bus_reg_dataout_1665_port, 
      DataPath_RF_bus_reg_dataout_1666_port, 
      DataPath_RF_bus_reg_dataout_1667_port, 
      DataPath_RF_bus_reg_dataout_1668_port, 
      DataPath_RF_bus_reg_dataout_1669_port, 
      DataPath_RF_bus_reg_dataout_1670_port, 
      DataPath_RF_bus_reg_dataout_1671_port, 
      DataPath_RF_bus_reg_dataout_1672_port, 
      DataPath_RF_bus_reg_dataout_1673_port, 
      DataPath_RF_bus_reg_dataout_1674_port, 
      DataPath_RF_bus_reg_dataout_1675_port, 
      DataPath_RF_bus_reg_dataout_1676_port, 
      DataPath_RF_bus_reg_dataout_1677_port, 
      DataPath_RF_bus_reg_dataout_1678_port, 
      DataPath_RF_bus_reg_dataout_1679_port, 
      DataPath_RF_bus_reg_dataout_1680_port, 
      DataPath_RF_bus_reg_dataout_1681_port, 
      DataPath_RF_bus_reg_dataout_1682_port, 
      DataPath_RF_bus_reg_dataout_1683_port, 
      DataPath_RF_bus_reg_dataout_1684_port, 
      DataPath_RF_bus_reg_dataout_1685_port, 
      DataPath_RF_bus_reg_dataout_1686_port, 
      DataPath_RF_bus_reg_dataout_1687_port, 
      DataPath_RF_bus_reg_dataout_1688_port, 
      DataPath_RF_bus_reg_dataout_1689_port, 
      DataPath_RF_bus_reg_dataout_1690_port, 
      DataPath_RF_bus_reg_dataout_1691_port, 
      DataPath_RF_bus_reg_dataout_1692_port, 
      DataPath_RF_bus_reg_dataout_1693_port, 
      DataPath_RF_bus_reg_dataout_1694_port, 
      DataPath_RF_bus_reg_dataout_1695_port, 
      DataPath_RF_bus_reg_dataout_1696_port, 
      DataPath_RF_bus_reg_dataout_1697_port, 
      DataPath_RF_bus_reg_dataout_1698_port, 
      DataPath_RF_bus_reg_dataout_1699_port, 
      DataPath_RF_bus_reg_dataout_1700_port, 
      DataPath_RF_bus_reg_dataout_1701_port, 
      DataPath_RF_bus_reg_dataout_1702_port, 
      DataPath_RF_bus_reg_dataout_1703_port, 
      DataPath_RF_bus_reg_dataout_1704_port, 
      DataPath_RF_bus_reg_dataout_1705_port, 
      DataPath_RF_bus_reg_dataout_1706_port, 
      DataPath_RF_bus_reg_dataout_1707_port, 
      DataPath_RF_bus_reg_dataout_1708_port, 
      DataPath_RF_bus_reg_dataout_1709_port, 
      DataPath_RF_bus_reg_dataout_1710_port, 
      DataPath_RF_bus_reg_dataout_1711_port, 
      DataPath_RF_bus_reg_dataout_1712_port, 
      DataPath_RF_bus_reg_dataout_1713_port, 
      DataPath_RF_bus_reg_dataout_1714_port, 
      DataPath_RF_bus_reg_dataout_1715_port, 
      DataPath_RF_bus_reg_dataout_1716_port, 
      DataPath_RF_bus_reg_dataout_1717_port, 
      DataPath_RF_bus_reg_dataout_1718_port, 
      DataPath_RF_bus_reg_dataout_1719_port, 
      DataPath_RF_bus_reg_dataout_1720_port, 
      DataPath_RF_bus_reg_dataout_1721_port, 
      DataPath_RF_bus_reg_dataout_1722_port, 
      DataPath_RF_bus_reg_dataout_1723_port, 
      DataPath_RF_bus_reg_dataout_1724_port, 
      DataPath_RF_bus_reg_dataout_1725_port, 
      DataPath_RF_bus_reg_dataout_1726_port, 
      DataPath_RF_bus_reg_dataout_1727_port, 
      DataPath_RF_bus_reg_dataout_1728_port, 
      DataPath_RF_bus_reg_dataout_1729_port, 
      DataPath_RF_bus_reg_dataout_1730_port, 
      DataPath_RF_bus_reg_dataout_1731_port, 
      DataPath_RF_bus_reg_dataout_1732_port, 
      DataPath_RF_bus_reg_dataout_1733_port, 
      DataPath_RF_bus_reg_dataout_1734_port, 
      DataPath_RF_bus_reg_dataout_1735_port, 
      DataPath_RF_bus_reg_dataout_1736_port, 
      DataPath_RF_bus_reg_dataout_1737_port, 
      DataPath_RF_bus_reg_dataout_1738_port, 
      DataPath_RF_bus_reg_dataout_1739_port, 
      DataPath_RF_bus_reg_dataout_1740_port, 
      DataPath_RF_bus_reg_dataout_1741_port, 
      DataPath_RF_bus_reg_dataout_1742_port, 
      DataPath_RF_bus_reg_dataout_1743_port, 
      DataPath_RF_bus_reg_dataout_1744_port, 
      DataPath_RF_bus_reg_dataout_1745_port, 
      DataPath_RF_bus_reg_dataout_1746_port, 
      DataPath_RF_bus_reg_dataout_1747_port, 
      DataPath_RF_bus_reg_dataout_1748_port, 
      DataPath_RF_bus_reg_dataout_1749_port, 
      DataPath_RF_bus_reg_dataout_1750_port, 
      DataPath_RF_bus_reg_dataout_1751_port, 
      DataPath_RF_bus_reg_dataout_1752_port, 
      DataPath_RF_bus_reg_dataout_1753_port, 
      DataPath_RF_bus_reg_dataout_1754_port, 
      DataPath_RF_bus_reg_dataout_1755_port, 
      DataPath_RF_bus_reg_dataout_1756_port, 
      DataPath_RF_bus_reg_dataout_1757_port, 
      DataPath_RF_bus_reg_dataout_1758_port, 
      DataPath_RF_bus_reg_dataout_1759_port, 
      DataPath_RF_bus_reg_dataout_1760_port, 
      DataPath_RF_bus_reg_dataout_1761_port, 
      DataPath_RF_bus_reg_dataout_1762_port, 
      DataPath_RF_bus_reg_dataout_1763_port, 
      DataPath_RF_bus_reg_dataout_1764_port, 
      DataPath_RF_bus_reg_dataout_1765_port, 
      DataPath_RF_bus_reg_dataout_1766_port, 
      DataPath_RF_bus_reg_dataout_1767_port, 
      DataPath_RF_bus_reg_dataout_1768_port, 
      DataPath_RF_bus_reg_dataout_1769_port, 
      DataPath_RF_bus_reg_dataout_1770_port, 
      DataPath_RF_bus_reg_dataout_1771_port, 
      DataPath_RF_bus_reg_dataout_1772_port, 
      DataPath_RF_bus_reg_dataout_1773_port, 
      DataPath_RF_bus_reg_dataout_1774_port, 
      DataPath_RF_bus_reg_dataout_1775_port, 
      DataPath_RF_bus_reg_dataout_1776_port, 
      DataPath_RF_bus_reg_dataout_1777_port, 
      DataPath_RF_bus_reg_dataout_1778_port, 
      DataPath_RF_bus_reg_dataout_1779_port, 
      DataPath_RF_bus_reg_dataout_1780_port, 
      DataPath_RF_bus_reg_dataout_1781_port, 
      DataPath_RF_bus_reg_dataout_1782_port, 
      DataPath_RF_bus_reg_dataout_1783_port, 
      DataPath_RF_bus_reg_dataout_1784_port, 
      DataPath_RF_bus_reg_dataout_1785_port, 
      DataPath_RF_bus_reg_dataout_1786_port, 
      DataPath_RF_bus_reg_dataout_1787_port, 
      DataPath_RF_bus_reg_dataout_1788_port, 
      DataPath_RF_bus_reg_dataout_1789_port, 
      DataPath_RF_bus_reg_dataout_1790_port, 
      DataPath_RF_bus_reg_dataout_1791_port, 
      DataPath_RF_bus_reg_dataout_1792_port, 
      DataPath_RF_bus_reg_dataout_1793_port, 
      DataPath_RF_bus_reg_dataout_1794_port, 
      DataPath_RF_bus_reg_dataout_1795_port, 
      DataPath_RF_bus_reg_dataout_1796_port, 
      DataPath_RF_bus_reg_dataout_1797_port, 
      DataPath_RF_bus_reg_dataout_1798_port, 
      DataPath_RF_bus_reg_dataout_1799_port, 
      DataPath_RF_bus_reg_dataout_1800_port, 
      DataPath_RF_bus_reg_dataout_1801_port, 
      DataPath_RF_bus_reg_dataout_1802_port, 
      DataPath_RF_bus_reg_dataout_1803_port, 
      DataPath_RF_bus_reg_dataout_1804_port, 
      DataPath_RF_bus_reg_dataout_1805_port, 
      DataPath_RF_bus_reg_dataout_1806_port, 
      DataPath_RF_bus_reg_dataout_1807_port, 
      DataPath_RF_bus_reg_dataout_1808_port, 
      DataPath_RF_bus_reg_dataout_1809_port, 
      DataPath_RF_bus_reg_dataout_1810_port, 
      DataPath_RF_bus_reg_dataout_1811_port, 
      DataPath_RF_bus_reg_dataout_1812_port, 
      DataPath_RF_bus_reg_dataout_1813_port, 
      DataPath_RF_bus_reg_dataout_1814_port, 
      DataPath_RF_bus_reg_dataout_1815_port, 
      DataPath_RF_bus_reg_dataout_1816_port, 
      DataPath_RF_bus_reg_dataout_1817_port, 
      DataPath_RF_bus_reg_dataout_1818_port, 
      DataPath_RF_bus_reg_dataout_1819_port, 
      DataPath_RF_bus_reg_dataout_1820_port, 
      DataPath_RF_bus_reg_dataout_1821_port, 
      DataPath_RF_bus_reg_dataout_1822_port, 
      DataPath_RF_bus_reg_dataout_1823_port, 
      DataPath_RF_bus_reg_dataout_1824_port, 
      DataPath_RF_bus_reg_dataout_1825_port, 
      DataPath_RF_bus_reg_dataout_1826_port, 
      DataPath_RF_bus_reg_dataout_1827_port, 
      DataPath_RF_bus_reg_dataout_1828_port, 
      DataPath_RF_bus_reg_dataout_1829_port, 
      DataPath_RF_bus_reg_dataout_1830_port, 
      DataPath_RF_bus_reg_dataout_1831_port, 
      DataPath_RF_bus_reg_dataout_1832_port, 
      DataPath_RF_bus_reg_dataout_1833_port, 
      DataPath_RF_bus_reg_dataout_1834_port, 
      DataPath_RF_bus_reg_dataout_1835_port, 
      DataPath_RF_bus_reg_dataout_1836_port, 
      DataPath_RF_bus_reg_dataout_1837_port, 
      DataPath_RF_bus_reg_dataout_1838_port, 
      DataPath_RF_bus_reg_dataout_1839_port, 
      DataPath_RF_bus_reg_dataout_1840_port, 
      DataPath_RF_bus_reg_dataout_1841_port, 
      DataPath_RF_bus_reg_dataout_1842_port, 
      DataPath_RF_bus_reg_dataout_1843_port, 
      DataPath_RF_bus_reg_dataout_1844_port, 
      DataPath_RF_bus_reg_dataout_1845_port, 
      DataPath_RF_bus_reg_dataout_1846_port, 
      DataPath_RF_bus_reg_dataout_1847_port, 
      DataPath_RF_bus_reg_dataout_1848_port, 
      DataPath_RF_bus_reg_dataout_1849_port, 
      DataPath_RF_bus_reg_dataout_1850_port, 
      DataPath_RF_bus_reg_dataout_1851_port, 
      DataPath_RF_bus_reg_dataout_1852_port, 
      DataPath_RF_bus_reg_dataout_1853_port, 
      DataPath_RF_bus_reg_dataout_1854_port, 
      DataPath_RF_bus_reg_dataout_1855_port, 
      DataPath_RF_bus_reg_dataout_1856_port, 
      DataPath_RF_bus_reg_dataout_1857_port, 
      DataPath_RF_bus_reg_dataout_1858_port, 
      DataPath_RF_bus_reg_dataout_1859_port, 
      DataPath_RF_bus_reg_dataout_1860_port, 
      DataPath_RF_bus_reg_dataout_1861_port, 
      DataPath_RF_bus_reg_dataout_1862_port, 
      DataPath_RF_bus_reg_dataout_1863_port, 
      DataPath_RF_bus_reg_dataout_1864_port, 
      DataPath_RF_bus_reg_dataout_1865_port, 
      DataPath_RF_bus_reg_dataout_1866_port, 
      DataPath_RF_bus_reg_dataout_1867_port, 
      DataPath_RF_bus_reg_dataout_1868_port, 
      DataPath_RF_bus_reg_dataout_1869_port, 
      DataPath_RF_bus_reg_dataout_1870_port, 
      DataPath_RF_bus_reg_dataout_1871_port, 
      DataPath_RF_bus_reg_dataout_1872_port, 
      DataPath_RF_bus_reg_dataout_1873_port, 
      DataPath_RF_bus_reg_dataout_1874_port, 
      DataPath_RF_bus_reg_dataout_1875_port, 
      DataPath_RF_bus_reg_dataout_1876_port, 
      DataPath_RF_bus_reg_dataout_1877_port, 
      DataPath_RF_bus_reg_dataout_1878_port, 
      DataPath_RF_bus_reg_dataout_1879_port, 
      DataPath_RF_bus_reg_dataout_1880_port, 
      DataPath_RF_bus_reg_dataout_1881_port, 
      DataPath_RF_bus_reg_dataout_1882_port, 
      DataPath_RF_bus_reg_dataout_1883_port, 
      DataPath_RF_bus_reg_dataout_1884_port, 
      DataPath_RF_bus_reg_dataout_1885_port, 
      DataPath_RF_bus_reg_dataout_1886_port, 
      DataPath_RF_bus_reg_dataout_1887_port, 
      DataPath_RF_bus_reg_dataout_1888_port, 
      DataPath_RF_bus_reg_dataout_1889_port, 
      DataPath_RF_bus_reg_dataout_1890_port, 
      DataPath_RF_bus_reg_dataout_1891_port, 
      DataPath_RF_bus_reg_dataout_1892_port, 
      DataPath_RF_bus_reg_dataout_1893_port, 
      DataPath_RF_bus_reg_dataout_1894_port, 
      DataPath_RF_bus_reg_dataout_1895_port, 
      DataPath_RF_bus_reg_dataout_1896_port, 
      DataPath_RF_bus_reg_dataout_1897_port, 
      DataPath_RF_bus_reg_dataout_1898_port, 
      DataPath_RF_bus_reg_dataout_1899_port, 
      DataPath_RF_bus_reg_dataout_1900_port, 
      DataPath_RF_bus_reg_dataout_1901_port, 
      DataPath_RF_bus_reg_dataout_1902_port, 
      DataPath_RF_bus_reg_dataout_1903_port, 
      DataPath_RF_bus_reg_dataout_1904_port, 
      DataPath_RF_bus_reg_dataout_1905_port, 
      DataPath_RF_bus_reg_dataout_1906_port, 
      DataPath_RF_bus_reg_dataout_1907_port, 
      DataPath_RF_bus_reg_dataout_1908_port, 
      DataPath_RF_bus_reg_dataout_1909_port, 
      DataPath_RF_bus_reg_dataout_1910_port, 
      DataPath_RF_bus_reg_dataout_1911_port, 
      DataPath_RF_bus_reg_dataout_1912_port, 
      DataPath_RF_bus_reg_dataout_1913_port, 
      DataPath_RF_bus_reg_dataout_1914_port, 
      DataPath_RF_bus_reg_dataout_1915_port, 
      DataPath_RF_bus_reg_dataout_1916_port, 
      DataPath_RF_bus_reg_dataout_1917_port, 
      DataPath_RF_bus_reg_dataout_1918_port, 
      DataPath_RF_bus_reg_dataout_1919_port, 
      DataPath_RF_bus_reg_dataout_1920_port, 
      DataPath_RF_bus_reg_dataout_1921_port, 
      DataPath_RF_bus_reg_dataout_1922_port, 
      DataPath_RF_bus_reg_dataout_1923_port, 
      DataPath_RF_bus_reg_dataout_1924_port, 
      DataPath_RF_bus_reg_dataout_1925_port, 
      DataPath_RF_bus_reg_dataout_1926_port, 
      DataPath_RF_bus_reg_dataout_1927_port, 
      DataPath_RF_bus_reg_dataout_1928_port, 
      DataPath_RF_bus_reg_dataout_1929_port, 
      DataPath_RF_bus_reg_dataout_1930_port, 
      DataPath_RF_bus_reg_dataout_1931_port, 
      DataPath_RF_bus_reg_dataout_1932_port, 
      DataPath_RF_bus_reg_dataout_1933_port, 
      DataPath_RF_bus_reg_dataout_1934_port, 
      DataPath_RF_bus_reg_dataout_1935_port, 
      DataPath_RF_bus_reg_dataout_1936_port, 
      DataPath_RF_bus_reg_dataout_1937_port, 
      DataPath_RF_bus_reg_dataout_1938_port, 
      DataPath_RF_bus_reg_dataout_1939_port, 
      DataPath_RF_bus_reg_dataout_1940_port, 
      DataPath_RF_bus_reg_dataout_1941_port, 
      DataPath_RF_bus_reg_dataout_1942_port, 
      DataPath_RF_bus_reg_dataout_1943_port, 
      DataPath_RF_bus_reg_dataout_1944_port, 
      DataPath_RF_bus_reg_dataout_1945_port, 
      DataPath_RF_bus_reg_dataout_1946_port, 
      DataPath_RF_bus_reg_dataout_1947_port, 
      DataPath_RF_bus_reg_dataout_1948_port, 
      DataPath_RF_bus_reg_dataout_1949_port, 
      DataPath_RF_bus_reg_dataout_1950_port, 
      DataPath_RF_bus_reg_dataout_1951_port, 
      DataPath_RF_bus_reg_dataout_1952_port, 
      DataPath_RF_bus_reg_dataout_1953_port, 
      DataPath_RF_bus_reg_dataout_1954_port, 
      DataPath_RF_bus_reg_dataout_1955_port, 
      DataPath_RF_bus_reg_dataout_1956_port, 
      DataPath_RF_bus_reg_dataout_1957_port, 
      DataPath_RF_bus_reg_dataout_1958_port, 
      DataPath_RF_bus_reg_dataout_1959_port, 
      DataPath_RF_bus_reg_dataout_1960_port, 
      DataPath_RF_bus_reg_dataout_1961_port, 
      DataPath_RF_bus_reg_dataout_1962_port, 
      DataPath_RF_bus_reg_dataout_1963_port, 
      DataPath_RF_bus_reg_dataout_1964_port, 
      DataPath_RF_bus_reg_dataout_1965_port, 
      DataPath_RF_bus_reg_dataout_1966_port, 
      DataPath_RF_bus_reg_dataout_1967_port, 
      DataPath_RF_bus_reg_dataout_1968_port, 
      DataPath_RF_bus_reg_dataout_1969_port, 
      DataPath_RF_bus_reg_dataout_1970_port, 
      DataPath_RF_bus_reg_dataout_1971_port, 
      DataPath_RF_bus_reg_dataout_1972_port, 
      DataPath_RF_bus_reg_dataout_1973_port, 
      DataPath_RF_bus_reg_dataout_1974_port, 
      DataPath_RF_bus_reg_dataout_1975_port, 
      DataPath_RF_bus_reg_dataout_1976_port, 
      DataPath_RF_bus_reg_dataout_1977_port, 
      DataPath_RF_bus_reg_dataout_1978_port, 
      DataPath_RF_bus_reg_dataout_1979_port, 
      DataPath_RF_bus_reg_dataout_1980_port, 
      DataPath_RF_bus_reg_dataout_1981_port, 
      DataPath_RF_bus_reg_dataout_1982_port, 
      DataPath_RF_bus_reg_dataout_1983_port, 
      DataPath_RF_bus_reg_dataout_1984_port, 
      DataPath_RF_bus_reg_dataout_1985_port, 
      DataPath_RF_bus_reg_dataout_1986_port, 
      DataPath_RF_bus_reg_dataout_1987_port, 
      DataPath_RF_bus_reg_dataout_1988_port, 
      DataPath_RF_bus_reg_dataout_1989_port, 
      DataPath_RF_bus_reg_dataout_1990_port, 
      DataPath_RF_bus_reg_dataout_1991_port, 
      DataPath_RF_bus_reg_dataout_1992_port, 
      DataPath_RF_bus_reg_dataout_1993_port, 
      DataPath_RF_bus_reg_dataout_1994_port, 
      DataPath_RF_bus_reg_dataout_1995_port, 
      DataPath_RF_bus_reg_dataout_1996_port, 
      DataPath_RF_bus_reg_dataout_1997_port, 
      DataPath_RF_bus_reg_dataout_1998_port, 
      DataPath_RF_bus_reg_dataout_1999_port, 
      DataPath_RF_bus_reg_dataout_2000_port, 
      DataPath_RF_bus_reg_dataout_2001_port, 
      DataPath_RF_bus_reg_dataout_2002_port, 
      DataPath_RF_bus_reg_dataout_2003_port, 
      DataPath_RF_bus_reg_dataout_2004_port, 
      DataPath_RF_bus_reg_dataout_2005_port, 
      DataPath_RF_bus_reg_dataout_2006_port, 
      DataPath_RF_bus_reg_dataout_2007_port, 
      DataPath_RF_bus_reg_dataout_2008_port, 
      DataPath_RF_bus_reg_dataout_2009_port, 
      DataPath_RF_bus_reg_dataout_2010_port, 
      DataPath_RF_bus_reg_dataout_2011_port, 
      DataPath_RF_bus_reg_dataout_2012_port, 
      DataPath_RF_bus_reg_dataout_2013_port, 
      DataPath_RF_bus_reg_dataout_2014_port, 
      DataPath_RF_bus_reg_dataout_2015_port, 
      DataPath_RF_bus_reg_dataout_2016_port, 
      DataPath_RF_bus_reg_dataout_2017_port, 
      DataPath_RF_bus_reg_dataout_2018_port, 
      DataPath_RF_bus_reg_dataout_2019_port, 
      DataPath_RF_bus_reg_dataout_2020_port, 
      DataPath_RF_bus_reg_dataout_2021_port, 
      DataPath_RF_bus_reg_dataout_2022_port, 
      DataPath_RF_bus_reg_dataout_2023_port, 
      DataPath_RF_bus_reg_dataout_2024_port, 
      DataPath_RF_bus_reg_dataout_2025_port, 
      DataPath_RF_bus_reg_dataout_2026_port, 
      DataPath_RF_bus_reg_dataout_2027_port, 
      DataPath_RF_bus_reg_dataout_2028_port, 
      DataPath_RF_bus_reg_dataout_2029_port, 
      DataPath_RF_bus_reg_dataout_2030_port, 
      DataPath_RF_bus_reg_dataout_2031_port, 
      DataPath_RF_bus_reg_dataout_2032_port, 
      DataPath_RF_bus_reg_dataout_2033_port, 
      DataPath_RF_bus_reg_dataout_2034_port, 
      DataPath_RF_bus_reg_dataout_2035_port, 
      DataPath_RF_bus_reg_dataout_2036_port, 
      DataPath_RF_bus_reg_dataout_2037_port, 
      DataPath_RF_bus_reg_dataout_2038_port, 
      DataPath_RF_bus_reg_dataout_2039_port, 
      DataPath_RF_bus_reg_dataout_2040_port, 
      DataPath_RF_bus_reg_dataout_2041_port, 
      DataPath_RF_bus_reg_dataout_2042_port, 
      DataPath_RF_bus_reg_dataout_2043_port, 
      DataPath_RF_bus_reg_dataout_2044_port, 
      DataPath_RF_bus_reg_dataout_2045_port, 
      DataPath_RF_bus_reg_dataout_2046_port, 
      DataPath_RF_bus_reg_dataout_2047_port, 
      DataPath_RF_bus_reg_dataout_2048_port, 
      DataPath_RF_bus_reg_dataout_2049_port, 
      DataPath_RF_bus_reg_dataout_2050_port, 
      DataPath_RF_bus_reg_dataout_2051_port, 
      DataPath_RF_bus_reg_dataout_2052_port, 
      DataPath_RF_bus_reg_dataout_2053_port, 
      DataPath_RF_bus_reg_dataout_2054_port, 
      DataPath_RF_bus_reg_dataout_2055_port, 
      DataPath_RF_bus_reg_dataout_2056_port, 
      DataPath_RF_bus_reg_dataout_2057_port, 
      DataPath_RF_bus_reg_dataout_2058_port, 
      DataPath_RF_bus_reg_dataout_2059_port, 
      DataPath_RF_bus_reg_dataout_2060_port, 
      DataPath_RF_bus_reg_dataout_2061_port, 
      DataPath_RF_bus_reg_dataout_2062_port, 
      DataPath_RF_bus_reg_dataout_2063_port, 
      DataPath_RF_bus_reg_dataout_2064_port, 
      DataPath_RF_bus_reg_dataout_2065_port, 
      DataPath_RF_bus_reg_dataout_2066_port, 
      DataPath_RF_bus_reg_dataout_2067_port, 
      DataPath_RF_bus_reg_dataout_2068_port, 
      DataPath_RF_bus_reg_dataout_2069_port, 
      DataPath_RF_bus_reg_dataout_2070_port, 
      DataPath_RF_bus_reg_dataout_2071_port, 
      DataPath_RF_bus_reg_dataout_2072_port, 
      DataPath_RF_bus_reg_dataout_2073_port, 
      DataPath_RF_bus_reg_dataout_2074_port, 
      DataPath_RF_bus_reg_dataout_2075_port, 
      DataPath_RF_bus_reg_dataout_2076_port, 
      DataPath_RF_bus_reg_dataout_2077_port, 
      DataPath_RF_bus_reg_dataout_2078_port, 
      DataPath_RF_bus_reg_dataout_2079_port, 
      DataPath_RF_bus_reg_dataout_2080_port, 
      DataPath_RF_bus_reg_dataout_2081_port, 
      DataPath_RF_bus_reg_dataout_2082_port, 
      DataPath_RF_bus_reg_dataout_2083_port, 
      DataPath_RF_bus_reg_dataout_2084_port, 
      DataPath_RF_bus_reg_dataout_2085_port, 
      DataPath_RF_bus_reg_dataout_2086_port, 
      DataPath_RF_bus_reg_dataout_2087_port, 
      DataPath_RF_bus_reg_dataout_2088_port, 
      DataPath_RF_bus_reg_dataout_2089_port, 
      DataPath_RF_bus_reg_dataout_2090_port, 
      DataPath_RF_bus_reg_dataout_2091_port, 
      DataPath_RF_bus_reg_dataout_2092_port, 
      DataPath_RF_bus_reg_dataout_2093_port, 
      DataPath_RF_bus_reg_dataout_2094_port, 
      DataPath_RF_bus_reg_dataout_2095_port, 
      DataPath_RF_bus_reg_dataout_2096_port, 
      DataPath_RF_bus_reg_dataout_2097_port, 
      DataPath_RF_bus_reg_dataout_2098_port, 
      DataPath_RF_bus_reg_dataout_2099_port, 
      DataPath_RF_bus_reg_dataout_2100_port, 
      DataPath_RF_bus_reg_dataout_2101_port, 
      DataPath_RF_bus_reg_dataout_2102_port, 
      DataPath_RF_bus_reg_dataout_2103_port, 
      DataPath_RF_bus_reg_dataout_2104_port, 
      DataPath_RF_bus_reg_dataout_2105_port, 
      DataPath_RF_bus_reg_dataout_2106_port, 
      DataPath_RF_bus_reg_dataout_2107_port, 
      DataPath_RF_bus_reg_dataout_2108_port, 
      DataPath_RF_bus_reg_dataout_2109_port, 
      DataPath_RF_bus_reg_dataout_2110_port, 
      DataPath_RF_bus_reg_dataout_2111_port, 
      DataPath_RF_bus_reg_dataout_2112_port, 
      DataPath_RF_bus_reg_dataout_2113_port, 
      DataPath_RF_bus_reg_dataout_2114_port, 
      DataPath_RF_bus_reg_dataout_2115_port, 
      DataPath_RF_bus_reg_dataout_2116_port, 
      DataPath_RF_bus_reg_dataout_2117_port, 
      DataPath_RF_bus_reg_dataout_2118_port, 
      DataPath_RF_bus_reg_dataout_2119_port, 
      DataPath_RF_bus_reg_dataout_2120_port, 
      DataPath_RF_bus_reg_dataout_2121_port, 
      DataPath_RF_bus_reg_dataout_2122_port, 
      DataPath_RF_bus_reg_dataout_2123_port, 
      DataPath_RF_bus_reg_dataout_2124_port, 
      DataPath_RF_bus_reg_dataout_2125_port, 
      DataPath_RF_bus_reg_dataout_2126_port, 
      DataPath_RF_bus_reg_dataout_2127_port, 
      DataPath_RF_bus_reg_dataout_2128_port, 
      DataPath_RF_bus_reg_dataout_2129_port, 
      DataPath_RF_bus_reg_dataout_2130_port, 
      DataPath_RF_bus_reg_dataout_2131_port, 
      DataPath_RF_bus_reg_dataout_2132_port, 
      DataPath_RF_bus_reg_dataout_2133_port, 
      DataPath_RF_bus_reg_dataout_2134_port, 
      DataPath_RF_bus_reg_dataout_2135_port, 
      DataPath_RF_bus_reg_dataout_2136_port, 
      DataPath_RF_bus_reg_dataout_2137_port, 
      DataPath_RF_bus_reg_dataout_2138_port, 
      DataPath_RF_bus_reg_dataout_2139_port, 
      DataPath_RF_bus_reg_dataout_2140_port, 
      DataPath_RF_bus_reg_dataout_2141_port, 
      DataPath_RF_bus_reg_dataout_2142_port, 
      DataPath_RF_bus_reg_dataout_2143_port, 
      DataPath_RF_bus_reg_dataout_2144_port, 
      DataPath_RF_bus_reg_dataout_2145_port, 
      DataPath_RF_bus_reg_dataout_2146_port, 
      DataPath_RF_bus_reg_dataout_2147_port, 
      DataPath_RF_bus_reg_dataout_2148_port, 
      DataPath_RF_bus_reg_dataout_2149_port, 
      DataPath_RF_bus_reg_dataout_2150_port, 
      DataPath_RF_bus_reg_dataout_2151_port, 
      DataPath_RF_bus_reg_dataout_2152_port, 
      DataPath_RF_bus_reg_dataout_2153_port, 
      DataPath_RF_bus_reg_dataout_2154_port, 
      DataPath_RF_bus_reg_dataout_2155_port, 
      DataPath_RF_bus_reg_dataout_2156_port, 
      DataPath_RF_bus_reg_dataout_2157_port, 
      DataPath_RF_bus_reg_dataout_2158_port, 
      DataPath_RF_bus_reg_dataout_2159_port, 
      DataPath_RF_bus_reg_dataout_2160_port, 
      DataPath_RF_bus_reg_dataout_2161_port, 
      DataPath_RF_bus_reg_dataout_2162_port, 
      DataPath_RF_bus_reg_dataout_2163_port, 
      DataPath_RF_bus_reg_dataout_2164_port, 
      DataPath_RF_bus_reg_dataout_2165_port, 
      DataPath_RF_bus_reg_dataout_2166_port, 
      DataPath_RF_bus_reg_dataout_2167_port, 
      DataPath_RF_bus_reg_dataout_2168_port, 
      DataPath_RF_bus_reg_dataout_2169_port, 
      DataPath_RF_bus_reg_dataout_2170_port, 
      DataPath_RF_bus_reg_dataout_2171_port, 
      DataPath_RF_bus_reg_dataout_2172_port, 
      DataPath_RF_bus_reg_dataout_2173_port, 
      DataPath_RF_bus_reg_dataout_2174_port, 
      DataPath_RF_bus_reg_dataout_2175_port, 
      DataPath_RF_bus_reg_dataout_2176_port, 
      DataPath_RF_bus_reg_dataout_2177_port, 
      DataPath_RF_bus_reg_dataout_2178_port, 
      DataPath_RF_bus_reg_dataout_2179_port, 
      DataPath_RF_bus_reg_dataout_2180_port, 
      DataPath_RF_bus_reg_dataout_2181_port, 
      DataPath_RF_bus_reg_dataout_2182_port, 
      DataPath_RF_bus_reg_dataout_2183_port, 
      DataPath_RF_bus_reg_dataout_2184_port, 
      DataPath_RF_bus_reg_dataout_2185_port, 
      DataPath_RF_bus_reg_dataout_2186_port, 
      DataPath_RF_bus_reg_dataout_2187_port, 
      DataPath_RF_bus_reg_dataout_2188_port, 
      DataPath_RF_bus_reg_dataout_2189_port, 
      DataPath_RF_bus_reg_dataout_2190_port, 
      DataPath_RF_bus_reg_dataout_2191_port, 
      DataPath_RF_bus_reg_dataout_2192_port, 
      DataPath_RF_bus_reg_dataout_2193_port, 
      DataPath_RF_bus_reg_dataout_2194_port, 
      DataPath_RF_bus_reg_dataout_2195_port, 
      DataPath_RF_bus_reg_dataout_2196_port, 
      DataPath_RF_bus_reg_dataout_2197_port, 
      DataPath_RF_bus_reg_dataout_2198_port, 
      DataPath_RF_bus_reg_dataout_2199_port, 
      DataPath_RF_bus_reg_dataout_2200_port, 
      DataPath_RF_bus_reg_dataout_2201_port, 
      DataPath_RF_bus_reg_dataout_2202_port, 
      DataPath_RF_bus_reg_dataout_2203_port, 
      DataPath_RF_bus_reg_dataout_2204_port, 
      DataPath_RF_bus_reg_dataout_2205_port, 
      DataPath_RF_bus_reg_dataout_2206_port, 
      DataPath_RF_bus_reg_dataout_2207_port, 
      DataPath_RF_bus_reg_dataout_2208_port, 
      DataPath_RF_bus_reg_dataout_2209_port, 
      DataPath_RF_bus_reg_dataout_2210_port, 
      DataPath_RF_bus_reg_dataout_2211_port, 
      DataPath_RF_bus_reg_dataout_2212_port, 
      DataPath_RF_bus_reg_dataout_2213_port, 
      DataPath_RF_bus_reg_dataout_2214_port, 
      DataPath_RF_bus_reg_dataout_2215_port, 
      DataPath_RF_bus_reg_dataout_2216_port, 
      DataPath_RF_bus_reg_dataout_2217_port, 
      DataPath_RF_bus_reg_dataout_2218_port, 
      DataPath_RF_bus_reg_dataout_2219_port, 
      DataPath_RF_bus_reg_dataout_2220_port, 
      DataPath_RF_bus_reg_dataout_2221_port, 
      DataPath_RF_bus_reg_dataout_2222_port, 
      DataPath_RF_bus_reg_dataout_2223_port, 
      DataPath_RF_bus_reg_dataout_2224_port, 
      DataPath_RF_bus_reg_dataout_2225_port, 
      DataPath_RF_bus_reg_dataout_2226_port, 
      DataPath_RF_bus_reg_dataout_2227_port, 
      DataPath_RF_bus_reg_dataout_2228_port, 
      DataPath_RF_bus_reg_dataout_2229_port, 
      DataPath_RF_bus_reg_dataout_2230_port, 
      DataPath_RF_bus_reg_dataout_2231_port, 
      DataPath_RF_bus_reg_dataout_2232_port, 
      DataPath_RF_bus_reg_dataout_2233_port, 
      DataPath_RF_bus_reg_dataout_2234_port, 
      DataPath_RF_bus_reg_dataout_2235_port, 
      DataPath_RF_bus_reg_dataout_2236_port, 
      DataPath_RF_bus_reg_dataout_2237_port, 
      DataPath_RF_bus_reg_dataout_2238_port, 
      DataPath_RF_bus_reg_dataout_2239_port, 
      DataPath_RF_bus_reg_dataout_2240_port, 
      DataPath_RF_bus_reg_dataout_2241_port, 
      DataPath_RF_bus_reg_dataout_2242_port, 
      DataPath_RF_bus_reg_dataout_2243_port, 
      DataPath_RF_bus_reg_dataout_2244_port, 
      DataPath_RF_bus_reg_dataout_2245_port, 
      DataPath_RF_bus_reg_dataout_2246_port, 
      DataPath_RF_bus_reg_dataout_2247_port, 
      DataPath_RF_bus_reg_dataout_2248_port, 
      DataPath_RF_bus_reg_dataout_2249_port, 
      DataPath_RF_bus_reg_dataout_2250_port, 
      DataPath_RF_bus_reg_dataout_2251_port, 
      DataPath_RF_bus_reg_dataout_2252_port, 
      DataPath_RF_bus_reg_dataout_2253_port, 
      DataPath_RF_bus_reg_dataout_2254_port, 
      DataPath_RF_bus_reg_dataout_2255_port, 
      DataPath_RF_bus_reg_dataout_2256_port, 
      DataPath_RF_bus_reg_dataout_2257_port, 
      DataPath_RF_bus_reg_dataout_2258_port, 
      DataPath_RF_bus_reg_dataout_2259_port, 
      DataPath_RF_bus_reg_dataout_2260_port, 
      DataPath_RF_bus_reg_dataout_2261_port, 
      DataPath_RF_bus_reg_dataout_2262_port, 
      DataPath_RF_bus_reg_dataout_2263_port, 
      DataPath_RF_bus_reg_dataout_2264_port, 
      DataPath_RF_bus_reg_dataout_2265_port, 
      DataPath_RF_bus_reg_dataout_2266_port, 
      DataPath_RF_bus_reg_dataout_2267_port, 
      DataPath_RF_bus_reg_dataout_2268_port, 
      DataPath_RF_bus_reg_dataout_2269_port, 
      DataPath_RF_bus_reg_dataout_2270_port, 
      DataPath_RF_bus_reg_dataout_2271_port, 
      DataPath_RF_bus_reg_dataout_2272_port, 
      DataPath_RF_bus_reg_dataout_2273_port, 
      DataPath_RF_bus_reg_dataout_2274_port, 
      DataPath_RF_bus_reg_dataout_2275_port, 
      DataPath_RF_bus_reg_dataout_2276_port, 
      DataPath_RF_bus_reg_dataout_2277_port, 
      DataPath_RF_bus_reg_dataout_2278_port, 
      DataPath_RF_bus_reg_dataout_2279_port, 
      DataPath_RF_bus_reg_dataout_2280_port, 
      DataPath_RF_bus_reg_dataout_2281_port, 
      DataPath_RF_bus_reg_dataout_2282_port, 
      DataPath_RF_bus_reg_dataout_2283_port, 
      DataPath_RF_bus_reg_dataout_2284_port, 
      DataPath_RF_bus_reg_dataout_2285_port, 
      DataPath_RF_bus_reg_dataout_2286_port, 
      DataPath_RF_bus_reg_dataout_2287_port, 
      DataPath_RF_bus_reg_dataout_2288_port, 
      DataPath_RF_bus_reg_dataout_2289_port, 
      DataPath_RF_bus_reg_dataout_2290_port, 
      DataPath_RF_bus_reg_dataout_2291_port, 
      DataPath_RF_bus_reg_dataout_2292_port, 
      DataPath_RF_bus_reg_dataout_2293_port, 
      DataPath_RF_bus_reg_dataout_2294_port, 
      DataPath_RF_bus_reg_dataout_2295_port, 
      DataPath_RF_bus_reg_dataout_2296_port, 
      DataPath_RF_bus_reg_dataout_2297_port, 
      DataPath_RF_bus_reg_dataout_2298_port, 
      DataPath_RF_bus_reg_dataout_2299_port, 
      DataPath_RF_bus_reg_dataout_2300_port, 
      DataPath_RF_bus_reg_dataout_2301_port, 
      DataPath_RF_bus_reg_dataout_2302_port, 
      DataPath_RF_bus_reg_dataout_2303_port, 
      DataPath_RF_bus_reg_dataout_2304_port, 
      DataPath_RF_bus_reg_dataout_2305_port, 
      DataPath_RF_bus_reg_dataout_2306_port, 
      DataPath_RF_bus_reg_dataout_2307_port, 
      DataPath_RF_bus_reg_dataout_2308_port, 
      DataPath_RF_bus_reg_dataout_2309_port, 
      DataPath_RF_bus_reg_dataout_2310_port, 
      DataPath_RF_bus_reg_dataout_2311_port, 
      DataPath_RF_bus_reg_dataout_2312_port, 
      DataPath_RF_bus_reg_dataout_2313_port, 
      DataPath_RF_bus_reg_dataout_2314_port, 
      DataPath_RF_bus_reg_dataout_2315_port, 
      DataPath_RF_bus_reg_dataout_2316_port, 
      DataPath_RF_bus_reg_dataout_2317_port, 
      DataPath_RF_bus_reg_dataout_2318_port, 
      DataPath_RF_bus_reg_dataout_2319_port, 
      DataPath_RF_bus_reg_dataout_2320_port, 
      DataPath_RF_bus_reg_dataout_2321_port, 
      DataPath_RF_bus_reg_dataout_2322_port, 
      DataPath_RF_bus_reg_dataout_2323_port, 
      DataPath_RF_bus_reg_dataout_2324_port, 
      DataPath_RF_bus_reg_dataout_2325_port, 
      DataPath_RF_bus_reg_dataout_2326_port, 
      DataPath_RF_bus_reg_dataout_2327_port, 
      DataPath_RF_bus_reg_dataout_2328_port, 
      DataPath_RF_bus_reg_dataout_2329_port, 
      DataPath_RF_bus_reg_dataout_2330_port, 
      DataPath_RF_bus_reg_dataout_2331_port, 
      DataPath_RF_bus_reg_dataout_2332_port, 
      DataPath_RF_bus_reg_dataout_2333_port, 
      DataPath_RF_bus_reg_dataout_2334_port, 
      DataPath_RF_bus_reg_dataout_2335_port, 
      DataPath_RF_bus_reg_dataout_2336_port, 
      DataPath_RF_bus_reg_dataout_2337_port, 
      DataPath_RF_bus_reg_dataout_2338_port, 
      DataPath_RF_bus_reg_dataout_2339_port, 
      DataPath_RF_bus_reg_dataout_2340_port, 
      DataPath_RF_bus_reg_dataout_2341_port, 
      DataPath_RF_bus_reg_dataout_2342_port, 
      DataPath_RF_bus_reg_dataout_2343_port, 
      DataPath_RF_bus_reg_dataout_2344_port, 
      DataPath_RF_bus_reg_dataout_2345_port, 
      DataPath_RF_bus_reg_dataout_2346_port, 
      DataPath_RF_bus_reg_dataout_2347_port, 
      DataPath_RF_bus_reg_dataout_2348_port, 
      DataPath_RF_bus_reg_dataout_2349_port, 
      DataPath_RF_bus_reg_dataout_2350_port, 
      DataPath_RF_bus_reg_dataout_2351_port, 
      DataPath_RF_bus_reg_dataout_2352_port, 
      DataPath_RF_bus_reg_dataout_2353_port, 
      DataPath_RF_bus_reg_dataout_2354_port, 
      DataPath_RF_bus_reg_dataout_2355_port, 
      DataPath_RF_bus_reg_dataout_2356_port, 
      DataPath_RF_bus_reg_dataout_2357_port, 
      DataPath_RF_bus_reg_dataout_2358_port, 
      DataPath_RF_bus_reg_dataout_2359_port, 
      DataPath_RF_bus_reg_dataout_2360_port, 
      DataPath_RF_bus_reg_dataout_2361_port, 
      DataPath_RF_bus_reg_dataout_2362_port, 
      DataPath_RF_bus_reg_dataout_2363_port, 
      DataPath_RF_bus_reg_dataout_2364_port, 
      DataPath_RF_bus_reg_dataout_2365_port, 
      DataPath_RF_bus_reg_dataout_2366_port, 
      DataPath_RF_bus_reg_dataout_2367_port, 
      DataPath_RF_bus_reg_dataout_2368_port, 
      DataPath_RF_bus_reg_dataout_2369_port, 
      DataPath_RF_bus_reg_dataout_2370_port, 
      DataPath_RF_bus_reg_dataout_2371_port, 
      DataPath_RF_bus_reg_dataout_2372_port, 
      DataPath_RF_bus_reg_dataout_2373_port, 
      DataPath_RF_bus_reg_dataout_2374_port, 
      DataPath_RF_bus_reg_dataout_2375_port, 
      DataPath_RF_bus_reg_dataout_2376_port, 
      DataPath_RF_bus_reg_dataout_2377_port, 
      DataPath_RF_bus_reg_dataout_2378_port, 
      DataPath_RF_bus_reg_dataout_2379_port, 
      DataPath_RF_bus_reg_dataout_2380_port, 
      DataPath_RF_bus_reg_dataout_2381_port, 
      DataPath_RF_bus_reg_dataout_2382_port, 
      DataPath_RF_bus_reg_dataout_2383_port, 
      DataPath_RF_bus_reg_dataout_2384_port, 
      DataPath_RF_bus_reg_dataout_2385_port, 
      DataPath_RF_bus_reg_dataout_2386_port, 
      DataPath_RF_bus_reg_dataout_2387_port, 
      DataPath_RF_bus_reg_dataout_2388_port, 
      DataPath_RF_bus_reg_dataout_2389_port, 
      DataPath_RF_bus_reg_dataout_2390_port, 
      DataPath_RF_bus_reg_dataout_2391_port, 
      DataPath_RF_bus_reg_dataout_2392_port, 
      DataPath_RF_bus_reg_dataout_2393_port, 
      DataPath_RF_bus_reg_dataout_2394_port, 
      DataPath_RF_bus_reg_dataout_2395_port, 
      DataPath_RF_bus_reg_dataout_2396_port, 
      DataPath_RF_bus_reg_dataout_2397_port, 
      DataPath_RF_bus_reg_dataout_2398_port, 
      DataPath_RF_bus_reg_dataout_2399_port, 
      DataPath_RF_bus_reg_dataout_2400_port, 
      DataPath_RF_bus_reg_dataout_2401_port, 
      DataPath_RF_bus_reg_dataout_2402_port, 
      DataPath_RF_bus_reg_dataout_2403_port, 
      DataPath_RF_bus_reg_dataout_2404_port, 
      DataPath_RF_bus_reg_dataout_2405_port, 
      DataPath_RF_bus_reg_dataout_2406_port, 
      DataPath_RF_bus_reg_dataout_2407_port, 
      DataPath_RF_bus_reg_dataout_2408_port, 
      DataPath_RF_bus_reg_dataout_2409_port, 
      DataPath_RF_bus_reg_dataout_2410_port, 
      DataPath_RF_bus_reg_dataout_2411_port, 
      DataPath_RF_bus_reg_dataout_2412_port, 
      DataPath_RF_bus_reg_dataout_2413_port, 
      DataPath_RF_bus_reg_dataout_2414_port, 
      DataPath_RF_bus_reg_dataout_2415_port, 
      DataPath_RF_bus_reg_dataout_2416_port, 
      DataPath_RF_bus_reg_dataout_2417_port, 
      DataPath_RF_bus_reg_dataout_2418_port, 
      DataPath_RF_bus_reg_dataout_2419_port, 
      DataPath_RF_bus_reg_dataout_2420_port, 
      DataPath_RF_bus_reg_dataout_2421_port, 
      DataPath_RF_bus_reg_dataout_2422_port, 
      DataPath_RF_bus_reg_dataout_2423_port, 
      DataPath_RF_bus_reg_dataout_2424_port, 
      DataPath_RF_bus_reg_dataout_2425_port, 
      DataPath_RF_bus_reg_dataout_2426_port, 
      DataPath_RF_bus_reg_dataout_2427_port, 
      DataPath_RF_bus_reg_dataout_2428_port, 
      DataPath_RF_bus_reg_dataout_2429_port, 
      DataPath_RF_bus_reg_dataout_2430_port, 
      DataPath_RF_bus_reg_dataout_2431_port, 
      DataPath_RF_bus_reg_dataout_2432_port, 
      DataPath_RF_bus_reg_dataout_2433_port, 
      DataPath_RF_bus_reg_dataout_2434_port, 
      DataPath_RF_bus_reg_dataout_2435_port, 
      DataPath_RF_bus_reg_dataout_2436_port, 
      DataPath_RF_bus_reg_dataout_2437_port, 
      DataPath_RF_bus_reg_dataout_2438_port, 
      DataPath_RF_bus_reg_dataout_2439_port, 
      DataPath_RF_bus_reg_dataout_2440_port, 
      DataPath_RF_bus_reg_dataout_2441_port, 
      DataPath_RF_bus_reg_dataout_2442_port, 
      DataPath_RF_bus_reg_dataout_2443_port, 
      DataPath_RF_bus_reg_dataout_2444_port, 
      DataPath_RF_bus_reg_dataout_2445_port, 
      DataPath_RF_bus_reg_dataout_2446_port, 
      DataPath_RF_bus_reg_dataout_2447_port, 
      DataPath_RF_bus_reg_dataout_2448_port, 
      DataPath_RF_bus_reg_dataout_2449_port, 
      DataPath_RF_bus_reg_dataout_2450_port, 
      DataPath_RF_bus_reg_dataout_2451_port, 
      DataPath_RF_bus_reg_dataout_2452_port, 
      DataPath_RF_bus_reg_dataout_2453_port, 
      DataPath_RF_bus_reg_dataout_2454_port, 
      DataPath_RF_bus_reg_dataout_2455_port, 
      DataPath_RF_bus_reg_dataout_2456_port, 
      DataPath_RF_bus_reg_dataout_2457_port, 
      DataPath_RF_bus_reg_dataout_2458_port, 
      DataPath_RF_bus_reg_dataout_2459_port, 
      DataPath_RF_bus_reg_dataout_2460_port, 
      DataPath_RF_bus_reg_dataout_2461_port, 
      DataPath_RF_bus_reg_dataout_2462_port, 
      DataPath_RF_bus_reg_dataout_2463_port, 
      DataPath_RF_bus_reg_dataout_2464_port, 
      DataPath_RF_bus_reg_dataout_2465_port, 
      DataPath_RF_bus_reg_dataout_2466_port, 
      DataPath_RF_bus_reg_dataout_2467_port, 
      DataPath_RF_bus_reg_dataout_2468_port, 
      DataPath_RF_bus_reg_dataout_2469_port, 
      DataPath_RF_bus_reg_dataout_2470_port, 
      DataPath_RF_bus_reg_dataout_2471_port, 
      DataPath_RF_bus_reg_dataout_2472_port, 
      DataPath_RF_bus_reg_dataout_2473_port, 
      DataPath_RF_bus_reg_dataout_2474_port, 
      DataPath_RF_bus_reg_dataout_2475_port, 
      DataPath_RF_bus_reg_dataout_2476_port, 
      DataPath_RF_bus_reg_dataout_2477_port, 
      DataPath_RF_bus_reg_dataout_2478_port, 
      DataPath_RF_bus_reg_dataout_2479_port, 
      DataPath_RF_bus_reg_dataout_2480_port, 
      DataPath_RF_bus_reg_dataout_2481_port, 
      DataPath_RF_bus_reg_dataout_2482_port, 
      DataPath_RF_bus_reg_dataout_2483_port, 
      DataPath_RF_bus_reg_dataout_2484_port, 
      DataPath_RF_bus_reg_dataout_2485_port, 
      DataPath_RF_bus_reg_dataout_2486_port, 
      DataPath_RF_bus_reg_dataout_2487_port, 
      DataPath_RF_bus_reg_dataout_2488_port, 
      DataPath_RF_bus_reg_dataout_2489_port, 
      DataPath_RF_bus_reg_dataout_2490_port, 
      DataPath_RF_bus_reg_dataout_2491_port, 
      DataPath_RF_bus_reg_dataout_2492_port, 
      DataPath_RF_bus_reg_dataout_2493_port, 
      DataPath_RF_bus_reg_dataout_2494_port, 
      DataPath_RF_bus_reg_dataout_2495_port, 
      DataPath_RF_bus_reg_dataout_2496_port, 
      DataPath_RF_bus_reg_dataout_2497_port, 
      DataPath_RF_bus_reg_dataout_2498_port, 
      DataPath_RF_bus_reg_dataout_2499_port, 
      DataPath_RF_bus_reg_dataout_2500_port, 
      DataPath_RF_bus_reg_dataout_2501_port, 
      DataPath_RF_bus_reg_dataout_2502_port, 
      DataPath_RF_bus_reg_dataout_2503_port, 
      DataPath_RF_bus_reg_dataout_2504_port, 
      DataPath_RF_bus_reg_dataout_2505_port, 
      DataPath_RF_bus_reg_dataout_2506_port, 
      DataPath_RF_bus_reg_dataout_2507_port, 
      DataPath_RF_bus_reg_dataout_2508_port, 
      DataPath_RF_bus_reg_dataout_2509_port, 
      DataPath_RF_bus_reg_dataout_2510_port, 
      DataPath_RF_bus_reg_dataout_2511_port, 
      DataPath_RF_bus_reg_dataout_2512_port, 
      DataPath_RF_bus_reg_dataout_2513_port, 
      DataPath_RF_bus_reg_dataout_2514_port, 
      DataPath_RF_bus_reg_dataout_2515_port, 
      DataPath_RF_bus_reg_dataout_2516_port, 
      DataPath_RF_bus_reg_dataout_2517_port, 
      DataPath_RF_bus_reg_dataout_2518_port, 
      DataPath_RF_bus_reg_dataout_2519_port, 
      DataPath_RF_bus_reg_dataout_2520_port, 
      DataPath_RF_bus_reg_dataout_2521_port, 
      DataPath_RF_bus_reg_dataout_2522_port, 
      DataPath_RF_bus_reg_dataout_2523_port, 
      DataPath_RF_bus_reg_dataout_2524_port, 
      DataPath_RF_bus_reg_dataout_2525_port, 
      DataPath_RF_bus_reg_dataout_2526_port, 
      DataPath_RF_bus_reg_dataout_2527_port, 
      DataPath_RF_bus_reg_dataout_2528_port, 
      DataPath_RF_bus_reg_dataout_2529_port, 
      DataPath_RF_bus_reg_dataout_2530_port, 
      DataPath_RF_bus_reg_dataout_2531_port, 
      DataPath_RF_bus_reg_dataout_2532_port, 
      DataPath_RF_bus_reg_dataout_2533_port, 
      DataPath_RF_bus_reg_dataout_2534_port, 
      DataPath_RF_bus_reg_dataout_2535_port, 
      DataPath_RF_bus_reg_dataout_2536_port, 
      DataPath_RF_bus_reg_dataout_2537_port, 
      DataPath_RF_bus_reg_dataout_2538_port, 
      DataPath_RF_bus_reg_dataout_2539_port, 
      DataPath_RF_bus_reg_dataout_2540_port, 
      DataPath_RF_bus_reg_dataout_2541_port, 
      DataPath_RF_bus_reg_dataout_2542_port, 
      DataPath_RF_bus_reg_dataout_2543_port, 
      DataPath_RF_bus_reg_dataout_2544_port, 
      DataPath_RF_bus_reg_dataout_2545_port, 
      DataPath_RF_bus_reg_dataout_2546_port, 
      DataPath_RF_bus_reg_dataout_2547_port, 
      DataPath_RF_bus_reg_dataout_2548_port, 
      DataPath_RF_bus_reg_dataout_2549_port, 
      DataPath_RF_bus_reg_dataout_2550_port, 
      DataPath_RF_bus_reg_dataout_2551_port, 
      DataPath_RF_bus_reg_dataout_2552_port, 
      DataPath_RF_bus_reg_dataout_2553_port, 
      DataPath_RF_bus_reg_dataout_2554_port, 
      DataPath_RF_bus_reg_dataout_2555_port, 
      DataPath_RF_bus_reg_dataout_2556_port, 
      DataPath_RF_bus_reg_dataout_2557_port, 
      DataPath_RF_bus_reg_dataout_2558_port, 
      DataPath_RF_bus_reg_dataout_2559_port, DataPath_RF_c_win_0_port, 
      DataPath_RF_c_win_1_port, DataPath_RF_c_win_2_port, 
      DataPath_RF_c_win_3_port, DataPath_RF_c_win_4_port, 
      DataPath_WRF_CUhw_N145, DataPath_WRF_CUhw_curr_addr_2_port, 
      DataPath_WRF_CUhw_curr_addr_3_port, DataPath_WRF_CUhw_curr_addr_4_port, 
      DataPath_WRF_CUhw_curr_addr_5_port, DataPath_WRF_CUhw_curr_addr_6_port, 
      DataPath_WRF_CUhw_curr_addr_7_port, DataPath_WRF_CUhw_curr_addr_8_port, 
      DataPath_WRF_CUhw_curr_addr_9_port, DataPath_WRF_CUhw_curr_addr_10_port, 
      DataPath_WRF_CUhw_curr_addr_11_port, DataPath_WRF_CUhw_curr_addr_12_port,
      DataPath_WRF_CUhw_curr_addr_13_port, DataPath_WRF_CUhw_curr_addr_14_port,
      DataPath_WRF_CUhw_curr_addr_15_port, DataPath_WRF_CUhw_curr_addr_16_port,
      DataPath_WRF_CUhw_curr_addr_17_port, DataPath_WRF_CUhw_curr_addr_18_port,
      DataPath_WRF_CUhw_curr_addr_19_port, DataPath_WRF_CUhw_curr_addr_20_port,
      DataPath_WRF_CUhw_curr_addr_21_port, DataPath_WRF_CUhw_curr_addr_22_port,
      DataPath_WRF_CUhw_curr_addr_23_port, DataPath_WRF_CUhw_curr_addr_24_port,
      DataPath_WRF_CUhw_curr_addr_25_port, DataPath_WRF_CUhw_curr_addr_26_port,
      DataPath_WRF_CUhw_curr_addr_27_port, DataPath_WRF_CUhw_curr_addr_28_port,
      DataPath_WRF_CUhw_curr_addr_29_port, DataPath_WRF_CUhw_curr_addr_30_port,
      DataPath_WRF_CUhw_curr_addr_31_port, DataPath_WRF_CUhw_curr_data_0_port, 
      DataPath_WRF_CUhw_curr_data_1_port, DataPath_WRF_CUhw_curr_data_2_port, 
      DataPath_WRF_CUhw_curr_data_3_port, DataPath_WRF_CUhw_curr_data_4_port, 
      DataPath_WRF_CUhw_curr_data_5_port, DataPath_WRF_CUhw_curr_data_6_port, 
      DataPath_WRF_CUhw_curr_data_7_port, DataPath_WRF_CUhw_curr_data_8_port, 
      DataPath_WRF_CUhw_curr_data_9_port, DataPath_WRF_CUhw_curr_data_10_port, 
      DataPath_WRF_CUhw_curr_data_11_port, DataPath_WRF_CUhw_curr_data_12_port,
      DataPath_WRF_CUhw_curr_data_13_port, DataPath_WRF_CUhw_curr_data_14_port,
      DataPath_WRF_CUhw_curr_data_15_port, DataPath_WRF_CUhw_curr_data_16_port,
      DataPath_WRF_CUhw_curr_data_17_port, DataPath_WRF_CUhw_curr_data_18_port,
      DataPath_WRF_CUhw_curr_data_19_port, DataPath_WRF_CUhw_curr_data_20_port,
      DataPath_WRF_CUhw_curr_data_21_port, DataPath_WRF_CUhw_curr_data_22_port,
      DataPath_WRF_CUhw_curr_data_23_port, DataPath_WRF_CUhw_curr_data_24_port,
      DataPath_WRF_CUhw_curr_data_25_port, DataPath_WRF_CUhw_curr_data_26_port,
      DataPath_WRF_CUhw_curr_data_27_port, DataPath_WRF_CUhw_curr_data_28_port,
      DataPath_WRF_CUhw_curr_data_29_port, DataPath_WRF_CUhw_curr_data_30_port,
      DataPath_WRF_CUhw_curr_data_31_port, DataPath_ALUhw_i_Q_EXTENDED_34_port,
      DataPath_ALUhw_i_Q_EXTENDED_41_port, DataPath_ALUhw_i_Q_EXTENDED_42_port,
      DataPath_ALUhw_i_Q_EXTENDED_44_port, DataPath_ALUhw_i_Q_EXTENDED_45_port,
      DataPath_ALUhw_i_Q_EXTENDED_47_port, DataPath_ALUhw_i_Q_EXTENDED_48_port,
      DataPath_ALUhw_i_Q_EXTENDED_49_port, DataPath_ALUhw_i_Q_EXTENDED_50_port,
      DataPath_ALUhw_i_Q_EXTENDED_51_port, DataPath_ALUhw_i_Q_EXTENDED_52_port,
      DataPath_ALUhw_i_Q_EXTENDED_53_port, DataPath_ALUhw_i_Q_EXTENDED_54_port,
      DataPath_ALUhw_i_Q_EXTENDED_55_port, DataPath_ALUhw_i_Q_EXTENDED_56_port,
      DataPath_ALUhw_i_Q_EXTENDED_57_port, DataPath_ALUhw_i_Q_EXTENDED_58_port,
      DataPath_ALUhw_i_Q_EXTENDED_59_port, DataPath_ALUhw_i_Q_EXTENDED_60_port,
      DataPath_RF_RDPORT0_OUTLATCH_N35, DataPath_RF_RDPORT0_OUTLATCH_N34, 
      DataPath_RF_RDPORT0_OUTLATCH_N33, DataPath_RF_RDPORT0_OUTLATCH_N32, 
      DataPath_RF_RDPORT0_OUTLATCH_N31, DataPath_RF_RDPORT0_OUTLATCH_N30, 
      DataPath_RF_RDPORT0_OUTLATCH_N29, DataPath_RF_RDPORT0_OUTLATCH_N28, 
      DataPath_RF_RDPORT0_OUTLATCH_N27, DataPath_RF_RDPORT0_OUTLATCH_N26, 
      DataPath_RF_RDPORT0_OUTLATCH_N25, DataPath_RF_RDPORT0_OUTLATCH_N24, 
      DataPath_RF_RDPORT0_OUTLATCH_N23, DataPath_RF_RDPORT0_OUTLATCH_N22, 
      DataPath_RF_RDPORT0_OUTLATCH_N21, DataPath_RF_RDPORT0_OUTLATCH_N20, 
      DataPath_RF_RDPORT0_OUTLATCH_N19, DataPath_RF_RDPORT0_OUTLATCH_N18, 
      DataPath_RF_RDPORT0_OUTLATCH_N17, DataPath_RF_RDPORT0_OUTLATCH_N16, 
      DataPath_RF_RDPORT0_OUTLATCH_N15, DataPath_RF_RDPORT0_OUTLATCH_N14, 
      DataPath_RF_RDPORT0_OUTLATCH_N13, DataPath_RF_RDPORT0_OUTLATCH_N12, 
      DataPath_RF_RDPORT0_OUTLATCH_N11, DataPath_RF_RDPORT0_OUTLATCH_N10, 
      DataPath_RF_RDPORT0_OUTLATCH_N9, DataPath_RF_RDPORT0_OUTLATCH_N8, 
      DataPath_RF_RDPORT0_OUTLATCH_N7, DataPath_RF_RDPORT0_OUTLATCH_N6, 
      DataPath_RF_RDPORT0_OUTLATCH_N5, DataPath_RF_RDPORT0_OUTLATCH_N4, 
      DataPath_RF_RDPORT0_OUTLATCH_N3, DataPath_RF_RDPORT1_OUTLATCH_N35, 
      DataPath_RF_RDPORT1_OUTLATCH_N34, DataPath_RF_RDPORT1_OUTLATCH_N33, 
      DataPath_RF_RDPORT1_OUTLATCH_N32, DataPath_RF_RDPORT1_OUTLATCH_N31, 
      DataPath_RF_RDPORT1_OUTLATCH_N30, DataPath_RF_RDPORT1_OUTLATCH_N29, 
      DataPath_RF_RDPORT1_OUTLATCH_N28, DataPath_RF_RDPORT1_OUTLATCH_N27, 
      DataPath_RF_RDPORT1_OUTLATCH_N26, DataPath_RF_RDPORT1_OUTLATCH_N25, 
      DataPath_RF_RDPORT1_OUTLATCH_N24, DataPath_RF_RDPORT1_OUTLATCH_N23, 
      DataPath_RF_RDPORT1_OUTLATCH_N22, DataPath_RF_RDPORT1_OUTLATCH_N21, 
      DataPath_RF_RDPORT1_OUTLATCH_N20, DataPath_RF_RDPORT1_OUTLATCH_N19, 
      DataPath_RF_RDPORT1_OUTLATCH_N18, DataPath_RF_RDPORT1_OUTLATCH_N17, 
      DataPath_RF_RDPORT1_OUTLATCH_N16, DataPath_RF_RDPORT1_OUTLATCH_N15, 
      DataPath_RF_RDPORT1_OUTLATCH_N14, DataPath_RF_RDPORT1_OUTLATCH_N13, 
      DataPath_RF_RDPORT1_OUTLATCH_N12, DataPath_RF_RDPORT1_OUTLATCH_N11, 
      DataPath_RF_RDPORT1_OUTLATCH_N10, DataPath_RF_RDPORT1_OUTLATCH_N9, 
      DataPath_RF_RDPORT1_OUTLATCH_N8, DataPath_RF_RDPORT1_OUTLATCH_N7, 
      DataPath_RF_RDPORT1_OUTLATCH_N6, DataPath_RF_RDPORT1_OUTLATCH_N5, 
      DataPath_RF_RDPORT1_OUTLATCH_N4, DataPath_RF_RDPORT1_OUTLATCH_N3, 
      DataPath_RF_PUSH_ADDRGEN_N61, DataPath_RF_PUSH_ADDRGEN_N60, 
      DataPath_RF_PUSH_ADDRGEN_N59, DataPath_RF_PUSH_ADDRGEN_N58, 
      DataPath_RF_PUSH_ADDRGEN_N57, DataPath_RF_PUSH_ADDRGEN_N56, 
      DataPath_RF_PUSH_ADDRGEN_N55, DataPath_RF_PUSH_ADDRGEN_N54, 
      DataPath_RF_PUSH_ADDRGEN_N53, DataPath_RF_PUSH_ADDRGEN_N52, 
      DataPath_RF_PUSH_ADDRGEN_N51, DataPath_RF_PUSH_ADDRGEN_N50, 
      DataPath_RF_PUSH_ADDRGEN_N49, DataPath_RF_PUSH_ADDRGEN_N48, 
      DataPath_RF_PUSH_ADDRGEN_N47, DataPath_RF_PUSH_ADDRGEN_N46, 
      DataPath_RF_PUSH_ADDRGEN_curr_state_0_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_14_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_15_port, DataPath_RF_POP_ADDRGEN_N61, 
      DataPath_RF_POP_ADDRGEN_N46, DataPath_RF_POP_ADDRGEN_curr_state_0_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_15_port, 
      DataPath_ALUhw_MULT_mux_out_15_30_port, 
      DataPath_ALUhw_MULT_mux_out_14_28_port, 
      DataPath_ALUhw_MULT_mux_out_14_29_port, 
      DataPath_ALUhw_MULT_mux_out_14_30_port, 
      DataPath_ALUhw_MULT_mux_out_14_31_port, 
      DataPath_ALUhw_MULT_mux_out_13_26_port, 
      DataPath_ALUhw_MULT_mux_out_13_27_port, 
      DataPath_ALUhw_MULT_mux_out_13_28_port, 
      DataPath_ALUhw_MULT_mux_out_13_29_port, 
      DataPath_ALUhw_MULT_mux_out_13_30_port, 
      DataPath_ALUhw_MULT_mux_out_13_31_port, 
      DataPath_ALUhw_MULT_mux_out_12_24_port, 
      DataPath_ALUhw_MULT_mux_out_12_25_port, 
      DataPath_ALUhw_MULT_mux_out_12_26_port, 
      DataPath_ALUhw_MULT_mux_out_12_27_port, 
      DataPath_ALUhw_MULT_mux_out_12_28_port, 
      DataPath_ALUhw_MULT_mux_out_12_29_port, 
      DataPath_ALUhw_MULT_mux_out_12_30_port, 
      DataPath_ALUhw_MULT_mux_out_12_31_port, 
      DataPath_ALUhw_MULT_mux_out_11_22_port, 
      DataPath_ALUhw_MULT_mux_out_11_23_port, 
      DataPath_ALUhw_MULT_mux_out_11_24_port, 
      DataPath_ALUhw_MULT_mux_out_11_25_port, 
      DataPath_ALUhw_MULT_mux_out_11_26_port, 
      DataPath_ALUhw_MULT_mux_out_11_27_port, 
      DataPath_ALUhw_MULT_mux_out_11_28_port, 
      DataPath_ALUhw_MULT_mux_out_11_29_port, 
      DataPath_ALUhw_MULT_mux_out_11_30_port, 
      DataPath_ALUhw_MULT_mux_out_11_31_port, 
      DataPath_ALUhw_MULT_mux_out_10_20_port, 
      DataPath_ALUhw_MULT_mux_out_10_21_port, 
      DataPath_ALUhw_MULT_mux_out_10_22_port, 
      DataPath_ALUhw_MULT_mux_out_10_23_port, 
      DataPath_ALUhw_MULT_mux_out_10_24_port, 
      DataPath_ALUhw_MULT_mux_out_10_25_port, 
      DataPath_ALUhw_MULT_mux_out_10_26_port, 
      DataPath_ALUhw_MULT_mux_out_10_27_port, 
      DataPath_ALUhw_MULT_mux_out_10_28_port, 
      DataPath_ALUhw_MULT_mux_out_10_29_port, 
      DataPath_ALUhw_MULT_mux_out_10_30_port, 
      DataPath_ALUhw_MULT_mux_out_10_31_port, 
      DataPath_ALUhw_MULT_mux_out_9_19_port, 
      DataPath_ALUhw_MULT_mux_out_9_20_port, 
      DataPath_ALUhw_MULT_mux_out_9_21_port, 
      DataPath_ALUhw_MULT_mux_out_9_22_port, 
      DataPath_ALUhw_MULT_mux_out_9_23_port, 
      DataPath_ALUhw_MULT_mux_out_9_24_port, 
      DataPath_ALUhw_MULT_mux_out_9_25_port, 
      DataPath_ALUhw_MULT_mux_out_9_26_port, 
      DataPath_ALUhw_MULT_mux_out_9_27_port, 
      DataPath_ALUhw_MULT_mux_out_9_28_port, 
      DataPath_ALUhw_MULT_mux_out_9_29_port, 
      DataPath_ALUhw_MULT_mux_out_9_30_port, 
      DataPath_ALUhw_MULT_mux_out_9_31_port, 
      DataPath_ALUhw_MULT_mux_out_8_16_port, 
      DataPath_ALUhw_MULT_mux_out_8_17_port, 
      DataPath_ALUhw_MULT_mux_out_8_18_port, 
      DataPath_ALUhw_MULT_mux_out_8_19_port, 
      DataPath_ALUhw_MULT_mux_out_8_20_port, 
      DataPath_ALUhw_MULT_mux_out_8_21_port, 
      DataPath_ALUhw_MULT_mux_out_8_22_port, 
      DataPath_ALUhw_MULT_mux_out_8_23_port, 
      DataPath_ALUhw_MULT_mux_out_8_24_port, 
      DataPath_ALUhw_MULT_mux_out_8_25_port, 
      DataPath_ALUhw_MULT_mux_out_8_26_port, 
      DataPath_ALUhw_MULT_mux_out_8_27_port, 
      DataPath_ALUhw_MULT_mux_out_8_28_port, 
      DataPath_ALUhw_MULT_mux_out_8_29_port, 
      DataPath_ALUhw_MULT_mux_out_8_30_port, 
      DataPath_ALUhw_MULT_mux_out_8_31_port, 
      DataPath_ALUhw_MULT_mux_out_7_15_port, 
      DataPath_ALUhw_MULT_mux_out_7_16_port, 
      DataPath_ALUhw_MULT_mux_out_7_17_port, 
      DataPath_ALUhw_MULT_mux_out_7_18_port, 
      DataPath_ALUhw_MULT_mux_out_7_19_port, 
      DataPath_ALUhw_MULT_mux_out_7_20_port, 
      DataPath_ALUhw_MULT_mux_out_7_21_port, 
      DataPath_ALUhw_MULT_mux_out_7_22_port, 
      DataPath_ALUhw_MULT_mux_out_7_23_port, 
      DataPath_ALUhw_MULT_mux_out_7_24_port, 
      DataPath_ALUhw_MULT_mux_out_7_25_port, 
      DataPath_ALUhw_MULT_mux_out_7_26_port, 
      DataPath_ALUhw_MULT_mux_out_7_27_port, 
      DataPath_ALUhw_MULT_mux_out_7_28_port, 
      DataPath_ALUhw_MULT_mux_out_7_29_port, 
      DataPath_ALUhw_MULT_mux_out_7_30_port, 
      DataPath_ALUhw_MULT_mux_out_7_31_port, 
      DataPath_ALUhw_MULT_mux_out_6_13_port, 
      DataPath_ALUhw_MULT_mux_out_6_14_port, 
      DataPath_ALUhw_MULT_mux_out_6_15_port, 
      DataPath_ALUhw_MULT_mux_out_6_16_port, 
      DataPath_ALUhw_MULT_mux_out_6_17_port, 
      DataPath_ALUhw_MULT_mux_out_6_18_port, 
      DataPath_ALUhw_MULT_mux_out_6_19_port, 
      DataPath_ALUhw_MULT_mux_out_6_20_port, 
      DataPath_ALUhw_MULT_mux_out_6_21_port, 
      DataPath_ALUhw_MULT_mux_out_6_22_port, 
      DataPath_ALUhw_MULT_mux_out_6_23_port, 
      DataPath_ALUhw_MULT_mux_out_6_24_port, 
      DataPath_ALUhw_MULT_mux_out_6_25_port, 
      DataPath_ALUhw_MULT_mux_out_6_26_port, 
      DataPath_ALUhw_MULT_mux_out_6_27_port, 
      DataPath_ALUhw_MULT_mux_out_6_28_port, 
      DataPath_ALUhw_MULT_mux_out_6_29_port, 
      DataPath_ALUhw_MULT_mux_out_6_30_port, 
      DataPath_ALUhw_MULT_mux_out_6_31_port, 
      DataPath_ALUhw_MULT_mux_out_5_10_port, 
      DataPath_ALUhw_MULT_mux_out_5_11_port, 
      DataPath_ALUhw_MULT_mux_out_5_12_port, 
      DataPath_ALUhw_MULT_mux_out_5_13_port, 
      DataPath_ALUhw_MULT_mux_out_5_14_port, 
      DataPath_ALUhw_MULT_mux_out_5_15_port, 
      DataPath_ALUhw_MULT_mux_out_5_16_port, 
      DataPath_ALUhw_MULT_mux_out_5_17_port, 
      DataPath_ALUhw_MULT_mux_out_5_18_port, 
      DataPath_ALUhw_MULT_mux_out_5_19_port, 
      DataPath_ALUhw_MULT_mux_out_5_20_port, 
      DataPath_ALUhw_MULT_mux_out_5_21_port, 
      DataPath_ALUhw_MULT_mux_out_5_22_port, 
      DataPath_ALUhw_MULT_mux_out_5_23_port, 
      DataPath_ALUhw_MULT_mux_out_5_24_port, 
      DataPath_ALUhw_MULT_mux_out_5_25_port, 
      DataPath_ALUhw_MULT_mux_out_5_26_port, 
      DataPath_ALUhw_MULT_mux_out_5_27_port, 
      DataPath_ALUhw_MULT_mux_out_5_28_port, 
      DataPath_ALUhw_MULT_mux_out_5_29_port, 
      DataPath_ALUhw_MULT_mux_out_5_30_port, 
      DataPath_ALUhw_MULT_mux_out_5_31_port, 
      DataPath_ALUhw_MULT_mux_out_4_9_port, 
      DataPath_ALUhw_MULT_mux_out_4_10_port, 
      DataPath_ALUhw_MULT_mux_out_4_11_port, 
      DataPath_ALUhw_MULT_mux_out_4_12_port, 
      DataPath_ALUhw_MULT_mux_out_4_13_port, 
      DataPath_ALUhw_MULT_mux_out_4_14_port, 
      DataPath_ALUhw_MULT_mux_out_4_15_port, 
      DataPath_ALUhw_MULT_mux_out_4_16_port, 
      DataPath_ALUhw_MULT_mux_out_4_17_port, 
      DataPath_ALUhw_MULT_mux_out_4_18_port, 
      DataPath_ALUhw_MULT_mux_out_4_19_port, 
      DataPath_ALUhw_MULT_mux_out_4_20_port, 
      DataPath_ALUhw_MULT_mux_out_4_21_port, 
      DataPath_ALUhw_MULT_mux_out_4_22_port, 
      DataPath_ALUhw_MULT_mux_out_4_23_port, 
      DataPath_ALUhw_MULT_mux_out_4_24_port, 
      DataPath_ALUhw_MULT_mux_out_4_25_port, 
      DataPath_ALUhw_MULT_mux_out_4_26_port, 
      DataPath_ALUhw_MULT_mux_out_4_27_port, 
      DataPath_ALUhw_MULT_mux_out_4_28_port, 
      DataPath_ALUhw_MULT_mux_out_4_29_port, 
      DataPath_ALUhw_MULT_mux_out_4_30_port, 
      DataPath_ALUhw_MULT_mux_out_4_31_port, 
      DataPath_ALUhw_MULT_mux_out_3_7_port, 
      DataPath_ALUhw_MULT_mux_out_3_8_port, 
      DataPath_ALUhw_MULT_mux_out_3_9_port, 
      DataPath_ALUhw_MULT_mux_out_3_10_port, 
      DataPath_ALUhw_MULT_mux_out_3_11_port, 
      DataPath_ALUhw_MULT_mux_out_3_12_port, 
      DataPath_ALUhw_MULT_mux_out_3_13_port, 
      DataPath_ALUhw_MULT_mux_out_3_14_port, 
      DataPath_ALUhw_MULT_mux_out_3_15_port, 
      DataPath_ALUhw_MULT_mux_out_3_16_port, 
      DataPath_ALUhw_MULT_mux_out_3_17_port, 
      DataPath_ALUhw_MULT_mux_out_3_18_port, 
      DataPath_ALUhw_MULT_mux_out_3_19_port, 
      DataPath_ALUhw_MULT_mux_out_3_20_port, 
      DataPath_ALUhw_MULT_mux_out_3_21_port, 
      DataPath_ALUhw_MULT_mux_out_3_22_port, 
      DataPath_ALUhw_MULT_mux_out_3_23_port, 
      DataPath_ALUhw_MULT_mux_out_3_24_port, 
      DataPath_ALUhw_MULT_mux_out_3_26_port, 
      DataPath_ALUhw_MULT_mux_out_3_27_port, 
      DataPath_ALUhw_MULT_mux_out_3_28_port, 
      DataPath_ALUhw_MULT_mux_out_3_29_port, 
      DataPath_ALUhw_MULT_mux_out_3_30_port, 
      DataPath_ALUhw_MULT_mux_out_3_31_port, 
      DataPath_ALUhw_MULT_mux_out_2_5_port, 
      DataPath_ALUhw_MULT_mux_out_2_6_port, 
      DataPath_ALUhw_MULT_mux_out_2_7_port, 
      DataPath_ALUhw_MULT_mux_out_2_8_port, 
      DataPath_ALUhw_MULT_mux_out_2_9_port, 
      DataPath_ALUhw_MULT_mux_out_2_10_port, 
      DataPath_ALUhw_MULT_mux_out_2_11_port, 
      DataPath_ALUhw_MULT_mux_out_2_12_port, 
      DataPath_ALUhw_MULT_mux_out_2_13_port, 
      DataPath_ALUhw_MULT_mux_out_2_14_port, 
      DataPath_ALUhw_MULT_mux_out_2_15_port, 
      DataPath_ALUhw_MULT_mux_out_2_16_port, 
      DataPath_ALUhw_MULT_mux_out_2_17_port, 
      DataPath_ALUhw_MULT_mux_out_2_18_port, 
      DataPath_ALUhw_MULT_mux_out_2_19_port, 
      DataPath_ALUhw_MULT_mux_out_2_20_port, 
      DataPath_ALUhw_MULT_mux_out_2_21_port, 
      DataPath_ALUhw_MULT_mux_out_2_22_port, 
      DataPath_ALUhw_MULT_mux_out_2_23_port, 
      DataPath_ALUhw_MULT_mux_out_2_24_port, 
      DataPath_ALUhw_MULT_mux_out_2_25_port, 
      DataPath_ALUhw_MULT_mux_out_2_26_port, 
      DataPath_ALUhw_MULT_mux_out_2_27_port, 
      DataPath_ALUhw_MULT_mux_out_2_28_port, 
      DataPath_ALUhw_MULT_mux_out_2_29_port, 
      DataPath_ALUhw_MULT_mux_out_2_30_port, 
      DataPath_ALUhw_MULT_mux_out_2_31_port, 
      DataPath_ALUhw_MULT_mux_out_1_2_port, 
      DataPath_ALUhw_MULT_mux_out_1_3_port, 
      DataPath_ALUhw_MULT_mux_out_1_6_port, 
      DataPath_ALUhw_MULT_mux_out_1_7_port, 
      DataPath_ALUhw_MULT_mux_out_1_8_port, 
      DataPath_ALUhw_MULT_mux_out_1_12_port, 
      DataPath_ALUhw_MULT_mux_out_1_13_port, 
      DataPath_ALUhw_MULT_mux_out_1_14_port, 
      DataPath_ALUhw_MULT_mux_out_1_15_port, 
      DataPath_ALUhw_MULT_mux_out_1_16_port, 
      DataPath_ALUhw_MULT_mux_out_1_17_port, 
      DataPath_ALUhw_MULT_mux_out_1_18_port, 
      DataPath_ALUhw_MULT_mux_out_1_19_port, 
      DataPath_ALUhw_MULT_mux_out_1_20_port, 
      DataPath_ALUhw_MULT_mux_out_1_26_port, 
      DataPath_ALUhw_MULT_mux_out_1_28_port, 
      DataPath_ALUhw_MULT_mux_out_1_31_port, 
      DataPath_ALUhw_MULT_mux_out_0_0_port, 
      DataPath_ALUhw_MULT_mux_out_0_1_port, 
      DataPath_ALUhw_MULT_mux_out_0_10_port, 
      DataPath_ALUhw_MULT_mux_out_0_11_port, 
      DataPath_ALUhw_MULT_mux_out_0_13_port, 
      DataPath_ALUhw_MULT_mux_out_0_14_port, 
      DataPath_ALUhw_MULT_mux_out_0_15_port, 
      DataPath_ALUhw_MULT_mux_out_0_16_port, 
      DataPath_ALUhw_MULT_mux_out_0_17_port, 
      DataPath_ALUhw_MULT_mux_out_0_18_port, 
      DataPath_ALUhw_MULT_mux_out_0_19_port, 
      DataPath_ALUhw_MULT_mux_out_0_20_port, 
      DataPath_ALUhw_MULT_mux_out_0_22_port, 
      DataPath_ALUhw_MULT_mux_out_0_27_port, 
      DataPath_ALUhw_MULT_mux_out_0_29_port, 
      DataPath_ALUhw_MULT_mux_out_0_31_port, C620_DATA2_2, C620_DATA2_3, 
      C620_DATA2_4, C620_DATA2_5, C620_DATA2_6, C620_DATA2_7, C620_DATA2_8, 
      C620_DATA2_9, C620_DATA2_10, C620_DATA2_11, C620_DATA2_12, C620_DATA2_13,
      C620_DATA2_14, C620_DATA2_15, C620_DATA2_20, C620_DATA2_21, C620_DATA2_27
      , C620_DATA2_29, C620_DATA2_30, C620_DATA2_31, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n104, n116, n171, n176, n181, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n210, 
      n220, n222, n224, n226, n230, n235, n368, n372, n373, n374, n375, n376, 
      n382, n383, n384, n385, n392, n393, n411, n415, n417, n472, n473, n476, 
      n477, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
      n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, 
      n525, n526, n527, n543, n544, n546, n548, n550, n552, n554, n556, n558, 
      n560, n562, n564, n566, n568, n570, n571, n572, n577, n596, n597, n598, 
      n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, 
      n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, 
      n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, 
      n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, 
      n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, 
      n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, 
      n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, 
      n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, 
      n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, 
      n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, 
      n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, 
      n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, 
      n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, 
      n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, 
      n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, 
      n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, 
      n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, 
      n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, 
      n815, n816, n817, n818, n819, n821, n822, n823, n824, n838, n851, n852, 
      n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, 
      n865, n866, n879, n883, n885, n887, n889, n891, n893, n895, n897, n899, 
      n901, n903, n905, n907, n909, n911, n913, n917, n919, n921, n923, n925, 
      n927, n929, n931, n933, n935, n937, n939, n941, n943, n945, n947, n948, 
      n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, 
      n961, n962, n966, n969, n970, n971, n972, n973, n974, n975, n976, n977, 
      n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, 
      n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1003, n1006,
      n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, 
      n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, 
      n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, 
      n1040, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, 
      n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, 
      n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, 
      n1072, n1073, n1077, n1080, n1081, n1082, n1083, n1084, n1085, n1086, 
      n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, 
      n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, 
      n1107, n1108, n1109, n1110, n1114, n1117, n1118, n1119, n1120, n1121, 
      n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, 
      n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, 
      n1142, n1143, n1144, n1145, n1146, n1147, n1151, n1154, n1155, n1156, 
      n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, 
      n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, 
      n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1188, n1191, 
      n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, 
      n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, 
      n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, 
      n1225, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, 
      n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, 
      n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, 
      n1257, n1258, n2106, n2228, n2260, n2287, n2288, n2289, n2290, n2291, 
      n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, 
      n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, 
      n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2441, n2443, n2445, 
      n2447, n2449, n2451, n2453, n2455, n2457, n2459, n2461, n2463, n2465, 
      n2467, n2469, n2474, n2478, n2480, n2483, n2486, n2489, n2491, n2494, 
      n2496, n2498, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, 
      n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, 
      n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, 
      n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, 
      n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, 
      n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, 
      n2871, n2872, n2873, n2874, n2876, n2882, n2883, n2884, n2885, n2886, 
      n2887, n2953, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, 
      n2963, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, 
      n2974, n2975, n2976, n2977, n2981, n2982, n2986, n2987, n2988, n2989, 
      n2990, n2992, n3006, n3009, n3010, n3274, n3280, n3324, n3327, n3328, 
      n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, 
      n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, 
      n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, 
      n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, 
      n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, 
      n3379, n3380, n3381, n3382, n3383, n3432, n3434, n3436, n3438, n3440, 
      n3442, n3444, n3446, n3448, n3450, n3452, n3454, n3456, n3458, n3460, 
      n3462, n3464, n3466, n3468, n3470, n3472, n3474, n3476, n3478, n3480, 
      n3482, n3484, n3486, n3488, n3490, n3492, n3499, n3502, n3503, n3504, 
      n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, 
      n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, 
      n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3537, n3540, 
      n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, 
      n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, 
      n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, 
      n3575, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, 
      n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, 
      n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, 
      n3607, n3608, n3613, n3616, n3617, n3618, n3619, n3620, n3621, n3622, 
      n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, 
      n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, 
      n3643, n3644, n3645, n3646, n3651, n3654, n3655, n3656, n3657, n3658, 
      n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, 
      n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, 
      n3679, n3680, n3681, n3682, n3683, n3684, n3689, n3692, n3693, n3694, 
      n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, 
      n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, 
      n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3727, n3730, 
      n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, 
      n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, 
      n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, 
      n3765, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, 
      n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, 
      n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, 
      n3797, n3798, n3800, n3803, n3804, n3805, n3806, n3807, n3808, n3809, 
      n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, 
      n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, 
      n3830, n3831, n3832, n3833, n3835, n3838, n3839, n3840, n3841, n3842, 
      n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, 
      n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, 
      n3863, n3864, n3865, n3866, n3867, n3868, n3870, n3873, n3874, n3875, 
      n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, 
      n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, 
      n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3905, n3908, 
      n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, 
      n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, 
      n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, 
      n3940, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, 
      n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, 
      n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, 
      n3972, n3973, n3975, n3978, n3979, n3980, n3981, n3982, n3983, n3984, 
      n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, 
      n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, 
      n4005, n4006, n4007, n4008, n4010, n4014, n4016, n4018, n4020, n4022, 
      n4024, n4026, n4028, n4030, n4032, n4034, n4036, n4038, n4040, n4042, 
      n4044, n4046, n4048, n4050, n4052, n4054, n4056, n4058, n4060, n4062, 
      n4064, n4066, n4068, n4070, n4072, n4074, n4077, n4081, n4083, n4085, 
      n4087, n4089, n4091, n4093, n4095, n4097, n4099, n4101, n4103, n4105, 
      n4107, n4109, n4111, n4113, n4115, n4117, n4119, n4121, n4123, n4125, 
      n4127, n4129, n4131, n4133, n4135, n4137, n4139, n4141, n4145, n4148, 
      n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, 
      n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, 
      n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, 
      n4180, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, 
      n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, 
      n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, 
      n4212, n4213, n4215, n4218, n4219, n4220, n4221, n4222, n4223, n4224, 
      n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, 
      n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, 
      n4245, n4246, n4247, n4248, n4250, n4253, n4254, n4255, n4256, n4257, 
      n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, 
      n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, 
      n4278, n4279, n4280, n4281, n4282, n4283, n4285, n4288, n4289, n4290, 
      n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, 
      n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, 
      n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4320, n4323, 
      n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, 
      n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, 
      n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, 
      n4355, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, 
      n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, 
      n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, 
      n4387, n4388, n4390, n4393, n4394, n4395, n4396, n4397, n4398, n4399, 
      n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, 
      n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, 
      n4420, n4421, n4422, n4423, n4425, n4428, n4429, n4430, n4431, n4432, 
      n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, 
      n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, 
      n4453, n4454, n4455, n4456, n4457, n4458, n4460, n4463, n4464, n4465, 
      n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, 
      n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, 
      n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4495, n4498, 
      n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, 
      n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, 
      n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, 
      n4530, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, 
      n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, 
      n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, 
      n4562, n4563, n4565, n4568, n4569, n4570, n4571, n4572, n4573, n4574, 
      n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, 
      n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, 
      n4595, n4596, n4597, n4598, n4600, n4603, n4604, n4605, n4606, n4607, 
      n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, 
      n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, 
      n4628, n4629, n4630, n4631, n4632, n4633, n4635, n4638, n4639, n4640, 
      n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, 
      n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, 
      n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4670, n4674, 
      n4676, n4678, n4680, n4682, n4684, n4686, n4688, n4690, n4692, n4694, 
      n4696, n4698, n4700, n4702, n4704, n4706, n4708, n4710, n4712, n4714, 
      n4716, n4718, n4720, n4722, n4724, n4726, n4728, n4730, n4732, n4734, 
      n4738, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, 
      n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, 
      n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, 
      n4770, n4771, n4773, n4776, n4777, n4778, n4779, n4780, n4781, n4782, 
      n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, 
      n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, 
      n4803, n4804, n4805, n4806, n4808, n4811, n4812, n4813, n4814, n4815, 
      n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, 
      n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, 
      n4836, n4837, n4838, n4839, n4840, n4841, n4843, n4846, n4847, n4848, 
      n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, 
      n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, 
      n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4878, n4881, 
      n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, 
      n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, 
      n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, 
      n4913, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, 
      n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, 
      n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, 
      n4945, n4946, n4948, n4951, n4952, n4953, n4954, n4955, n4956, n4957, 
      n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, 
      n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, 
      n4978, n4979, n4980, n4981, n4983, n4986, n4987, n4988, n4989, n4990, 
      n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, 
      n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, 
      n5011, n5012, n5013, n5014, n5015, n5016, n5018, n5021, n5022, n5023, 
      n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, 
      n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, 
      n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5053, n5056, 
      n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, 
      n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, 
      n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, 
      n5088, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, 
      n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, 
      n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, 
      n5120, n5121, n5123, n5126, n5127, n5128, n5129, n5130, n5131, n5132, 
      n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, 
      n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, 
      n5153, n5154, n5155, n5156, n5158, n5161, n5162, n5163, n5164, n5165, 
      n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, 
      n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, 
      n5186, n5187, n5188, n5189, n5190, n5191, n5193, n5196, n5197, n5198, 
      n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, 
      n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, 
      n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5228, n5231, 
      n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, 
      n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, 
      n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, 
      n5263, n5267, n5269, n5271, n5273, n5275, n5277, n5279, n5281, n5283, 
      n5285, n5287, n5289, n5291, n5293, n5295, n5297, n5299, n5301, n5303, 
      n5305, n5307, n5309, n5311, n5313, n5315, n5317, n5319, n5321, n5323, 
      n5325, n5327, n5331, n5334, n5335, n5336, n5337, n5338, n5339, n5340, 
      n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, 
      n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, 
      n5361, n5362, n5363, n5364, n5366, n5369, n5370, n5371, n5372, n5373, 
      n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, 
      n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, 
      n5394, n5395, n5396, n5397, n5398, n5399, n5401, n5404, n5405, n5406, 
      n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, 
      n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, 
      n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5436, n5439, 
      n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, 
      n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, 
      n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, 
      n5471, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, 
      n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, 
      n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, 
      n5503, n5504, n5506, n5509, n5510, n5511, n5512, n5513, n5514, n5515, 
      n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, 
      n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, 
      n5536, n5537, n5538, n5539, n5541, n5544, n5545, n5546, n5547, n5548, 
      n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, 
      n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, 
      n5569, n5570, n5571, n5572, n5573, n5574, n5576, n5579, n5580, n5581, 
      n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, 
      n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, 
      n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5614, n5615, 
      n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, 
      n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, 
      n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, 
      n5648, n5650, n5651, n5654, n5655, n5656, n5657, n5658, n5659, n5660, 
      n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, 
      n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, 
      n5681, n5682, n5683, n5684, n5686, n5687, n5690, n5691, n5692, n5693, 
      n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, 
      n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, 
      n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5722, n5723, n5726, 
      n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, 
      n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, 
      n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, 
      n5758, n5759, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, 
      n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, 
      n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, 
      n5790, n5791, n5792, n5794, n5795, n5798, n5799, n5800, n5801, n5802, 
      n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, 
      n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, 
      n5823, n5824, n5825, n5826, n5827, n5828, n5830, n5831, n5834, n5835, 
      n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, 
      n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, 
      n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5867, 
      n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, 
      n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, 
      n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, 
      n5900, n5905, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, 
      n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, 
      n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, 
      n5936, n5937, n5938, n5941, n5942, n5945, n5946, n5947, n5948, n5949, 
      n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, 
      n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, 
      n5970, n5971, n5972, n5973, n5974, n5975, n5978, n5979, n5982, n5983, 
      n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, 
      n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, 
      n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6015, 
      n6016, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, 
      n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, 
      n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, 
      n6048, n6049, n6052, n6053, n6056, n6057, n6058, n6059, n6060, n6061, 
      n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, 
      n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, 
      n6082, n6083, n6084, n6085, n6086, n6089, n6090, n6093, n6094, n6095, 
      n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, 
      n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, 
      n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6126, n6127, 
      n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, 
      n6138, n6139, n6140, n6141, n6142, n6146, n6730, n6731, n6732, n6733, 
      n6734, n6735, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, 
      n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, 
      n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, 
      n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805, 
      n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, 
      n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, 
      n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, 
      n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, 
      n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, 
      n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, 
      n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, 
      n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885, 
      n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895, 
      n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905, 
      n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915, 
      n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925, 
      n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935, 
      n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, 
      n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955, 
      n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, 
      n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, 
      n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, 
      n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995, 
      n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, 
      n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, 
      n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, 
      n7026, n7027, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, 
      n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, 
      n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, 
      n7059, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, 
      n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, 
      n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7104, n7105, 
      n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, 
      n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, 
      n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, 
      n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, 
      n7147, n7148, n7149, n7151, n7152, n7153, intadd_0_A_0_port, 
      intadd_1_A_1_port, intadd_1_A_0_port, DP_OP_1090J1_126_7243_n75, 
      DP_OP_1090J1_126_7243_n72, DP_OP_1090J1_126_7243_n37, 
      DP_OP_1090J1_126_7243_n30, DP_OP_1090J1_126_7243_n29, 
      DP_OP_1090J1_126_7243_n28, DP_OP_1090J1_126_7243_n27, 
      DP_OP_1090J1_126_7243_n26, DP_OP_1090J1_126_7243_n25, 
      DP_OP_1090J1_126_7243_n24, DP_OP_1090J1_126_7243_n23, 
      DP_OP_1090J1_126_7243_n22, DP_OP_1090J1_126_7243_n21, 
      DP_OP_1090J1_126_7243_n20, DP_OP_1090J1_126_7243_n19, 
      DP_OP_1090J1_126_7243_n18, DP_OP_1090J1_126_7243_n17, 
      DP_OP_1090J1_126_7243_n16, DP_OP_1090J1_126_7243_n14, 
      DP_OP_1090J1_126_7243_n13, DP_OP_1090J1_126_7243_n12, 
      DP_OP_1090J1_126_7243_n11, DP_OP_1090J1_126_7243_n9, 
      DP_OP_1090J1_126_7243_n1, DP_OP_751_130_5637_I2, DP_OP_751_130_5637_n1828
      , DP_OP_751_130_5637_n1816, DP_OP_751_130_5637_n1815, 
      DP_OP_751_130_5637_n1814, DP_OP_751_130_5637_n1813, 
      DP_OP_751_130_5637_n1812, DP_OP_751_130_5637_n1811, 
      DP_OP_751_130_5637_n1810, DP_OP_751_130_5637_n1809, 
      DP_OP_751_130_5637_n1807, DP_OP_751_130_5637_n1798, 
      DP_OP_751_130_5637_n1795, DP_OP_751_130_5637_n1794, 
      DP_OP_751_130_5637_n1792, DP_OP_751_130_5637_n1781, 
      DP_OP_751_130_5637_n1780, DP_OP_751_130_5637_n1779, 
      DP_OP_751_130_5637_n1778, DP_OP_751_130_5637_n1777, 
      DP_OP_751_130_5637_n1776, DP_OP_751_130_5637_n1775, 
      DP_OP_751_130_5637_n1774, DP_OP_751_130_5637_n1773, 
      DP_OP_751_130_5637_n1772, DP_OP_751_130_5637_n1771, 
      DP_OP_751_130_5637_n1770, DP_OP_751_130_5637_n1769, 
      DP_OP_751_130_5637_n1768, DP_OP_751_130_5637_n1767, 
      DP_OP_751_130_5637_n1765, DP_OP_751_130_5637_n1764, 
      DP_OP_751_130_5637_n1763, DP_OP_751_130_5637_n1761, 
      DP_OP_751_130_5637_n1760, DP_OP_751_130_5637_n1750, 
      DP_OP_751_130_5637_n1749, DP_OP_751_130_5637_n1748, 
      DP_OP_751_130_5637_n1747, DP_OP_751_130_5637_n1746, 
      DP_OP_751_130_5637_n1745, DP_OP_751_130_5637_n1743, 
      DP_OP_751_130_5637_n1742, DP_OP_751_130_5637_n1740, 
      DP_OP_751_130_5637_n1739, DP_OP_751_130_5637_n1738, 
      DP_OP_751_130_5637_n1737, DP_OP_751_130_5637_n1736, 
      DP_OP_751_130_5637_n1734, DP_OP_751_130_5637_n1733, 
      DP_OP_751_130_5637_n1732, DP_OP_751_130_5637_n1727, 
      DP_OP_751_130_5637_n1726, DP_OP_751_130_5637_n1725, 
      DP_OP_751_130_5637_n1724, DP_OP_751_130_5637_n1723, 
      DP_OP_751_130_5637_n1722, DP_OP_751_130_5637_n1721, 
      DP_OP_751_130_5637_n1720, DP_OP_751_130_5637_n1719, 
      DP_OP_751_130_5637_n1718, DP_OP_751_130_5637_n1717, 
      DP_OP_751_130_5637_n1716, DP_OP_751_130_5637_n1715, 
      DP_OP_751_130_5637_n1714, DP_OP_751_130_5637_n1713, 
      DP_OP_751_130_5637_n1712, DP_OP_751_130_5637_n1711, 
      DP_OP_751_130_5637_n1710, DP_OP_751_130_5637_n1709, 
      DP_OP_751_130_5637_n1708, DP_OP_751_130_5637_n1707, 
      DP_OP_751_130_5637_n1706, DP_OP_751_130_5637_n1705, 
      DP_OP_751_130_5637_n1704, DP_OP_751_130_5637_n1703, 
      DP_OP_751_130_5637_n1702, DP_OP_751_130_5637_n1701, 
      DP_OP_751_130_5637_n1700, DP_OP_751_130_5637_n1699, 
      DP_OP_751_130_5637_n1698, DP_OP_751_130_5637_n1697, 
      DP_OP_751_130_5637_n1696, DP_OP_751_130_5637_n1695, 
      DP_OP_751_130_5637_n1694, DP_OP_751_130_5637_n1693, 
      DP_OP_751_130_5637_n1692, DP_OP_751_130_5637_n1691, 
      DP_OP_751_130_5637_n1690, DP_OP_751_130_5637_n1689, 
      DP_OP_751_130_5637_n1688, DP_OP_751_130_5637_n1687, 
      DP_OP_751_130_5637_n1686, DP_OP_751_130_5637_n1685, 
      DP_OP_751_130_5637_n1684, DP_OP_751_130_5637_n1683, 
      DP_OP_751_130_5637_n1682, DP_OP_751_130_5637_n1681, 
      DP_OP_751_130_5637_n1680, DP_OP_751_130_5637_n1679, 
      DP_OP_751_130_5637_n1678, DP_OP_751_130_5637_n1677, 
      DP_OP_751_130_5637_n1676, DP_OP_751_130_5637_n1675, 
      DP_OP_751_130_5637_n1674, DP_OP_751_130_5637_n1673, 
      DP_OP_751_130_5637_n1672, DP_OP_751_130_5637_n1671, 
      DP_OP_751_130_5637_n1670, DP_OP_751_130_5637_n1669, 
      DP_OP_751_130_5637_n1668, DP_OP_751_130_5637_n1659, 
      DP_OP_751_130_5637_n1657, DP_OP_751_130_5637_n1656, 
      DP_OP_751_130_5637_n1655, DP_OP_751_130_5637_n1654, 
      DP_OP_751_130_5637_n1653, DP_OP_751_130_5637_n1652, 
      DP_OP_751_130_5637_n1651, DP_OP_751_130_5637_n1650, 
      DP_OP_751_130_5637_n1649, DP_OP_751_130_5637_n1648, 
      DP_OP_751_130_5637_n1647, DP_OP_751_130_5637_n1646, 
      DP_OP_751_130_5637_n1645, DP_OP_751_130_5637_n1644, 
      DP_OP_751_130_5637_n1643, DP_OP_751_130_5637_n1642, 
      DP_OP_751_130_5637_n1641, DP_OP_751_130_5637_n1640, 
      DP_OP_751_130_5637_n1639, DP_OP_751_130_5637_n1638, 
      DP_OP_751_130_5637_n1637, DP_OP_751_130_5637_n1636, 
      DP_OP_751_130_5637_n1635, DP_OP_751_130_5637_n1634, 
      DP_OP_751_130_5637_n1633, DP_OP_751_130_5637_n1632, 
      DP_OP_751_130_5637_n1631, DP_OP_751_130_5637_n1624, 
      DP_OP_751_130_5637_n1623, DP_OP_751_130_5637_n1622, 
      DP_OP_751_130_5637_n1621, DP_OP_751_130_5637_n1620, 
      DP_OP_751_130_5637_n1619, DP_OP_751_130_5637_n1618, 
      DP_OP_751_130_5637_n1617, DP_OP_751_130_5637_n1616, 
      DP_OP_751_130_5637_n1615, DP_OP_751_130_5637_n1614, 
      DP_OP_751_130_5637_n1613, DP_OP_751_130_5637_n1612, 
      DP_OP_751_130_5637_n1611, DP_OP_751_130_5637_n1610, 
      DP_OP_751_130_5637_n1609, DP_OP_751_130_5637_n1608, 
      DP_OP_751_130_5637_n1607, DP_OP_751_130_5637_n1606, 
      DP_OP_751_130_5637_n1605, DP_OP_751_130_5637_n1604, 
      DP_OP_751_130_5637_n1603, DP_OP_751_130_5637_n1602, 
      DP_OP_751_130_5637_n1601, DP_OP_751_130_5637_n1600, 
      DP_OP_751_130_5637_n1599, DP_OP_751_130_5637_n1598, 
      DP_OP_751_130_5637_n1597, DP_OP_751_130_5637_n1596, 
      DP_OP_751_130_5637_n1595, DP_OP_751_130_5637_n1594, 
      DP_OP_751_130_5637_n1593, DP_OP_751_130_5637_n1592, 
      DP_OP_751_130_5637_n1591, DP_OP_751_130_5637_n1589, 
      DP_OP_751_130_5637_n1588, DP_OP_751_130_5637_n1587, 
      DP_OP_751_130_5637_n1584, DP_OP_751_130_5637_n1583, 
      DP_OP_751_130_5637_n1581, DP_OP_751_130_5637_n1580, 
      DP_OP_751_130_5637_n1579, DP_OP_751_130_5637_n1577, 
      DP_OP_751_130_5637_n1576, DP_OP_751_130_5637_n1575, 
      DP_OP_751_130_5637_n1574, DP_OP_751_130_5637_n1573, 
      DP_OP_751_130_5637_n1572, DP_OP_751_130_5637_n1571, 
      DP_OP_751_130_5637_n1570, DP_OP_751_130_5637_n1557, 
      DP_OP_751_130_5637_n1555, DP_OP_751_130_5637_n1554, 
      DP_OP_751_130_5637_n1553, DP_OP_751_130_5637_n1552, 
      DP_OP_751_130_5637_n1551, DP_OP_751_130_5637_n1550, 
      DP_OP_751_130_5637_n1549, DP_OP_751_130_5637_n1548, 
      DP_OP_751_130_5637_n1547, DP_OP_751_130_5637_n1546, 
      DP_OP_751_130_5637_n1545, DP_OP_751_130_5637_n1544, 
      DP_OP_751_130_5637_n1543, DP_OP_751_130_5637_n1542, 
      DP_OP_751_130_5637_n1541, DP_OP_751_130_5637_n1540, 
      DP_OP_751_130_5637_n1539, DP_OP_751_130_5637_n1538, 
      DP_OP_751_130_5637_n1537, DP_OP_751_130_5637_n1536, 
      DP_OP_751_130_5637_n1535, DP_OP_751_130_5637_n1534, 
      DP_OP_751_130_5637_n1533, DP_OP_751_130_5637_n1532, 
      DP_OP_751_130_5637_n1531, DP_OP_751_130_5637_n1522, 
      DP_OP_751_130_5637_n1521, DP_OP_751_130_5637_n1520, 
      DP_OP_751_130_5637_n1519, DP_OP_751_130_5637_n1518, 
      DP_OP_751_130_5637_n1517, DP_OP_751_130_5637_n1516, 
      DP_OP_751_130_5637_n1515, DP_OP_751_130_5637_n1514, 
      DP_OP_751_130_5637_n1513, DP_OP_751_130_5637_n1512, 
      DP_OP_751_130_5637_n1511, DP_OP_751_130_5637_n1510, 
      DP_OP_751_130_5637_n1509, DP_OP_751_130_5637_n1508, 
      DP_OP_751_130_5637_n1507, DP_OP_751_130_5637_n1506, 
      DP_OP_751_130_5637_n1505, DP_OP_751_130_5637_n1504, 
      DP_OP_751_130_5637_n1503, DP_OP_751_130_5637_n1502, 
      DP_OP_751_130_5637_n1501, DP_OP_751_130_5637_n1500, 
      DP_OP_751_130_5637_n1499, DP_OP_751_130_5637_n1498, 
      DP_OP_751_130_5637_n1497, DP_OP_751_130_5637_n1496, 
      DP_OP_751_130_5637_n1495, DP_OP_751_130_5637_n1494, 
      DP_OP_751_130_5637_n1493, DP_OP_751_130_5637_n1492, 
      DP_OP_751_130_5637_n1491, DP_OP_751_130_5637_n1490, 
      DP_OP_751_130_5637_n1489, DP_OP_751_130_5637_n1488, 
      DP_OP_751_130_5637_n1487, DP_OP_751_130_5637_n1486, 
      DP_OP_751_130_5637_n1485, DP_OP_751_130_5637_n1484, 
      DP_OP_751_130_5637_n1483, DP_OP_751_130_5637_n1481, 
      DP_OP_751_130_5637_n1480, DP_OP_751_130_5637_n1479, 
      DP_OP_751_130_5637_n1477, DP_OP_751_130_5637_n1476, 
      DP_OP_751_130_5637_n1475, DP_OP_751_130_5637_n1473, 
      DP_OP_751_130_5637_n1472, DP_OP_751_130_5637_n1455, 
      DP_OP_751_130_5637_n1453, DP_OP_751_130_5637_n1452, 
      DP_OP_751_130_5637_n1451, DP_OP_751_130_5637_n1450, 
      DP_OP_751_130_5637_n1449, DP_OP_751_130_5637_n1448, 
      DP_OP_751_130_5637_n1447, DP_OP_751_130_5637_n1446, 
      DP_OP_751_130_5637_n1445, DP_OP_751_130_5637_n1444, 
      DP_OP_751_130_5637_n1443, DP_OP_751_130_5637_n1442, 
      DP_OP_751_130_5637_n1441, DP_OP_751_130_5637_n1440, 
      DP_OP_751_130_5637_n1439, DP_OP_751_130_5637_n1438, 
      DP_OP_751_130_5637_n1437, DP_OP_751_130_5637_n1436, 
      DP_OP_751_130_5637_n1435, DP_OP_751_130_5637_n1434, 
      DP_OP_751_130_5637_n1433, DP_OP_751_130_5637_n1432, 
      DP_OP_751_130_5637_n1431, DP_OP_751_130_5637_n1420, 
      DP_OP_751_130_5637_n1419, DP_OP_751_130_5637_n1418, 
      DP_OP_751_130_5637_n1417, DP_OP_751_130_5637_n1416, 
      DP_OP_751_130_5637_n1415, DP_OP_751_130_5637_n1414, 
      DP_OP_751_130_5637_n1413, DP_OP_751_130_5637_n1412, 
      DP_OP_751_130_5637_n1411, DP_OP_751_130_5637_n1410, 
      DP_OP_751_130_5637_n1409, DP_OP_751_130_5637_n1408, 
      DP_OP_751_130_5637_n1407, DP_OP_751_130_5637_n1406, 
      DP_OP_751_130_5637_n1405, DP_OP_751_130_5637_n1404, 
      DP_OP_751_130_5637_n1403, DP_OP_751_130_5637_n1402, 
      DP_OP_751_130_5637_n1401, DP_OP_751_130_5637_n1400, 
      DP_OP_751_130_5637_n1399, DP_OP_751_130_5637_n1398, 
      DP_OP_751_130_5637_n1397, DP_OP_751_130_5637_n1396, 
      DP_OP_751_130_5637_n1395, DP_OP_751_130_5637_n1394, 
      DP_OP_751_130_5637_n1393, DP_OP_751_130_5637_n1391, 
      DP_OP_751_130_5637_n1389, DP_OP_751_130_5637_n1388, 
      DP_OP_751_130_5637_n1387, DP_OP_751_130_5637_n1386, 
      DP_OP_751_130_5637_n1385, DP_OP_751_130_5637_n1384, 
      DP_OP_751_130_5637_n1381, DP_OP_751_130_5637_n1380, 
      DP_OP_751_130_5637_n1377, DP_OP_751_130_5637_n1376, 
      DP_OP_751_130_5637_n1375, DP_OP_751_130_5637_n1374, 
      DP_OP_751_130_5637_n1353, DP_OP_751_130_5637_n1352, 
      DP_OP_751_130_5637_n1351, DP_OP_751_130_5637_n1350, 
      DP_OP_751_130_5637_n1349, DP_OP_751_130_5637_n1348, 
      DP_OP_751_130_5637_n1347, DP_OP_751_130_5637_n1346, 
      DP_OP_751_130_5637_n1345, DP_OP_751_130_5637_n1344, 
      DP_OP_751_130_5637_n1343, DP_OP_751_130_5637_n1342, 
      DP_OP_751_130_5637_n1341, DP_OP_751_130_5637_n1340, 
      DP_OP_751_130_5637_n1339, DP_OP_751_130_5637_n1338, 
      DP_OP_751_130_5637_n1337, DP_OP_751_130_5637_n1336, 
      DP_OP_751_130_5637_n1335, DP_OP_751_130_5637_n1334, 
      DP_OP_751_130_5637_n1333, DP_OP_751_130_5637_n1332, 
      DP_OP_751_130_5637_n1331, DP_OP_751_130_5637_n1318, 
      DP_OP_751_130_5637_n1317, DP_OP_751_130_5637_n1316, 
      DP_OP_751_130_5637_n1315, DP_OP_751_130_5637_n1314, 
      DP_OP_751_130_5637_n1313, DP_OP_751_130_5637_n1312, 
      DP_OP_751_130_5637_n1311, DP_OP_751_130_5637_n1310, 
      DP_OP_751_130_5637_n1309, DP_OP_751_130_5637_n1308, 
      DP_OP_751_130_5637_n1307, DP_OP_751_130_5637_n1306, 
      DP_OP_751_130_5637_n1305, DP_OP_751_130_5637_n1304, 
      DP_OP_751_130_5637_n1303, DP_OP_751_130_5637_n1302, 
      DP_OP_751_130_5637_n1301, DP_OP_751_130_5637_n1300, 
      DP_OP_751_130_5637_n1299, DP_OP_751_130_5637_n1298, 
      DP_OP_751_130_5637_n1297, DP_OP_751_130_5637_n1296, 
      DP_OP_751_130_5637_n1295, DP_OP_751_130_5637_n1294, 
      DP_OP_751_130_5637_n1293, DP_OP_751_130_5637_n1292, 
      DP_OP_751_130_5637_n1291, DP_OP_751_130_5637_n1290, 
      DP_OP_751_130_5637_n1289, DP_OP_751_130_5637_n1288, 
      DP_OP_751_130_5637_n1287, DP_OP_751_130_5637_n1286, 
      DP_OP_751_130_5637_n1285, DP_OP_751_130_5637_n1284, 
      DP_OP_751_130_5637_n1283, DP_OP_751_130_5637_n1282, 
      DP_OP_751_130_5637_n1281, DP_OP_751_130_5637_n1280, 
      DP_OP_751_130_5637_n1279, DP_OP_751_130_5637_n1277, 
      DP_OP_751_130_5637_n1276, DP_OP_751_130_5637_n1251, 
      DP_OP_751_130_5637_n1249, DP_OP_751_130_5637_n1248, 
      DP_OP_751_130_5637_n1247, DP_OP_751_130_5637_n1246, 
      DP_OP_751_130_5637_n1245, DP_OP_751_130_5637_n1244, 
      DP_OP_751_130_5637_n1243, DP_OP_751_130_5637_n1242, 
      DP_OP_751_130_5637_n1241, DP_OP_751_130_5637_n1240, 
      DP_OP_751_130_5637_n1239, DP_OP_751_130_5637_n1238, 
      DP_OP_751_130_5637_n1237, DP_OP_751_130_5637_n1236, 
      DP_OP_751_130_5637_n1235, DP_OP_751_130_5637_n1234, 
      DP_OP_751_130_5637_n1233, DP_OP_751_130_5637_n1232, 
      DP_OP_751_130_5637_n1231, DP_OP_751_130_5637_n1216, 
      DP_OP_751_130_5637_n1215, DP_OP_751_130_5637_n1214, 
      DP_OP_751_130_5637_n1213, DP_OP_751_130_5637_n1212, 
      DP_OP_751_130_5637_n1211, DP_OP_751_130_5637_n1210, 
      DP_OP_751_130_5637_n1209, DP_OP_751_130_5637_n1208, 
      DP_OP_751_130_5637_n1207, DP_OP_751_130_5637_n1206, 
      DP_OP_751_130_5637_n1205, DP_OP_751_130_5637_n1204, 
      DP_OP_751_130_5637_n1203, DP_OP_751_130_5637_n1202, 
      DP_OP_751_130_5637_n1201, DP_OP_751_130_5637_n1200, 
      DP_OP_751_130_5637_n1199, DP_OP_751_130_5637_n1198, 
      DP_OP_751_130_5637_n1197, DP_OP_751_130_5637_n1196, 
      DP_OP_751_130_5637_n1195, DP_OP_751_130_5637_n1194, 
      DP_OP_751_130_5637_n1193, DP_OP_751_130_5637_n1192, 
      DP_OP_751_130_5637_n1191, DP_OP_751_130_5637_n1190, 
      DP_OP_751_130_5637_n1189, DP_OP_751_130_5637_n1188, 
      DP_OP_751_130_5637_n1187, DP_OP_751_130_5637_n1186, 
      DP_OP_751_130_5637_n1185, DP_OP_751_130_5637_n1184, 
      DP_OP_751_130_5637_n1183, DP_OP_751_130_5637_n1182, 
      DP_OP_751_130_5637_n1181, DP_OP_751_130_5637_n1180, 
      DP_OP_751_130_5637_n1178, DP_OP_751_130_5637_n1149, 
      DP_OP_751_130_5637_n1147, DP_OP_751_130_5637_n1146, 
      DP_OP_751_130_5637_n1145, DP_OP_751_130_5637_n1144, 
      DP_OP_751_130_5637_n1143, DP_OP_751_130_5637_n1142, 
      DP_OP_751_130_5637_n1141, DP_OP_751_130_5637_n1140, 
      DP_OP_751_130_5637_n1139, DP_OP_751_130_5637_n1138, 
      DP_OP_751_130_5637_n1137, DP_OP_751_130_5637_n1136, 
      DP_OP_751_130_5637_n1135, DP_OP_751_130_5637_n1134, 
      DP_OP_751_130_5637_n1133, DP_OP_751_130_5637_n1132, 
      DP_OP_751_130_5637_n1131, DP_OP_751_130_5637_n1114, 
      DP_OP_751_130_5637_n1113, DP_OP_751_130_5637_n1112, 
      DP_OP_751_130_5637_n1111, DP_OP_751_130_5637_n1110, 
      DP_OP_751_130_5637_n1109, DP_OP_751_130_5637_n1108, 
      DP_OP_751_130_5637_n1107, DP_OP_751_130_5637_n1106, 
      DP_OP_751_130_5637_n1105, DP_OP_751_130_5637_n1104, 
      DP_OP_751_130_5637_n1103, DP_OP_751_130_5637_n1102, 
      DP_OP_751_130_5637_n1101, DP_OP_751_130_5637_n1100, 
      DP_OP_751_130_5637_n1099, DP_OP_751_130_5637_n1098, 
      DP_OP_751_130_5637_n1097, DP_OP_751_130_5637_n1096, 
      DP_OP_751_130_5637_n1095, DP_OP_751_130_5637_n1094, 
      DP_OP_751_130_5637_n1093, DP_OP_751_130_5637_n1092, 
      DP_OP_751_130_5637_n1091, DP_OP_751_130_5637_n1090, 
      DP_OP_751_130_5637_n1089, DP_OP_751_130_5637_n1088, 
      DP_OP_751_130_5637_n1087, DP_OP_751_130_5637_n1086, 
      DP_OP_751_130_5637_n1085, DP_OP_751_130_5637_n1084, 
      DP_OP_751_130_5637_n1083, DP_OP_751_130_5637_n1082, 
      DP_OP_751_130_5637_n1081, DP_OP_751_130_5637_n1080, 
      DP_OP_751_130_5637_n1047, DP_OP_751_130_5637_n1046, 
      DP_OP_751_130_5637_n1045, DP_OP_751_130_5637_n1044, 
      DP_OP_751_130_5637_n1043, DP_OP_751_130_5637_n1042, 
      DP_OP_751_130_5637_n1041, DP_OP_751_130_5637_n1040, 
      DP_OP_751_130_5637_n1039, DP_OP_751_130_5637_n1038, 
      DP_OP_751_130_5637_n1037, DP_OP_751_130_5637_n1036, 
      DP_OP_751_130_5637_n1035, DP_OP_751_130_5637_n1034, 
      DP_OP_751_130_5637_n1033, DP_OP_751_130_5637_n1032, 
      DP_OP_751_130_5637_n1031, DP_OP_751_130_5637_n1012, 
      DP_OP_751_130_5637_n1011, DP_OP_751_130_5637_n1010, 
      DP_OP_751_130_5637_n1009, DP_OP_751_130_5637_n1008, 
      DP_OP_751_130_5637_n1007, DP_OP_751_130_5637_n1006, 
      DP_OP_751_130_5637_n1005, DP_OP_751_130_5637_n1004, 
      DP_OP_751_130_5637_n1003, DP_OP_751_130_5637_n1002, 
      DP_OP_751_130_5637_n1001, DP_OP_751_130_5637_n1000, 
      DP_OP_751_130_5637_n999, DP_OP_751_130_5637_n998, DP_OP_751_130_5637_n997
      , DP_OP_751_130_5637_n996, DP_OP_751_130_5637_n995, 
      DP_OP_751_130_5637_n994, DP_OP_751_130_5637_n993, DP_OP_751_130_5637_n992
      , DP_OP_751_130_5637_n991, DP_OP_751_130_5637_n990, 
      DP_OP_751_130_5637_n989, DP_OP_751_130_5637_n988, DP_OP_751_130_5637_n987
      , DP_OP_751_130_5637_n986, DP_OP_751_130_5637_n985, 
      DP_OP_751_130_5637_n984, DP_OP_751_130_5637_n983, DP_OP_751_130_5637_n982
      , DP_OP_751_130_5637_n945, DP_OP_751_130_5637_n943, 
      DP_OP_751_130_5637_n942, DP_OP_751_130_5637_n941, DP_OP_751_130_5637_n940
      , DP_OP_751_130_5637_n939, DP_OP_751_130_5637_n938, 
      DP_OP_751_130_5637_n937, DP_OP_751_130_5637_n936, DP_OP_751_130_5637_n935
      , DP_OP_751_130_5637_n934, DP_OP_751_130_5637_n933, 
      DP_OP_751_130_5637_n932, DP_OP_751_130_5637_n931, DP_OP_751_130_5637_n910
      , DP_OP_751_130_5637_n909, DP_OP_751_130_5637_n908, 
      DP_OP_751_130_5637_n907, DP_OP_751_130_5637_n906, DP_OP_751_130_5637_n905
      , DP_OP_751_130_5637_n904, DP_OP_751_130_5637_n903, 
      DP_OP_751_130_5637_n902, DP_OP_751_130_5637_n901, DP_OP_751_130_5637_n900
      , DP_OP_751_130_5637_n899, DP_OP_751_130_5637_n898, 
      DP_OP_751_130_5637_n897, DP_OP_751_130_5637_n896, DP_OP_751_130_5637_n895
      , DP_OP_751_130_5637_n894, DP_OP_751_130_5637_n893, 
      DP_OP_751_130_5637_n892, DP_OP_751_130_5637_n891, DP_OP_751_130_5637_n890
      , DP_OP_751_130_5637_n889, DP_OP_751_130_5637_n888, 
      DP_OP_751_130_5637_n887, DP_OP_751_130_5637_n886, DP_OP_751_130_5637_n885
      , DP_OP_751_130_5637_n884, DP_OP_751_130_5637_n843, 
      DP_OP_751_130_5637_n842, DP_OP_751_130_5637_n841, DP_OP_751_130_5637_n840
      , DP_OP_751_130_5637_n839, DP_OP_751_130_5637_n838, 
      DP_OP_751_130_5637_n837, DP_OP_751_130_5637_n836, DP_OP_751_130_5637_n835
      , DP_OP_751_130_5637_n834, DP_OP_751_130_5637_n833, 
      DP_OP_751_130_5637_n832, DP_OP_751_130_5637_n831, DP_OP_751_130_5637_n808
      , DP_OP_751_130_5637_n807, DP_OP_751_130_5637_n806, 
      DP_OP_751_130_5637_n805, DP_OP_751_130_5637_n804, DP_OP_751_130_5637_n803
      , DP_OP_751_130_5637_n802, DP_OP_751_130_5637_n801, 
      DP_OP_751_130_5637_n800, DP_OP_751_130_5637_n799, DP_OP_751_130_5637_n798
      , DP_OP_751_130_5637_n797, DP_OP_751_130_5637_n796, 
      DP_OP_751_130_5637_n795, DP_OP_751_130_5637_n794, DP_OP_751_130_5637_n793
      , DP_OP_751_130_5637_n792, DP_OP_751_130_5637_n791, 
      DP_OP_751_130_5637_n790, DP_OP_751_130_5637_n789, DP_OP_751_130_5637_n788
      , DP_OP_751_130_5637_n787, DP_OP_751_130_5637_n786, 
      DP_OP_751_130_5637_n741, DP_OP_751_130_5637_n740, DP_OP_751_130_5637_n739
      , DP_OP_751_130_5637_n738, DP_OP_751_130_5637_n737, 
      DP_OP_751_130_5637_n736, DP_OP_751_130_5637_n735, DP_OP_751_130_5637_n734
      , DP_OP_751_130_5637_n733, DP_OP_751_130_5637_n732, 
      DP_OP_751_130_5637_n731, DP_OP_751_130_5637_n706, DP_OP_751_130_5637_n705
      , DP_OP_751_130_5637_n704, DP_OP_751_130_5637_n703, 
      DP_OP_751_130_5637_n702, DP_OP_751_130_5637_n701, DP_OP_751_130_5637_n700
      , DP_OP_751_130_5637_n699, DP_OP_751_130_5637_n698, 
      DP_OP_751_130_5637_n697, DP_OP_751_130_5637_n696, DP_OP_751_130_5637_n695
      , DP_OP_751_130_5637_n694, DP_OP_751_130_5637_n693, 
      DP_OP_751_130_5637_n692, DP_OP_751_130_5637_n689, DP_OP_751_130_5637_n688
      , DP_OP_751_130_5637_n639, DP_OP_751_130_5637_n638, 
      DP_OP_751_130_5637_n637, DP_OP_751_130_5637_n636, DP_OP_751_130_5637_n635
      , DP_OP_751_130_5637_n634, DP_OP_751_130_5637_n633, 
      DP_OP_751_130_5637_n632, DP_OP_751_130_5637_n631, DP_OP_751_130_5637_n604
      , DP_OP_751_130_5637_n603, DP_OP_751_130_5637_n602, 
      DP_OP_751_130_5637_n601, DP_OP_751_130_5637_n600, DP_OP_751_130_5637_n599
      , DP_OP_751_130_5637_n598, DP_OP_751_130_5637_n597, 
      DP_OP_751_130_5637_n596, DP_OP_751_130_5637_n595, DP_OP_751_130_5637_n594
      , DP_OP_751_130_5637_n593, DP_OP_751_130_5637_n592, 
      DP_OP_751_130_5637_n591, DP_OP_751_130_5637_n590, DP_OP_751_130_5637_n537
      , DP_OP_751_130_5637_n536, DP_OP_751_130_5637_n535, 
      DP_OP_751_130_5637_n534, DP_OP_751_130_5637_n533, DP_OP_751_130_5637_n532
      , DP_OP_751_130_5637_n531, DP_OP_751_130_5637_n502, 
      DP_OP_751_130_5637_n501, DP_OP_751_130_5637_n500, DP_OP_751_130_5637_n499
      , DP_OP_751_130_5637_n498, DP_OP_751_130_5637_n497, 
      DP_OP_751_130_5637_n494, DP_OP_751_130_5637_n493, DP_OP_751_130_5637_n492
      , DP_OP_751_130_5637_n435, DP_OP_751_130_5637_n434, 
      DP_OP_751_130_5637_n433, DP_OP_751_130_5637_n432, DP_OP_751_130_5637_n431
      , DP_OP_751_130_5637_n400, DP_OP_751_130_5637_n399, 
      DP_OP_751_130_5637_n398, DP_OP_751_130_5637_n396, DP_OP_751_130_5637_n394
      , DP_OP_751_130_5637_n333, DP_OP_751_130_5637_n332, 
      DP_OP_751_130_5637_n298, DP_OP_751_130_5637_n297, DP_OP_751_130_5637_n218
      , DP_OP_751_130_5637_n216, DP_OP_751_130_5637_n215, 
      DP_OP_751_130_5637_n213, DP_OP_751_130_5637_n211, DP_OP_751_130_5637_n209
      , DP_OP_751_130_5637_n206, DP_OP_751_130_5637_n201, 
      DP_OP_751_130_5637_n198, DP_OP_751_130_5637_n196, DP_OP_751_130_5637_n194
      , DP_OP_751_130_5637_n191, DP_OP_751_130_5637_n189, 
      DP_OP_751_130_5637_n187, DP_OP_751_130_5637_n186, DP_OP_751_130_5637_n185
      , DP_OP_751_130_5637_n184, DP_OP_751_130_5637_n183, 
      DP_OP_751_130_5637_n178, DP_OP_751_130_5637_n177, DP_OP_751_130_5637_n175
      , DP_OP_751_130_5637_n173, DP_OP_751_130_5637_n172, 
      DP_OP_751_130_5637_n171, DP_OP_751_130_5637_n170, DP_OP_751_130_5637_n169
      , DP_OP_751_130_5637_n167, DP_OP_751_130_5637_n165, 
      DP_OP_751_130_5637_n164, DP_OP_751_130_5637_n163, DP_OP_751_130_5637_n162
      , DP_OP_751_130_5637_n161, DP_OP_751_130_5637_n156, 
      DP_OP_751_130_5637_n155, DP_OP_751_130_5637_n153, DP_OP_751_130_5637_n151
      , DP_OP_751_130_5637_n150, DP_OP_751_130_5637_n149, 
      DP_OP_751_130_5637_n148, DP_OP_751_130_5637_n147, DP_OP_751_130_5637_n145
      , DP_OP_751_130_5637_n143, DP_OP_751_130_5637_n142, 
      DP_OP_751_130_5637_n141, DP_OP_751_130_5637_n140, DP_OP_751_130_5637_n139
      , DP_OP_751_130_5637_n137, DP_OP_751_130_5637_n135, 
      DP_OP_751_130_5637_n134, DP_OP_751_130_5637_n133, DP_OP_751_130_5637_n131
      , DP_OP_751_130_5637_n130, DP_OP_751_130_5637_n129, 
      DP_OP_751_130_5637_n128, DP_OP_751_130_5637_n127, DP_OP_751_130_5637_n125
      , DP_OP_751_130_5637_n123, DP_OP_751_130_5637_n122, 
      DP_OP_751_130_5637_n121, DP_OP_751_130_5637_n120, DP_OP_751_130_5637_n119
      , DP_OP_751_130_5637_n117, DP_OP_751_130_5637_n115, 
      DP_OP_751_130_5637_n114, DP_OP_751_130_5637_n113, DP_OP_751_130_5637_n112
      , DP_OP_751_130_5637_n111, DP_OP_751_130_5637_n107, 
      DP_OP_751_130_5637_n106, DP_OP_751_130_5637_n105, DP_OP_751_130_5637_n104
      , DP_OP_751_130_5637_n101, DP_OP_751_130_5637_n98, DP_OP_751_130_5637_n97
      , DP_OP_751_130_5637_n93, DP_OP_751_130_5637_n92, DP_OP_751_130_5637_n91,
      DP_OP_751_130_5637_n90, DP_OP_751_130_5637_n89, DP_OP_751_130_5637_n85, 
      DP_OP_751_130_5637_n84, DP_OP_751_130_5637_n83, DP_OP_751_130_5637_n82, 
      DP_OP_751_130_5637_n79, DP_OP_751_130_5637_n77, DP_OP_751_130_5637_n76, 
      DP_OP_751_130_5637_n75, DP_OP_751_130_5637_n72, DP_OP_751_130_5637_n71, 
      DP_OP_751_130_5637_n69, DP_OP_751_130_5637_n31, DP_OP_751_130_5637_n24, 
      DP_OP_751_130_5637_n23, DP_OP_751_130_5637_n21, DP_OP_751_130_5637_n20, 
      DP_OP_751_130_5637_n18, DP_OP_751_130_5637_n17, DP_OP_751_130_5637_n16, 
      DP_OP_751_130_5637_n15, DP_OP_751_130_5637_n14, DP_OP_751_130_5637_n13, 
      DP_OP_751_130_5637_n12, DP_OP_751_130_5637_n11, DP_OP_751_130_5637_n10, 
      DP_OP_751_130_5637_n9, DP_OP_751_130_5637_n8, DP_OP_751_130_5637_n7, 
      DP_OP_751_130_5637_n6, DP_OP_751_130_5637_n5, n7174, n7175, n7176, n7177,
      n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, 
      n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, 
      n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, 
      n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, 
      n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, 
      n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, 
      n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, 
      n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, 
      n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, 
      n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, 
      n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, 
      n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, 
      n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, 
      n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, 
      n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, 
      n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, 
      n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, 
      n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, 
      n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, 
      n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, 
      n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, 
      n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, 
      n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, 
      n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, 
      n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, 
      n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, 
      n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, 
      n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, 
      n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, 
      n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, 
      n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, 
      n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, 
      n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, 
      n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, 
      n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, 
      n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, 
      n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, 
      n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, 
      n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, 
      n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, 
      n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, 
      n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, 
      n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, 
      n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, 
      n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, 
      n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, 
      n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, 
      n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, 
      n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, 
      n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, 
      n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, 
      n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, 
      n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, 
      n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, 
      n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, 
      n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, 
      n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, 
      n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, 
      n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, 
      n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, 
      n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, 
      n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, 
      n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, 
      n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, 
      n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, 
      n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, 
      n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, 
      n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, 
      n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, 
      n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, 
      n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, 
      n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, 
      n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, 
      n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, 
      n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, 
      n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, 
      n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, 
      n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, 
      n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, 
      n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, 
      n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, 
      n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, 
      n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, 
      n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, 
      n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, 
      n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, 
      n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, 
      n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, 
      n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, 
      n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, 
      n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, 
      n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, 
      n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, 
      n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, 
      n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, 
      n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, 
      n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, 
      n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, 
      n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, 
      n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, 
      n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, 
      n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, 
      n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, 
      n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, 
      n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, 
      n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, 
      n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, 
      n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, 
      n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, 
      n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, 
      n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, 
      n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, 
      n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, 
      n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, 
      n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, 
      n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, 
      n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, 
      n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, 
      n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, 
      n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, 
      n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, 
      n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, 
      n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, 
      n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, 
      n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, 
      n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, 
      n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, 
      n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, 
      n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, 
      n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, 
      n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, 
      n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, 
      n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, 
      n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, 
      n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, 
      n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, 
      n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, 
      n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, 
      n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, 
      n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, 
      n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, 
      n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, 
      n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, 
      n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, 
      n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, 
      n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, 
      n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, 
      n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, 
      n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, 
      n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, 
      n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, 
      n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, 
      n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, 
      n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, 
      n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, 
      n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, 
      n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, 
      n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, 
      n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, 
      n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, 
      n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, 
      n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, 
      n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, 
      n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, 
      n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, 
      n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, 
      n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, 
      n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, 
      n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, 
      n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, 
      n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, 
      n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, 
      n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, 
      n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, 
      n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, 
      n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, 
      n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, 
      n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, 
      n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, 
      n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, 
      n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, 
      n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, 
      n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, 
      n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, 
      n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, 
      n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, 
      n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, 
      n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, 
      n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, 
      n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, 
      n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, 
      n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, 
      n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, 
      n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, 
      n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, 
      n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, 
      n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, 
      n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, 
      n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, 
      n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, 
      n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, 
      n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, 
      n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, 
      n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, 
      n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, 
      n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, 
      n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, 
      n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, 
      n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, 
      n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, 
      n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, 
      n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, 
      n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, 
      n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, 
      n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, 
      n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, 
      n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, 
      n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, 
      n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, 
      n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, 
      n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, 
      n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, 
      n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, 
      n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, 
      n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, 
      n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, 
      n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, 
      n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, 
      n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, 
      n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, 
      n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, 
      n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, 
      n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, 
      n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, 
      n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, 
      n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, 
      n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, 
      n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, 
      n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, 
      n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, 
      n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, 
      n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, 
      n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, 
      n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, 
      n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, 
      n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, 
      n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, 
      n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, 
      n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, 
      n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, 
      n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, 
      n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, 
      n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, 
      n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, 
      n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, 
      n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, 
      n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, 
      n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, 
      n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, 
      n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, 
      n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, 
      n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, 
      n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, 
      n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, 
      n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, 
      n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, 
      n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, 
      n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, 
      n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, 
      n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, 
      n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, 
      n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, 
      n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, 
      n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, 
      n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, 
      n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, 
      n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, 
      n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, 
      n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, 
      n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, 
      n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, 
      n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, 
      n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, 
      n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015, 
      n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024, 
      n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033, 
      n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042, 
      n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051, 
      n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060, 
      n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069, 
      n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078, 
      n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087, 
      n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096, 
      n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105, 
      n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114, 
      n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, 
      n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132, 
      n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141, 
      n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150, 
      n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159, 
      n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168, 
      n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177, 
      n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186, 
      n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195, 
      n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204, 
      n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213, 
      n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222, 
      n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231, 
      n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240, 
      n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249, 
      n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, 
      n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267, 
      n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276, 
      n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285, 
      n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294, 
      n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303, 
      n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312, 
      n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321, 
      n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330, 
      n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339, 
      n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348, 
      n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357, 
      n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, 
      n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375, 
      n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384, 
      n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393, 
      n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, 
      n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, 
      n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, 
      n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, 
      n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, 
      n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, 
      n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, 
      n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, 
      n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, 
      n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, 
      n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, 
      n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, 
      n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, 
      n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, 
      n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, 
      n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, 
      n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, 
      n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, 
      n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, 
      n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, 
      n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, 
      n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, 
      n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, 
      n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, 
      n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, 
      n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, 
      n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, 
      n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, 
      n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, 
      n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, 
      n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672, 
      n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681, 
      n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690, 
      n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699, 
      n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708, 
      n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717, 
      n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, 
      n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735, 
      n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744, 
      n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753, 
      n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762, 
      n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771, 
      n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780, 
      n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789, 
      n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798, 
      n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807, 
      n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, 
      n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825, 
      n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834, 
      n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843, 
      n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852, 
      n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861, 
      n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870, 
      n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879, 
      n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888, 
      n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897, 
      n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906, 
      n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915, 
      n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924, 
      n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, 
      n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, 
      n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951, 
      n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960, 
      n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969, 
      n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978, 
      n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987, 
      n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996, 
      n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005, 
      n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014, 
      n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023, 
      n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032, 
      n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041, 
      n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050, 
      n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059, 
      n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068, 
      n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077, 
      n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086, 
      n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095, 
      n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104, 
      n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113, 
      n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122, 
      n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131, 
      n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140, 
      n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149, 
      n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158, 
      n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167, 
      n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176, 
      n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185, 
      n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194, 
      n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203, 
      n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212, 
      n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221, 
      n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230, 
      n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, 
      n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, 
      n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, 
      n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, 
      n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, 
      n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, 
      n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, 
      n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, 
      n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, 
      n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, 
      n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, 
      n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, 
      n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, 
      n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356, 
      n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365, 
      n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374, 
      n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383, 
      n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392, 
      n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401, 
      n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410, 
      n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419, 
      n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428, 
      n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437, 
      n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446, 
      n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455, 
      n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464, 
      n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473, 
      n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482, 
      n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491, 
      n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500, 
      n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509, 
      n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518, 
      n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527, 
      n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536, 
      n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545, 
      n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, 
      n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563, 
      n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572, 
      n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581, 
      n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590, 
      n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599, 
      n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608, 
      n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617, 
      n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626, 
      n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635, 
      n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644, 
      n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, 
      n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, 
      n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, 
      n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, 
      n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, 
      n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698, 
      n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, 
      n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, 
      n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725, 
      n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734, 
      n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743, 
      n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752, 
      n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761, 
      n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770, 
      n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779, 
      n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788, 
      n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797, 
      n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, 
      n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, 
      n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824, 
      n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833, 
      n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842, 
      n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851, 
      n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, 
      n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869, 
      n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878, 
      n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887, 
      n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896, 
      n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905, 
      n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914, 
      n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923, 
      n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932, 
      n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941, 
      n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950, 
      n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959, 
      n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968, 
      n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977, 
      n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986, 
      n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995, 
      n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004, 
      n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013, 
      n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022, 
      n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031, 
      n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040, 
      n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049, 
      n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058, 
      n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067, 
      n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, 
      n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, 
      n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, 
      n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, 
      n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112, 
      n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121, 
      n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130, 
      n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139, 
      n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, 
      n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, 
      n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, 
      n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, 
      n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184, 
      n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193, 
      n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202, 
      n12203, n12204, n12205, n12206, n12207, n12208, n_1064, n_1065, n_1066, 
      n_1067, n_1068, n_1069, n_1070, n_1071, n_1072, n_1073, n_1074, n_1075, 
      n_1076, n_1077, n_1078, n_1079, n_1080, n_1081, n_1082, n_1083, n_1084, 
      n_1085, n_1086, n_1087, n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, 
      n_1094, n_1095, n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, 
      n_1103, n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111, 
      n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119, n_1120, 
      n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127, n_1128, n_1129, 
      n_1130, n_1131, n_1132, n_1133, n_1134, n_1135, n_1136, n_1137, n_1138, 
      n_1139, n_1140, n_1141, n_1142, n_1143, n_1144, n_1145, n_1146, n_1147, 
      n_1148, n_1149, n_1150, n_1151, n_1152, n_1153, n_1154, n_1155, n_1156, 
      n_1157, n_1158, n_1159, n_1160, n_1161, n_1162, n_1163, n_1164, n_1165, 
      n_1166, n_1167, n_1168, n_1169, n_1170, n_1171, n_1172, n_1173, n_1174, 
      n_1175, n_1176, n_1177, n_1178, n_1179, n_1180, n_1181, n_1182, n_1183, 
      n_1184, n_1185, n_1186, n_1187, n_1188, n_1189, n_1190, n_1191, n_1192, 
      n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199, n_1200, n_1201, 
      n_1202, n_1203, n_1204, n_1205, n_1206, n_1207, n_1208, n_1209, n_1210, 
      n_1211, n_1212, n_1213, n_1214, n_1215, n_1216, n_1217, n_1218, n_1219, 
      n_1220, n_1221, n_1222, n_1223, n_1224, n_1225, n_1226, n_1227, n_1228, 
      n_1229, n_1230, n_1231, n_1232, n_1233, n_1234, n_1235, n_1236, n_1237, 
      n_1238, n_1239, n_1240, n_1241, n_1242, n_1243, n_1244, n_1245, n_1246, 
      n_1247, n_1248, n_1249, n_1250, n_1251, n_1252, n_1253, n_1254, n_1255, 
      n_1256, n_1257, n_1258, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, 
      n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, 
      n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, 
      n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, 
      n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, 
      n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, 
      n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, 
      n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, 
      n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, 
      n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, 
      n_1346, n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, 
      n_1355, n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, 
      n_1364, n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, 
      n_1373, n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, 
      n_1382, n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, 
      n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, 
      n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, 
      n_1409, n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, 
      n_1418, n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, 
      n_1427, n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, 
      n_1436, n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, 
      n_1445, n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, 
      n_1454, n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, 
      n_1463, n_1464, n_1465, n_1466, n_1467, n_1468, n_1469, n_1470, n_1471, 
      n_1472, n_1473, n_1474, n_1475, n_1476, n_1477, n_1478, n_1479, n_1480, 
      n_1481, n_1482, n_1483, n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, 
      n_1490, n_1491, n_1492, n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, 
      n_1499, n_1500, n_1501, n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, 
      n_1508, n_1509, n_1510, n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, 
      n_1517, n_1518, n_1519, n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, 
      n_1526, n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534, 
      n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542, n_1543, 
      n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550, n_1551, n_1552, 
      n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559, n_1560, n_1561, 
      n_1562, n_1563, n_1564, n_1565, n_1566, n_1567, n_1568, n_1569, n_1570, 
      n_1571, n_1572, n_1573, n_1574, n_1575, n_1576, n_1577, n_1578, n_1579, 
      n_1580, n_1581, n_1582, n_1583, n_1584, n_1585, n_1586, n_1587, n_1588, 
      n_1589, n_1590, n_1591, n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, 
      n_1598, n_1599, n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, 
      n_1607, n_1608, n_1609, n_1610, n_1611, n_1612, n_1613, n_1614, n_1615, 
      n_1616, n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624, 
      n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, 
      n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, 
      n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, 
      n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, 
      n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, 
      n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, 
      n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, 
      n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, 
      n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, 
      n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, 
      n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, 
      n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, 
      n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, 
      n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, 
      n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, 
      n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, 
      n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, 
      n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, 
      n_1787, n_1788, n_1789, n_1790, n_1791, n_1792, n_1793, n_1794, n_1795, 
      n_1796, n_1797, n_1798, n_1799, n_1800, n_1801, n_1802, n_1803, n_1804, 
      n_1805, n_1806, n_1807, n_1808, n_1809, n_1810, n_1811, n_1812, n_1813, 
      n_1814, n_1815, n_1816, n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, 
      n_1823, n_1824, n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, 
      n_1832, n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840, 
      n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848, n_1849, 
      n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856, n_1857, n_1858, 
      n_1859, n_1860, n_1861, n_1862, n_1863, n_1864, n_1865, n_1866, n_1867, 
      n_1868, n_1869, n_1870, n_1871, n_1872, n_1873, n_1874, n_1875, n_1876, 
      n_1877, n_1878, n_1879, n_1880, n_1881, n_1882, n_1883, n_1884, n_1885, 
      n_1886, n_1887, n_1888, n_1889, n_1890, n_1891, n_1892, n_1893, n_1894, 
      n_1895, n_1896, n_1897, n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, 
      n_1904, n_1905, n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, 
      n_1913, n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921, 
      n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929, n_1930, 
      n_1931, n_1932, n_1933, n_1934, n_1935, n_1936, n_1937, n_1938, n_1939, 
      n_1940, n_1941, n_1942, n_1943, n_1944, n_1945, n_1946, n_1947, n_1948, 
      n_1949, n_1950, n_1951, n_1952, n_1953, n_1954, n_1955, n_1956, n_1957, 
      n_1958, n_1959, n_1960, n_1961, n_1962, n_1963, n_1964, n_1965, n_1966, 
      n_1967, n_1968, n_1969, n_1970, n_1971, n_1972, n_1973, n_1974, n_1975, 
      n_1976, n_1977, n_1978, n_1979, n_1980, n_1981, n_1982, n_1983, n_1984, 
      n_1985, n_1986, n_1987, n_1988, n_1989, n_1990, n_1991, n_1992, n_1993, 
      n_1994, n_1995, n_1996, n_1997, n_1998, n_1999, n_2000, n_2001, n_2002, 
      n_2003, n_2004, n_2005, n_2006, n_2007, n_2008, n_2009, n_2010, n_2011, 
      n_2012, n_2013, n_2014, n_2015, n_2016, n_2017, n_2018, n_2019, n_2020, 
      n_2021, n_2022, n_2023, n_2024, n_2025, n_2026, n_2027, n_2028, n_2029, 
      n_2030, n_2031, n_2032, n_2033, n_2034, n_2035, n_2036, n_2037, n_2038, 
      n_2039, n_2040, n_2041, n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, 
      n_2048, n_2049, n_2050, n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, 
      n_2057, n_2058, n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, 
      n_2066, n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074, 
      n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082, n_2083, 
      n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090, n_2091, n_2092, 
      n_2093, n_2094, n_2095, n_2096, n_2097, n_2098, n_2099, n_2100, n_2101, 
      n_2102, n_2103, n_2104, n_2105, n_2106, n_2107, n_2108, n_2109, n_2110, 
      n_2111, n_2112, n_2113, n_2114, n_2115, n_2116, n_2117, n_2118, n_2119, 
      n_2120, n_2121, n_2122, n_2123, n_2124, n_2125, n_2126, n_2127, n_2128, 
      n_2129, n_2130, n_2131, n_2132, n_2133, n_2134, n_2135, n_2136, n_2137, 
      n_2138, n_2139, n_2140, n_2141, n_2142, n_2143, n_2144, n_2145, n_2146, 
      n_2147, n_2148, n_2149, n_2150, n_2151, n_2152, n_2153, n_2154, n_2155, 
      n_2156, n_2157, n_2158, n_2159, n_2160, n_2161, n_2162, n_2163, n_2164, 
      n_2165, n_2166, n_2167, n_2168, n_2169, n_2170, n_2171, n_2172, n_2173, 
      n_2174, n_2175, n_2176, n_2177, n_2178, n_2179, n_2180, n_2181, n_2182, 
      n_2183, n_2184, n_2185, n_2186, n_2187, n_2188, n_2189, n_2190, n_2191, 
      n_2192, n_2193, n_2194, n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, 
      n_2201, n_2202, n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, 
      n_2210, n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218, 
      n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226, n_2227, 
      n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234, n_2235, n_2236, 
      n_2237, n_2238, n_2239, n_2240, n_2241, n_2242, n_2243, n_2244, n_2245, 
      n_2246, n_2247, n_2248, n_2249, n_2250, n_2251, n_2252, n_2253, n_2254, 
      n_2255, n_2256, n_2257, n_2258, n_2259, n_2260, n_2261, n_2262, n_2263, 
      n_2264, n_2265, n_2266, n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, 
      n_2273, n_2274, n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, 
      n_2282, n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290, 
      n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298, n_2299, 
      n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306, n_2307, n_2308, 
      n_2309, n_2310, n_2311, n_2312, n_2313, n_2314, n_2315, n_2316, n_2317, 
      n_2318, n_2319, n_2320, n_2321, n_2322, n_2323, n_2324, n_2325, n_2326, 
      n_2327, n_2328, n_2329, n_2330, n_2331, n_2332, n_2333, n_2334, n_2335, 
      n_2336, n_2337, n_2338, n_2339, n_2340, n_2341, n_2342, n_2343, n_2344, 
      n_2345, n_2346, n_2347, n_2348, n_2349, n_2350, n_2351, n_2352, n_2353, 
      n_2354, n_2355, n_2356, n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, 
      n_2363, n_2364, n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, 
      n_2372, n_2373, n_2374, n_2375, n_2376, n_2377, n_2378, n_2379, n_2380, 
      n_2381, n_2382, n_2383, n_2384, n_2385, n_2386, n_2387, n_2388, n_2389, 
      n_2390, n_2391, n_2392, n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, 
      n_2399, n_2400, n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, 
      n_2408, n_2409, n_2410, n_2411, n_2412, n_2413, n_2414, n_2415, n_2416, 
      n_2417, n_2418, n_2419, n_2420, n_2421, n_2422, n_2423, n_2424, n_2425, 
      n_2426, n_2427, n_2428, n_2429, n_2430, n_2431, n_2432, n_2433, n_2434, 
      n_2435, n_2436, n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, 
      n_2444, n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452, 
      n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460, n_2461, 
      n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468, n_2469, n_2470, 
      n_2471, n_2472, n_2473, n_2474, n_2475, n_2476, n_2477, n_2478, n_2479, 
      n_2480, n_2481, n_2482, n_2483, n_2484, n_2485, n_2486, n_2487, n_2488, 
      n_2489, n_2490, n_2491, n_2492, n_2493, n_2494, n_2495, n_2496, n_2497, 
      n_2498, n_2499, n_2500, n_2501, n_2502, n_2503, n_2504, n_2505, n_2506, 
      n_2507, n_2508, n_2509, n_2510, n_2511, n_2512, n_2513, n_2514, n_2515, 
      n_2516, n_2517, n_2518, n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, 
      n_2525, n_2526, n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, 
      n_2534, n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542, 
      n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550, n_2551, 
      n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558, n_2559, n_2560, 
      n_2561, n_2562, n_2563, n_2564, n_2565, n_2566, n_2567, n_2568, n_2569, 
      n_2570, n_2571, n_2572, n_2573, n_2574, n_2575, n_2576, n_2577, n_2578, 
      n_2579, n_2580, n_2581, n_2582, n_2583, n_2584, n_2585, n_2586, n_2587, 
      n_2588, n_2589, n_2590, n_2591, n_2592, n_2593, n_2594, n_2595, n_2596, 
      n_2597, n_2598, n_2599, n_2600, n_2601, n_2602, n_2603, n_2604, n_2605, 
      n_2606, n_2607, n_2608, n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, 
      n_2615, n_2616, n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, 
      n_2624, n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632, 
      n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640, n_2641, 
      n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648, n_2649, n_2650, 
      n_2651, n_2652, n_2653, n_2654, n_2655, n_2656, n_2657, n_2658, n_2659, 
      n_2660, n_2661, n_2662, n_2663, n_2664, n_2665, n_2666, n_2667, n_2668, 
      n_2669, n_2670, n_2671, n_2672, n_2673, n_2674, n_2675, n_2676, n_2677, 
      n_2678, n_2679, n_2680, n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, 
      n_2687, n_2688, n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, 
      n_2696, n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704, 
      n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712, n_2713, 
      n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720, n_2721, n_2722, 
      n_2723, n_2724, n_2725, n_2726, n_2727, n_2728, n_2729, n_2730, n_2731, 
      n_2732, n_2733, n_2734, n_2735, n_2736, n_2737, n_2738, n_2739, n_2740, 
      n_2741, n_2742, n_2743, n_2744, n_2745, n_2746, n_2747, n_2748, n_2749, 
      n_2750, n_2751, n_2752, n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, 
      n_2759, n_2760, n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, 
      n_2768, n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776, 
      n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784, n_2785, 
      n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792, n_2793, n_2794, 
      n_2795, n_2796, n_2797, n_2798, n_2799, n_2800, n_2801, n_2802, n_2803, 
      n_2804, n_2805, n_2806, n_2807, n_2808, n_2809, n_2810, n_2811, n_2812, 
      n_2813, n_2814, n_2815, n_2816, n_2817, n_2818, n_2819, n_2820, n_2821, 
      n_2822, n_2823, n_2824, n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, 
      n_2831, n_2832, n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839, 
      n_2840, n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848, 
      n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856, n_2857, 
      n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864, n_2865, n_2866, 
      n_2867, n_2868, n_2869, n_2870, n_2871, n_2872, n_2873, n_2874, n_2875, 
      n_2876, n_2877, n_2878, n_2879, n_2880, n_2881, n_2882, n_2883, n_2884, 
      n_2885, n_2886, n_2887, n_2888, n_2889, n_2890, n_2891, n_2892, n_2893, 
      n_2894, n_2895, n_2896, n_2897, n_2898, n_2899, n_2900, n_2901, n_2902, 
      n_2903, n_2904, n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, 
      n_2912, n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920, 
      n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928, n_2929, 
      n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936, n_2937, n_2938, 
      n_2939, n_2940, n_2941, n_2942, n_2943, n_2944, n_2945, n_2946, n_2947, 
      n_2948, n_2949, n_2950, n_2951, n_2952, n_2953, n_2954, n_2955, n_2956, 
      n_2957, n_2958, n_2959, n_2960, n_2961, n_2962, n_2963, n_2964, n_2965, 
      n_2966, n_2967, n_2968, n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, 
      n_2975, n_2976, n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, 
      n_2984, n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992, 
      n_2993, n_2994, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001, 
      n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009, n_3010, 
      n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017, n_3018, n_3019, 
      n_3020, n_3021, n_3022, n_3023, n_3024, n_3025, n_3026, n_3027, n_3028, 
      n_3029, n_3030, n_3031, n_3032, n_3033, n_3034, n_3035, n_3036, n_3037, 
      n_3038, n_3039, n_3040, n_3041, n_3042, n_3043, n_3044, n_3045, n_3046, 
      n_3047, n_3048, n_3049, n_3050, n_3051, n_3052, n_3053, n_3054, n_3055, 
      n_3056, n_3057, n_3058, n_3059, n_3060, n_3061, n_3062, n_3063, n_3064, 
      n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071, n_3072, n_3073, 
      n_3074, n_3075, n_3076, n_3077, n_3078, n_3079, n_3080, n_3081, n_3082, 
      n_3083, n_3084, n_3085, n_3086, n_3087, n_3088, n_3089, n_3090, n_3091, 
      n_3092, n_3093, n_3094, n_3095, n_3096, n_3097, n_3098, n_3099, n_3100, 
      n_3101, n_3102, n_3103, n_3104, n_3105, n_3106, n_3107, n_3108, n_3109, 
      n_3110, n_3111, n_3112, n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, 
      n_3119, n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127, 
      n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135, n_3136, 
      n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143, n_3144, n_3145, 
      n_3146, n_3147, n_3148, n_3149, n_3150, n_3151, n_3152, n_3153, n_3154, 
      n_3155, n_3156, n_3157, n_3158, n_3159, n_3160, n_3161, n_3162, n_3163, 
      n_3164, n_3165, n_3166, n_3167, n_3168, n_3169, n_3170, n_3171, n_3172, 
      n_3173, n_3174, n_3175, n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, 
      n_3182, n_3183, n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, 
      n_3191, n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199, 
      n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207, n_3208, 
      n_3209, n_3210, n_3211, n_3212, n_3213, n_3214, n_3215, n_3216, n_3217, 
      n_3218, n_3219, n_3220, n_3221, n_3222, n_3223, n_3224, n_3225, n_3226, 
      n_3227, n_3228, n_3229, n_3230, n_3231, n_3232, n_3233, n_3234, n_3235, 
      n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242, n_3243, n_3244, 
      n_3245, n_3246, n_3247, n_3248, n_3249, n_3250, n_3251, n_3252, n_3253, 
      n_3254, n_3255, n_3256, n_3257, n_3258, n_3259, n_3260, n_3261, n_3262, 
      n_3263, n_3264, n_3265, n_3266, n_3267, n_3268, n_3269, n_3270, n_3271, 
      n_3272, n_3273, n_3274, n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, 
      n_3281, n_3282, n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, 
      n_3290, n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298, 
      n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306, n_3307, 
      n_3308, n_3309, n_3310, n_3311, n_3312, n_3313, n_3314, n_3315, n_3316, 
      n_3317, n_3318, n_3319, n_3320, n_3321, n_3322, n_3323, n_3324, n_3325, 
      n_3326, n_3327, n_3328, n_3329, n_3330, n_3331, n_3332, n_3333, n_3334, 
      n_3335, n_3336, n_3337, n_3338, n_3339, n_3340, n_3341, n_3342, n_3343, 
      n_3344, n_3345, n_3346, n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, 
      n_3353, n_3354, n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, 
      n_3362, n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370, 
      n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378, n_3379, 
      n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386, n_3387, n_3388, 
      n_3389, n_3390, n_3391, n_3392, n_3393, n_3394, n_3395, n_3396, n_3397, 
      n_3398, n_3399, n_3400, n_3401, n_3402, n_3403, n_3404, n_3405, n_3406, 
      n_3407, n_3408, n_3409, n_3410, n_3411, n_3412, n_3413, n_3414, n_3415, 
      n_3416, n_3417, n_3418, n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, 
      n_3425, n_3426, n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433, 
      n_3434, n_3435, n_3436, n_3437, n_3438, n_3439, n_3440, n_3441, n_3442, 
      n_3443, n_3444, n_3445, n_3446, n_3447, n_3448, n_3449, n_3450, n_3451, 
      n_3452, n_3453, n_3454, n_3455, n_3456, n_3457, n_3458, n_3459, n_3460, 
      n_3461, n_3462, n_3463, n_3464, n_3465, n_3466, n_3467, n_3468, n_3469, 
      n_3470, n_3471, n_3472, n_3473, n_3474, n_3475, n_3476, n_3477, n_3478, 
      n_3479, n_3480, n_3481, n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, 
      n_3488, n_3489, n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, 
      n_3497, n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505, 
      n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513, n_3514, 
      n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521, n_3522, n_3523, 
      n_3524, n_3525, n_3526, n_3527, n_3528, n_3529, n_3530, n_3531, n_3532, 
      n_3533, n_3534, n_3535, n_3536, n_3537, n_3538, n_3539, n_3540, n_3541, 
      n_3542, n_3543, n_3544, n_3545, n_3546, n_3547, n_3548, n_3549, n_3550, 
      n_3551, n_3552, n_3553, n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, 
      n_3560, n_3561, n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, 
      n_3569, n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577, 
      n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585, n_3586, 
      n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593, n_3594, n_3595, 
      n_3596, n_3597, n_3598, n_3599, n_3600, n_3601, n_3602, n_3603, n_3604, 
      n_3605, n_3606, n_3607, n_3608, n_3609, n_3610, n_3611, n_3612, n_3613, 
      n_3614, n_3615, n_3616, n_3617, n_3618, n_3619, n_3620, n_3621, n_3622, 
      n_3623, n_3624, n_3625, n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, 
      n_3632, n_3633, n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, 
      n_3641, n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649, 
      n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657, n_3658, 
      n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665, n_3666, n_3667, 
      n_3668, n_3669, n_3670, n_3671, n_3672, n_3673, n_3674, n_3675, n_3676, 
      n_3677, n_3678, n_3679, n_3680, n_3681, n_3682, n_3683, n_3684, n_3685, 
      n_3686, n_3687, n_3688, n_3689, n_3690, n_3691, n_3692, n_3693, n_3694, 
      n_3695, n_3696, n_3697, n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, 
      n_3704, n_3705, n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, 
      n_3713, n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721, 
      n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729, n_3730, 
      n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737, n_3738, n_3739, 
      n_3740, n_3741, n_3742, n_3743, n_3744, n_3745, n_3746, n_3747, n_3748, 
      n_3749, n_3750, n_3751, n_3752, n_3753, n_3754, n_3755, n_3756, n_3757, 
      n_3758, n_3759, n_3760, n_3761, n_3762, n_3763, n_3764, n_3765, n_3766, 
      n_3767, n_3768, n_3769, n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, 
      n_3776, n_3777, n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, n_3784, 
      n_3785, n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793, 
      n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801, n_3802, 
      n_3803, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809, n_3810, n_3811, 
      n_3812, n_3813, n_3814, n_3815, n_3816, n_3817, n_3818, n_3819, n_3820, 
      n_3821, n_3822, n_3823, n_3824, n_3825, n_3826, n_3827, n_3828, n_3829, 
      n_3830, n_3831, n_3832, n_3833, n_3834, n_3835, n_3836, n_3837, n_3838, 
      n_3839, n_3840, n_3841, n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, 
      n_3848, n_3849, n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, 
      n_3857, n_3858, n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865, 
      n_3866, n_3867, n_3868, n_3869, n_3870, n_3871, n_3872, n_3873, n_3874, 
      n_3875, n_3876, n_3877, n_3878, n_3879, n_3880, n_3881, n_3882, n_3883, 
      n_3884, n_3885, n_3886, n_3887, n_3888, n_3889, n_3890, n_3891, n_3892, 
      n_3893, n_3894, n_3895, n_3896, n_3897, n_3898, n_3899, n_3900, n_3901, 
      n_3902, n_3903, n_3904, n_3905, n_3906, n_3907, n_3908, n_3909, n_3910, 
      n_3911, n_3912, n_3913, n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, 
      n_3920, n_3921, n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, 
      n_3929, n_3930, n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937, 
      n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945, n_3946, 
      n_3947, n_3948, n_3949, n_3950 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port );
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, DRAM_ADDRESS_1_port, DRAM_ADDRESS_0_port );
   DRAM_DATA_OUT <= ( DRAM_DATA_OUT_31_port, DRAM_DATA_OUT_30_port, 
      DRAM_DATA_OUT_29_port, DRAM_DATA_OUT_28_port, DRAM_DATA_OUT_27_port, 
      DRAM_DATA_OUT_26_port, DRAM_DATA_OUT_25_port, DRAM_DATA_OUT_24_port, 
      DRAM_DATA_OUT_23_port, DRAM_DATA_OUT_22_port, DRAM_DATA_OUT_21_port, 
      DRAM_DATA_OUT_20_port, DRAM_DATA_OUT_19_port, DRAM_DATA_OUT_18_port, 
      DRAM_DATA_OUT_17_port, DRAM_DATA_OUT_16_port, DRAM_DATA_OUT_15_port, 
      DRAM_DATA_OUT_14_port, DRAM_DATA_OUT_13_port, DRAM_DATA_OUT_12_port, 
      DRAM_DATA_OUT_11_port, DRAM_DATA_OUT_10_port, DRAM_DATA_OUT_9_port, 
      DRAM_DATA_OUT_8_port, DRAM_DATA_OUT_7_port, DRAM_DATA_OUT_6_port, 
      DRAM_DATA_OUT_5_port, DRAM_DATA_OUT_4_port, DRAM_DATA_OUT_3_port, 
      DRAM_DATA_OUT_2_port, DRAM_DATA_OUT_1_port, DRAM_DATA_OUT_0_port );
   DATA_SIZE <= ( DATA_SIZE_1_port, DATA_SIZE_0_port );
   DRAMRF_ADDRESS <= ( DRAMRF_ADDRESS_31_port, DRAMRF_ADDRESS_30_port, 
      DRAMRF_ADDRESS_29_port, DRAMRF_ADDRESS_28_port, DRAMRF_ADDRESS_27_port, 
      DRAMRF_ADDRESS_26_port, DRAMRF_ADDRESS_25_port, DRAMRF_ADDRESS_24_port, 
      DRAMRF_ADDRESS_23_port, DRAMRF_ADDRESS_22_port, DRAMRF_ADDRESS_21_port, 
      DRAMRF_ADDRESS_20_port, DRAMRF_ADDRESS_19_port, DRAMRF_ADDRESS_18_port, 
      DRAMRF_ADDRESS_17_port, DRAMRF_ADDRESS_16_port, DRAMRF_ADDRESS_15_port, 
      DRAMRF_ADDRESS_14_port, DRAMRF_ADDRESS_13_port, DRAMRF_ADDRESS_12_port, 
      DRAMRF_ADDRESS_11_port, DRAMRF_ADDRESS_10_port, DRAMRF_ADDRESS_9_port, 
      DRAMRF_ADDRESS_8_port, DRAMRF_ADDRESS_7_port, DRAMRF_ADDRESS_6_port, 
      DRAMRF_ADDRESS_5_port, DRAMRF_ADDRESS_4_port, DRAMRF_ADDRESS_3_port, 
      DRAMRF_ADDRESS_2_port, DRAMRF_ADDRESS_1_port, DRAMRF_ADDRESS_0_port );
   DRAMRF_READNOTWRITE <= DRAMRF_READNOTWRITE_port;
   DATA_SIZE_RF <= ( DataPath_RF_bus_complete_win_data_0_port, 
      DataPath_RF_bus_complete_win_data_0_port );
   
   DECODEhw_HAZARD_CTRL : hazard_table_N_REGS_LOG5 port map( CLK => CLK, RST =>
                           RST, WR1 => DECODEhw_i_WR1, WR2 => i_WF, ADD_WR1(4) 
                           => i_ADD_WS1_4_port, ADD_WR1(3) => i_ADD_WS1_3_port,
                           ADD_WR1(2) => i_ADD_WS1_2_port, ADD_WR1(1) => 
                           i_ADD_WS1_1_port, ADD_WR1(0) => i_ADD_WS1_0_port, 
                           ADD_WR2(4) => i_ADD_WB_4_port, ADD_WR2(3) => 
                           i_ADD_WB_3_port, ADD_WR2(2) => i_ADD_WB_2_port, 
                           ADD_WR2(1) => i_ADD_WB_1_port, ADD_WR2(0) => 
                           i_ADD_WB_0_port, ADD_CHECK1(4) => n10858, 
                           ADD_CHECK1(3) => n10859, ADD_CHECK1(2) => n10860, 
                           ADD_CHECK1(1) => n10861, ADD_CHECK1(0) => n10862, 
                           ADD_CHECK2(4) => n10863, ADD_CHECK2(3) => n10864, 
                           ADD_CHECK2(2) => n10865, ADD_CHECK2(1) => n10866, 
                           ADD_CHECK2(0) => n10867, BUSY => i_HAZARD_SIG_CU, 
                           BUSY_WINDOW => i_BUSY_WINDOW);
   DataPath_RF_SELBLOCK_INLOC : in_loc_selblock_NBIT_DATA32_N8_F5 port map( 
                           regs(2559) => DataPath_RF_bus_reg_dataout_2559_port,
                           regs(2558) => DataPath_RF_bus_reg_dataout_2558_port,
                           regs(2557) => DataPath_RF_bus_reg_dataout_2557_port,
                           regs(2556) => DataPath_RF_bus_reg_dataout_2556_port,
                           regs(2555) => DataPath_RF_bus_reg_dataout_2555_port,
                           regs(2554) => DataPath_RF_bus_reg_dataout_2554_port,
                           regs(2553) => DataPath_RF_bus_reg_dataout_2553_port,
                           regs(2552) => DataPath_RF_bus_reg_dataout_2552_port,
                           regs(2551) => DataPath_RF_bus_reg_dataout_2551_port,
                           regs(2550) => DataPath_RF_bus_reg_dataout_2550_port,
                           regs(2549) => DataPath_RF_bus_reg_dataout_2549_port,
                           regs(2548) => DataPath_RF_bus_reg_dataout_2548_port,
                           regs(2547) => DataPath_RF_bus_reg_dataout_2547_port,
                           regs(2546) => DataPath_RF_bus_reg_dataout_2546_port,
                           regs(2545) => DataPath_RF_bus_reg_dataout_2545_port,
                           regs(2544) => DataPath_RF_bus_reg_dataout_2544_port,
                           regs(2543) => DataPath_RF_bus_reg_dataout_2543_port,
                           regs(2542) => DataPath_RF_bus_reg_dataout_2542_port,
                           regs(2541) => DataPath_RF_bus_reg_dataout_2541_port,
                           regs(2540) => DataPath_RF_bus_reg_dataout_2540_port,
                           regs(2539) => DataPath_RF_bus_reg_dataout_2539_port,
                           regs(2538) => DataPath_RF_bus_reg_dataout_2538_port,
                           regs(2537) => DataPath_RF_bus_reg_dataout_2537_port,
                           regs(2536) => DataPath_RF_bus_reg_dataout_2536_port,
                           regs(2535) => DataPath_RF_bus_reg_dataout_2535_port,
                           regs(2534) => DataPath_RF_bus_reg_dataout_2534_port,
                           regs(2533) => DataPath_RF_bus_reg_dataout_2533_port,
                           regs(2532) => DataPath_RF_bus_reg_dataout_2532_port,
                           regs(2531) => DataPath_RF_bus_reg_dataout_2531_port,
                           regs(2530) => DataPath_RF_bus_reg_dataout_2530_port,
                           regs(2529) => DataPath_RF_bus_reg_dataout_2529_port,
                           regs(2528) => DataPath_RF_bus_reg_dataout_2528_port,
                           regs(2527) => DataPath_RF_bus_reg_dataout_2527_port,
                           regs(2526) => DataPath_RF_bus_reg_dataout_2526_port,
                           regs(2525) => DataPath_RF_bus_reg_dataout_2525_port,
                           regs(2524) => DataPath_RF_bus_reg_dataout_2524_port,
                           regs(2523) => DataPath_RF_bus_reg_dataout_2523_port,
                           regs(2522) => DataPath_RF_bus_reg_dataout_2522_port,
                           regs(2521) => DataPath_RF_bus_reg_dataout_2521_port,
                           regs(2520) => DataPath_RF_bus_reg_dataout_2520_port,
                           regs(2519) => DataPath_RF_bus_reg_dataout_2519_port,
                           regs(2518) => DataPath_RF_bus_reg_dataout_2518_port,
                           regs(2517) => DataPath_RF_bus_reg_dataout_2517_port,
                           regs(2516) => DataPath_RF_bus_reg_dataout_2516_port,
                           regs(2515) => DataPath_RF_bus_reg_dataout_2515_port,
                           regs(2514) => DataPath_RF_bus_reg_dataout_2514_port,
                           regs(2513) => DataPath_RF_bus_reg_dataout_2513_port,
                           regs(2512) => DataPath_RF_bus_reg_dataout_2512_port,
                           regs(2511) => DataPath_RF_bus_reg_dataout_2511_port,
                           regs(2510) => DataPath_RF_bus_reg_dataout_2510_port,
                           regs(2509) => DataPath_RF_bus_reg_dataout_2509_port,
                           regs(2508) => DataPath_RF_bus_reg_dataout_2508_port,
                           regs(2507) => DataPath_RF_bus_reg_dataout_2507_port,
                           regs(2506) => DataPath_RF_bus_reg_dataout_2506_port,
                           regs(2505) => DataPath_RF_bus_reg_dataout_2505_port,
                           regs(2504) => DataPath_RF_bus_reg_dataout_2504_port,
                           regs(2503) => DataPath_RF_bus_reg_dataout_2503_port,
                           regs(2502) => DataPath_RF_bus_reg_dataout_2502_port,
                           regs(2501) => DataPath_RF_bus_reg_dataout_2501_port,
                           regs(2500) => DataPath_RF_bus_reg_dataout_2500_port,
                           regs(2499) => DataPath_RF_bus_reg_dataout_2499_port,
                           regs(2498) => DataPath_RF_bus_reg_dataout_2498_port,
                           regs(2497) => DataPath_RF_bus_reg_dataout_2497_port,
                           regs(2496) => DataPath_RF_bus_reg_dataout_2496_port,
                           regs(2495) => DataPath_RF_bus_reg_dataout_2495_port,
                           regs(2494) => DataPath_RF_bus_reg_dataout_2494_port,
                           regs(2493) => DataPath_RF_bus_reg_dataout_2493_port,
                           regs(2492) => DataPath_RF_bus_reg_dataout_2492_port,
                           regs(2491) => DataPath_RF_bus_reg_dataout_2491_port,
                           regs(2490) => DataPath_RF_bus_reg_dataout_2490_port,
                           regs(2489) => DataPath_RF_bus_reg_dataout_2489_port,
                           regs(2488) => DataPath_RF_bus_reg_dataout_2488_port,
                           regs(2487) => DataPath_RF_bus_reg_dataout_2487_port,
                           regs(2486) => DataPath_RF_bus_reg_dataout_2486_port,
                           regs(2485) => DataPath_RF_bus_reg_dataout_2485_port,
                           regs(2484) => DataPath_RF_bus_reg_dataout_2484_port,
                           regs(2483) => DataPath_RF_bus_reg_dataout_2483_port,
                           regs(2482) => DataPath_RF_bus_reg_dataout_2482_port,
                           regs(2481) => DataPath_RF_bus_reg_dataout_2481_port,
                           regs(2480) => DataPath_RF_bus_reg_dataout_2480_port,
                           regs(2479) => DataPath_RF_bus_reg_dataout_2479_port,
                           regs(2478) => DataPath_RF_bus_reg_dataout_2478_port,
                           regs(2477) => DataPath_RF_bus_reg_dataout_2477_port,
                           regs(2476) => DataPath_RF_bus_reg_dataout_2476_port,
                           regs(2475) => DataPath_RF_bus_reg_dataout_2475_port,
                           regs(2474) => DataPath_RF_bus_reg_dataout_2474_port,
                           regs(2473) => DataPath_RF_bus_reg_dataout_2473_port,
                           regs(2472) => DataPath_RF_bus_reg_dataout_2472_port,
                           regs(2471) => DataPath_RF_bus_reg_dataout_2471_port,
                           regs(2470) => DataPath_RF_bus_reg_dataout_2470_port,
                           regs(2469) => DataPath_RF_bus_reg_dataout_2469_port,
                           regs(2468) => DataPath_RF_bus_reg_dataout_2468_port,
                           regs(2467) => DataPath_RF_bus_reg_dataout_2467_port,
                           regs(2466) => DataPath_RF_bus_reg_dataout_2466_port,
                           regs(2465) => DataPath_RF_bus_reg_dataout_2465_port,
                           regs(2464) => DataPath_RF_bus_reg_dataout_2464_port,
                           regs(2463) => DataPath_RF_bus_reg_dataout_2463_port,
                           regs(2462) => DataPath_RF_bus_reg_dataout_2462_port,
                           regs(2461) => DataPath_RF_bus_reg_dataout_2461_port,
                           regs(2460) => DataPath_RF_bus_reg_dataout_2460_port,
                           regs(2459) => DataPath_RF_bus_reg_dataout_2459_port,
                           regs(2458) => DataPath_RF_bus_reg_dataout_2458_port,
                           regs(2457) => DataPath_RF_bus_reg_dataout_2457_port,
                           regs(2456) => DataPath_RF_bus_reg_dataout_2456_port,
                           regs(2455) => DataPath_RF_bus_reg_dataout_2455_port,
                           regs(2454) => DataPath_RF_bus_reg_dataout_2454_port,
                           regs(2453) => DataPath_RF_bus_reg_dataout_2453_port,
                           regs(2452) => DataPath_RF_bus_reg_dataout_2452_port,
                           regs(2451) => DataPath_RF_bus_reg_dataout_2451_port,
                           regs(2450) => DataPath_RF_bus_reg_dataout_2450_port,
                           regs(2449) => DataPath_RF_bus_reg_dataout_2449_port,
                           regs(2448) => DataPath_RF_bus_reg_dataout_2448_port,
                           regs(2447) => DataPath_RF_bus_reg_dataout_2447_port,
                           regs(2446) => DataPath_RF_bus_reg_dataout_2446_port,
                           regs(2445) => DataPath_RF_bus_reg_dataout_2445_port,
                           regs(2444) => DataPath_RF_bus_reg_dataout_2444_port,
                           regs(2443) => DataPath_RF_bus_reg_dataout_2443_port,
                           regs(2442) => DataPath_RF_bus_reg_dataout_2442_port,
                           regs(2441) => DataPath_RF_bus_reg_dataout_2441_port,
                           regs(2440) => DataPath_RF_bus_reg_dataout_2440_port,
                           regs(2439) => DataPath_RF_bus_reg_dataout_2439_port,
                           regs(2438) => DataPath_RF_bus_reg_dataout_2438_port,
                           regs(2437) => DataPath_RF_bus_reg_dataout_2437_port,
                           regs(2436) => DataPath_RF_bus_reg_dataout_2436_port,
                           regs(2435) => DataPath_RF_bus_reg_dataout_2435_port,
                           regs(2434) => DataPath_RF_bus_reg_dataout_2434_port,
                           regs(2433) => DataPath_RF_bus_reg_dataout_2433_port,
                           regs(2432) => DataPath_RF_bus_reg_dataout_2432_port,
                           regs(2431) => DataPath_RF_bus_reg_dataout_2431_port,
                           regs(2430) => DataPath_RF_bus_reg_dataout_2430_port,
                           regs(2429) => DataPath_RF_bus_reg_dataout_2429_port,
                           regs(2428) => DataPath_RF_bus_reg_dataout_2428_port,
                           regs(2427) => DataPath_RF_bus_reg_dataout_2427_port,
                           regs(2426) => DataPath_RF_bus_reg_dataout_2426_port,
                           regs(2425) => DataPath_RF_bus_reg_dataout_2425_port,
                           regs(2424) => DataPath_RF_bus_reg_dataout_2424_port,
                           regs(2423) => DataPath_RF_bus_reg_dataout_2423_port,
                           regs(2422) => DataPath_RF_bus_reg_dataout_2422_port,
                           regs(2421) => DataPath_RF_bus_reg_dataout_2421_port,
                           regs(2420) => DataPath_RF_bus_reg_dataout_2420_port,
                           regs(2419) => DataPath_RF_bus_reg_dataout_2419_port,
                           regs(2418) => DataPath_RF_bus_reg_dataout_2418_port,
                           regs(2417) => DataPath_RF_bus_reg_dataout_2417_port,
                           regs(2416) => DataPath_RF_bus_reg_dataout_2416_port,
                           regs(2415) => DataPath_RF_bus_reg_dataout_2415_port,
                           regs(2414) => DataPath_RF_bus_reg_dataout_2414_port,
                           regs(2413) => DataPath_RF_bus_reg_dataout_2413_port,
                           regs(2412) => DataPath_RF_bus_reg_dataout_2412_port,
                           regs(2411) => DataPath_RF_bus_reg_dataout_2411_port,
                           regs(2410) => DataPath_RF_bus_reg_dataout_2410_port,
                           regs(2409) => DataPath_RF_bus_reg_dataout_2409_port,
                           regs(2408) => DataPath_RF_bus_reg_dataout_2408_port,
                           regs(2407) => DataPath_RF_bus_reg_dataout_2407_port,
                           regs(2406) => DataPath_RF_bus_reg_dataout_2406_port,
                           regs(2405) => DataPath_RF_bus_reg_dataout_2405_port,
                           regs(2404) => DataPath_RF_bus_reg_dataout_2404_port,
                           regs(2403) => DataPath_RF_bus_reg_dataout_2403_port,
                           regs(2402) => DataPath_RF_bus_reg_dataout_2402_port,
                           regs(2401) => DataPath_RF_bus_reg_dataout_2401_port,
                           regs(2400) => DataPath_RF_bus_reg_dataout_2400_port,
                           regs(2399) => DataPath_RF_bus_reg_dataout_2399_port,
                           regs(2398) => DataPath_RF_bus_reg_dataout_2398_port,
                           regs(2397) => DataPath_RF_bus_reg_dataout_2397_port,
                           regs(2396) => DataPath_RF_bus_reg_dataout_2396_port,
                           regs(2395) => DataPath_RF_bus_reg_dataout_2395_port,
                           regs(2394) => DataPath_RF_bus_reg_dataout_2394_port,
                           regs(2393) => DataPath_RF_bus_reg_dataout_2393_port,
                           regs(2392) => DataPath_RF_bus_reg_dataout_2392_port,
                           regs(2391) => DataPath_RF_bus_reg_dataout_2391_port,
                           regs(2390) => DataPath_RF_bus_reg_dataout_2390_port,
                           regs(2389) => DataPath_RF_bus_reg_dataout_2389_port,
                           regs(2388) => DataPath_RF_bus_reg_dataout_2388_port,
                           regs(2387) => DataPath_RF_bus_reg_dataout_2387_port,
                           regs(2386) => DataPath_RF_bus_reg_dataout_2386_port,
                           regs(2385) => DataPath_RF_bus_reg_dataout_2385_port,
                           regs(2384) => DataPath_RF_bus_reg_dataout_2384_port,
                           regs(2383) => DataPath_RF_bus_reg_dataout_2383_port,
                           regs(2382) => DataPath_RF_bus_reg_dataout_2382_port,
                           regs(2381) => DataPath_RF_bus_reg_dataout_2381_port,
                           regs(2380) => DataPath_RF_bus_reg_dataout_2380_port,
                           regs(2379) => DataPath_RF_bus_reg_dataout_2379_port,
                           regs(2378) => DataPath_RF_bus_reg_dataout_2378_port,
                           regs(2377) => DataPath_RF_bus_reg_dataout_2377_port,
                           regs(2376) => DataPath_RF_bus_reg_dataout_2376_port,
                           regs(2375) => DataPath_RF_bus_reg_dataout_2375_port,
                           regs(2374) => DataPath_RF_bus_reg_dataout_2374_port,
                           regs(2373) => DataPath_RF_bus_reg_dataout_2373_port,
                           regs(2372) => DataPath_RF_bus_reg_dataout_2372_port,
                           regs(2371) => DataPath_RF_bus_reg_dataout_2371_port,
                           regs(2370) => DataPath_RF_bus_reg_dataout_2370_port,
                           regs(2369) => DataPath_RF_bus_reg_dataout_2369_port,
                           regs(2368) => DataPath_RF_bus_reg_dataout_2368_port,
                           regs(2367) => DataPath_RF_bus_reg_dataout_2367_port,
                           regs(2366) => DataPath_RF_bus_reg_dataout_2366_port,
                           regs(2365) => DataPath_RF_bus_reg_dataout_2365_port,
                           regs(2364) => DataPath_RF_bus_reg_dataout_2364_port,
                           regs(2363) => DataPath_RF_bus_reg_dataout_2363_port,
                           regs(2362) => DataPath_RF_bus_reg_dataout_2362_port,
                           regs(2361) => DataPath_RF_bus_reg_dataout_2361_port,
                           regs(2360) => DataPath_RF_bus_reg_dataout_2360_port,
                           regs(2359) => DataPath_RF_bus_reg_dataout_2359_port,
                           regs(2358) => DataPath_RF_bus_reg_dataout_2358_port,
                           regs(2357) => DataPath_RF_bus_reg_dataout_2357_port,
                           regs(2356) => DataPath_RF_bus_reg_dataout_2356_port,
                           regs(2355) => DataPath_RF_bus_reg_dataout_2355_port,
                           regs(2354) => DataPath_RF_bus_reg_dataout_2354_port,
                           regs(2353) => DataPath_RF_bus_reg_dataout_2353_port,
                           regs(2352) => DataPath_RF_bus_reg_dataout_2352_port,
                           regs(2351) => DataPath_RF_bus_reg_dataout_2351_port,
                           regs(2350) => DataPath_RF_bus_reg_dataout_2350_port,
                           regs(2349) => DataPath_RF_bus_reg_dataout_2349_port,
                           regs(2348) => DataPath_RF_bus_reg_dataout_2348_port,
                           regs(2347) => DataPath_RF_bus_reg_dataout_2347_port,
                           regs(2346) => DataPath_RF_bus_reg_dataout_2346_port,
                           regs(2345) => DataPath_RF_bus_reg_dataout_2345_port,
                           regs(2344) => DataPath_RF_bus_reg_dataout_2344_port,
                           regs(2343) => DataPath_RF_bus_reg_dataout_2343_port,
                           regs(2342) => DataPath_RF_bus_reg_dataout_2342_port,
                           regs(2341) => DataPath_RF_bus_reg_dataout_2341_port,
                           regs(2340) => DataPath_RF_bus_reg_dataout_2340_port,
                           regs(2339) => DataPath_RF_bus_reg_dataout_2339_port,
                           regs(2338) => DataPath_RF_bus_reg_dataout_2338_port,
                           regs(2337) => DataPath_RF_bus_reg_dataout_2337_port,
                           regs(2336) => DataPath_RF_bus_reg_dataout_2336_port,
                           regs(2335) => DataPath_RF_bus_reg_dataout_2335_port,
                           regs(2334) => DataPath_RF_bus_reg_dataout_2334_port,
                           regs(2333) => DataPath_RF_bus_reg_dataout_2333_port,
                           regs(2332) => DataPath_RF_bus_reg_dataout_2332_port,
                           regs(2331) => DataPath_RF_bus_reg_dataout_2331_port,
                           regs(2330) => DataPath_RF_bus_reg_dataout_2330_port,
                           regs(2329) => DataPath_RF_bus_reg_dataout_2329_port,
                           regs(2328) => DataPath_RF_bus_reg_dataout_2328_port,
                           regs(2327) => DataPath_RF_bus_reg_dataout_2327_port,
                           regs(2326) => DataPath_RF_bus_reg_dataout_2326_port,
                           regs(2325) => DataPath_RF_bus_reg_dataout_2325_port,
                           regs(2324) => DataPath_RF_bus_reg_dataout_2324_port,
                           regs(2323) => DataPath_RF_bus_reg_dataout_2323_port,
                           regs(2322) => DataPath_RF_bus_reg_dataout_2322_port,
                           regs(2321) => DataPath_RF_bus_reg_dataout_2321_port,
                           regs(2320) => DataPath_RF_bus_reg_dataout_2320_port,
                           regs(2319) => DataPath_RF_bus_reg_dataout_2319_port,
                           regs(2318) => DataPath_RF_bus_reg_dataout_2318_port,
                           regs(2317) => DataPath_RF_bus_reg_dataout_2317_port,
                           regs(2316) => DataPath_RF_bus_reg_dataout_2316_port,
                           regs(2315) => DataPath_RF_bus_reg_dataout_2315_port,
                           regs(2314) => DataPath_RF_bus_reg_dataout_2314_port,
                           regs(2313) => DataPath_RF_bus_reg_dataout_2313_port,
                           regs(2312) => DataPath_RF_bus_reg_dataout_2312_port,
                           regs(2311) => DataPath_RF_bus_reg_dataout_2311_port,
                           regs(2310) => DataPath_RF_bus_reg_dataout_2310_port,
                           regs(2309) => DataPath_RF_bus_reg_dataout_2309_port,
                           regs(2308) => DataPath_RF_bus_reg_dataout_2308_port,
                           regs(2307) => DataPath_RF_bus_reg_dataout_2307_port,
                           regs(2306) => DataPath_RF_bus_reg_dataout_2306_port,
                           regs(2305) => DataPath_RF_bus_reg_dataout_2305_port,
                           regs(2304) => DataPath_RF_bus_reg_dataout_2304_port,
                           regs(2303) => DataPath_RF_bus_reg_dataout_2303_port,
                           regs(2302) => DataPath_RF_bus_reg_dataout_2302_port,
                           regs(2301) => DataPath_RF_bus_reg_dataout_2301_port,
                           regs(2300) => DataPath_RF_bus_reg_dataout_2300_port,
                           regs(2299) => DataPath_RF_bus_reg_dataout_2299_port,
                           regs(2298) => DataPath_RF_bus_reg_dataout_2298_port,
                           regs(2297) => DataPath_RF_bus_reg_dataout_2297_port,
                           regs(2296) => DataPath_RF_bus_reg_dataout_2296_port,
                           regs(2295) => DataPath_RF_bus_reg_dataout_2295_port,
                           regs(2294) => DataPath_RF_bus_reg_dataout_2294_port,
                           regs(2293) => DataPath_RF_bus_reg_dataout_2293_port,
                           regs(2292) => DataPath_RF_bus_reg_dataout_2292_port,
                           regs(2291) => DataPath_RF_bus_reg_dataout_2291_port,
                           regs(2290) => DataPath_RF_bus_reg_dataout_2290_port,
                           regs(2289) => DataPath_RF_bus_reg_dataout_2289_port,
                           regs(2288) => DataPath_RF_bus_reg_dataout_2288_port,
                           regs(2287) => DataPath_RF_bus_reg_dataout_2287_port,
                           regs(2286) => DataPath_RF_bus_reg_dataout_2286_port,
                           regs(2285) => DataPath_RF_bus_reg_dataout_2285_port,
                           regs(2284) => DataPath_RF_bus_reg_dataout_2284_port,
                           regs(2283) => DataPath_RF_bus_reg_dataout_2283_port,
                           regs(2282) => DataPath_RF_bus_reg_dataout_2282_port,
                           regs(2281) => DataPath_RF_bus_reg_dataout_2281_port,
                           regs(2280) => DataPath_RF_bus_reg_dataout_2280_port,
                           regs(2279) => DataPath_RF_bus_reg_dataout_2279_port,
                           regs(2278) => DataPath_RF_bus_reg_dataout_2278_port,
                           regs(2277) => DataPath_RF_bus_reg_dataout_2277_port,
                           regs(2276) => DataPath_RF_bus_reg_dataout_2276_port,
                           regs(2275) => DataPath_RF_bus_reg_dataout_2275_port,
                           regs(2274) => DataPath_RF_bus_reg_dataout_2274_port,
                           regs(2273) => DataPath_RF_bus_reg_dataout_2273_port,
                           regs(2272) => DataPath_RF_bus_reg_dataout_2272_port,
                           regs(2271) => DataPath_RF_bus_reg_dataout_2271_port,
                           regs(2270) => DataPath_RF_bus_reg_dataout_2270_port,
                           regs(2269) => DataPath_RF_bus_reg_dataout_2269_port,
                           regs(2268) => DataPath_RF_bus_reg_dataout_2268_port,
                           regs(2267) => DataPath_RF_bus_reg_dataout_2267_port,
                           regs(2266) => DataPath_RF_bus_reg_dataout_2266_port,
                           regs(2265) => DataPath_RF_bus_reg_dataout_2265_port,
                           regs(2264) => DataPath_RF_bus_reg_dataout_2264_port,
                           regs(2263) => DataPath_RF_bus_reg_dataout_2263_port,
                           regs(2262) => DataPath_RF_bus_reg_dataout_2262_port,
                           regs(2261) => DataPath_RF_bus_reg_dataout_2261_port,
                           regs(2260) => DataPath_RF_bus_reg_dataout_2260_port,
                           regs(2259) => DataPath_RF_bus_reg_dataout_2259_port,
                           regs(2258) => DataPath_RF_bus_reg_dataout_2258_port,
                           regs(2257) => DataPath_RF_bus_reg_dataout_2257_port,
                           regs(2256) => DataPath_RF_bus_reg_dataout_2256_port,
                           regs(2255) => DataPath_RF_bus_reg_dataout_2255_port,
                           regs(2254) => DataPath_RF_bus_reg_dataout_2254_port,
                           regs(2253) => DataPath_RF_bus_reg_dataout_2253_port,
                           regs(2252) => DataPath_RF_bus_reg_dataout_2252_port,
                           regs(2251) => DataPath_RF_bus_reg_dataout_2251_port,
                           regs(2250) => DataPath_RF_bus_reg_dataout_2250_port,
                           regs(2249) => DataPath_RF_bus_reg_dataout_2249_port,
                           regs(2248) => DataPath_RF_bus_reg_dataout_2248_port,
                           regs(2247) => DataPath_RF_bus_reg_dataout_2247_port,
                           regs(2246) => DataPath_RF_bus_reg_dataout_2246_port,
                           regs(2245) => DataPath_RF_bus_reg_dataout_2245_port,
                           regs(2244) => DataPath_RF_bus_reg_dataout_2244_port,
                           regs(2243) => DataPath_RF_bus_reg_dataout_2243_port,
                           regs(2242) => DataPath_RF_bus_reg_dataout_2242_port,
                           regs(2241) => DataPath_RF_bus_reg_dataout_2241_port,
                           regs(2240) => DataPath_RF_bus_reg_dataout_2240_port,
                           regs(2239) => DataPath_RF_bus_reg_dataout_2239_port,
                           regs(2238) => DataPath_RF_bus_reg_dataout_2238_port,
                           regs(2237) => DataPath_RF_bus_reg_dataout_2237_port,
                           regs(2236) => DataPath_RF_bus_reg_dataout_2236_port,
                           regs(2235) => DataPath_RF_bus_reg_dataout_2235_port,
                           regs(2234) => DataPath_RF_bus_reg_dataout_2234_port,
                           regs(2233) => DataPath_RF_bus_reg_dataout_2233_port,
                           regs(2232) => DataPath_RF_bus_reg_dataout_2232_port,
                           regs(2231) => DataPath_RF_bus_reg_dataout_2231_port,
                           regs(2230) => DataPath_RF_bus_reg_dataout_2230_port,
                           regs(2229) => DataPath_RF_bus_reg_dataout_2229_port,
                           regs(2228) => DataPath_RF_bus_reg_dataout_2228_port,
                           regs(2227) => DataPath_RF_bus_reg_dataout_2227_port,
                           regs(2226) => DataPath_RF_bus_reg_dataout_2226_port,
                           regs(2225) => DataPath_RF_bus_reg_dataout_2225_port,
                           regs(2224) => DataPath_RF_bus_reg_dataout_2224_port,
                           regs(2223) => DataPath_RF_bus_reg_dataout_2223_port,
                           regs(2222) => DataPath_RF_bus_reg_dataout_2222_port,
                           regs(2221) => DataPath_RF_bus_reg_dataout_2221_port,
                           regs(2220) => DataPath_RF_bus_reg_dataout_2220_port,
                           regs(2219) => DataPath_RF_bus_reg_dataout_2219_port,
                           regs(2218) => DataPath_RF_bus_reg_dataout_2218_port,
                           regs(2217) => DataPath_RF_bus_reg_dataout_2217_port,
                           regs(2216) => DataPath_RF_bus_reg_dataout_2216_port,
                           regs(2215) => DataPath_RF_bus_reg_dataout_2215_port,
                           regs(2214) => DataPath_RF_bus_reg_dataout_2214_port,
                           regs(2213) => DataPath_RF_bus_reg_dataout_2213_port,
                           regs(2212) => DataPath_RF_bus_reg_dataout_2212_port,
                           regs(2211) => DataPath_RF_bus_reg_dataout_2211_port,
                           regs(2210) => DataPath_RF_bus_reg_dataout_2210_port,
                           regs(2209) => DataPath_RF_bus_reg_dataout_2209_port,
                           regs(2208) => DataPath_RF_bus_reg_dataout_2208_port,
                           regs(2207) => DataPath_RF_bus_reg_dataout_2207_port,
                           regs(2206) => DataPath_RF_bus_reg_dataout_2206_port,
                           regs(2205) => DataPath_RF_bus_reg_dataout_2205_port,
                           regs(2204) => DataPath_RF_bus_reg_dataout_2204_port,
                           regs(2203) => DataPath_RF_bus_reg_dataout_2203_port,
                           regs(2202) => DataPath_RF_bus_reg_dataout_2202_port,
                           regs(2201) => DataPath_RF_bus_reg_dataout_2201_port,
                           regs(2200) => DataPath_RF_bus_reg_dataout_2200_port,
                           regs(2199) => DataPath_RF_bus_reg_dataout_2199_port,
                           regs(2198) => DataPath_RF_bus_reg_dataout_2198_port,
                           regs(2197) => DataPath_RF_bus_reg_dataout_2197_port,
                           regs(2196) => DataPath_RF_bus_reg_dataout_2196_port,
                           regs(2195) => DataPath_RF_bus_reg_dataout_2195_port,
                           regs(2194) => DataPath_RF_bus_reg_dataout_2194_port,
                           regs(2193) => DataPath_RF_bus_reg_dataout_2193_port,
                           regs(2192) => DataPath_RF_bus_reg_dataout_2192_port,
                           regs(2191) => DataPath_RF_bus_reg_dataout_2191_port,
                           regs(2190) => DataPath_RF_bus_reg_dataout_2190_port,
                           regs(2189) => DataPath_RF_bus_reg_dataout_2189_port,
                           regs(2188) => DataPath_RF_bus_reg_dataout_2188_port,
                           regs(2187) => DataPath_RF_bus_reg_dataout_2187_port,
                           regs(2186) => DataPath_RF_bus_reg_dataout_2186_port,
                           regs(2185) => DataPath_RF_bus_reg_dataout_2185_port,
                           regs(2184) => DataPath_RF_bus_reg_dataout_2184_port,
                           regs(2183) => DataPath_RF_bus_reg_dataout_2183_port,
                           regs(2182) => DataPath_RF_bus_reg_dataout_2182_port,
                           regs(2181) => DataPath_RF_bus_reg_dataout_2181_port,
                           regs(2180) => DataPath_RF_bus_reg_dataout_2180_port,
                           regs(2179) => DataPath_RF_bus_reg_dataout_2179_port,
                           regs(2178) => DataPath_RF_bus_reg_dataout_2178_port,
                           regs(2177) => DataPath_RF_bus_reg_dataout_2177_port,
                           regs(2176) => DataPath_RF_bus_reg_dataout_2176_port,
                           regs(2175) => DataPath_RF_bus_reg_dataout_2175_port,
                           regs(2174) => DataPath_RF_bus_reg_dataout_2174_port,
                           regs(2173) => DataPath_RF_bus_reg_dataout_2173_port,
                           regs(2172) => DataPath_RF_bus_reg_dataout_2172_port,
                           regs(2171) => DataPath_RF_bus_reg_dataout_2171_port,
                           regs(2170) => DataPath_RF_bus_reg_dataout_2170_port,
                           regs(2169) => DataPath_RF_bus_reg_dataout_2169_port,
                           regs(2168) => DataPath_RF_bus_reg_dataout_2168_port,
                           regs(2167) => DataPath_RF_bus_reg_dataout_2167_port,
                           regs(2166) => DataPath_RF_bus_reg_dataout_2166_port,
                           regs(2165) => DataPath_RF_bus_reg_dataout_2165_port,
                           regs(2164) => DataPath_RF_bus_reg_dataout_2164_port,
                           regs(2163) => DataPath_RF_bus_reg_dataout_2163_port,
                           regs(2162) => DataPath_RF_bus_reg_dataout_2162_port,
                           regs(2161) => DataPath_RF_bus_reg_dataout_2161_port,
                           regs(2160) => DataPath_RF_bus_reg_dataout_2160_port,
                           regs(2159) => DataPath_RF_bus_reg_dataout_2159_port,
                           regs(2158) => DataPath_RF_bus_reg_dataout_2158_port,
                           regs(2157) => DataPath_RF_bus_reg_dataout_2157_port,
                           regs(2156) => DataPath_RF_bus_reg_dataout_2156_port,
                           regs(2155) => DataPath_RF_bus_reg_dataout_2155_port,
                           regs(2154) => DataPath_RF_bus_reg_dataout_2154_port,
                           regs(2153) => DataPath_RF_bus_reg_dataout_2153_port,
                           regs(2152) => DataPath_RF_bus_reg_dataout_2152_port,
                           regs(2151) => DataPath_RF_bus_reg_dataout_2151_port,
                           regs(2150) => DataPath_RF_bus_reg_dataout_2150_port,
                           regs(2149) => DataPath_RF_bus_reg_dataout_2149_port,
                           regs(2148) => DataPath_RF_bus_reg_dataout_2148_port,
                           regs(2147) => DataPath_RF_bus_reg_dataout_2147_port,
                           regs(2146) => DataPath_RF_bus_reg_dataout_2146_port,
                           regs(2145) => DataPath_RF_bus_reg_dataout_2145_port,
                           regs(2144) => DataPath_RF_bus_reg_dataout_2144_port,
                           regs(2143) => DataPath_RF_bus_reg_dataout_2143_port,
                           regs(2142) => DataPath_RF_bus_reg_dataout_2142_port,
                           regs(2141) => DataPath_RF_bus_reg_dataout_2141_port,
                           regs(2140) => DataPath_RF_bus_reg_dataout_2140_port,
                           regs(2139) => DataPath_RF_bus_reg_dataout_2139_port,
                           regs(2138) => DataPath_RF_bus_reg_dataout_2138_port,
                           regs(2137) => DataPath_RF_bus_reg_dataout_2137_port,
                           regs(2136) => DataPath_RF_bus_reg_dataout_2136_port,
                           regs(2135) => DataPath_RF_bus_reg_dataout_2135_port,
                           regs(2134) => DataPath_RF_bus_reg_dataout_2134_port,
                           regs(2133) => DataPath_RF_bus_reg_dataout_2133_port,
                           regs(2132) => DataPath_RF_bus_reg_dataout_2132_port,
                           regs(2131) => DataPath_RF_bus_reg_dataout_2131_port,
                           regs(2130) => DataPath_RF_bus_reg_dataout_2130_port,
                           regs(2129) => DataPath_RF_bus_reg_dataout_2129_port,
                           regs(2128) => DataPath_RF_bus_reg_dataout_2128_port,
                           regs(2127) => DataPath_RF_bus_reg_dataout_2127_port,
                           regs(2126) => DataPath_RF_bus_reg_dataout_2126_port,
                           regs(2125) => DataPath_RF_bus_reg_dataout_2125_port,
                           regs(2124) => DataPath_RF_bus_reg_dataout_2124_port,
                           regs(2123) => DataPath_RF_bus_reg_dataout_2123_port,
                           regs(2122) => DataPath_RF_bus_reg_dataout_2122_port,
                           regs(2121) => DataPath_RF_bus_reg_dataout_2121_port,
                           regs(2120) => DataPath_RF_bus_reg_dataout_2120_port,
                           regs(2119) => DataPath_RF_bus_reg_dataout_2119_port,
                           regs(2118) => DataPath_RF_bus_reg_dataout_2118_port,
                           regs(2117) => DataPath_RF_bus_reg_dataout_2117_port,
                           regs(2116) => DataPath_RF_bus_reg_dataout_2116_port,
                           regs(2115) => DataPath_RF_bus_reg_dataout_2115_port,
                           regs(2114) => DataPath_RF_bus_reg_dataout_2114_port,
                           regs(2113) => DataPath_RF_bus_reg_dataout_2113_port,
                           regs(2112) => DataPath_RF_bus_reg_dataout_2112_port,
                           regs(2111) => DataPath_RF_bus_reg_dataout_2111_port,
                           regs(2110) => DataPath_RF_bus_reg_dataout_2110_port,
                           regs(2109) => DataPath_RF_bus_reg_dataout_2109_port,
                           regs(2108) => DataPath_RF_bus_reg_dataout_2108_port,
                           regs(2107) => DataPath_RF_bus_reg_dataout_2107_port,
                           regs(2106) => DataPath_RF_bus_reg_dataout_2106_port,
                           regs(2105) => DataPath_RF_bus_reg_dataout_2105_port,
                           regs(2104) => DataPath_RF_bus_reg_dataout_2104_port,
                           regs(2103) => DataPath_RF_bus_reg_dataout_2103_port,
                           regs(2102) => DataPath_RF_bus_reg_dataout_2102_port,
                           regs(2101) => DataPath_RF_bus_reg_dataout_2101_port,
                           regs(2100) => DataPath_RF_bus_reg_dataout_2100_port,
                           regs(2099) => DataPath_RF_bus_reg_dataout_2099_port,
                           regs(2098) => DataPath_RF_bus_reg_dataout_2098_port,
                           regs(2097) => DataPath_RF_bus_reg_dataout_2097_port,
                           regs(2096) => DataPath_RF_bus_reg_dataout_2096_port,
                           regs(2095) => DataPath_RF_bus_reg_dataout_2095_port,
                           regs(2094) => DataPath_RF_bus_reg_dataout_2094_port,
                           regs(2093) => DataPath_RF_bus_reg_dataout_2093_port,
                           regs(2092) => DataPath_RF_bus_reg_dataout_2092_port,
                           regs(2091) => DataPath_RF_bus_reg_dataout_2091_port,
                           regs(2090) => DataPath_RF_bus_reg_dataout_2090_port,
                           regs(2089) => DataPath_RF_bus_reg_dataout_2089_port,
                           regs(2088) => DataPath_RF_bus_reg_dataout_2088_port,
                           regs(2087) => DataPath_RF_bus_reg_dataout_2087_port,
                           regs(2086) => DataPath_RF_bus_reg_dataout_2086_port,
                           regs(2085) => DataPath_RF_bus_reg_dataout_2085_port,
                           regs(2084) => DataPath_RF_bus_reg_dataout_2084_port,
                           regs(2083) => DataPath_RF_bus_reg_dataout_2083_port,
                           regs(2082) => DataPath_RF_bus_reg_dataout_2082_port,
                           regs(2081) => DataPath_RF_bus_reg_dataout_2081_port,
                           regs(2080) => DataPath_RF_bus_reg_dataout_2080_port,
                           regs(2079) => DataPath_RF_bus_reg_dataout_2079_port,
                           regs(2078) => DataPath_RF_bus_reg_dataout_2078_port,
                           regs(2077) => DataPath_RF_bus_reg_dataout_2077_port,
                           regs(2076) => DataPath_RF_bus_reg_dataout_2076_port,
                           regs(2075) => DataPath_RF_bus_reg_dataout_2075_port,
                           regs(2074) => DataPath_RF_bus_reg_dataout_2074_port,
                           regs(2073) => DataPath_RF_bus_reg_dataout_2073_port,
                           regs(2072) => DataPath_RF_bus_reg_dataout_2072_port,
                           regs(2071) => DataPath_RF_bus_reg_dataout_2071_port,
                           regs(2070) => DataPath_RF_bus_reg_dataout_2070_port,
                           regs(2069) => DataPath_RF_bus_reg_dataout_2069_port,
                           regs(2068) => DataPath_RF_bus_reg_dataout_2068_port,
                           regs(2067) => DataPath_RF_bus_reg_dataout_2067_port,
                           regs(2066) => DataPath_RF_bus_reg_dataout_2066_port,
                           regs(2065) => DataPath_RF_bus_reg_dataout_2065_port,
                           regs(2064) => DataPath_RF_bus_reg_dataout_2064_port,
                           regs(2063) => DataPath_RF_bus_reg_dataout_2063_port,
                           regs(2062) => DataPath_RF_bus_reg_dataout_2062_port,
                           regs(2061) => DataPath_RF_bus_reg_dataout_2061_port,
                           regs(2060) => DataPath_RF_bus_reg_dataout_2060_port,
                           regs(2059) => DataPath_RF_bus_reg_dataout_2059_port,
                           regs(2058) => DataPath_RF_bus_reg_dataout_2058_port,
                           regs(2057) => DataPath_RF_bus_reg_dataout_2057_port,
                           regs(2056) => DataPath_RF_bus_reg_dataout_2056_port,
                           regs(2055) => DataPath_RF_bus_reg_dataout_2055_port,
                           regs(2054) => DataPath_RF_bus_reg_dataout_2054_port,
                           regs(2053) => DataPath_RF_bus_reg_dataout_2053_port,
                           regs(2052) => DataPath_RF_bus_reg_dataout_2052_port,
                           regs(2051) => DataPath_RF_bus_reg_dataout_2051_port,
                           regs(2050) => DataPath_RF_bus_reg_dataout_2050_port,
                           regs(2049) => DataPath_RF_bus_reg_dataout_2049_port,
                           regs(2048) => DataPath_RF_bus_reg_dataout_2048_port,
                           regs(2047) => DataPath_RF_bus_reg_dataout_2047_port,
                           regs(2046) => DataPath_RF_bus_reg_dataout_2046_port,
                           regs(2045) => DataPath_RF_bus_reg_dataout_2045_port,
                           regs(2044) => DataPath_RF_bus_reg_dataout_2044_port,
                           regs(2043) => DataPath_RF_bus_reg_dataout_2043_port,
                           regs(2042) => DataPath_RF_bus_reg_dataout_2042_port,
                           regs(2041) => DataPath_RF_bus_reg_dataout_2041_port,
                           regs(2040) => DataPath_RF_bus_reg_dataout_2040_port,
                           regs(2039) => DataPath_RF_bus_reg_dataout_2039_port,
                           regs(2038) => DataPath_RF_bus_reg_dataout_2038_port,
                           regs(2037) => DataPath_RF_bus_reg_dataout_2037_port,
                           regs(2036) => DataPath_RF_bus_reg_dataout_2036_port,
                           regs(2035) => DataPath_RF_bus_reg_dataout_2035_port,
                           regs(2034) => DataPath_RF_bus_reg_dataout_2034_port,
                           regs(2033) => DataPath_RF_bus_reg_dataout_2033_port,
                           regs(2032) => DataPath_RF_bus_reg_dataout_2032_port,
                           regs(2031) => DataPath_RF_bus_reg_dataout_2031_port,
                           regs(2030) => DataPath_RF_bus_reg_dataout_2030_port,
                           regs(2029) => DataPath_RF_bus_reg_dataout_2029_port,
                           regs(2028) => DataPath_RF_bus_reg_dataout_2028_port,
                           regs(2027) => DataPath_RF_bus_reg_dataout_2027_port,
                           regs(2026) => DataPath_RF_bus_reg_dataout_2026_port,
                           regs(2025) => DataPath_RF_bus_reg_dataout_2025_port,
                           regs(2024) => DataPath_RF_bus_reg_dataout_2024_port,
                           regs(2023) => DataPath_RF_bus_reg_dataout_2023_port,
                           regs(2022) => DataPath_RF_bus_reg_dataout_2022_port,
                           regs(2021) => DataPath_RF_bus_reg_dataout_2021_port,
                           regs(2020) => DataPath_RF_bus_reg_dataout_2020_port,
                           regs(2019) => DataPath_RF_bus_reg_dataout_2019_port,
                           regs(2018) => DataPath_RF_bus_reg_dataout_2018_port,
                           regs(2017) => DataPath_RF_bus_reg_dataout_2017_port,
                           regs(2016) => DataPath_RF_bus_reg_dataout_2016_port,
                           regs(2015) => DataPath_RF_bus_reg_dataout_2015_port,
                           regs(2014) => DataPath_RF_bus_reg_dataout_2014_port,
                           regs(2013) => DataPath_RF_bus_reg_dataout_2013_port,
                           regs(2012) => DataPath_RF_bus_reg_dataout_2012_port,
                           regs(2011) => DataPath_RF_bus_reg_dataout_2011_port,
                           regs(2010) => DataPath_RF_bus_reg_dataout_2010_port,
                           regs(2009) => DataPath_RF_bus_reg_dataout_2009_port,
                           regs(2008) => DataPath_RF_bus_reg_dataout_2008_port,
                           regs(2007) => DataPath_RF_bus_reg_dataout_2007_port,
                           regs(2006) => DataPath_RF_bus_reg_dataout_2006_port,
                           regs(2005) => DataPath_RF_bus_reg_dataout_2005_port,
                           regs(2004) => DataPath_RF_bus_reg_dataout_2004_port,
                           regs(2003) => DataPath_RF_bus_reg_dataout_2003_port,
                           regs(2002) => DataPath_RF_bus_reg_dataout_2002_port,
                           regs(2001) => DataPath_RF_bus_reg_dataout_2001_port,
                           regs(2000) => DataPath_RF_bus_reg_dataout_2000_port,
                           regs(1999) => DataPath_RF_bus_reg_dataout_1999_port,
                           regs(1998) => DataPath_RF_bus_reg_dataout_1998_port,
                           regs(1997) => DataPath_RF_bus_reg_dataout_1997_port,
                           regs(1996) => DataPath_RF_bus_reg_dataout_1996_port,
                           regs(1995) => DataPath_RF_bus_reg_dataout_1995_port,
                           regs(1994) => DataPath_RF_bus_reg_dataout_1994_port,
                           regs(1993) => DataPath_RF_bus_reg_dataout_1993_port,
                           regs(1992) => DataPath_RF_bus_reg_dataout_1992_port,
                           regs(1991) => DataPath_RF_bus_reg_dataout_1991_port,
                           regs(1990) => DataPath_RF_bus_reg_dataout_1990_port,
                           regs(1989) => DataPath_RF_bus_reg_dataout_1989_port,
                           regs(1988) => DataPath_RF_bus_reg_dataout_1988_port,
                           regs(1987) => DataPath_RF_bus_reg_dataout_1987_port,
                           regs(1986) => DataPath_RF_bus_reg_dataout_1986_port,
                           regs(1985) => DataPath_RF_bus_reg_dataout_1985_port,
                           regs(1984) => DataPath_RF_bus_reg_dataout_1984_port,
                           regs(1983) => DataPath_RF_bus_reg_dataout_1983_port,
                           regs(1982) => DataPath_RF_bus_reg_dataout_1982_port,
                           regs(1981) => DataPath_RF_bus_reg_dataout_1981_port,
                           regs(1980) => DataPath_RF_bus_reg_dataout_1980_port,
                           regs(1979) => DataPath_RF_bus_reg_dataout_1979_port,
                           regs(1978) => DataPath_RF_bus_reg_dataout_1978_port,
                           regs(1977) => DataPath_RF_bus_reg_dataout_1977_port,
                           regs(1976) => DataPath_RF_bus_reg_dataout_1976_port,
                           regs(1975) => DataPath_RF_bus_reg_dataout_1975_port,
                           regs(1974) => DataPath_RF_bus_reg_dataout_1974_port,
                           regs(1973) => DataPath_RF_bus_reg_dataout_1973_port,
                           regs(1972) => DataPath_RF_bus_reg_dataout_1972_port,
                           regs(1971) => DataPath_RF_bus_reg_dataout_1971_port,
                           regs(1970) => DataPath_RF_bus_reg_dataout_1970_port,
                           regs(1969) => DataPath_RF_bus_reg_dataout_1969_port,
                           regs(1968) => DataPath_RF_bus_reg_dataout_1968_port,
                           regs(1967) => DataPath_RF_bus_reg_dataout_1967_port,
                           regs(1966) => DataPath_RF_bus_reg_dataout_1966_port,
                           regs(1965) => DataPath_RF_bus_reg_dataout_1965_port,
                           regs(1964) => DataPath_RF_bus_reg_dataout_1964_port,
                           regs(1963) => DataPath_RF_bus_reg_dataout_1963_port,
                           regs(1962) => DataPath_RF_bus_reg_dataout_1962_port,
                           regs(1961) => DataPath_RF_bus_reg_dataout_1961_port,
                           regs(1960) => DataPath_RF_bus_reg_dataout_1960_port,
                           regs(1959) => DataPath_RF_bus_reg_dataout_1959_port,
                           regs(1958) => DataPath_RF_bus_reg_dataout_1958_port,
                           regs(1957) => DataPath_RF_bus_reg_dataout_1957_port,
                           regs(1956) => DataPath_RF_bus_reg_dataout_1956_port,
                           regs(1955) => DataPath_RF_bus_reg_dataout_1955_port,
                           regs(1954) => DataPath_RF_bus_reg_dataout_1954_port,
                           regs(1953) => DataPath_RF_bus_reg_dataout_1953_port,
                           regs(1952) => DataPath_RF_bus_reg_dataout_1952_port,
                           regs(1951) => DataPath_RF_bus_reg_dataout_1951_port,
                           regs(1950) => DataPath_RF_bus_reg_dataout_1950_port,
                           regs(1949) => DataPath_RF_bus_reg_dataout_1949_port,
                           regs(1948) => DataPath_RF_bus_reg_dataout_1948_port,
                           regs(1947) => DataPath_RF_bus_reg_dataout_1947_port,
                           regs(1946) => DataPath_RF_bus_reg_dataout_1946_port,
                           regs(1945) => DataPath_RF_bus_reg_dataout_1945_port,
                           regs(1944) => DataPath_RF_bus_reg_dataout_1944_port,
                           regs(1943) => DataPath_RF_bus_reg_dataout_1943_port,
                           regs(1942) => DataPath_RF_bus_reg_dataout_1942_port,
                           regs(1941) => DataPath_RF_bus_reg_dataout_1941_port,
                           regs(1940) => DataPath_RF_bus_reg_dataout_1940_port,
                           regs(1939) => DataPath_RF_bus_reg_dataout_1939_port,
                           regs(1938) => DataPath_RF_bus_reg_dataout_1938_port,
                           regs(1937) => DataPath_RF_bus_reg_dataout_1937_port,
                           regs(1936) => DataPath_RF_bus_reg_dataout_1936_port,
                           regs(1935) => DataPath_RF_bus_reg_dataout_1935_port,
                           regs(1934) => DataPath_RF_bus_reg_dataout_1934_port,
                           regs(1933) => DataPath_RF_bus_reg_dataout_1933_port,
                           regs(1932) => DataPath_RF_bus_reg_dataout_1932_port,
                           regs(1931) => DataPath_RF_bus_reg_dataout_1931_port,
                           regs(1930) => DataPath_RF_bus_reg_dataout_1930_port,
                           regs(1929) => DataPath_RF_bus_reg_dataout_1929_port,
                           regs(1928) => DataPath_RF_bus_reg_dataout_1928_port,
                           regs(1927) => DataPath_RF_bus_reg_dataout_1927_port,
                           regs(1926) => DataPath_RF_bus_reg_dataout_1926_port,
                           regs(1925) => DataPath_RF_bus_reg_dataout_1925_port,
                           regs(1924) => DataPath_RF_bus_reg_dataout_1924_port,
                           regs(1923) => DataPath_RF_bus_reg_dataout_1923_port,
                           regs(1922) => DataPath_RF_bus_reg_dataout_1922_port,
                           regs(1921) => DataPath_RF_bus_reg_dataout_1921_port,
                           regs(1920) => DataPath_RF_bus_reg_dataout_1920_port,
                           regs(1919) => DataPath_RF_bus_reg_dataout_1919_port,
                           regs(1918) => DataPath_RF_bus_reg_dataout_1918_port,
                           regs(1917) => DataPath_RF_bus_reg_dataout_1917_port,
                           regs(1916) => DataPath_RF_bus_reg_dataout_1916_port,
                           regs(1915) => DataPath_RF_bus_reg_dataout_1915_port,
                           regs(1914) => DataPath_RF_bus_reg_dataout_1914_port,
                           regs(1913) => DataPath_RF_bus_reg_dataout_1913_port,
                           regs(1912) => DataPath_RF_bus_reg_dataout_1912_port,
                           regs(1911) => DataPath_RF_bus_reg_dataout_1911_port,
                           regs(1910) => DataPath_RF_bus_reg_dataout_1910_port,
                           regs(1909) => DataPath_RF_bus_reg_dataout_1909_port,
                           regs(1908) => DataPath_RF_bus_reg_dataout_1908_port,
                           regs(1907) => DataPath_RF_bus_reg_dataout_1907_port,
                           regs(1906) => DataPath_RF_bus_reg_dataout_1906_port,
                           regs(1905) => DataPath_RF_bus_reg_dataout_1905_port,
                           regs(1904) => DataPath_RF_bus_reg_dataout_1904_port,
                           regs(1903) => DataPath_RF_bus_reg_dataout_1903_port,
                           regs(1902) => DataPath_RF_bus_reg_dataout_1902_port,
                           regs(1901) => DataPath_RF_bus_reg_dataout_1901_port,
                           regs(1900) => DataPath_RF_bus_reg_dataout_1900_port,
                           regs(1899) => DataPath_RF_bus_reg_dataout_1899_port,
                           regs(1898) => DataPath_RF_bus_reg_dataout_1898_port,
                           regs(1897) => DataPath_RF_bus_reg_dataout_1897_port,
                           regs(1896) => DataPath_RF_bus_reg_dataout_1896_port,
                           regs(1895) => DataPath_RF_bus_reg_dataout_1895_port,
                           regs(1894) => DataPath_RF_bus_reg_dataout_1894_port,
                           regs(1893) => DataPath_RF_bus_reg_dataout_1893_port,
                           regs(1892) => DataPath_RF_bus_reg_dataout_1892_port,
                           regs(1891) => DataPath_RF_bus_reg_dataout_1891_port,
                           regs(1890) => DataPath_RF_bus_reg_dataout_1890_port,
                           regs(1889) => DataPath_RF_bus_reg_dataout_1889_port,
                           regs(1888) => DataPath_RF_bus_reg_dataout_1888_port,
                           regs(1887) => DataPath_RF_bus_reg_dataout_1887_port,
                           regs(1886) => DataPath_RF_bus_reg_dataout_1886_port,
                           regs(1885) => DataPath_RF_bus_reg_dataout_1885_port,
                           regs(1884) => DataPath_RF_bus_reg_dataout_1884_port,
                           regs(1883) => DataPath_RF_bus_reg_dataout_1883_port,
                           regs(1882) => DataPath_RF_bus_reg_dataout_1882_port,
                           regs(1881) => DataPath_RF_bus_reg_dataout_1881_port,
                           regs(1880) => DataPath_RF_bus_reg_dataout_1880_port,
                           regs(1879) => DataPath_RF_bus_reg_dataout_1879_port,
                           regs(1878) => DataPath_RF_bus_reg_dataout_1878_port,
                           regs(1877) => DataPath_RF_bus_reg_dataout_1877_port,
                           regs(1876) => DataPath_RF_bus_reg_dataout_1876_port,
                           regs(1875) => DataPath_RF_bus_reg_dataout_1875_port,
                           regs(1874) => DataPath_RF_bus_reg_dataout_1874_port,
                           regs(1873) => DataPath_RF_bus_reg_dataout_1873_port,
                           regs(1872) => DataPath_RF_bus_reg_dataout_1872_port,
                           regs(1871) => DataPath_RF_bus_reg_dataout_1871_port,
                           regs(1870) => DataPath_RF_bus_reg_dataout_1870_port,
                           regs(1869) => DataPath_RF_bus_reg_dataout_1869_port,
                           regs(1868) => DataPath_RF_bus_reg_dataout_1868_port,
                           regs(1867) => DataPath_RF_bus_reg_dataout_1867_port,
                           regs(1866) => DataPath_RF_bus_reg_dataout_1866_port,
                           regs(1865) => DataPath_RF_bus_reg_dataout_1865_port,
                           regs(1864) => DataPath_RF_bus_reg_dataout_1864_port,
                           regs(1863) => DataPath_RF_bus_reg_dataout_1863_port,
                           regs(1862) => DataPath_RF_bus_reg_dataout_1862_port,
                           regs(1861) => DataPath_RF_bus_reg_dataout_1861_port,
                           regs(1860) => DataPath_RF_bus_reg_dataout_1860_port,
                           regs(1859) => DataPath_RF_bus_reg_dataout_1859_port,
                           regs(1858) => DataPath_RF_bus_reg_dataout_1858_port,
                           regs(1857) => DataPath_RF_bus_reg_dataout_1857_port,
                           regs(1856) => DataPath_RF_bus_reg_dataout_1856_port,
                           regs(1855) => DataPath_RF_bus_reg_dataout_1855_port,
                           regs(1854) => DataPath_RF_bus_reg_dataout_1854_port,
                           regs(1853) => DataPath_RF_bus_reg_dataout_1853_port,
                           regs(1852) => DataPath_RF_bus_reg_dataout_1852_port,
                           regs(1851) => DataPath_RF_bus_reg_dataout_1851_port,
                           regs(1850) => DataPath_RF_bus_reg_dataout_1850_port,
                           regs(1849) => DataPath_RF_bus_reg_dataout_1849_port,
                           regs(1848) => DataPath_RF_bus_reg_dataout_1848_port,
                           regs(1847) => DataPath_RF_bus_reg_dataout_1847_port,
                           regs(1846) => DataPath_RF_bus_reg_dataout_1846_port,
                           regs(1845) => DataPath_RF_bus_reg_dataout_1845_port,
                           regs(1844) => DataPath_RF_bus_reg_dataout_1844_port,
                           regs(1843) => DataPath_RF_bus_reg_dataout_1843_port,
                           regs(1842) => DataPath_RF_bus_reg_dataout_1842_port,
                           regs(1841) => DataPath_RF_bus_reg_dataout_1841_port,
                           regs(1840) => DataPath_RF_bus_reg_dataout_1840_port,
                           regs(1839) => DataPath_RF_bus_reg_dataout_1839_port,
                           regs(1838) => DataPath_RF_bus_reg_dataout_1838_port,
                           regs(1837) => DataPath_RF_bus_reg_dataout_1837_port,
                           regs(1836) => DataPath_RF_bus_reg_dataout_1836_port,
                           regs(1835) => DataPath_RF_bus_reg_dataout_1835_port,
                           regs(1834) => DataPath_RF_bus_reg_dataout_1834_port,
                           regs(1833) => DataPath_RF_bus_reg_dataout_1833_port,
                           regs(1832) => DataPath_RF_bus_reg_dataout_1832_port,
                           regs(1831) => DataPath_RF_bus_reg_dataout_1831_port,
                           regs(1830) => DataPath_RF_bus_reg_dataout_1830_port,
                           regs(1829) => DataPath_RF_bus_reg_dataout_1829_port,
                           regs(1828) => DataPath_RF_bus_reg_dataout_1828_port,
                           regs(1827) => DataPath_RF_bus_reg_dataout_1827_port,
                           regs(1826) => DataPath_RF_bus_reg_dataout_1826_port,
                           regs(1825) => DataPath_RF_bus_reg_dataout_1825_port,
                           regs(1824) => DataPath_RF_bus_reg_dataout_1824_port,
                           regs(1823) => DataPath_RF_bus_reg_dataout_1823_port,
                           regs(1822) => DataPath_RF_bus_reg_dataout_1822_port,
                           regs(1821) => DataPath_RF_bus_reg_dataout_1821_port,
                           regs(1820) => DataPath_RF_bus_reg_dataout_1820_port,
                           regs(1819) => DataPath_RF_bus_reg_dataout_1819_port,
                           regs(1818) => DataPath_RF_bus_reg_dataout_1818_port,
                           regs(1817) => DataPath_RF_bus_reg_dataout_1817_port,
                           regs(1816) => DataPath_RF_bus_reg_dataout_1816_port,
                           regs(1815) => DataPath_RF_bus_reg_dataout_1815_port,
                           regs(1814) => DataPath_RF_bus_reg_dataout_1814_port,
                           regs(1813) => DataPath_RF_bus_reg_dataout_1813_port,
                           regs(1812) => DataPath_RF_bus_reg_dataout_1812_port,
                           regs(1811) => DataPath_RF_bus_reg_dataout_1811_port,
                           regs(1810) => DataPath_RF_bus_reg_dataout_1810_port,
                           regs(1809) => DataPath_RF_bus_reg_dataout_1809_port,
                           regs(1808) => DataPath_RF_bus_reg_dataout_1808_port,
                           regs(1807) => DataPath_RF_bus_reg_dataout_1807_port,
                           regs(1806) => DataPath_RF_bus_reg_dataout_1806_port,
                           regs(1805) => DataPath_RF_bus_reg_dataout_1805_port,
                           regs(1804) => DataPath_RF_bus_reg_dataout_1804_port,
                           regs(1803) => DataPath_RF_bus_reg_dataout_1803_port,
                           regs(1802) => DataPath_RF_bus_reg_dataout_1802_port,
                           regs(1801) => DataPath_RF_bus_reg_dataout_1801_port,
                           regs(1800) => DataPath_RF_bus_reg_dataout_1800_port,
                           regs(1799) => DataPath_RF_bus_reg_dataout_1799_port,
                           regs(1798) => DataPath_RF_bus_reg_dataout_1798_port,
                           regs(1797) => DataPath_RF_bus_reg_dataout_1797_port,
                           regs(1796) => DataPath_RF_bus_reg_dataout_1796_port,
                           regs(1795) => DataPath_RF_bus_reg_dataout_1795_port,
                           regs(1794) => DataPath_RF_bus_reg_dataout_1794_port,
                           regs(1793) => DataPath_RF_bus_reg_dataout_1793_port,
                           regs(1792) => DataPath_RF_bus_reg_dataout_1792_port,
                           regs(1791) => DataPath_RF_bus_reg_dataout_1791_port,
                           regs(1790) => DataPath_RF_bus_reg_dataout_1790_port,
                           regs(1789) => DataPath_RF_bus_reg_dataout_1789_port,
                           regs(1788) => DataPath_RF_bus_reg_dataout_1788_port,
                           regs(1787) => DataPath_RF_bus_reg_dataout_1787_port,
                           regs(1786) => DataPath_RF_bus_reg_dataout_1786_port,
                           regs(1785) => DataPath_RF_bus_reg_dataout_1785_port,
                           regs(1784) => DataPath_RF_bus_reg_dataout_1784_port,
                           regs(1783) => DataPath_RF_bus_reg_dataout_1783_port,
                           regs(1782) => DataPath_RF_bus_reg_dataout_1782_port,
                           regs(1781) => DataPath_RF_bus_reg_dataout_1781_port,
                           regs(1780) => DataPath_RF_bus_reg_dataout_1780_port,
                           regs(1779) => DataPath_RF_bus_reg_dataout_1779_port,
                           regs(1778) => DataPath_RF_bus_reg_dataout_1778_port,
                           regs(1777) => DataPath_RF_bus_reg_dataout_1777_port,
                           regs(1776) => DataPath_RF_bus_reg_dataout_1776_port,
                           regs(1775) => DataPath_RF_bus_reg_dataout_1775_port,
                           regs(1774) => DataPath_RF_bus_reg_dataout_1774_port,
                           regs(1773) => DataPath_RF_bus_reg_dataout_1773_port,
                           regs(1772) => DataPath_RF_bus_reg_dataout_1772_port,
                           regs(1771) => DataPath_RF_bus_reg_dataout_1771_port,
                           regs(1770) => DataPath_RF_bus_reg_dataout_1770_port,
                           regs(1769) => DataPath_RF_bus_reg_dataout_1769_port,
                           regs(1768) => DataPath_RF_bus_reg_dataout_1768_port,
                           regs(1767) => DataPath_RF_bus_reg_dataout_1767_port,
                           regs(1766) => DataPath_RF_bus_reg_dataout_1766_port,
                           regs(1765) => DataPath_RF_bus_reg_dataout_1765_port,
                           regs(1764) => DataPath_RF_bus_reg_dataout_1764_port,
                           regs(1763) => DataPath_RF_bus_reg_dataout_1763_port,
                           regs(1762) => DataPath_RF_bus_reg_dataout_1762_port,
                           regs(1761) => DataPath_RF_bus_reg_dataout_1761_port,
                           regs(1760) => DataPath_RF_bus_reg_dataout_1760_port,
                           regs(1759) => DataPath_RF_bus_reg_dataout_1759_port,
                           regs(1758) => DataPath_RF_bus_reg_dataout_1758_port,
                           regs(1757) => DataPath_RF_bus_reg_dataout_1757_port,
                           regs(1756) => DataPath_RF_bus_reg_dataout_1756_port,
                           regs(1755) => DataPath_RF_bus_reg_dataout_1755_port,
                           regs(1754) => DataPath_RF_bus_reg_dataout_1754_port,
                           regs(1753) => DataPath_RF_bus_reg_dataout_1753_port,
                           regs(1752) => DataPath_RF_bus_reg_dataout_1752_port,
                           regs(1751) => DataPath_RF_bus_reg_dataout_1751_port,
                           regs(1750) => DataPath_RF_bus_reg_dataout_1750_port,
                           regs(1749) => DataPath_RF_bus_reg_dataout_1749_port,
                           regs(1748) => DataPath_RF_bus_reg_dataout_1748_port,
                           regs(1747) => DataPath_RF_bus_reg_dataout_1747_port,
                           regs(1746) => DataPath_RF_bus_reg_dataout_1746_port,
                           regs(1745) => DataPath_RF_bus_reg_dataout_1745_port,
                           regs(1744) => DataPath_RF_bus_reg_dataout_1744_port,
                           regs(1743) => DataPath_RF_bus_reg_dataout_1743_port,
                           regs(1742) => DataPath_RF_bus_reg_dataout_1742_port,
                           regs(1741) => DataPath_RF_bus_reg_dataout_1741_port,
                           regs(1740) => DataPath_RF_bus_reg_dataout_1740_port,
                           regs(1739) => DataPath_RF_bus_reg_dataout_1739_port,
                           regs(1738) => DataPath_RF_bus_reg_dataout_1738_port,
                           regs(1737) => DataPath_RF_bus_reg_dataout_1737_port,
                           regs(1736) => DataPath_RF_bus_reg_dataout_1736_port,
                           regs(1735) => DataPath_RF_bus_reg_dataout_1735_port,
                           regs(1734) => DataPath_RF_bus_reg_dataout_1734_port,
                           regs(1733) => DataPath_RF_bus_reg_dataout_1733_port,
                           regs(1732) => DataPath_RF_bus_reg_dataout_1732_port,
                           regs(1731) => DataPath_RF_bus_reg_dataout_1731_port,
                           regs(1730) => DataPath_RF_bus_reg_dataout_1730_port,
                           regs(1729) => DataPath_RF_bus_reg_dataout_1729_port,
                           regs(1728) => DataPath_RF_bus_reg_dataout_1728_port,
                           regs(1727) => DataPath_RF_bus_reg_dataout_1727_port,
                           regs(1726) => DataPath_RF_bus_reg_dataout_1726_port,
                           regs(1725) => DataPath_RF_bus_reg_dataout_1725_port,
                           regs(1724) => DataPath_RF_bus_reg_dataout_1724_port,
                           regs(1723) => DataPath_RF_bus_reg_dataout_1723_port,
                           regs(1722) => DataPath_RF_bus_reg_dataout_1722_port,
                           regs(1721) => DataPath_RF_bus_reg_dataout_1721_port,
                           regs(1720) => DataPath_RF_bus_reg_dataout_1720_port,
                           regs(1719) => DataPath_RF_bus_reg_dataout_1719_port,
                           regs(1718) => DataPath_RF_bus_reg_dataout_1718_port,
                           regs(1717) => DataPath_RF_bus_reg_dataout_1717_port,
                           regs(1716) => DataPath_RF_bus_reg_dataout_1716_port,
                           regs(1715) => DataPath_RF_bus_reg_dataout_1715_port,
                           regs(1714) => DataPath_RF_bus_reg_dataout_1714_port,
                           regs(1713) => DataPath_RF_bus_reg_dataout_1713_port,
                           regs(1712) => DataPath_RF_bus_reg_dataout_1712_port,
                           regs(1711) => DataPath_RF_bus_reg_dataout_1711_port,
                           regs(1710) => DataPath_RF_bus_reg_dataout_1710_port,
                           regs(1709) => DataPath_RF_bus_reg_dataout_1709_port,
                           regs(1708) => DataPath_RF_bus_reg_dataout_1708_port,
                           regs(1707) => DataPath_RF_bus_reg_dataout_1707_port,
                           regs(1706) => DataPath_RF_bus_reg_dataout_1706_port,
                           regs(1705) => DataPath_RF_bus_reg_dataout_1705_port,
                           regs(1704) => DataPath_RF_bus_reg_dataout_1704_port,
                           regs(1703) => DataPath_RF_bus_reg_dataout_1703_port,
                           regs(1702) => DataPath_RF_bus_reg_dataout_1702_port,
                           regs(1701) => DataPath_RF_bus_reg_dataout_1701_port,
                           regs(1700) => DataPath_RF_bus_reg_dataout_1700_port,
                           regs(1699) => DataPath_RF_bus_reg_dataout_1699_port,
                           regs(1698) => DataPath_RF_bus_reg_dataout_1698_port,
                           regs(1697) => DataPath_RF_bus_reg_dataout_1697_port,
                           regs(1696) => DataPath_RF_bus_reg_dataout_1696_port,
                           regs(1695) => DataPath_RF_bus_reg_dataout_1695_port,
                           regs(1694) => DataPath_RF_bus_reg_dataout_1694_port,
                           regs(1693) => DataPath_RF_bus_reg_dataout_1693_port,
                           regs(1692) => DataPath_RF_bus_reg_dataout_1692_port,
                           regs(1691) => DataPath_RF_bus_reg_dataout_1691_port,
                           regs(1690) => DataPath_RF_bus_reg_dataout_1690_port,
                           regs(1689) => DataPath_RF_bus_reg_dataout_1689_port,
                           regs(1688) => DataPath_RF_bus_reg_dataout_1688_port,
                           regs(1687) => DataPath_RF_bus_reg_dataout_1687_port,
                           regs(1686) => DataPath_RF_bus_reg_dataout_1686_port,
                           regs(1685) => DataPath_RF_bus_reg_dataout_1685_port,
                           regs(1684) => DataPath_RF_bus_reg_dataout_1684_port,
                           regs(1683) => DataPath_RF_bus_reg_dataout_1683_port,
                           regs(1682) => DataPath_RF_bus_reg_dataout_1682_port,
                           regs(1681) => DataPath_RF_bus_reg_dataout_1681_port,
                           regs(1680) => DataPath_RF_bus_reg_dataout_1680_port,
                           regs(1679) => DataPath_RF_bus_reg_dataout_1679_port,
                           regs(1678) => DataPath_RF_bus_reg_dataout_1678_port,
                           regs(1677) => DataPath_RF_bus_reg_dataout_1677_port,
                           regs(1676) => DataPath_RF_bus_reg_dataout_1676_port,
                           regs(1675) => DataPath_RF_bus_reg_dataout_1675_port,
                           regs(1674) => DataPath_RF_bus_reg_dataout_1674_port,
                           regs(1673) => DataPath_RF_bus_reg_dataout_1673_port,
                           regs(1672) => DataPath_RF_bus_reg_dataout_1672_port,
                           regs(1671) => DataPath_RF_bus_reg_dataout_1671_port,
                           regs(1670) => DataPath_RF_bus_reg_dataout_1670_port,
                           regs(1669) => DataPath_RF_bus_reg_dataout_1669_port,
                           regs(1668) => DataPath_RF_bus_reg_dataout_1668_port,
                           regs(1667) => DataPath_RF_bus_reg_dataout_1667_port,
                           regs(1666) => DataPath_RF_bus_reg_dataout_1666_port,
                           regs(1665) => DataPath_RF_bus_reg_dataout_1665_port,
                           regs(1664) => DataPath_RF_bus_reg_dataout_1664_port,
                           regs(1663) => DataPath_RF_bus_reg_dataout_1663_port,
                           regs(1662) => DataPath_RF_bus_reg_dataout_1662_port,
                           regs(1661) => DataPath_RF_bus_reg_dataout_1661_port,
                           regs(1660) => DataPath_RF_bus_reg_dataout_1660_port,
                           regs(1659) => DataPath_RF_bus_reg_dataout_1659_port,
                           regs(1658) => DataPath_RF_bus_reg_dataout_1658_port,
                           regs(1657) => DataPath_RF_bus_reg_dataout_1657_port,
                           regs(1656) => DataPath_RF_bus_reg_dataout_1656_port,
                           regs(1655) => DataPath_RF_bus_reg_dataout_1655_port,
                           regs(1654) => DataPath_RF_bus_reg_dataout_1654_port,
                           regs(1653) => DataPath_RF_bus_reg_dataout_1653_port,
                           regs(1652) => DataPath_RF_bus_reg_dataout_1652_port,
                           regs(1651) => DataPath_RF_bus_reg_dataout_1651_port,
                           regs(1650) => DataPath_RF_bus_reg_dataout_1650_port,
                           regs(1649) => DataPath_RF_bus_reg_dataout_1649_port,
                           regs(1648) => DataPath_RF_bus_reg_dataout_1648_port,
                           regs(1647) => DataPath_RF_bus_reg_dataout_1647_port,
                           regs(1646) => DataPath_RF_bus_reg_dataout_1646_port,
                           regs(1645) => DataPath_RF_bus_reg_dataout_1645_port,
                           regs(1644) => DataPath_RF_bus_reg_dataout_1644_port,
                           regs(1643) => DataPath_RF_bus_reg_dataout_1643_port,
                           regs(1642) => DataPath_RF_bus_reg_dataout_1642_port,
                           regs(1641) => DataPath_RF_bus_reg_dataout_1641_port,
                           regs(1640) => DataPath_RF_bus_reg_dataout_1640_port,
                           regs(1639) => DataPath_RF_bus_reg_dataout_1639_port,
                           regs(1638) => DataPath_RF_bus_reg_dataout_1638_port,
                           regs(1637) => DataPath_RF_bus_reg_dataout_1637_port,
                           regs(1636) => DataPath_RF_bus_reg_dataout_1636_port,
                           regs(1635) => DataPath_RF_bus_reg_dataout_1635_port,
                           regs(1634) => DataPath_RF_bus_reg_dataout_1634_port,
                           regs(1633) => DataPath_RF_bus_reg_dataout_1633_port,
                           regs(1632) => DataPath_RF_bus_reg_dataout_1632_port,
                           regs(1631) => DataPath_RF_bus_reg_dataout_1631_port,
                           regs(1630) => DataPath_RF_bus_reg_dataout_1630_port,
                           regs(1629) => DataPath_RF_bus_reg_dataout_1629_port,
                           regs(1628) => DataPath_RF_bus_reg_dataout_1628_port,
                           regs(1627) => DataPath_RF_bus_reg_dataout_1627_port,
                           regs(1626) => DataPath_RF_bus_reg_dataout_1626_port,
                           regs(1625) => DataPath_RF_bus_reg_dataout_1625_port,
                           regs(1624) => DataPath_RF_bus_reg_dataout_1624_port,
                           regs(1623) => DataPath_RF_bus_reg_dataout_1623_port,
                           regs(1622) => DataPath_RF_bus_reg_dataout_1622_port,
                           regs(1621) => DataPath_RF_bus_reg_dataout_1621_port,
                           regs(1620) => DataPath_RF_bus_reg_dataout_1620_port,
                           regs(1619) => DataPath_RF_bus_reg_dataout_1619_port,
                           regs(1618) => DataPath_RF_bus_reg_dataout_1618_port,
                           regs(1617) => DataPath_RF_bus_reg_dataout_1617_port,
                           regs(1616) => DataPath_RF_bus_reg_dataout_1616_port,
                           regs(1615) => DataPath_RF_bus_reg_dataout_1615_port,
                           regs(1614) => DataPath_RF_bus_reg_dataout_1614_port,
                           regs(1613) => DataPath_RF_bus_reg_dataout_1613_port,
                           regs(1612) => DataPath_RF_bus_reg_dataout_1612_port,
                           regs(1611) => DataPath_RF_bus_reg_dataout_1611_port,
                           regs(1610) => DataPath_RF_bus_reg_dataout_1610_port,
                           regs(1609) => DataPath_RF_bus_reg_dataout_1609_port,
                           regs(1608) => DataPath_RF_bus_reg_dataout_1608_port,
                           regs(1607) => DataPath_RF_bus_reg_dataout_1607_port,
                           regs(1606) => DataPath_RF_bus_reg_dataout_1606_port,
                           regs(1605) => DataPath_RF_bus_reg_dataout_1605_port,
                           regs(1604) => DataPath_RF_bus_reg_dataout_1604_port,
                           regs(1603) => DataPath_RF_bus_reg_dataout_1603_port,
                           regs(1602) => DataPath_RF_bus_reg_dataout_1602_port,
                           regs(1601) => DataPath_RF_bus_reg_dataout_1601_port,
                           regs(1600) => DataPath_RF_bus_reg_dataout_1600_port,
                           regs(1599) => DataPath_RF_bus_reg_dataout_1599_port,
                           regs(1598) => DataPath_RF_bus_reg_dataout_1598_port,
                           regs(1597) => DataPath_RF_bus_reg_dataout_1597_port,
                           regs(1596) => DataPath_RF_bus_reg_dataout_1596_port,
                           regs(1595) => DataPath_RF_bus_reg_dataout_1595_port,
                           regs(1594) => DataPath_RF_bus_reg_dataout_1594_port,
                           regs(1593) => DataPath_RF_bus_reg_dataout_1593_port,
                           regs(1592) => DataPath_RF_bus_reg_dataout_1592_port,
                           regs(1591) => DataPath_RF_bus_reg_dataout_1591_port,
                           regs(1590) => DataPath_RF_bus_reg_dataout_1590_port,
                           regs(1589) => DataPath_RF_bus_reg_dataout_1589_port,
                           regs(1588) => DataPath_RF_bus_reg_dataout_1588_port,
                           regs(1587) => DataPath_RF_bus_reg_dataout_1587_port,
                           regs(1586) => DataPath_RF_bus_reg_dataout_1586_port,
                           regs(1585) => DataPath_RF_bus_reg_dataout_1585_port,
                           regs(1584) => DataPath_RF_bus_reg_dataout_1584_port,
                           regs(1583) => DataPath_RF_bus_reg_dataout_1583_port,
                           regs(1582) => DataPath_RF_bus_reg_dataout_1582_port,
                           regs(1581) => DataPath_RF_bus_reg_dataout_1581_port,
                           regs(1580) => DataPath_RF_bus_reg_dataout_1580_port,
                           regs(1579) => DataPath_RF_bus_reg_dataout_1579_port,
                           regs(1578) => DataPath_RF_bus_reg_dataout_1578_port,
                           regs(1577) => DataPath_RF_bus_reg_dataout_1577_port,
                           regs(1576) => DataPath_RF_bus_reg_dataout_1576_port,
                           regs(1575) => DataPath_RF_bus_reg_dataout_1575_port,
                           regs(1574) => DataPath_RF_bus_reg_dataout_1574_port,
                           regs(1573) => DataPath_RF_bus_reg_dataout_1573_port,
                           regs(1572) => DataPath_RF_bus_reg_dataout_1572_port,
                           regs(1571) => DataPath_RF_bus_reg_dataout_1571_port,
                           regs(1570) => DataPath_RF_bus_reg_dataout_1570_port,
                           regs(1569) => DataPath_RF_bus_reg_dataout_1569_port,
                           regs(1568) => DataPath_RF_bus_reg_dataout_1568_port,
                           regs(1567) => DataPath_RF_bus_reg_dataout_1567_port,
                           regs(1566) => DataPath_RF_bus_reg_dataout_1566_port,
                           regs(1565) => DataPath_RF_bus_reg_dataout_1565_port,
                           regs(1564) => DataPath_RF_bus_reg_dataout_1564_port,
                           regs(1563) => DataPath_RF_bus_reg_dataout_1563_port,
                           regs(1562) => DataPath_RF_bus_reg_dataout_1562_port,
                           regs(1561) => DataPath_RF_bus_reg_dataout_1561_port,
                           regs(1560) => DataPath_RF_bus_reg_dataout_1560_port,
                           regs(1559) => DataPath_RF_bus_reg_dataout_1559_port,
                           regs(1558) => DataPath_RF_bus_reg_dataout_1558_port,
                           regs(1557) => DataPath_RF_bus_reg_dataout_1557_port,
                           regs(1556) => DataPath_RF_bus_reg_dataout_1556_port,
                           regs(1555) => DataPath_RF_bus_reg_dataout_1555_port,
                           regs(1554) => DataPath_RF_bus_reg_dataout_1554_port,
                           regs(1553) => DataPath_RF_bus_reg_dataout_1553_port,
                           regs(1552) => DataPath_RF_bus_reg_dataout_1552_port,
                           regs(1551) => DataPath_RF_bus_reg_dataout_1551_port,
                           regs(1550) => DataPath_RF_bus_reg_dataout_1550_port,
                           regs(1549) => DataPath_RF_bus_reg_dataout_1549_port,
                           regs(1548) => DataPath_RF_bus_reg_dataout_1548_port,
                           regs(1547) => DataPath_RF_bus_reg_dataout_1547_port,
                           regs(1546) => DataPath_RF_bus_reg_dataout_1546_port,
                           regs(1545) => DataPath_RF_bus_reg_dataout_1545_port,
                           regs(1544) => DataPath_RF_bus_reg_dataout_1544_port,
                           regs(1543) => DataPath_RF_bus_reg_dataout_1543_port,
                           regs(1542) => DataPath_RF_bus_reg_dataout_1542_port,
                           regs(1541) => DataPath_RF_bus_reg_dataout_1541_port,
                           regs(1540) => DataPath_RF_bus_reg_dataout_1540_port,
                           regs(1539) => DataPath_RF_bus_reg_dataout_1539_port,
                           regs(1538) => DataPath_RF_bus_reg_dataout_1538_port,
                           regs(1537) => DataPath_RF_bus_reg_dataout_1537_port,
                           regs(1536) => DataPath_RF_bus_reg_dataout_1536_port,
                           regs(1535) => DataPath_RF_bus_reg_dataout_1535_port,
                           regs(1534) => DataPath_RF_bus_reg_dataout_1534_port,
                           regs(1533) => DataPath_RF_bus_reg_dataout_1533_port,
                           regs(1532) => DataPath_RF_bus_reg_dataout_1532_port,
                           regs(1531) => DataPath_RF_bus_reg_dataout_1531_port,
                           regs(1530) => DataPath_RF_bus_reg_dataout_1530_port,
                           regs(1529) => DataPath_RF_bus_reg_dataout_1529_port,
                           regs(1528) => DataPath_RF_bus_reg_dataout_1528_port,
                           regs(1527) => DataPath_RF_bus_reg_dataout_1527_port,
                           regs(1526) => DataPath_RF_bus_reg_dataout_1526_port,
                           regs(1525) => DataPath_RF_bus_reg_dataout_1525_port,
                           regs(1524) => DataPath_RF_bus_reg_dataout_1524_port,
                           regs(1523) => DataPath_RF_bus_reg_dataout_1523_port,
                           regs(1522) => DataPath_RF_bus_reg_dataout_1522_port,
                           regs(1521) => DataPath_RF_bus_reg_dataout_1521_port,
                           regs(1520) => DataPath_RF_bus_reg_dataout_1520_port,
                           regs(1519) => DataPath_RF_bus_reg_dataout_1519_port,
                           regs(1518) => DataPath_RF_bus_reg_dataout_1518_port,
                           regs(1517) => DataPath_RF_bus_reg_dataout_1517_port,
                           regs(1516) => DataPath_RF_bus_reg_dataout_1516_port,
                           regs(1515) => DataPath_RF_bus_reg_dataout_1515_port,
                           regs(1514) => DataPath_RF_bus_reg_dataout_1514_port,
                           regs(1513) => DataPath_RF_bus_reg_dataout_1513_port,
                           regs(1512) => DataPath_RF_bus_reg_dataout_1512_port,
                           regs(1511) => DataPath_RF_bus_reg_dataout_1511_port,
                           regs(1510) => DataPath_RF_bus_reg_dataout_1510_port,
                           regs(1509) => DataPath_RF_bus_reg_dataout_1509_port,
                           regs(1508) => DataPath_RF_bus_reg_dataout_1508_port,
                           regs(1507) => DataPath_RF_bus_reg_dataout_1507_port,
                           regs(1506) => DataPath_RF_bus_reg_dataout_1506_port,
                           regs(1505) => DataPath_RF_bus_reg_dataout_1505_port,
                           regs(1504) => DataPath_RF_bus_reg_dataout_1504_port,
                           regs(1503) => DataPath_RF_bus_reg_dataout_1503_port,
                           regs(1502) => DataPath_RF_bus_reg_dataout_1502_port,
                           regs(1501) => DataPath_RF_bus_reg_dataout_1501_port,
                           regs(1500) => DataPath_RF_bus_reg_dataout_1500_port,
                           regs(1499) => DataPath_RF_bus_reg_dataout_1499_port,
                           regs(1498) => DataPath_RF_bus_reg_dataout_1498_port,
                           regs(1497) => DataPath_RF_bus_reg_dataout_1497_port,
                           regs(1496) => DataPath_RF_bus_reg_dataout_1496_port,
                           regs(1495) => DataPath_RF_bus_reg_dataout_1495_port,
                           regs(1494) => DataPath_RF_bus_reg_dataout_1494_port,
                           regs(1493) => DataPath_RF_bus_reg_dataout_1493_port,
                           regs(1492) => DataPath_RF_bus_reg_dataout_1492_port,
                           regs(1491) => DataPath_RF_bus_reg_dataout_1491_port,
                           regs(1490) => DataPath_RF_bus_reg_dataout_1490_port,
                           regs(1489) => DataPath_RF_bus_reg_dataout_1489_port,
                           regs(1488) => DataPath_RF_bus_reg_dataout_1488_port,
                           regs(1487) => DataPath_RF_bus_reg_dataout_1487_port,
                           regs(1486) => DataPath_RF_bus_reg_dataout_1486_port,
                           regs(1485) => DataPath_RF_bus_reg_dataout_1485_port,
                           regs(1484) => DataPath_RF_bus_reg_dataout_1484_port,
                           regs(1483) => DataPath_RF_bus_reg_dataout_1483_port,
                           regs(1482) => DataPath_RF_bus_reg_dataout_1482_port,
                           regs(1481) => DataPath_RF_bus_reg_dataout_1481_port,
                           regs(1480) => DataPath_RF_bus_reg_dataout_1480_port,
                           regs(1479) => DataPath_RF_bus_reg_dataout_1479_port,
                           regs(1478) => DataPath_RF_bus_reg_dataout_1478_port,
                           regs(1477) => DataPath_RF_bus_reg_dataout_1477_port,
                           regs(1476) => DataPath_RF_bus_reg_dataout_1476_port,
                           regs(1475) => DataPath_RF_bus_reg_dataout_1475_port,
                           regs(1474) => DataPath_RF_bus_reg_dataout_1474_port,
                           regs(1473) => DataPath_RF_bus_reg_dataout_1473_port,
                           regs(1472) => DataPath_RF_bus_reg_dataout_1472_port,
                           regs(1471) => DataPath_RF_bus_reg_dataout_1471_port,
                           regs(1470) => DataPath_RF_bus_reg_dataout_1470_port,
                           regs(1469) => DataPath_RF_bus_reg_dataout_1469_port,
                           regs(1468) => DataPath_RF_bus_reg_dataout_1468_port,
                           regs(1467) => DataPath_RF_bus_reg_dataout_1467_port,
                           regs(1466) => DataPath_RF_bus_reg_dataout_1466_port,
                           regs(1465) => DataPath_RF_bus_reg_dataout_1465_port,
                           regs(1464) => DataPath_RF_bus_reg_dataout_1464_port,
                           regs(1463) => DataPath_RF_bus_reg_dataout_1463_port,
                           regs(1462) => DataPath_RF_bus_reg_dataout_1462_port,
                           regs(1461) => DataPath_RF_bus_reg_dataout_1461_port,
                           regs(1460) => DataPath_RF_bus_reg_dataout_1460_port,
                           regs(1459) => DataPath_RF_bus_reg_dataout_1459_port,
                           regs(1458) => DataPath_RF_bus_reg_dataout_1458_port,
                           regs(1457) => DataPath_RF_bus_reg_dataout_1457_port,
                           regs(1456) => DataPath_RF_bus_reg_dataout_1456_port,
                           regs(1455) => DataPath_RF_bus_reg_dataout_1455_port,
                           regs(1454) => DataPath_RF_bus_reg_dataout_1454_port,
                           regs(1453) => DataPath_RF_bus_reg_dataout_1453_port,
                           regs(1452) => DataPath_RF_bus_reg_dataout_1452_port,
                           regs(1451) => DataPath_RF_bus_reg_dataout_1451_port,
                           regs(1450) => DataPath_RF_bus_reg_dataout_1450_port,
                           regs(1449) => DataPath_RF_bus_reg_dataout_1449_port,
                           regs(1448) => DataPath_RF_bus_reg_dataout_1448_port,
                           regs(1447) => DataPath_RF_bus_reg_dataout_1447_port,
                           regs(1446) => DataPath_RF_bus_reg_dataout_1446_port,
                           regs(1445) => DataPath_RF_bus_reg_dataout_1445_port,
                           regs(1444) => DataPath_RF_bus_reg_dataout_1444_port,
                           regs(1443) => DataPath_RF_bus_reg_dataout_1443_port,
                           regs(1442) => DataPath_RF_bus_reg_dataout_1442_port,
                           regs(1441) => DataPath_RF_bus_reg_dataout_1441_port,
                           regs(1440) => DataPath_RF_bus_reg_dataout_1440_port,
                           regs(1439) => DataPath_RF_bus_reg_dataout_1439_port,
                           regs(1438) => DataPath_RF_bus_reg_dataout_1438_port,
                           regs(1437) => DataPath_RF_bus_reg_dataout_1437_port,
                           regs(1436) => DataPath_RF_bus_reg_dataout_1436_port,
                           regs(1435) => DataPath_RF_bus_reg_dataout_1435_port,
                           regs(1434) => DataPath_RF_bus_reg_dataout_1434_port,
                           regs(1433) => DataPath_RF_bus_reg_dataout_1433_port,
                           regs(1432) => DataPath_RF_bus_reg_dataout_1432_port,
                           regs(1431) => DataPath_RF_bus_reg_dataout_1431_port,
                           regs(1430) => DataPath_RF_bus_reg_dataout_1430_port,
                           regs(1429) => DataPath_RF_bus_reg_dataout_1429_port,
                           regs(1428) => DataPath_RF_bus_reg_dataout_1428_port,
                           regs(1427) => DataPath_RF_bus_reg_dataout_1427_port,
                           regs(1426) => DataPath_RF_bus_reg_dataout_1426_port,
                           regs(1425) => DataPath_RF_bus_reg_dataout_1425_port,
                           regs(1424) => DataPath_RF_bus_reg_dataout_1424_port,
                           regs(1423) => DataPath_RF_bus_reg_dataout_1423_port,
                           regs(1422) => DataPath_RF_bus_reg_dataout_1422_port,
                           regs(1421) => DataPath_RF_bus_reg_dataout_1421_port,
                           regs(1420) => DataPath_RF_bus_reg_dataout_1420_port,
                           regs(1419) => DataPath_RF_bus_reg_dataout_1419_port,
                           regs(1418) => DataPath_RF_bus_reg_dataout_1418_port,
                           regs(1417) => DataPath_RF_bus_reg_dataout_1417_port,
                           regs(1416) => DataPath_RF_bus_reg_dataout_1416_port,
                           regs(1415) => DataPath_RF_bus_reg_dataout_1415_port,
                           regs(1414) => DataPath_RF_bus_reg_dataout_1414_port,
                           regs(1413) => DataPath_RF_bus_reg_dataout_1413_port,
                           regs(1412) => DataPath_RF_bus_reg_dataout_1412_port,
                           regs(1411) => DataPath_RF_bus_reg_dataout_1411_port,
                           regs(1410) => DataPath_RF_bus_reg_dataout_1410_port,
                           regs(1409) => DataPath_RF_bus_reg_dataout_1409_port,
                           regs(1408) => DataPath_RF_bus_reg_dataout_1408_port,
                           regs(1407) => DataPath_RF_bus_reg_dataout_1407_port,
                           regs(1406) => DataPath_RF_bus_reg_dataout_1406_port,
                           regs(1405) => DataPath_RF_bus_reg_dataout_1405_port,
                           regs(1404) => DataPath_RF_bus_reg_dataout_1404_port,
                           regs(1403) => DataPath_RF_bus_reg_dataout_1403_port,
                           regs(1402) => DataPath_RF_bus_reg_dataout_1402_port,
                           regs(1401) => DataPath_RF_bus_reg_dataout_1401_port,
                           regs(1400) => DataPath_RF_bus_reg_dataout_1400_port,
                           regs(1399) => DataPath_RF_bus_reg_dataout_1399_port,
                           regs(1398) => DataPath_RF_bus_reg_dataout_1398_port,
                           regs(1397) => DataPath_RF_bus_reg_dataout_1397_port,
                           regs(1396) => DataPath_RF_bus_reg_dataout_1396_port,
                           regs(1395) => DataPath_RF_bus_reg_dataout_1395_port,
                           regs(1394) => DataPath_RF_bus_reg_dataout_1394_port,
                           regs(1393) => DataPath_RF_bus_reg_dataout_1393_port,
                           regs(1392) => DataPath_RF_bus_reg_dataout_1392_port,
                           regs(1391) => DataPath_RF_bus_reg_dataout_1391_port,
                           regs(1390) => DataPath_RF_bus_reg_dataout_1390_port,
                           regs(1389) => DataPath_RF_bus_reg_dataout_1389_port,
                           regs(1388) => DataPath_RF_bus_reg_dataout_1388_port,
                           regs(1387) => DataPath_RF_bus_reg_dataout_1387_port,
                           regs(1386) => DataPath_RF_bus_reg_dataout_1386_port,
                           regs(1385) => DataPath_RF_bus_reg_dataout_1385_port,
                           regs(1384) => DataPath_RF_bus_reg_dataout_1384_port,
                           regs(1383) => DataPath_RF_bus_reg_dataout_1383_port,
                           regs(1382) => DataPath_RF_bus_reg_dataout_1382_port,
                           regs(1381) => DataPath_RF_bus_reg_dataout_1381_port,
                           regs(1380) => DataPath_RF_bus_reg_dataout_1380_port,
                           regs(1379) => DataPath_RF_bus_reg_dataout_1379_port,
                           regs(1378) => DataPath_RF_bus_reg_dataout_1378_port,
                           regs(1377) => DataPath_RF_bus_reg_dataout_1377_port,
                           regs(1376) => DataPath_RF_bus_reg_dataout_1376_port,
                           regs(1375) => DataPath_RF_bus_reg_dataout_1375_port,
                           regs(1374) => DataPath_RF_bus_reg_dataout_1374_port,
                           regs(1373) => DataPath_RF_bus_reg_dataout_1373_port,
                           regs(1372) => DataPath_RF_bus_reg_dataout_1372_port,
                           regs(1371) => DataPath_RF_bus_reg_dataout_1371_port,
                           regs(1370) => DataPath_RF_bus_reg_dataout_1370_port,
                           regs(1369) => DataPath_RF_bus_reg_dataout_1369_port,
                           regs(1368) => DataPath_RF_bus_reg_dataout_1368_port,
                           regs(1367) => DataPath_RF_bus_reg_dataout_1367_port,
                           regs(1366) => DataPath_RF_bus_reg_dataout_1366_port,
                           regs(1365) => DataPath_RF_bus_reg_dataout_1365_port,
                           regs(1364) => DataPath_RF_bus_reg_dataout_1364_port,
                           regs(1363) => DataPath_RF_bus_reg_dataout_1363_port,
                           regs(1362) => DataPath_RF_bus_reg_dataout_1362_port,
                           regs(1361) => DataPath_RF_bus_reg_dataout_1361_port,
                           regs(1360) => DataPath_RF_bus_reg_dataout_1360_port,
                           regs(1359) => DataPath_RF_bus_reg_dataout_1359_port,
                           regs(1358) => DataPath_RF_bus_reg_dataout_1358_port,
                           regs(1357) => DataPath_RF_bus_reg_dataout_1357_port,
                           regs(1356) => DataPath_RF_bus_reg_dataout_1356_port,
                           regs(1355) => DataPath_RF_bus_reg_dataout_1355_port,
                           regs(1354) => DataPath_RF_bus_reg_dataout_1354_port,
                           regs(1353) => DataPath_RF_bus_reg_dataout_1353_port,
                           regs(1352) => DataPath_RF_bus_reg_dataout_1352_port,
                           regs(1351) => DataPath_RF_bus_reg_dataout_1351_port,
                           regs(1350) => DataPath_RF_bus_reg_dataout_1350_port,
                           regs(1349) => DataPath_RF_bus_reg_dataout_1349_port,
                           regs(1348) => DataPath_RF_bus_reg_dataout_1348_port,
                           regs(1347) => DataPath_RF_bus_reg_dataout_1347_port,
                           regs(1346) => DataPath_RF_bus_reg_dataout_1346_port,
                           regs(1345) => DataPath_RF_bus_reg_dataout_1345_port,
                           regs(1344) => DataPath_RF_bus_reg_dataout_1344_port,
                           regs(1343) => DataPath_RF_bus_reg_dataout_1343_port,
                           regs(1342) => DataPath_RF_bus_reg_dataout_1342_port,
                           regs(1341) => DataPath_RF_bus_reg_dataout_1341_port,
                           regs(1340) => DataPath_RF_bus_reg_dataout_1340_port,
                           regs(1339) => DataPath_RF_bus_reg_dataout_1339_port,
                           regs(1338) => DataPath_RF_bus_reg_dataout_1338_port,
                           regs(1337) => DataPath_RF_bus_reg_dataout_1337_port,
                           regs(1336) => DataPath_RF_bus_reg_dataout_1336_port,
                           regs(1335) => DataPath_RF_bus_reg_dataout_1335_port,
                           regs(1334) => DataPath_RF_bus_reg_dataout_1334_port,
                           regs(1333) => DataPath_RF_bus_reg_dataout_1333_port,
                           regs(1332) => DataPath_RF_bus_reg_dataout_1332_port,
                           regs(1331) => DataPath_RF_bus_reg_dataout_1331_port,
                           regs(1330) => DataPath_RF_bus_reg_dataout_1330_port,
                           regs(1329) => DataPath_RF_bus_reg_dataout_1329_port,
                           regs(1328) => DataPath_RF_bus_reg_dataout_1328_port,
                           regs(1327) => DataPath_RF_bus_reg_dataout_1327_port,
                           regs(1326) => DataPath_RF_bus_reg_dataout_1326_port,
                           regs(1325) => DataPath_RF_bus_reg_dataout_1325_port,
                           regs(1324) => DataPath_RF_bus_reg_dataout_1324_port,
                           regs(1323) => DataPath_RF_bus_reg_dataout_1323_port,
                           regs(1322) => DataPath_RF_bus_reg_dataout_1322_port,
                           regs(1321) => DataPath_RF_bus_reg_dataout_1321_port,
                           regs(1320) => DataPath_RF_bus_reg_dataout_1320_port,
                           regs(1319) => DataPath_RF_bus_reg_dataout_1319_port,
                           regs(1318) => DataPath_RF_bus_reg_dataout_1318_port,
                           regs(1317) => DataPath_RF_bus_reg_dataout_1317_port,
                           regs(1316) => DataPath_RF_bus_reg_dataout_1316_port,
                           regs(1315) => DataPath_RF_bus_reg_dataout_1315_port,
                           regs(1314) => DataPath_RF_bus_reg_dataout_1314_port,
                           regs(1313) => DataPath_RF_bus_reg_dataout_1313_port,
                           regs(1312) => DataPath_RF_bus_reg_dataout_1312_port,
                           regs(1311) => DataPath_RF_bus_reg_dataout_1311_port,
                           regs(1310) => DataPath_RF_bus_reg_dataout_1310_port,
                           regs(1309) => DataPath_RF_bus_reg_dataout_1309_port,
                           regs(1308) => DataPath_RF_bus_reg_dataout_1308_port,
                           regs(1307) => DataPath_RF_bus_reg_dataout_1307_port,
                           regs(1306) => DataPath_RF_bus_reg_dataout_1306_port,
                           regs(1305) => DataPath_RF_bus_reg_dataout_1305_port,
                           regs(1304) => DataPath_RF_bus_reg_dataout_1304_port,
                           regs(1303) => DataPath_RF_bus_reg_dataout_1303_port,
                           regs(1302) => DataPath_RF_bus_reg_dataout_1302_port,
                           regs(1301) => DataPath_RF_bus_reg_dataout_1301_port,
                           regs(1300) => DataPath_RF_bus_reg_dataout_1300_port,
                           regs(1299) => DataPath_RF_bus_reg_dataout_1299_port,
                           regs(1298) => DataPath_RF_bus_reg_dataout_1298_port,
                           regs(1297) => DataPath_RF_bus_reg_dataout_1297_port,
                           regs(1296) => DataPath_RF_bus_reg_dataout_1296_port,
                           regs(1295) => DataPath_RF_bus_reg_dataout_1295_port,
                           regs(1294) => DataPath_RF_bus_reg_dataout_1294_port,
                           regs(1293) => DataPath_RF_bus_reg_dataout_1293_port,
                           regs(1292) => DataPath_RF_bus_reg_dataout_1292_port,
                           regs(1291) => DataPath_RF_bus_reg_dataout_1291_port,
                           regs(1290) => DataPath_RF_bus_reg_dataout_1290_port,
                           regs(1289) => DataPath_RF_bus_reg_dataout_1289_port,
                           regs(1288) => DataPath_RF_bus_reg_dataout_1288_port,
                           regs(1287) => DataPath_RF_bus_reg_dataout_1287_port,
                           regs(1286) => DataPath_RF_bus_reg_dataout_1286_port,
                           regs(1285) => DataPath_RF_bus_reg_dataout_1285_port,
                           regs(1284) => DataPath_RF_bus_reg_dataout_1284_port,
                           regs(1283) => DataPath_RF_bus_reg_dataout_1283_port,
                           regs(1282) => DataPath_RF_bus_reg_dataout_1282_port,
                           regs(1281) => DataPath_RF_bus_reg_dataout_1281_port,
                           regs(1280) => DataPath_RF_bus_reg_dataout_1280_port,
                           regs(1279) => DataPath_RF_bus_reg_dataout_1279_port,
                           regs(1278) => DataPath_RF_bus_reg_dataout_1278_port,
                           regs(1277) => DataPath_RF_bus_reg_dataout_1277_port,
                           regs(1276) => DataPath_RF_bus_reg_dataout_1276_port,
                           regs(1275) => DataPath_RF_bus_reg_dataout_1275_port,
                           regs(1274) => DataPath_RF_bus_reg_dataout_1274_port,
                           regs(1273) => DataPath_RF_bus_reg_dataout_1273_port,
                           regs(1272) => DataPath_RF_bus_reg_dataout_1272_port,
                           regs(1271) => DataPath_RF_bus_reg_dataout_1271_port,
                           regs(1270) => DataPath_RF_bus_reg_dataout_1270_port,
                           regs(1269) => DataPath_RF_bus_reg_dataout_1269_port,
                           regs(1268) => DataPath_RF_bus_reg_dataout_1268_port,
                           regs(1267) => DataPath_RF_bus_reg_dataout_1267_port,
                           regs(1266) => DataPath_RF_bus_reg_dataout_1266_port,
                           regs(1265) => DataPath_RF_bus_reg_dataout_1265_port,
                           regs(1264) => DataPath_RF_bus_reg_dataout_1264_port,
                           regs(1263) => DataPath_RF_bus_reg_dataout_1263_port,
                           regs(1262) => DataPath_RF_bus_reg_dataout_1262_port,
                           regs(1261) => DataPath_RF_bus_reg_dataout_1261_port,
                           regs(1260) => DataPath_RF_bus_reg_dataout_1260_port,
                           regs(1259) => DataPath_RF_bus_reg_dataout_1259_port,
                           regs(1258) => DataPath_RF_bus_reg_dataout_1258_port,
                           regs(1257) => DataPath_RF_bus_reg_dataout_1257_port,
                           regs(1256) => DataPath_RF_bus_reg_dataout_1256_port,
                           regs(1255) => DataPath_RF_bus_reg_dataout_1255_port,
                           regs(1254) => DataPath_RF_bus_reg_dataout_1254_port,
                           regs(1253) => DataPath_RF_bus_reg_dataout_1253_port,
                           regs(1252) => DataPath_RF_bus_reg_dataout_1252_port,
                           regs(1251) => DataPath_RF_bus_reg_dataout_1251_port,
                           regs(1250) => DataPath_RF_bus_reg_dataout_1250_port,
                           regs(1249) => DataPath_RF_bus_reg_dataout_1249_port,
                           regs(1248) => DataPath_RF_bus_reg_dataout_1248_port,
                           regs(1247) => DataPath_RF_bus_reg_dataout_1247_port,
                           regs(1246) => DataPath_RF_bus_reg_dataout_1246_port,
                           regs(1245) => DataPath_RF_bus_reg_dataout_1245_port,
                           regs(1244) => DataPath_RF_bus_reg_dataout_1244_port,
                           regs(1243) => DataPath_RF_bus_reg_dataout_1243_port,
                           regs(1242) => DataPath_RF_bus_reg_dataout_1242_port,
                           regs(1241) => DataPath_RF_bus_reg_dataout_1241_port,
                           regs(1240) => DataPath_RF_bus_reg_dataout_1240_port,
                           regs(1239) => DataPath_RF_bus_reg_dataout_1239_port,
                           regs(1238) => DataPath_RF_bus_reg_dataout_1238_port,
                           regs(1237) => DataPath_RF_bus_reg_dataout_1237_port,
                           regs(1236) => DataPath_RF_bus_reg_dataout_1236_port,
                           regs(1235) => DataPath_RF_bus_reg_dataout_1235_port,
                           regs(1234) => DataPath_RF_bus_reg_dataout_1234_port,
                           regs(1233) => DataPath_RF_bus_reg_dataout_1233_port,
                           regs(1232) => DataPath_RF_bus_reg_dataout_1232_port,
                           regs(1231) => DataPath_RF_bus_reg_dataout_1231_port,
                           regs(1230) => DataPath_RF_bus_reg_dataout_1230_port,
                           regs(1229) => DataPath_RF_bus_reg_dataout_1229_port,
                           regs(1228) => DataPath_RF_bus_reg_dataout_1228_port,
                           regs(1227) => DataPath_RF_bus_reg_dataout_1227_port,
                           regs(1226) => DataPath_RF_bus_reg_dataout_1226_port,
                           regs(1225) => DataPath_RF_bus_reg_dataout_1225_port,
                           regs(1224) => DataPath_RF_bus_reg_dataout_1224_port,
                           regs(1223) => DataPath_RF_bus_reg_dataout_1223_port,
                           regs(1222) => DataPath_RF_bus_reg_dataout_1222_port,
                           regs(1221) => DataPath_RF_bus_reg_dataout_1221_port,
                           regs(1220) => DataPath_RF_bus_reg_dataout_1220_port,
                           regs(1219) => DataPath_RF_bus_reg_dataout_1219_port,
                           regs(1218) => DataPath_RF_bus_reg_dataout_1218_port,
                           regs(1217) => DataPath_RF_bus_reg_dataout_1217_port,
                           regs(1216) => DataPath_RF_bus_reg_dataout_1216_port,
                           regs(1215) => DataPath_RF_bus_reg_dataout_1215_port,
                           regs(1214) => DataPath_RF_bus_reg_dataout_1214_port,
                           regs(1213) => DataPath_RF_bus_reg_dataout_1213_port,
                           regs(1212) => DataPath_RF_bus_reg_dataout_1212_port,
                           regs(1211) => DataPath_RF_bus_reg_dataout_1211_port,
                           regs(1210) => DataPath_RF_bus_reg_dataout_1210_port,
                           regs(1209) => DataPath_RF_bus_reg_dataout_1209_port,
                           regs(1208) => DataPath_RF_bus_reg_dataout_1208_port,
                           regs(1207) => DataPath_RF_bus_reg_dataout_1207_port,
                           regs(1206) => DataPath_RF_bus_reg_dataout_1206_port,
                           regs(1205) => DataPath_RF_bus_reg_dataout_1205_port,
                           regs(1204) => DataPath_RF_bus_reg_dataout_1204_port,
                           regs(1203) => DataPath_RF_bus_reg_dataout_1203_port,
                           regs(1202) => DataPath_RF_bus_reg_dataout_1202_port,
                           regs(1201) => DataPath_RF_bus_reg_dataout_1201_port,
                           regs(1200) => DataPath_RF_bus_reg_dataout_1200_port,
                           regs(1199) => DataPath_RF_bus_reg_dataout_1199_port,
                           regs(1198) => DataPath_RF_bus_reg_dataout_1198_port,
                           regs(1197) => DataPath_RF_bus_reg_dataout_1197_port,
                           regs(1196) => DataPath_RF_bus_reg_dataout_1196_port,
                           regs(1195) => DataPath_RF_bus_reg_dataout_1195_port,
                           regs(1194) => DataPath_RF_bus_reg_dataout_1194_port,
                           regs(1193) => DataPath_RF_bus_reg_dataout_1193_port,
                           regs(1192) => DataPath_RF_bus_reg_dataout_1192_port,
                           regs(1191) => DataPath_RF_bus_reg_dataout_1191_port,
                           regs(1190) => DataPath_RF_bus_reg_dataout_1190_port,
                           regs(1189) => DataPath_RF_bus_reg_dataout_1189_port,
                           regs(1188) => DataPath_RF_bus_reg_dataout_1188_port,
                           regs(1187) => DataPath_RF_bus_reg_dataout_1187_port,
                           regs(1186) => DataPath_RF_bus_reg_dataout_1186_port,
                           regs(1185) => DataPath_RF_bus_reg_dataout_1185_port,
                           regs(1184) => DataPath_RF_bus_reg_dataout_1184_port,
                           regs(1183) => DataPath_RF_bus_reg_dataout_1183_port,
                           regs(1182) => DataPath_RF_bus_reg_dataout_1182_port,
                           regs(1181) => DataPath_RF_bus_reg_dataout_1181_port,
                           regs(1180) => DataPath_RF_bus_reg_dataout_1180_port,
                           regs(1179) => DataPath_RF_bus_reg_dataout_1179_port,
                           regs(1178) => DataPath_RF_bus_reg_dataout_1178_port,
                           regs(1177) => DataPath_RF_bus_reg_dataout_1177_port,
                           regs(1176) => DataPath_RF_bus_reg_dataout_1176_port,
                           regs(1175) => DataPath_RF_bus_reg_dataout_1175_port,
                           regs(1174) => DataPath_RF_bus_reg_dataout_1174_port,
                           regs(1173) => DataPath_RF_bus_reg_dataout_1173_port,
                           regs(1172) => DataPath_RF_bus_reg_dataout_1172_port,
                           regs(1171) => DataPath_RF_bus_reg_dataout_1171_port,
                           regs(1170) => DataPath_RF_bus_reg_dataout_1170_port,
                           regs(1169) => DataPath_RF_bus_reg_dataout_1169_port,
                           regs(1168) => DataPath_RF_bus_reg_dataout_1168_port,
                           regs(1167) => DataPath_RF_bus_reg_dataout_1167_port,
                           regs(1166) => DataPath_RF_bus_reg_dataout_1166_port,
                           regs(1165) => DataPath_RF_bus_reg_dataout_1165_port,
                           regs(1164) => DataPath_RF_bus_reg_dataout_1164_port,
                           regs(1163) => DataPath_RF_bus_reg_dataout_1163_port,
                           regs(1162) => DataPath_RF_bus_reg_dataout_1162_port,
                           regs(1161) => DataPath_RF_bus_reg_dataout_1161_port,
                           regs(1160) => DataPath_RF_bus_reg_dataout_1160_port,
                           regs(1159) => DataPath_RF_bus_reg_dataout_1159_port,
                           regs(1158) => DataPath_RF_bus_reg_dataout_1158_port,
                           regs(1157) => DataPath_RF_bus_reg_dataout_1157_port,
                           regs(1156) => DataPath_RF_bus_reg_dataout_1156_port,
                           regs(1155) => DataPath_RF_bus_reg_dataout_1155_port,
                           regs(1154) => DataPath_RF_bus_reg_dataout_1154_port,
                           regs(1153) => DataPath_RF_bus_reg_dataout_1153_port,
                           regs(1152) => DataPath_RF_bus_reg_dataout_1152_port,
                           regs(1151) => DataPath_RF_bus_reg_dataout_1151_port,
                           regs(1150) => DataPath_RF_bus_reg_dataout_1150_port,
                           regs(1149) => DataPath_RF_bus_reg_dataout_1149_port,
                           regs(1148) => DataPath_RF_bus_reg_dataout_1148_port,
                           regs(1147) => DataPath_RF_bus_reg_dataout_1147_port,
                           regs(1146) => DataPath_RF_bus_reg_dataout_1146_port,
                           regs(1145) => DataPath_RF_bus_reg_dataout_1145_port,
                           regs(1144) => DataPath_RF_bus_reg_dataout_1144_port,
                           regs(1143) => DataPath_RF_bus_reg_dataout_1143_port,
                           regs(1142) => DataPath_RF_bus_reg_dataout_1142_port,
                           regs(1141) => DataPath_RF_bus_reg_dataout_1141_port,
                           regs(1140) => DataPath_RF_bus_reg_dataout_1140_port,
                           regs(1139) => DataPath_RF_bus_reg_dataout_1139_port,
                           regs(1138) => DataPath_RF_bus_reg_dataout_1138_port,
                           regs(1137) => DataPath_RF_bus_reg_dataout_1137_port,
                           regs(1136) => DataPath_RF_bus_reg_dataout_1136_port,
                           regs(1135) => DataPath_RF_bus_reg_dataout_1135_port,
                           regs(1134) => DataPath_RF_bus_reg_dataout_1134_port,
                           regs(1133) => DataPath_RF_bus_reg_dataout_1133_port,
                           regs(1132) => DataPath_RF_bus_reg_dataout_1132_port,
                           regs(1131) => DataPath_RF_bus_reg_dataout_1131_port,
                           regs(1130) => DataPath_RF_bus_reg_dataout_1130_port,
                           regs(1129) => DataPath_RF_bus_reg_dataout_1129_port,
                           regs(1128) => DataPath_RF_bus_reg_dataout_1128_port,
                           regs(1127) => DataPath_RF_bus_reg_dataout_1127_port,
                           regs(1126) => DataPath_RF_bus_reg_dataout_1126_port,
                           regs(1125) => DataPath_RF_bus_reg_dataout_1125_port,
                           regs(1124) => DataPath_RF_bus_reg_dataout_1124_port,
                           regs(1123) => DataPath_RF_bus_reg_dataout_1123_port,
                           regs(1122) => DataPath_RF_bus_reg_dataout_1122_port,
                           regs(1121) => DataPath_RF_bus_reg_dataout_1121_port,
                           regs(1120) => DataPath_RF_bus_reg_dataout_1120_port,
                           regs(1119) => DataPath_RF_bus_reg_dataout_1119_port,
                           regs(1118) => DataPath_RF_bus_reg_dataout_1118_port,
                           regs(1117) => DataPath_RF_bus_reg_dataout_1117_port,
                           regs(1116) => DataPath_RF_bus_reg_dataout_1116_port,
                           regs(1115) => DataPath_RF_bus_reg_dataout_1115_port,
                           regs(1114) => DataPath_RF_bus_reg_dataout_1114_port,
                           regs(1113) => DataPath_RF_bus_reg_dataout_1113_port,
                           regs(1112) => DataPath_RF_bus_reg_dataout_1112_port,
                           regs(1111) => DataPath_RF_bus_reg_dataout_1111_port,
                           regs(1110) => DataPath_RF_bus_reg_dataout_1110_port,
                           regs(1109) => DataPath_RF_bus_reg_dataout_1109_port,
                           regs(1108) => DataPath_RF_bus_reg_dataout_1108_port,
                           regs(1107) => DataPath_RF_bus_reg_dataout_1107_port,
                           regs(1106) => DataPath_RF_bus_reg_dataout_1106_port,
                           regs(1105) => DataPath_RF_bus_reg_dataout_1105_port,
                           regs(1104) => DataPath_RF_bus_reg_dataout_1104_port,
                           regs(1103) => DataPath_RF_bus_reg_dataout_1103_port,
                           regs(1102) => DataPath_RF_bus_reg_dataout_1102_port,
                           regs(1101) => DataPath_RF_bus_reg_dataout_1101_port,
                           regs(1100) => DataPath_RF_bus_reg_dataout_1100_port,
                           regs(1099) => DataPath_RF_bus_reg_dataout_1099_port,
                           regs(1098) => DataPath_RF_bus_reg_dataout_1098_port,
                           regs(1097) => DataPath_RF_bus_reg_dataout_1097_port,
                           regs(1096) => DataPath_RF_bus_reg_dataout_1096_port,
                           regs(1095) => DataPath_RF_bus_reg_dataout_1095_port,
                           regs(1094) => DataPath_RF_bus_reg_dataout_1094_port,
                           regs(1093) => DataPath_RF_bus_reg_dataout_1093_port,
                           regs(1092) => DataPath_RF_bus_reg_dataout_1092_port,
                           regs(1091) => DataPath_RF_bus_reg_dataout_1091_port,
                           regs(1090) => DataPath_RF_bus_reg_dataout_1090_port,
                           regs(1089) => DataPath_RF_bus_reg_dataout_1089_port,
                           regs(1088) => DataPath_RF_bus_reg_dataout_1088_port,
                           regs(1087) => DataPath_RF_bus_reg_dataout_1087_port,
                           regs(1086) => DataPath_RF_bus_reg_dataout_1086_port,
                           regs(1085) => DataPath_RF_bus_reg_dataout_1085_port,
                           regs(1084) => DataPath_RF_bus_reg_dataout_1084_port,
                           regs(1083) => DataPath_RF_bus_reg_dataout_1083_port,
                           regs(1082) => DataPath_RF_bus_reg_dataout_1082_port,
                           regs(1081) => DataPath_RF_bus_reg_dataout_1081_port,
                           regs(1080) => DataPath_RF_bus_reg_dataout_1080_port,
                           regs(1079) => DataPath_RF_bus_reg_dataout_1079_port,
                           regs(1078) => DataPath_RF_bus_reg_dataout_1078_port,
                           regs(1077) => DataPath_RF_bus_reg_dataout_1077_port,
                           regs(1076) => DataPath_RF_bus_reg_dataout_1076_port,
                           regs(1075) => DataPath_RF_bus_reg_dataout_1075_port,
                           regs(1074) => DataPath_RF_bus_reg_dataout_1074_port,
                           regs(1073) => DataPath_RF_bus_reg_dataout_1073_port,
                           regs(1072) => DataPath_RF_bus_reg_dataout_1072_port,
                           regs(1071) => DataPath_RF_bus_reg_dataout_1071_port,
                           regs(1070) => DataPath_RF_bus_reg_dataout_1070_port,
                           regs(1069) => DataPath_RF_bus_reg_dataout_1069_port,
                           regs(1068) => DataPath_RF_bus_reg_dataout_1068_port,
                           regs(1067) => DataPath_RF_bus_reg_dataout_1067_port,
                           regs(1066) => DataPath_RF_bus_reg_dataout_1066_port,
                           regs(1065) => DataPath_RF_bus_reg_dataout_1065_port,
                           regs(1064) => DataPath_RF_bus_reg_dataout_1064_port,
                           regs(1063) => DataPath_RF_bus_reg_dataout_1063_port,
                           regs(1062) => DataPath_RF_bus_reg_dataout_1062_port,
                           regs(1061) => DataPath_RF_bus_reg_dataout_1061_port,
                           regs(1060) => DataPath_RF_bus_reg_dataout_1060_port,
                           regs(1059) => DataPath_RF_bus_reg_dataout_1059_port,
                           regs(1058) => DataPath_RF_bus_reg_dataout_1058_port,
                           regs(1057) => DataPath_RF_bus_reg_dataout_1057_port,
                           regs(1056) => DataPath_RF_bus_reg_dataout_1056_port,
                           regs(1055) => DataPath_RF_bus_reg_dataout_1055_port,
                           regs(1054) => DataPath_RF_bus_reg_dataout_1054_port,
                           regs(1053) => DataPath_RF_bus_reg_dataout_1053_port,
                           regs(1052) => DataPath_RF_bus_reg_dataout_1052_port,
                           regs(1051) => DataPath_RF_bus_reg_dataout_1051_port,
                           regs(1050) => DataPath_RF_bus_reg_dataout_1050_port,
                           regs(1049) => DataPath_RF_bus_reg_dataout_1049_port,
                           regs(1048) => DataPath_RF_bus_reg_dataout_1048_port,
                           regs(1047) => DataPath_RF_bus_reg_dataout_1047_port,
                           regs(1046) => DataPath_RF_bus_reg_dataout_1046_port,
                           regs(1045) => DataPath_RF_bus_reg_dataout_1045_port,
                           regs(1044) => DataPath_RF_bus_reg_dataout_1044_port,
                           regs(1043) => DataPath_RF_bus_reg_dataout_1043_port,
                           regs(1042) => DataPath_RF_bus_reg_dataout_1042_port,
                           regs(1041) => DataPath_RF_bus_reg_dataout_1041_port,
                           regs(1040) => DataPath_RF_bus_reg_dataout_1040_port,
                           regs(1039) => DataPath_RF_bus_reg_dataout_1039_port,
                           regs(1038) => DataPath_RF_bus_reg_dataout_1038_port,
                           regs(1037) => DataPath_RF_bus_reg_dataout_1037_port,
                           regs(1036) => DataPath_RF_bus_reg_dataout_1036_port,
                           regs(1035) => DataPath_RF_bus_reg_dataout_1035_port,
                           regs(1034) => DataPath_RF_bus_reg_dataout_1034_port,
                           regs(1033) => DataPath_RF_bus_reg_dataout_1033_port,
                           regs(1032) => DataPath_RF_bus_reg_dataout_1032_port,
                           regs(1031) => DataPath_RF_bus_reg_dataout_1031_port,
                           regs(1030) => DataPath_RF_bus_reg_dataout_1030_port,
                           regs(1029) => DataPath_RF_bus_reg_dataout_1029_port,
                           regs(1028) => DataPath_RF_bus_reg_dataout_1028_port,
                           regs(1027) => DataPath_RF_bus_reg_dataout_1027_port,
                           regs(1026) => DataPath_RF_bus_reg_dataout_1026_port,
                           regs(1025) => DataPath_RF_bus_reg_dataout_1025_port,
                           regs(1024) => DataPath_RF_bus_reg_dataout_1024_port,
                           regs(1023) => DataPath_RF_bus_reg_dataout_1023_port,
                           regs(1022) => DataPath_RF_bus_reg_dataout_1022_port,
                           regs(1021) => DataPath_RF_bus_reg_dataout_1021_port,
                           regs(1020) => DataPath_RF_bus_reg_dataout_1020_port,
                           regs(1019) => DataPath_RF_bus_reg_dataout_1019_port,
                           regs(1018) => DataPath_RF_bus_reg_dataout_1018_port,
                           regs(1017) => DataPath_RF_bus_reg_dataout_1017_port,
                           regs(1016) => DataPath_RF_bus_reg_dataout_1016_port,
                           regs(1015) => DataPath_RF_bus_reg_dataout_1015_port,
                           regs(1014) => DataPath_RF_bus_reg_dataout_1014_port,
                           regs(1013) => DataPath_RF_bus_reg_dataout_1013_port,
                           regs(1012) => DataPath_RF_bus_reg_dataout_1012_port,
                           regs(1011) => DataPath_RF_bus_reg_dataout_1011_port,
                           regs(1010) => DataPath_RF_bus_reg_dataout_1010_port,
                           regs(1009) => DataPath_RF_bus_reg_dataout_1009_port,
                           regs(1008) => DataPath_RF_bus_reg_dataout_1008_port,
                           regs(1007) => DataPath_RF_bus_reg_dataout_1007_port,
                           regs(1006) => DataPath_RF_bus_reg_dataout_1006_port,
                           regs(1005) => DataPath_RF_bus_reg_dataout_1005_port,
                           regs(1004) => DataPath_RF_bus_reg_dataout_1004_port,
                           regs(1003) => DataPath_RF_bus_reg_dataout_1003_port,
                           regs(1002) => DataPath_RF_bus_reg_dataout_1002_port,
                           regs(1001) => DataPath_RF_bus_reg_dataout_1001_port,
                           regs(1000) => DataPath_RF_bus_reg_dataout_1000_port,
                           regs(999) => DataPath_RF_bus_reg_dataout_999_port, 
                           regs(998) => DataPath_RF_bus_reg_dataout_998_port, 
                           regs(997) => DataPath_RF_bus_reg_dataout_997_port, 
                           regs(996) => DataPath_RF_bus_reg_dataout_996_port, 
                           regs(995) => DataPath_RF_bus_reg_dataout_995_port, 
                           regs(994) => DataPath_RF_bus_reg_dataout_994_port, 
                           regs(993) => DataPath_RF_bus_reg_dataout_993_port, 
                           regs(992) => DataPath_RF_bus_reg_dataout_992_port, 
                           regs(991) => DataPath_RF_bus_reg_dataout_991_port, 
                           regs(990) => DataPath_RF_bus_reg_dataout_990_port, 
                           regs(989) => DataPath_RF_bus_reg_dataout_989_port, 
                           regs(988) => DataPath_RF_bus_reg_dataout_988_port, 
                           regs(987) => DataPath_RF_bus_reg_dataout_987_port, 
                           regs(986) => DataPath_RF_bus_reg_dataout_986_port, 
                           regs(985) => DataPath_RF_bus_reg_dataout_985_port, 
                           regs(984) => DataPath_RF_bus_reg_dataout_984_port, 
                           regs(983) => DataPath_RF_bus_reg_dataout_983_port, 
                           regs(982) => DataPath_RF_bus_reg_dataout_982_port, 
                           regs(981) => DataPath_RF_bus_reg_dataout_981_port, 
                           regs(980) => DataPath_RF_bus_reg_dataout_980_port, 
                           regs(979) => DataPath_RF_bus_reg_dataout_979_port, 
                           regs(978) => DataPath_RF_bus_reg_dataout_978_port, 
                           regs(977) => DataPath_RF_bus_reg_dataout_977_port, 
                           regs(976) => DataPath_RF_bus_reg_dataout_976_port, 
                           regs(975) => DataPath_RF_bus_reg_dataout_975_port, 
                           regs(974) => DataPath_RF_bus_reg_dataout_974_port, 
                           regs(973) => DataPath_RF_bus_reg_dataout_973_port, 
                           regs(972) => DataPath_RF_bus_reg_dataout_972_port, 
                           regs(971) => DataPath_RF_bus_reg_dataout_971_port, 
                           regs(970) => DataPath_RF_bus_reg_dataout_970_port, 
                           regs(969) => DataPath_RF_bus_reg_dataout_969_port, 
                           regs(968) => DataPath_RF_bus_reg_dataout_968_port, 
                           regs(967) => DataPath_RF_bus_reg_dataout_967_port, 
                           regs(966) => DataPath_RF_bus_reg_dataout_966_port, 
                           regs(965) => DataPath_RF_bus_reg_dataout_965_port, 
                           regs(964) => DataPath_RF_bus_reg_dataout_964_port, 
                           regs(963) => DataPath_RF_bus_reg_dataout_963_port, 
                           regs(962) => DataPath_RF_bus_reg_dataout_962_port, 
                           regs(961) => DataPath_RF_bus_reg_dataout_961_port, 
                           regs(960) => DataPath_RF_bus_reg_dataout_960_port, 
                           regs(959) => DataPath_RF_bus_reg_dataout_959_port, 
                           regs(958) => DataPath_RF_bus_reg_dataout_958_port, 
                           regs(957) => DataPath_RF_bus_reg_dataout_957_port, 
                           regs(956) => DataPath_RF_bus_reg_dataout_956_port, 
                           regs(955) => DataPath_RF_bus_reg_dataout_955_port, 
                           regs(954) => DataPath_RF_bus_reg_dataout_954_port, 
                           regs(953) => DataPath_RF_bus_reg_dataout_953_port, 
                           regs(952) => DataPath_RF_bus_reg_dataout_952_port, 
                           regs(951) => DataPath_RF_bus_reg_dataout_951_port, 
                           regs(950) => DataPath_RF_bus_reg_dataout_950_port, 
                           regs(949) => DataPath_RF_bus_reg_dataout_949_port, 
                           regs(948) => DataPath_RF_bus_reg_dataout_948_port, 
                           regs(947) => DataPath_RF_bus_reg_dataout_947_port, 
                           regs(946) => DataPath_RF_bus_reg_dataout_946_port, 
                           regs(945) => DataPath_RF_bus_reg_dataout_945_port, 
                           regs(944) => DataPath_RF_bus_reg_dataout_944_port, 
                           regs(943) => DataPath_RF_bus_reg_dataout_943_port, 
                           regs(942) => DataPath_RF_bus_reg_dataout_942_port, 
                           regs(941) => DataPath_RF_bus_reg_dataout_941_port, 
                           regs(940) => DataPath_RF_bus_reg_dataout_940_port, 
                           regs(939) => DataPath_RF_bus_reg_dataout_939_port, 
                           regs(938) => DataPath_RF_bus_reg_dataout_938_port, 
                           regs(937) => DataPath_RF_bus_reg_dataout_937_port, 
                           regs(936) => DataPath_RF_bus_reg_dataout_936_port, 
                           regs(935) => DataPath_RF_bus_reg_dataout_935_port, 
                           regs(934) => DataPath_RF_bus_reg_dataout_934_port, 
                           regs(933) => DataPath_RF_bus_reg_dataout_933_port, 
                           regs(932) => DataPath_RF_bus_reg_dataout_932_port, 
                           regs(931) => DataPath_RF_bus_reg_dataout_931_port, 
                           regs(930) => DataPath_RF_bus_reg_dataout_930_port, 
                           regs(929) => DataPath_RF_bus_reg_dataout_929_port, 
                           regs(928) => DataPath_RF_bus_reg_dataout_928_port, 
                           regs(927) => DataPath_RF_bus_reg_dataout_927_port, 
                           regs(926) => DataPath_RF_bus_reg_dataout_926_port, 
                           regs(925) => DataPath_RF_bus_reg_dataout_925_port, 
                           regs(924) => DataPath_RF_bus_reg_dataout_924_port, 
                           regs(923) => DataPath_RF_bus_reg_dataout_923_port, 
                           regs(922) => DataPath_RF_bus_reg_dataout_922_port, 
                           regs(921) => DataPath_RF_bus_reg_dataout_921_port, 
                           regs(920) => DataPath_RF_bus_reg_dataout_920_port, 
                           regs(919) => DataPath_RF_bus_reg_dataout_919_port, 
                           regs(918) => DataPath_RF_bus_reg_dataout_918_port, 
                           regs(917) => DataPath_RF_bus_reg_dataout_917_port, 
                           regs(916) => DataPath_RF_bus_reg_dataout_916_port, 
                           regs(915) => DataPath_RF_bus_reg_dataout_915_port, 
                           regs(914) => DataPath_RF_bus_reg_dataout_914_port, 
                           regs(913) => DataPath_RF_bus_reg_dataout_913_port, 
                           regs(912) => DataPath_RF_bus_reg_dataout_912_port, 
                           regs(911) => DataPath_RF_bus_reg_dataout_911_port, 
                           regs(910) => DataPath_RF_bus_reg_dataout_910_port, 
                           regs(909) => DataPath_RF_bus_reg_dataout_909_port, 
                           regs(908) => DataPath_RF_bus_reg_dataout_908_port, 
                           regs(907) => DataPath_RF_bus_reg_dataout_907_port, 
                           regs(906) => DataPath_RF_bus_reg_dataout_906_port, 
                           regs(905) => DataPath_RF_bus_reg_dataout_905_port, 
                           regs(904) => DataPath_RF_bus_reg_dataout_904_port, 
                           regs(903) => DataPath_RF_bus_reg_dataout_903_port, 
                           regs(902) => DataPath_RF_bus_reg_dataout_902_port, 
                           regs(901) => DataPath_RF_bus_reg_dataout_901_port, 
                           regs(900) => DataPath_RF_bus_reg_dataout_900_port, 
                           regs(899) => DataPath_RF_bus_reg_dataout_899_port, 
                           regs(898) => DataPath_RF_bus_reg_dataout_898_port, 
                           regs(897) => DataPath_RF_bus_reg_dataout_897_port, 
                           regs(896) => DataPath_RF_bus_reg_dataout_896_port, 
                           regs(895) => DataPath_RF_bus_reg_dataout_895_port, 
                           regs(894) => DataPath_RF_bus_reg_dataout_894_port, 
                           regs(893) => DataPath_RF_bus_reg_dataout_893_port, 
                           regs(892) => DataPath_RF_bus_reg_dataout_892_port, 
                           regs(891) => DataPath_RF_bus_reg_dataout_891_port, 
                           regs(890) => DataPath_RF_bus_reg_dataout_890_port, 
                           regs(889) => DataPath_RF_bus_reg_dataout_889_port, 
                           regs(888) => DataPath_RF_bus_reg_dataout_888_port, 
                           regs(887) => DataPath_RF_bus_reg_dataout_887_port, 
                           regs(886) => DataPath_RF_bus_reg_dataout_886_port, 
                           regs(885) => DataPath_RF_bus_reg_dataout_885_port, 
                           regs(884) => DataPath_RF_bus_reg_dataout_884_port, 
                           regs(883) => DataPath_RF_bus_reg_dataout_883_port, 
                           regs(882) => DataPath_RF_bus_reg_dataout_882_port, 
                           regs(881) => DataPath_RF_bus_reg_dataout_881_port, 
                           regs(880) => DataPath_RF_bus_reg_dataout_880_port, 
                           regs(879) => DataPath_RF_bus_reg_dataout_879_port, 
                           regs(878) => DataPath_RF_bus_reg_dataout_878_port, 
                           regs(877) => DataPath_RF_bus_reg_dataout_877_port, 
                           regs(876) => DataPath_RF_bus_reg_dataout_876_port, 
                           regs(875) => DataPath_RF_bus_reg_dataout_875_port, 
                           regs(874) => DataPath_RF_bus_reg_dataout_874_port, 
                           regs(873) => DataPath_RF_bus_reg_dataout_873_port, 
                           regs(872) => DataPath_RF_bus_reg_dataout_872_port, 
                           regs(871) => DataPath_RF_bus_reg_dataout_871_port, 
                           regs(870) => DataPath_RF_bus_reg_dataout_870_port, 
                           regs(869) => DataPath_RF_bus_reg_dataout_869_port, 
                           regs(868) => DataPath_RF_bus_reg_dataout_868_port, 
                           regs(867) => DataPath_RF_bus_reg_dataout_867_port, 
                           regs(866) => DataPath_RF_bus_reg_dataout_866_port, 
                           regs(865) => DataPath_RF_bus_reg_dataout_865_port, 
                           regs(864) => DataPath_RF_bus_reg_dataout_864_port, 
                           regs(863) => DataPath_RF_bus_reg_dataout_863_port, 
                           regs(862) => DataPath_RF_bus_reg_dataout_862_port, 
                           regs(861) => DataPath_RF_bus_reg_dataout_861_port, 
                           regs(860) => DataPath_RF_bus_reg_dataout_860_port, 
                           regs(859) => DataPath_RF_bus_reg_dataout_859_port, 
                           regs(858) => DataPath_RF_bus_reg_dataout_858_port, 
                           regs(857) => DataPath_RF_bus_reg_dataout_857_port, 
                           regs(856) => DataPath_RF_bus_reg_dataout_856_port, 
                           regs(855) => DataPath_RF_bus_reg_dataout_855_port, 
                           regs(854) => DataPath_RF_bus_reg_dataout_854_port, 
                           regs(853) => DataPath_RF_bus_reg_dataout_853_port, 
                           regs(852) => DataPath_RF_bus_reg_dataout_852_port, 
                           regs(851) => DataPath_RF_bus_reg_dataout_851_port, 
                           regs(850) => DataPath_RF_bus_reg_dataout_850_port, 
                           regs(849) => DataPath_RF_bus_reg_dataout_849_port, 
                           regs(848) => DataPath_RF_bus_reg_dataout_848_port, 
                           regs(847) => DataPath_RF_bus_reg_dataout_847_port, 
                           regs(846) => DataPath_RF_bus_reg_dataout_846_port, 
                           regs(845) => DataPath_RF_bus_reg_dataout_845_port, 
                           regs(844) => DataPath_RF_bus_reg_dataout_844_port, 
                           regs(843) => DataPath_RF_bus_reg_dataout_843_port, 
                           regs(842) => DataPath_RF_bus_reg_dataout_842_port, 
                           regs(841) => DataPath_RF_bus_reg_dataout_841_port, 
                           regs(840) => DataPath_RF_bus_reg_dataout_840_port, 
                           regs(839) => DataPath_RF_bus_reg_dataout_839_port, 
                           regs(838) => DataPath_RF_bus_reg_dataout_838_port, 
                           regs(837) => DataPath_RF_bus_reg_dataout_837_port, 
                           regs(836) => DataPath_RF_bus_reg_dataout_836_port, 
                           regs(835) => DataPath_RF_bus_reg_dataout_835_port, 
                           regs(834) => DataPath_RF_bus_reg_dataout_834_port, 
                           regs(833) => DataPath_RF_bus_reg_dataout_833_port, 
                           regs(832) => DataPath_RF_bus_reg_dataout_832_port, 
                           regs(831) => DataPath_RF_bus_reg_dataout_831_port, 
                           regs(830) => DataPath_RF_bus_reg_dataout_830_port, 
                           regs(829) => DataPath_RF_bus_reg_dataout_829_port, 
                           regs(828) => DataPath_RF_bus_reg_dataout_828_port, 
                           regs(827) => DataPath_RF_bus_reg_dataout_827_port, 
                           regs(826) => DataPath_RF_bus_reg_dataout_826_port, 
                           regs(825) => DataPath_RF_bus_reg_dataout_825_port, 
                           regs(824) => DataPath_RF_bus_reg_dataout_824_port, 
                           regs(823) => DataPath_RF_bus_reg_dataout_823_port, 
                           regs(822) => DataPath_RF_bus_reg_dataout_822_port, 
                           regs(821) => DataPath_RF_bus_reg_dataout_821_port, 
                           regs(820) => DataPath_RF_bus_reg_dataout_820_port, 
                           regs(819) => DataPath_RF_bus_reg_dataout_819_port, 
                           regs(818) => DataPath_RF_bus_reg_dataout_818_port, 
                           regs(817) => DataPath_RF_bus_reg_dataout_817_port, 
                           regs(816) => DataPath_RF_bus_reg_dataout_816_port, 
                           regs(815) => DataPath_RF_bus_reg_dataout_815_port, 
                           regs(814) => DataPath_RF_bus_reg_dataout_814_port, 
                           regs(813) => DataPath_RF_bus_reg_dataout_813_port, 
                           regs(812) => DataPath_RF_bus_reg_dataout_812_port, 
                           regs(811) => DataPath_RF_bus_reg_dataout_811_port, 
                           regs(810) => DataPath_RF_bus_reg_dataout_810_port, 
                           regs(809) => DataPath_RF_bus_reg_dataout_809_port, 
                           regs(808) => DataPath_RF_bus_reg_dataout_808_port, 
                           regs(807) => DataPath_RF_bus_reg_dataout_807_port, 
                           regs(806) => DataPath_RF_bus_reg_dataout_806_port, 
                           regs(805) => DataPath_RF_bus_reg_dataout_805_port, 
                           regs(804) => DataPath_RF_bus_reg_dataout_804_port, 
                           regs(803) => DataPath_RF_bus_reg_dataout_803_port, 
                           regs(802) => DataPath_RF_bus_reg_dataout_802_port, 
                           regs(801) => DataPath_RF_bus_reg_dataout_801_port, 
                           regs(800) => DataPath_RF_bus_reg_dataout_800_port, 
                           regs(799) => DataPath_RF_bus_reg_dataout_799_port, 
                           regs(798) => DataPath_RF_bus_reg_dataout_798_port, 
                           regs(797) => DataPath_RF_bus_reg_dataout_797_port, 
                           regs(796) => DataPath_RF_bus_reg_dataout_796_port, 
                           regs(795) => DataPath_RF_bus_reg_dataout_795_port, 
                           regs(794) => DataPath_RF_bus_reg_dataout_794_port, 
                           regs(793) => DataPath_RF_bus_reg_dataout_793_port, 
                           regs(792) => DataPath_RF_bus_reg_dataout_792_port, 
                           regs(791) => DataPath_RF_bus_reg_dataout_791_port, 
                           regs(790) => DataPath_RF_bus_reg_dataout_790_port, 
                           regs(789) => DataPath_RF_bus_reg_dataout_789_port, 
                           regs(788) => DataPath_RF_bus_reg_dataout_788_port, 
                           regs(787) => DataPath_RF_bus_reg_dataout_787_port, 
                           regs(786) => DataPath_RF_bus_reg_dataout_786_port, 
                           regs(785) => DataPath_RF_bus_reg_dataout_785_port, 
                           regs(784) => DataPath_RF_bus_reg_dataout_784_port, 
                           regs(783) => DataPath_RF_bus_reg_dataout_783_port, 
                           regs(782) => DataPath_RF_bus_reg_dataout_782_port, 
                           regs(781) => DataPath_RF_bus_reg_dataout_781_port, 
                           regs(780) => DataPath_RF_bus_reg_dataout_780_port, 
                           regs(779) => DataPath_RF_bus_reg_dataout_779_port, 
                           regs(778) => DataPath_RF_bus_reg_dataout_778_port, 
                           regs(777) => DataPath_RF_bus_reg_dataout_777_port, 
                           regs(776) => DataPath_RF_bus_reg_dataout_776_port, 
                           regs(775) => DataPath_RF_bus_reg_dataout_775_port, 
                           regs(774) => DataPath_RF_bus_reg_dataout_774_port, 
                           regs(773) => DataPath_RF_bus_reg_dataout_773_port, 
                           regs(772) => DataPath_RF_bus_reg_dataout_772_port, 
                           regs(771) => DataPath_RF_bus_reg_dataout_771_port, 
                           regs(770) => DataPath_RF_bus_reg_dataout_770_port, 
                           regs(769) => DataPath_RF_bus_reg_dataout_769_port, 
                           regs(768) => DataPath_RF_bus_reg_dataout_768_port, 
                           regs(767) => DataPath_RF_bus_reg_dataout_767_port, 
                           regs(766) => DataPath_RF_bus_reg_dataout_766_port, 
                           regs(765) => DataPath_RF_bus_reg_dataout_765_port, 
                           regs(764) => DataPath_RF_bus_reg_dataout_764_port, 
                           regs(763) => DataPath_RF_bus_reg_dataout_763_port, 
                           regs(762) => DataPath_RF_bus_reg_dataout_762_port, 
                           regs(761) => DataPath_RF_bus_reg_dataout_761_port, 
                           regs(760) => DataPath_RF_bus_reg_dataout_760_port, 
                           regs(759) => DataPath_RF_bus_reg_dataout_759_port, 
                           regs(758) => DataPath_RF_bus_reg_dataout_758_port, 
                           regs(757) => DataPath_RF_bus_reg_dataout_757_port, 
                           regs(756) => DataPath_RF_bus_reg_dataout_756_port, 
                           regs(755) => DataPath_RF_bus_reg_dataout_755_port, 
                           regs(754) => DataPath_RF_bus_reg_dataout_754_port, 
                           regs(753) => DataPath_RF_bus_reg_dataout_753_port, 
                           regs(752) => DataPath_RF_bus_reg_dataout_752_port, 
                           regs(751) => DataPath_RF_bus_reg_dataout_751_port, 
                           regs(750) => DataPath_RF_bus_reg_dataout_750_port, 
                           regs(749) => DataPath_RF_bus_reg_dataout_749_port, 
                           regs(748) => DataPath_RF_bus_reg_dataout_748_port, 
                           regs(747) => DataPath_RF_bus_reg_dataout_747_port, 
                           regs(746) => DataPath_RF_bus_reg_dataout_746_port, 
                           regs(745) => DataPath_RF_bus_reg_dataout_745_port, 
                           regs(744) => DataPath_RF_bus_reg_dataout_744_port, 
                           regs(743) => DataPath_RF_bus_reg_dataout_743_port, 
                           regs(742) => DataPath_RF_bus_reg_dataout_742_port, 
                           regs(741) => DataPath_RF_bus_reg_dataout_741_port, 
                           regs(740) => DataPath_RF_bus_reg_dataout_740_port, 
                           regs(739) => DataPath_RF_bus_reg_dataout_739_port, 
                           regs(738) => DataPath_RF_bus_reg_dataout_738_port, 
                           regs(737) => DataPath_RF_bus_reg_dataout_737_port, 
                           regs(736) => DataPath_RF_bus_reg_dataout_736_port, 
                           regs(735) => DataPath_RF_bus_reg_dataout_735_port, 
                           regs(734) => DataPath_RF_bus_reg_dataout_734_port, 
                           regs(733) => DataPath_RF_bus_reg_dataout_733_port, 
                           regs(732) => DataPath_RF_bus_reg_dataout_732_port, 
                           regs(731) => DataPath_RF_bus_reg_dataout_731_port, 
                           regs(730) => DataPath_RF_bus_reg_dataout_730_port, 
                           regs(729) => DataPath_RF_bus_reg_dataout_729_port, 
                           regs(728) => DataPath_RF_bus_reg_dataout_728_port, 
                           regs(727) => DataPath_RF_bus_reg_dataout_727_port, 
                           regs(726) => DataPath_RF_bus_reg_dataout_726_port, 
                           regs(725) => DataPath_RF_bus_reg_dataout_725_port, 
                           regs(724) => DataPath_RF_bus_reg_dataout_724_port, 
                           regs(723) => DataPath_RF_bus_reg_dataout_723_port, 
                           regs(722) => DataPath_RF_bus_reg_dataout_722_port, 
                           regs(721) => DataPath_RF_bus_reg_dataout_721_port, 
                           regs(720) => DataPath_RF_bus_reg_dataout_720_port, 
                           regs(719) => DataPath_RF_bus_reg_dataout_719_port, 
                           regs(718) => DataPath_RF_bus_reg_dataout_718_port, 
                           regs(717) => DataPath_RF_bus_reg_dataout_717_port, 
                           regs(716) => DataPath_RF_bus_reg_dataout_716_port, 
                           regs(715) => DataPath_RF_bus_reg_dataout_715_port, 
                           regs(714) => DataPath_RF_bus_reg_dataout_714_port, 
                           regs(713) => DataPath_RF_bus_reg_dataout_713_port, 
                           regs(712) => DataPath_RF_bus_reg_dataout_712_port, 
                           regs(711) => DataPath_RF_bus_reg_dataout_711_port, 
                           regs(710) => DataPath_RF_bus_reg_dataout_710_port, 
                           regs(709) => DataPath_RF_bus_reg_dataout_709_port, 
                           regs(708) => DataPath_RF_bus_reg_dataout_708_port, 
                           regs(707) => DataPath_RF_bus_reg_dataout_707_port, 
                           regs(706) => DataPath_RF_bus_reg_dataout_706_port, 
                           regs(705) => DataPath_RF_bus_reg_dataout_705_port, 
                           regs(704) => DataPath_RF_bus_reg_dataout_704_port, 
                           regs(703) => DataPath_RF_bus_reg_dataout_703_port, 
                           regs(702) => DataPath_RF_bus_reg_dataout_702_port, 
                           regs(701) => DataPath_RF_bus_reg_dataout_701_port, 
                           regs(700) => DataPath_RF_bus_reg_dataout_700_port, 
                           regs(699) => DataPath_RF_bus_reg_dataout_699_port, 
                           regs(698) => DataPath_RF_bus_reg_dataout_698_port, 
                           regs(697) => DataPath_RF_bus_reg_dataout_697_port, 
                           regs(696) => DataPath_RF_bus_reg_dataout_696_port, 
                           regs(695) => DataPath_RF_bus_reg_dataout_695_port, 
                           regs(694) => DataPath_RF_bus_reg_dataout_694_port, 
                           regs(693) => DataPath_RF_bus_reg_dataout_693_port, 
                           regs(692) => DataPath_RF_bus_reg_dataout_692_port, 
                           regs(691) => DataPath_RF_bus_reg_dataout_691_port, 
                           regs(690) => DataPath_RF_bus_reg_dataout_690_port, 
                           regs(689) => DataPath_RF_bus_reg_dataout_689_port, 
                           regs(688) => DataPath_RF_bus_reg_dataout_688_port, 
                           regs(687) => DataPath_RF_bus_reg_dataout_687_port, 
                           regs(686) => DataPath_RF_bus_reg_dataout_686_port, 
                           regs(685) => DataPath_RF_bus_reg_dataout_685_port, 
                           regs(684) => DataPath_RF_bus_reg_dataout_684_port, 
                           regs(683) => DataPath_RF_bus_reg_dataout_683_port, 
                           regs(682) => DataPath_RF_bus_reg_dataout_682_port, 
                           regs(681) => DataPath_RF_bus_reg_dataout_681_port, 
                           regs(680) => DataPath_RF_bus_reg_dataout_680_port, 
                           regs(679) => DataPath_RF_bus_reg_dataout_679_port, 
                           regs(678) => DataPath_RF_bus_reg_dataout_678_port, 
                           regs(677) => DataPath_RF_bus_reg_dataout_677_port, 
                           regs(676) => DataPath_RF_bus_reg_dataout_676_port, 
                           regs(675) => DataPath_RF_bus_reg_dataout_675_port, 
                           regs(674) => DataPath_RF_bus_reg_dataout_674_port, 
                           regs(673) => DataPath_RF_bus_reg_dataout_673_port, 
                           regs(672) => DataPath_RF_bus_reg_dataout_672_port, 
                           regs(671) => DataPath_RF_bus_reg_dataout_671_port, 
                           regs(670) => DataPath_RF_bus_reg_dataout_670_port, 
                           regs(669) => DataPath_RF_bus_reg_dataout_669_port, 
                           regs(668) => DataPath_RF_bus_reg_dataout_668_port, 
                           regs(667) => DataPath_RF_bus_reg_dataout_667_port, 
                           regs(666) => DataPath_RF_bus_reg_dataout_666_port, 
                           regs(665) => DataPath_RF_bus_reg_dataout_665_port, 
                           regs(664) => DataPath_RF_bus_reg_dataout_664_port, 
                           regs(663) => DataPath_RF_bus_reg_dataout_663_port, 
                           regs(662) => DataPath_RF_bus_reg_dataout_662_port, 
                           regs(661) => DataPath_RF_bus_reg_dataout_661_port, 
                           regs(660) => DataPath_RF_bus_reg_dataout_660_port, 
                           regs(659) => DataPath_RF_bus_reg_dataout_659_port, 
                           regs(658) => DataPath_RF_bus_reg_dataout_658_port, 
                           regs(657) => DataPath_RF_bus_reg_dataout_657_port, 
                           regs(656) => DataPath_RF_bus_reg_dataout_656_port, 
                           regs(655) => DataPath_RF_bus_reg_dataout_655_port, 
                           regs(654) => DataPath_RF_bus_reg_dataout_654_port, 
                           regs(653) => DataPath_RF_bus_reg_dataout_653_port, 
                           regs(652) => DataPath_RF_bus_reg_dataout_652_port, 
                           regs(651) => DataPath_RF_bus_reg_dataout_651_port, 
                           regs(650) => DataPath_RF_bus_reg_dataout_650_port, 
                           regs(649) => DataPath_RF_bus_reg_dataout_649_port, 
                           regs(648) => DataPath_RF_bus_reg_dataout_648_port, 
                           regs(647) => DataPath_RF_bus_reg_dataout_647_port, 
                           regs(646) => DataPath_RF_bus_reg_dataout_646_port, 
                           regs(645) => DataPath_RF_bus_reg_dataout_645_port, 
                           regs(644) => DataPath_RF_bus_reg_dataout_644_port, 
                           regs(643) => DataPath_RF_bus_reg_dataout_643_port, 
                           regs(642) => DataPath_RF_bus_reg_dataout_642_port, 
                           regs(641) => DataPath_RF_bus_reg_dataout_641_port, 
                           regs(640) => DataPath_RF_bus_reg_dataout_640_port, 
                           regs(639) => DataPath_RF_bus_reg_dataout_639_port, 
                           regs(638) => DataPath_RF_bus_reg_dataout_638_port, 
                           regs(637) => DataPath_RF_bus_reg_dataout_637_port, 
                           regs(636) => DataPath_RF_bus_reg_dataout_636_port, 
                           regs(635) => DataPath_RF_bus_reg_dataout_635_port, 
                           regs(634) => DataPath_RF_bus_reg_dataout_634_port, 
                           regs(633) => DataPath_RF_bus_reg_dataout_633_port, 
                           regs(632) => DataPath_RF_bus_reg_dataout_632_port, 
                           regs(631) => DataPath_RF_bus_reg_dataout_631_port, 
                           regs(630) => DataPath_RF_bus_reg_dataout_630_port, 
                           regs(629) => DataPath_RF_bus_reg_dataout_629_port, 
                           regs(628) => DataPath_RF_bus_reg_dataout_628_port, 
                           regs(627) => DataPath_RF_bus_reg_dataout_627_port, 
                           regs(626) => DataPath_RF_bus_reg_dataout_626_port, 
                           regs(625) => DataPath_RF_bus_reg_dataout_625_port, 
                           regs(624) => DataPath_RF_bus_reg_dataout_624_port, 
                           regs(623) => DataPath_RF_bus_reg_dataout_623_port, 
                           regs(622) => DataPath_RF_bus_reg_dataout_622_port, 
                           regs(621) => DataPath_RF_bus_reg_dataout_621_port, 
                           regs(620) => DataPath_RF_bus_reg_dataout_620_port, 
                           regs(619) => DataPath_RF_bus_reg_dataout_619_port, 
                           regs(618) => DataPath_RF_bus_reg_dataout_618_port, 
                           regs(617) => DataPath_RF_bus_reg_dataout_617_port, 
                           regs(616) => DataPath_RF_bus_reg_dataout_616_port, 
                           regs(615) => DataPath_RF_bus_reg_dataout_615_port, 
                           regs(614) => DataPath_RF_bus_reg_dataout_614_port, 
                           regs(613) => DataPath_RF_bus_reg_dataout_613_port, 
                           regs(612) => DataPath_RF_bus_reg_dataout_612_port, 
                           regs(611) => DataPath_RF_bus_reg_dataout_611_port, 
                           regs(610) => DataPath_RF_bus_reg_dataout_610_port, 
                           regs(609) => DataPath_RF_bus_reg_dataout_609_port, 
                           regs(608) => DataPath_RF_bus_reg_dataout_608_port, 
                           regs(607) => DataPath_RF_bus_reg_dataout_607_port, 
                           regs(606) => DataPath_RF_bus_reg_dataout_606_port, 
                           regs(605) => DataPath_RF_bus_reg_dataout_605_port, 
                           regs(604) => DataPath_RF_bus_reg_dataout_604_port, 
                           regs(603) => DataPath_RF_bus_reg_dataout_603_port, 
                           regs(602) => DataPath_RF_bus_reg_dataout_602_port, 
                           regs(601) => DataPath_RF_bus_reg_dataout_601_port, 
                           regs(600) => DataPath_RF_bus_reg_dataout_600_port, 
                           regs(599) => DataPath_RF_bus_reg_dataout_599_port, 
                           regs(598) => DataPath_RF_bus_reg_dataout_598_port, 
                           regs(597) => DataPath_RF_bus_reg_dataout_597_port, 
                           regs(596) => DataPath_RF_bus_reg_dataout_596_port, 
                           regs(595) => DataPath_RF_bus_reg_dataout_595_port, 
                           regs(594) => DataPath_RF_bus_reg_dataout_594_port, 
                           regs(593) => DataPath_RF_bus_reg_dataout_593_port, 
                           regs(592) => DataPath_RF_bus_reg_dataout_592_port, 
                           regs(591) => DataPath_RF_bus_reg_dataout_591_port, 
                           regs(590) => DataPath_RF_bus_reg_dataout_590_port, 
                           regs(589) => DataPath_RF_bus_reg_dataout_589_port, 
                           regs(588) => DataPath_RF_bus_reg_dataout_588_port, 
                           regs(587) => DataPath_RF_bus_reg_dataout_587_port, 
                           regs(586) => DataPath_RF_bus_reg_dataout_586_port, 
                           regs(585) => DataPath_RF_bus_reg_dataout_585_port, 
                           regs(584) => DataPath_RF_bus_reg_dataout_584_port, 
                           regs(583) => DataPath_RF_bus_reg_dataout_583_port, 
                           regs(582) => DataPath_RF_bus_reg_dataout_582_port, 
                           regs(581) => DataPath_RF_bus_reg_dataout_581_port, 
                           regs(580) => DataPath_RF_bus_reg_dataout_580_port, 
                           regs(579) => DataPath_RF_bus_reg_dataout_579_port, 
                           regs(578) => DataPath_RF_bus_reg_dataout_578_port, 
                           regs(577) => DataPath_RF_bus_reg_dataout_577_port, 
                           regs(576) => DataPath_RF_bus_reg_dataout_576_port, 
                           regs(575) => DataPath_RF_bus_reg_dataout_575_port, 
                           regs(574) => DataPath_RF_bus_reg_dataout_574_port, 
                           regs(573) => DataPath_RF_bus_reg_dataout_573_port, 
                           regs(572) => DataPath_RF_bus_reg_dataout_572_port, 
                           regs(571) => DataPath_RF_bus_reg_dataout_571_port, 
                           regs(570) => DataPath_RF_bus_reg_dataout_570_port, 
                           regs(569) => DataPath_RF_bus_reg_dataout_569_port, 
                           regs(568) => DataPath_RF_bus_reg_dataout_568_port, 
                           regs(567) => DataPath_RF_bus_reg_dataout_567_port, 
                           regs(566) => DataPath_RF_bus_reg_dataout_566_port, 
                           regs(565) => DataPath_RF_bus_reg_dataout_565_port, 
                           regs(564) => DataPath_RF_bus_reg_dataout_564_port, 
                           regs(563) => DataPath_RF_bus_reg_dataout_563_port, 
                           regs(562) => DataPath_RF_bus_reg_dataout_562_port, 
                           regs(561) => DataPath_RF_bus_reg_dataout_561_port, 
                           regs(560) => DataPath_RF_bus_reg_dataout_560_port, 
                           regs(559) => DataPath_RF_bus_reg_dataout_559_port, 
                           regs(558) => DataPath_RF_bus_reg_dataout_558_port, 
                           regs(557) => DataPath_RF_bus_reg_dataout_557_port, 
                           regs(556) => DataPath_RF_bus_reg_dataout_556_port, 
                           regs(555) => DataPath_RF_bus_reg_dataout_555_port, 
                           regs(554) => DataPath_RF_bus_reg_dataout_554_port, 
                           regs(553) => DataPath_RF_bus_reg_dataout_553_port, 
                           regs(552) => DataPath_RF_bus_reg_dataout_552_port, 
                           regs(551) => DataPath_RF_bus_reg_dataout_551_port, 
                           regs(550) => DataPath_RF_bus_reg_dataout_550_port, 
                           regs(549) => DataPath_RF_bus_reg_dataout_549_port, 
                           regs(548) => DataPath_RF_bus_reg_dataout_548_port, 
                           regs(547) => DataPath_RF_bus_reg_dataout_547_port, 
                           regs(546) => DataPath_RF_bus_reg_dataout_546_port, 
                           regs(545) => DataPath_RF_bus_reg_dataout_545_port, 
                           regs(544) => DataPath_RF_bus_reg_dataout_544_port, 
                           regs(543) => DataPath_RF_bus_reg_dataout_543_port, 
                           regs(542) => DataPath_RF_bus_reg_dataout_542_port, 
                           regs(541) => DataPath_RF_bus_reg_dataout_541_port, 
                           regs(540) => DataPath_RF_bus_reg_dataout_540_port, 
                           regs(539) => DataPath_RF_bus_reg_dataout_539_port, 
                           regs(538) => DataPath_RF_bus_reg_dataout_538_port, 
                           regs(537) => DataPath_RF_bus_reg_dataout_537_port, 
                           regs(536) => DataPath_RF_bus_reg_dataout_536_port, 
                           regs(535) => DataPath_RF_bus_reg_dataout_535_port, 
                           regs(534) => DataPath_RF_bus_reg_dataout_534_port, 
                           regs(533) => DataPath_RF_bus_reg_dataout_533_port, 
                           regs(532) => DataPath_RF_bus_reg_dataout_532_port, 
                           regs(531) => DataPath_RF_bus_reg_dataout_531_port, 
                           regs(530) => DataPath_RF_bus_reg_dataout_530_port, 
                           regs(529) => DataPath_RF_bus_reg_dataout_529_port, 
                           regs(528) => DataPath_RF_bus_reg_dataout_528_port, 
                           regs(527) => DataPath_RF_bus_reg_dataout_527_port, 
                           regs(526) => DataPath_RF_bus_reg_dataout_526_port, 
                           regs(525) => DataPath_RF_bus_reg_dataout_525_port, 
                           regs(524) => DataPath_RF_bus_reg_dataout_524_port, 
                           regs(523) => DataPath_RF_bus_reg_dataout_523_port, 
                           regs(522) => DataPath_RF_bus_reg_dataout_522_port, 
                           regs(521) => DataPath_RF_bus_reg_dataout_521_port, 
                           regs(520) => DataPath_RF_bus_reg_dataout_520_port, 
                           regs(519) => DataPath_RF_bus_reg_dataout_519_port, 
                           regs(518) => DataPath_RF_bus_reg_dataout_518_port, 
                           regs(517) => DataPath_RF_bus_reg_dataout_517_port, 
                           regs(516) => DataPath_RF_bus_reg_dataout_516_port, 
                           regs(515) => DataPath_RF_bus_reg_dataout_515_port, 
                           regs(514) => DataPath_RF_bus_reg_dataout_514_port, 
                           regs(513) => DataPath_RF_bus_reg_dataout_513_port, 
                           regs(512) => DataPath_RF_bus_reg_dataout_512_port, 
                           regs(511) => DataPath_RF_bus_reg_dataout_511_port, 
                           regs(510) => DataPath_RF_bus_reg_dataout_510_port, 
                           regs(509) => DataPath_RF_bus_reg_dataout_509_port, 
                           regs(508) => DataPath_RF_bus_reg_dataout_508_port, 
                           regs(507) => DataPath_RF_bus_reg_dataout_507_port, 
                           regs(506) => DataPath_RF_bus_reg_dataout_506_port, 
                           regs(505) => DataPath_RF_bus_reg_dataout_505_port, 
                           regs(504) => DataPath_RF_bus_reg_dataout_504_port, 
                           regs(503) => DataPath_RF_bus_reg_dataout_503_port, 
                           regs(502) => DataPath_RF_bus_reg_dataout_502_port, 
                           regs(501) => DataPath_RF_bus_reg_dataout_501_port, 
                           regs(500) => DataPath_RF_bus_reg_dataout_500_port, 
                           regs(499) => DataPath_RF_bus_reg_dataout_499_port, 
                           regs(498) => DataPath_RF_bus_reg_dataout_498_port, 
                           regs(497) => DataPath_RF_bus_reg_dataout_497_port, 
                           regs(496) => DataPath_RF_bus_reg_dataout_496_port, 
                           regs(495) => DataPath_RF_bus_reg_dataout_495_port, 
                           regs(494) => DataPath_RF_bus_reg_dataout_494_port, 
                           regs(493) => DataPath_RF_bus_reg_dataout_493_port, 
                           regs(492) => DataPath_RF_bus_reg_dataout_492_port, 
                           regs(491) => DataPath_RF_bus_reg_dataout_491_port, 
                           regs(490) => DataPath_RF_bus_reg_dataout_490_port, 
                           regs(489) => DataPath_RF_bus_reg_dataout_489_port, 
                           regs(488) => DataPath_RF_bus_reg_dataout_488_port, 
                           regs(487) => DataPath_RF_bus_reg_dataout_487_port, 
                           regs(486) => DataPath_RF_bus_reg_dataout_486_port, 
                           regs(485) => DataPath_RF_bus_reg_dataout_485_port, 
                           regs(484) => DataPath_RF_bus_reg_dataout_484_port, 
                           regs(483) => DataPath_RF_bus_reg_dataout_483_port, 
                           regs(482) => DataPath_RF_bus_reg_dataout_482_port, 
                           regs(481) => DataPath_RF_bus_reg_dataout_481_port, 
                           regs(480) => DataPath_RF_bus_reg_dataout_480_port, 
                           regs(479) => DataPath_RF_bus_reg_dataout_479_port, 
                           regs(478) => DataPath_RF_bus_reg_dataout_478_port, 
                           regs(477) => DataPath_RF_bus_reg_dataout_477_port, 
                           regs(476) => DataPath_RF_bus_reg_dataout_476_port, 
                           regs(475) => DataPath_RF_bus_reg_dataout_475_port, 
                           regs(474) => DataPath_RF_bus_reg_dataout_474_port, 
                           regs(473) => DataPath_RF_bus_reg_dataout_473_port, 
                           regs(472) => DataPath_RF_bus_reg_dataout_472_port, 
                           regs(471) => DataPath_RF_bus_reg_dataout_471_port, 
                           regs(470) => DataPath_RF_bus_reg_dataout_470_port, 
                           regs(469) => DataPath_RF_bus_reg_dataout_469_port, 
                           regs(468) => DataPath_RF_bus_reg_dataout_468_port, 
                           regs(467) => DataPath_RF_bus_reg_dataout_467_port, 
                           regs(466) => DataPath_RF_bus_reg_dataout_466_port, 
                           regs(465) => DataPath_RF_bus_reg_dataout_465_port, 
                           regs(464) => DataPath_RF_bus_reg_dataout_464_port, 
                           regs(463) => DataPath_RF_bus_reg_dataout_463_port, 
                           regs(462) => DataPath_RF_bus_reg_dataout_462_port, 
                           regs(461) => DataPath_RF_bus_reg_dataout_461_port, 
                           regs(460) => DataPath_RF_bus_reg_dataout_460_port, 
                           regs(459) => DataPath_RF_bus_reg_dataout_459_port, 
                           regs(458) => DataPath_RF_bus_reg_dataout_458_port, 
                           regs(457) => DataPath_RF_bus_reg_dataout_457_port, 
                           regs(456) => DataPath_RF_bus_reg_dataout_456_port, 
                           regs(455) => DataPath_RF_bus_reg_dataout_455_port, 
                           regs(454) => DataPath_RF_bus_reg_dataout_454_port, 
                           regs(453) => DataPath_RF_bus_reg_dataout_453_port, 
                           regs(452) => DataPath_RF_bus_reg_dataout_452_port, 
                           regs(451) => DataPath_RF_bus_reg_dataout_451_port, 
                           regs(450) => DataPath_RF_bus_reg_dataout_450_port, 
                           regs(449) => DataPath_RF_bus_reg_dataout_449_port, 
                           regs(448) => DataPath_RF_bus_reg_dataout_448_port, 
                           regs(447) => DataPath_RF_bus_reg_dataout_447_port, 
                           regs(446) => DataPath_RF_bus_reg_dataout_446_port, 
                           regs(445) => DataPath_RF_bus_reg_dataout_445_port, 
                           regs(444) => DataPath_RF_bus_reg_dataout_444_port, 
                           regs(443) => DataPath_RF_bus_reg_dataout_443_port, 
                           regs(442) => DataPath_RF_bus_reg_dataout_442_port, 
                           regs(441) => DataPath_RF_bus_reg_dataout_441_port, 
                           regs(440) => DataPath_RF_bus_reg_dataout_440_port, 
                           regs(439) => DataPath_RF_bus_reg_dataout_439_port, 
                           regs(438) => DataPath_RF_bus_reg_dataout_438_port, 
                           regs(437) => DataPath_RF_bus_reg_dataout_437_port, 
                           regs(436) => DataPath_RF_bus_reg_dataout_436_port, 
                           regs(435) => DataPath_RF_bus_reg_dataout_435_port, 
                           regs(434) => DataPath_RF_bus_reg_dataout_434_port, 
                           regs(433) => DataPath_RF_bus_reg_dataout_433_port, 
                           regs(432) => DataPath_RF_bus_reg_dataout_432_port, 
                           regs(431) => DataPath_RF_bus_reg_dataout_431_port, 
                           regs(430) => DataPath_RF_bus_reg_dataout_430_port, 
                           regs(429) => DataPath_RF_bus_reg_dataout_429_port, 
                           regs(428) => DataPath_RF_bus_reg_dataout_428_port, 
                           regs(427) => DataPath_RF_bus_reg_dataout_427_port, 
                           regs(426) => DataPath_RF_bus_reg_dataout_426_port, 
                           regs(425) => DataPath_RF_bus_reg_dataout_425_port, 
                           regs(424) => DataPath_RF_bus_reg_dataout_424_port, 
                           regs(423) => DataPath_RF_bus_reg_dataout_423_port, 
                           regs(422) => DataPath_RF_bus_reg_dataout_422_port, 
                           regs(421) => DataPath_RF_bus_reg_dataout_421_port, 
                           regs(420) => DataPath_RF_bus_reg_dataout_420_port, 
                           regs(419) => DataPath_RF_bus_reg_dataout_419_port, 
                           regs(418) => DataPath_RF_bus_reg_dataout_418_port, 
                           regs(417) => DataPath_RF_bus_reg_dataout_417_port, 
                           regs(416) => DataPath_RF_bus_reg_dataout_416_port, 
                           regs(415) => DataPath_RF_bus_reg_dataout_415_port, 
                           regs(414) => DataPath_RF_bus_reg_dataout_414_port, 
                           regs(413) => DataPath_RF_bus_reg_dataout_413_port, 
                           regs(412) => DataPath_RF_bus_reg_dataout_412_port, 
                           regs(411) => DataPath_RF_bus_reg_dataout_411_port, 
                           regs(410) => DataPath_RF_bus_reg_dataout_410_port, 
                           regs(409) => DataPath_RF_bus_reg_dataout_409_port, 
                           regs(408) => DataPath_RF_bus_reg_dataout_408_port, 
                           regs(407) => DataPath_RF_bus_reg_dataout_407_port, 
                           regs(406) => DataPath_RF_bus_reg_dataout_406_port, 
                           regs(405) => DataPath_RF_bus_reg_dataout_405_port, 
                           regs(404) => DataPath_RF_bus_reg_dataout_404_port, 
                           regs(403) => DataPath_RF_bus_reg_dataout_403_port, 
                           regs(402) => DataPath_RF_bus_reg_dataout_402_port, 
                           regs(401) => DataPath_RF_bus_reg_dataout_401_port, 
                           regs(400) => DataPath_RF_bus_reg_dataout_400_port, 
                           regs(399) => DataPath_RF_bus_reg_dataout_399_port, 
                           regs(398) => DataPath_RF_bus_reg_dataout_398_port, 
                           regs(397) => DataPath_RF_bus_reg_dataout_397_port, 
                           regs(396) => DataPath_RF_bus_reg_dataout_396_port, 
                           regs(395) => DataPath_RF_bus_reg_dataout_395_port, 
                           regs(394) => DataPath_RF_bus_reg_dataout_394_port, 
                           regs(393) => DataPath_RF_bus_reg_dataout_393_port, 
                           regs(392) => DataPath_RF_bus_reg_dataout_392_port, 
                           regs(391) => DataPath_RF_bus_reg_dataout_391_port, 
                           regs(390) => DataPath_RF_bus_reg_dataout_390_port, 
                           regs(389) => DataPath_RF_bus_reg_dataout_389_port, 
                           regs(388) => DataPath_RF_bus_reg_dataout_388_port, 
                           regs(387) => DataPath_RF_bus_reg_dataout_387_port, 
                           regs(386) => DataPath_RF_bus_reg_dataout_386_port, 
                           regs(385) => DataPath_RF_bus_reg_dataout_385_port, 
                           regs(384) => DataPath_RF_bus_reg_dataout_384_port, 
                           regs(383) => DataPath_RF_bus_reg_dataout_383_port, 
                           regs(382) => DataPath_RF_bus_reg_dataout_382_port, 
                           regs(381) => DataPath_RF_bus_reg_dataout_381_port, 
                           regs(380) => DataPath_RF_bus_reg_dataout_380_port, 
                           regs(379) => DataPath_RF_bus_reg_dataout_379_port, 
                           regs(378) => DataPath_RF_bus_reg_dataout_378_port, 
                           regs(377) => DataPath_RF_bus_reg_dataout_377_port, 
                           regs(376) => DataPath_RF_bus_reg_dataout_376_port, 
                           regs(375) => DataPath_RF_bus_reg_dataout_375_port, 
                           regs(374) => DataPath_RF_bus_reg_dataout_374_port, 
                           regs(373) => DataPath_RF_bus_reg_dataout_373_port, 
                           regs(372) => DataPath_RF_bus_reg_dataout_372_port, 
                           regs(371) => DataPath_RF_bus_reg_dataout_371_port, 
                           regs(370) => DataPath_RF_bus_reg_dataout_370_port, 
                           regs(369) => DataPath_RF_bus_reg_dataout_369_port, 
                           regs(368) => DataPath_RF_bus_reg_dataout_368_port, 
                           regs(367) => DataPath_RF_bus_reg_dataout_367_port, 
                           regs(366) => DataPath_RF_bus_reg_dataout_366_port, 
                           regs(365) => DataPath_RF_bus_reg_dataout_365_port, 
                           regs(364) => DataPath_RF_bus_reg_dataout_364_port, 
                           regs(363) => DataPath_RF_bus_reg_dataout_363_port, 
                           regs(362) => DataPath_RF_bus_reg_dataout_362_port, 
                           regs(361) => DataPath_RF_bus_reg_dataout_361_port, 
                           regs(360) => DataPath_RF_bus_reg_dataout_360_port, 
                           regs(359) => DataPath_RF_bus_reg_dataout_359_port, 
                           regs(358) => DataPath_RF_bus_reg_dataout_358_port, 
                           regs(357) => DataPath_RF_bus_reg_dataout_357_port, 
                           regs(356) => DataPath_RF_bus_reg_dataout_356_port, 
                           regs(355) => DataPath_RF_bus_reg_dataout_355_port, 
                           regs(354) => DataPath_RF_bus_reg_dataout_354_port, 
                           regs(353) => DataPath_RF_bus_reg_dataout_353_port, 
                           regs(352) => DataPath_RF_bus_reg_dataout_352_port, 
                           regs(351) => DataPath_RF_bus_reg_dataout_351_port, 
                           regs(350) => DataPath_RF_bus_reg_dataout_350_port, 
                           regs(349) => DataPath_RF_bus_reg_dataout_349_port, 
                           regs(348) => DataPath_RF_bus_reg_dataout_348_port, 
                           regs(347) => DataPath_RF_bus_reg_dataout_347_port, 
                           regs(346) => DataPath_RF_bus_reg_dataout_346_port, 
                           regs(345) => DataPath_RF_bus_reg_dataout_345_port, 
                           regs(344) => DataPath_RF_bus_reg_dataout_344_port, 
                           regs(343) => DataPath_RF_bus_reg_dataout_343_port, 
                           regs(342) => DataPath_RF_bus_reg_dataout_342_port, 
                           regs(341) => DataPath_RF_bus_reg_dataout_341_port, 
                           regs(340) => DataPath_RF_bus_reg_dataout_340_port, 
                           regs(339) => DataPath_RF_bus_reg_dataout_339_port, 
                           regs(338) => DataPath_RF_bus_reg_dataout_338_port, 
                           regs(337) => DataPath_RF_bus_reg_dataout_337_port, 
                           regs(336) => DataPath_RF_bus_reg_dataout_336_port, 
                           regs(335) => DataPath_RF_bus_reg_dataout_335_port, 
                           regs(334) => DataPath_RF_bus_reg_dataout_334_port, 
                           regs(333) => DataPath_RF_bus_reg_dataout_333_port, 
                           regs(332) => DataPath_RF_bus_reg_dataout_332_port, 
                           regs(331) => DataPath_RF_bus_reg_dataout_331_port, 
                           regs(330) => DataPath_RF_bus_reg_dataout_330_port, 
                           regs(329) => DataPath_RF_bus_reg_dataout_329_port, 
                           regs(328) => DataPath_RF_bus_reg_dataout_328_port, 
                           regs(327) => DataPath_RF_bus_reg_dataout_327_port, 
                           regs(326) => DataPath_RF_bus_reg_dataout_326_port, 
                           regs(325) => DataPath_RF_bus_reg_dataout_325_port, 
                           regs(324) => DataPath_RF_bus_reg_dataout_324_port, 
                           regs(323) => DataPath_RF_bus_reg_dataout_323_port, 
                           regs(322) => DataPath_RF_bus_reg_dataout_322_port, 
                           regs(321) => DataPath_RF_bus_reg_dataout_321_port, 
                           regs(320) => DataPath_RF_bus_reg_dataout_320_port, 
                           regs(319) => DataPath_RF_bus_reg_dataout_319_port, 
                           regs(318) => DataPath_RF_bus_reg_dataout_318_port, 
                           regs(317) => DataPath_RF_bus_reg_dataout_317_port, 
                           regs(316) => DataPath_RF_bus_reg_dataout_316_port, 
                           regs(315) => DataPath_RF_bus_reg_dataout_315_port, 
                           regs(314) => DataPath_RF_bus_reg_dataout_314_port, 
                           regs(313) => DataPath_RF_bus_reg_dataout_313_port, 
                           regs(312) => DataPath_RF_bus_reg_dataout_312_port, 
                           regs(311) => DataPath_RF_bus_reg_dataout_311_port, 
                           regs(310) => DataPath_RF_bus_reg_dataout_310_port, 
                           regs(309) => DataPath_RF_bus_reg_dataout_309_port, 
                           regs(308) => DataPath_RF_bus_reg_dataout_308_port, 
                           regs(307) => DataPath_RF_bus_reg_dataout_307_port, 
                           regs(306) => DataPath_RF_bus_reg_dataout_306_port, 
                           regs(305) => DataPath_RF_bus_reg_dataout_305_port, 
                           regs(304) => DataPath_RF_bus_reg_dataout_304_port, 
                           regs(303) => DataPath_RF_bus_reg_dataout_303_port, 
                           regs(302) => DataPath_RF_bus_reg_dataout_302_port, 
                           regs(301) => DataPath_RF_bus_reg_dataout_301_port, 
                           regs(300) => DataPath_RF_bus_reg_dataout_300_port, 
                           regs(299) => DataPath_RF_bus_reg_dataout_299_port, 
                           regs(298) => DataPath_RF_bus_reg_dataout_298_port, 
                           regs(297) => DataPath_RF_bus_reg_dataout_297_port, 
                           regs(296) => DataPath_RF_bus_reg_dataout_296_port, 
                           regs(295) => DataPath_RF_bus_reg_dataout_295_port, 
                           regs(294) => DataPath_RF_bus_reg_dataout_294_port, 
                           regs(293) => DataPath_RF_bus_reg_dataout_293_port, 
                           regs(292) => DataPath_RF_bus_reg_dataout_292_port, 
                           regs(291) => DataPath_RF_bus_reg_dataout_291_port, 
                           regs(290) => DataPath_RF_bus_reg_dataout_290_port, 
                           regs(289) => DataPath_RF_bus_reg_dataout_289_port, 
                           regs(288) => DataPath_RF_bus_reg_dataout_288_port, 
                           regs(287) => DataPath_RF_bus_reg_dataout_287_port, 
                           regs(286) => DataPath_RF_bus_reg_dataout_286_port, 
                           regs(285) => DataPath_RF_bus_reg_dataout_285_port, 
                           regs(284) => DataPath_RF_bus_reg_dataout_284_port, 
                           regs(283) => DataPath_RF_bus_reg_dataout_283_port, 
                           regs(282) => DataPath_RF_bus_reg_dataout_282_port, 
                           regs(281) => DataPath_RF_bus_reg_dataout_281_port, 
                           regs(280) => DataPath_RF_bus_reg_dataout_280_port, 
                           regs(279) => DataPath_RF_bus_reg_dataout_279_port, 
                           regs(278) => DataPath_RF_bus_reg_dataout_278_port, 
                           regs(277) => DataPath_RF_bus_reg_dataout_277_port, 
                           regs(276) => DataPath_RF_bus_reg_dataout_276_port, 
                           regs(275) => DataPath_RF_bus_reg_dataout_275_port, 
                           regs(274) => DataPath_RF_bus_reg_dataout_274_port, 
                           regs(273) => DataPath_RF_bus_reg_dataout_273_port, 
                           regs(272) => DataPath_RF_bus_reg_dataout_272_port, 
                           regs(271) => DataPath_RF_bus_reg_dataout_271_port, 
                           regs(270) => DataPath_RF_bus_reg_dataout_270_port, 
                           regs(269) => DataPath_RF_bus_reg_dataout_269_port, 
                           regs(268) => DataPath_RF_bus_reg_dataout_268_port, 
                           regs(267) => DataPath_RF_bus_reg_dataout_267_port, 
                           regs(266) => DataPath_RF_bus_reg_dataout_266_port, 
                           regs(265) => DataPath_RF_bus_reg_dataout_265_port, 
                           regs(264) => DataPath_RF_bus_reg_dataout_264_port, 
                           regs(263) => DataPath_RF_bus_reg_dataout_263_port, 
                           regs(262) => DataPath_RF_bus_reg_dataout_262_port, 
                           regs(261) => DataPath_RF_bus_reg_dataout_261_port, 
                           regs(260) => DataPath_RF_bus_reg_dataout_260_port, 
                           regs(259) => DataPath_RF_bus_reg_dataout_259_port, 
                           regs(258) => DataPath_RF_bus_reg_dataout_258_port, 
                           regs(257) => DataPath_RF_bus_reg_dataout_257_port, 
                           regs(256) => DataPath_RF_bus_reg_dataout_256_port, 
                           regs(255) => DataPath_RF_bus_reg_dataout_255_port, 
                           regs(254) => DataPath_RF_bus_reg_dataout_254_port, 
                           regs(253) => DataPath_RF_bus_reg_dataout_253_port, 
                           regs(252) => DataPath_RF_bus_reg_dataout_252_port, 
                           regs(251) => DataPath_RF_bus_reg_dataout_251_port, 
                           regs(250) => DataPath_RF_bus_reg_dataout_250_port, 
                           regs(249) => DataPath_RF_bus_reg_dataout_249_port, 
                           regs(248) => DataPath_RF_bus_reg_dataout_248_port, 
                           regs(247) => DataPath_RF_bus_reg_dataout_247_port, 
                           regs(246) => DataPath_RF_bus_reg_dataout_246_port, 
                           regs(245) => DataPath_RF_bus_reg_dataout_245_port, 
                           regs(244) => DataPath_RF_bus_reg_dataout_244_port, 
                           regs(243) => DataPath_RF_bus_reg_dataout_243_port, 
                           regs(242) => DataPath_RF_bus_reg_dataout_242_port, 
                           regs(241) => DataPath_RF_bus_reg_dataout_241_port, 
                           regs(240) => DataPath_RF_bus_reg_dataout_240_port, 
                           regs(239) => DataPath_RF_bus_reg_dataout_239_port, 
                           regs(238) => DataPath_RF_bus_reg_dataout_238_port, 
                           regs(237) => DataPath_RF_bus_reg_dataout_237_port, 
                           regs(236) => DataPath_RF_bus_reg_dataout_236_port, 
                           regs(235) => DataPath_RF_bus_reg_dataout_235_port, 
                           regs(234) => DataPath_RF_bus_reg_dataout_234_port, 
                           regs(233) => DataPath_RF_bus_reg_dataout_233_port, 
                           regs(232) => DataPath_RF_bus_reg_dataout_232_port, 
                           regs(231) => DataPath_RF_bus_reg_dataout_231_port, 
                           regs(230) => DataPath_RF_bus_reg_dataout_230_port, 
                           regs(229) => DataPath_RF_bus_reg_dataout_229_port, 
                           regs(228) => DataPath_RF_bus_reg_dataout_228_port, 
                           regs(227) => DataPath_RF_bus_reg_dataout_227_port, 
                           regs(226) => DataPath_RF_bus_reg_dataout_226_port, 
                           regs(225) => DataPath_RF_bus_reg_dataout_225_port, 
                           regs(224) => DataPath_RF_bus_reg_dataout_224_port, 
                           regs(223) => DataPath_RF_bus_reg_dataout_223_port, 
                           regs(222) => DataPath_RF_bus_reg_dataout_222_port, 
                           regs(221) => DataPath_RF_bus_reg_dataout_221_port, 
                           regs(220) => DataPath_RF_bus_reg_dataout_220_port, 
                           regs(219) => DataPath_RF_bus_reg_dataout_219_port, 
                           regs(218) => DataPath_RF_bus_reg_dataout_218_port, 
                           regs(217) => DataPath_RF_bus_reg_dataout_217_port, 
                           regs(216) => DataPath_RF_bus_reg_dataout_216_port, 
                           regs(215) => DataPath_RF_bus_reg_dataout_215_port, 
                           regs(214) => DataPath_RF_bus_reg_dataout_214_port, 
                           regs(213) => DataPath_RF_bus_reg_dataout_213_port, 
                           regs(212) => DataPath_RF_bus_reg_dataout_212_port, 
                           regs(211) => DataPath_RF_bus_reg_dataout_211_port, 
                           regs(210) => DataPath_RF_bus_reg_dataout_210_port, 
                           regs(209) => DataPath_RF_bus_reg_dataout_209_port, 
                           regs(208) => DataPath_RF_bus_reg_dataout_208_port, 
                           regs(207) => DataPath_RF_bus_reg_dataout_207_port, 
                           regs(206) => DataPath_RF_bus_reg_dataout_206_port, 
                           regs(205) => DataPath_RF_bus_reg_dataout_205_port, 
                           regs(204) => DataPath_RF_bus_reg_dataout_204_port, 
                           regs(203) => DataPath_RF_bus_reg_dataout_203_port, 
                           regs(202) => DataPath_RF_bus_reg_dataout_202_port, 
                           regs(201) => DataPath_RF_bus_reg_dataout_201_port, 
                           regs(200) => DataPath_RF_bus_reg_dataout_200_port, 
                           regs(199) => DataPath_RF_bus_reg_dataout_199_port, 
                           regs(198) => DataPath_RF_bus_reg_dataout_198_port, 
                           regs(197) => DataPath_RF_bus_reg_dataout_197_port, 
                           regs(196) => DataPath_RF_bus_reg_dataout_196_port, 
                           regs(195) => DataPath_RF_bus_reg_dataout_195_port, 
                           regs(194) => DataPath_RF_bus_reg_dataout_194_port, 
                           regs(193) => DataPath_RF_bus_reg_dataout_193_port, 
                           regs(192) => DataPath_RF_bus_reg_dataout_192_port, 
                           regs(191) => DataPath_RF_bus_reg_dataout_191_port, 
                           regs(190) => DataPath_RF_bus_reg_dataout_190_port, 
                           regs(189) => DataPath_RF_bus_reg_dataout_189_port, 
                           regs(188) => DataPath_RF_bus_reg_dataout_188_port, 
                           regs(187) => DataPath_RF_bus_reg_dataout_187_port, 
                           regs(186) => DataPath_RF_bus_reg_dataout_186_port, 
                           regs(185) => DataPath_RF_bus_reg_dataout_185_port, 
                           regs(184) => DataPath_RF_bus_reg_dataout_184_port, 
                           regs(183) => DataPath_RF_bus_reg_dataout_183_port, 
                           regs(182) => DataPath_RF_bus_reg_dataout_182_port, 
                           regs(181) => DataPath_RF_bus_reg_dataout_181_port, 
                           regs(180) => DataPath_RF_bus_reg_dataout_180_port, 
                           regs(179) => DataPath_RF_bus_reg_dataout_179_port, 
                           regs(178) => DataPath_RF_bus_reg_dataout_178_port, 
                           regs(177) => DataPath_RF_bus_reg_dataout_177_port, 
                           regs(176) => DataPath_RF_bus_reg_dataout_176_port, 
                           regs(175) => DataPath_RF_bus_reg_dataout_175_port, 
                           regs(174) => DataPath_RF_bus_reg_dataout_174_port, 
                           regs(173) => DataPath_RF_bus_reg_dataout_173_port, 
                           regs(172) => DataPath_RF_bus_reg_dataout_172_port, 
                           regs(171) => DataPath_RF_bus_reg_dataout_171_port, 
                           regs(170) => DataPath_RF_bus_reg_dataout_170_port, 
                           regs(169) => DataPath_RF_bus_reg_dataout_169_port, 
                           regs(168) => DataPath_RF_bus_reg_dataout_168_port, 
                           regs(167) => DataPath_RF_bus_reg_dataout_167_port, 
                           regs(166) => DataPath_RF_bus_reg_dataout_166_port, 
                           regs(165) => DataPath_RF_bus_reg_dataout_165_port, 
                           regs(164) => DataPath_RF_bus_reg_dataout_164_port, 
                           regs(163) => DataPath_RF_bus_reg_dataout_163_port, 
                           regs(162) => DataPath_RF_bus_reg_dataout_162_port, 
                           regs(161) => DataPath_RF_bus_reg_dataout_161_port, 
                           regs(160) => DataPath_RF_bus_reg_dataout_160_port, 
                           regs(159) => DataPath_RF_bus_reg_dataout_159_port, 
                           regs(158) => DataPath_RF_bus_reg_dataout_158_port, 
                           regs(157) => DataPath_RF_bus_reg_dataout_157_port, 
                           regs(156) => DataPath_RF_bus_reg_dataout_156_port, 
                           regs(155) => DataPath_RF_bus_reg_dataout_155_port, 
                           regs(154) => DataPath_RF_bus_reg_dataout_154_port, 
                           regs(153) => DataPath_RF_bus_reg_dataout_153_port, 
                           regs(152) => DataPath_RF_bus_reg_dataout_152_port, 
                           regs(151) => DataPath_RF_bus_reg_dataout_151_port, 
                           regs(150) => DataPath_RF_bus_reg_dataout_150_port, 
                           regs(149) => DataPath_RF_bus_reg_dataout_149_port, 
                           regs(148) => DataPath_RF_bus_reg_dataout_148_port, 
                           regs(147) => DataPath_RF_bus_reg_dataout_147_port, 
                           regs(146) => DataPath_RF_bus_reg_dataout_146_port, 
                           regs(145) => DataPath_RF_bus_reg_dataout_145_port, 
                           regs(144) => DataPath_RF_bus_reg_dataout_144_port, 
                           regs(143) => DataPath_RF_bus_reg_dataout_143_port, 
                           regs(142) => DataPath_RF_bus_reg_dataout_142_port, 
                           regs(141) => DataPath_RF_bus_reg_dataout_141_port, 
                           regs(140) => DataPath_RF_bus_reg_dataout_140_port, 
                           regs(139) => DataPath_RF_bus_reg_dataout_139_port, 
                           regs(138) => DataPath_RF_bus_reg_dataout_138_port, 
                           regs(137) => DataPath_RF_bus_reg_dataout_137_port, 
                           regs(136) => DataPath_RF_bus_reg_dataout_136_port, 
                           regs(135) => DataPath_RF_bus_reg_dataout_135_port, 
                           regs(134) => DataPath_RF_bus_reg_dataout_134_port, 
                           regs(133) => DataPath_RF_bus_reg_dataout_133_port, 
                           regs(132) => DataPath_RF_bus_reg_dataout_132_port, 
                           regs(131) => DataPath_RF_bus_reg_dataout_131_port, 
                           regs(130) => DataPath_RF_bus_reg_dataout_130_port, 
                           regs(129) => DataPath_RF_bus_reg_dataout_129_port, 
                           regs(128) => DataPath_RF_bus_reg_dataout_128_port, 
                           regs(127) => DataPath_RF_bus_reg_dataout_127_port, 
                           regs(126) => DataPath_RF_bus_reg_dataout_126_port, 
                           regs(125) => DataPath_RF_bus_reg_dataout_125_port, 
                           regs(124) => DataPath_RF_bus_reg_dataout_124_port, 
                           regs(123) => DataPath_RF_bus_reg_dataout_123_port, 
                           regs(122) => DataPath_RF_bus_reg_dataout_122_port, 
                           regs(121) => DataPath_RF_bus_reg_dataout_121_port, 
                           regs(120) => DataPath_RF_bus_reg_dataout_120_port, 
                           regs(119) => DataPath_RF_bus_reg_dataout_119_port, 
                           regs(118) => DataPath_RF_bus_reg_dataout_118_port, 
                           regs(117) => DataPath_RF_bus_reg_dataout_117_port, 
                           regs(116) => DataPath_RF_bus_reg_dataout_116_port, 
                           regs(115) => DataPath_RF_bus_reg_dataout_115_port, 
                           regs(114) => DataPath_RF_bus_reg_dataout_114_port, 
                           regs(113) => DataPath_RF_bus_reg_dataout_113_port, 
                           regs(112) => DataPath_RF_bus_reg_dataout_112_port, 
                           regs(111) => DataPath_RF_bus_reg_dataout_111_port, 
                           regs(110) => DataPath_RF_bus_reg_dataout_110_port, 
                           regs(109) => DataPath_RF_bus_reg_dataout_109_port, 
                           regs(108) => DataPath_RF_bus_reg_dataout_108_port, 
                           regs(107) => DataPath_RF_bus_reg_dataout_107_port, 
                           regs(106) => DataPath_RF_bus_reg_dataout_106_port, 
                           regs(105) => DataPath_RF_bus_reg_dataout_105_port, 
                           regs(104) => DataPath_RF_bus_reg_dataout_104_port, 
                           regs(103) => DataPath_RF_bus_reg_dataout_103_port, 
                           regs(102) => DataPath_RF_bus_reg_dataout_102_port, 
                           regs(101) => DataPath_RF_bus_reg_dataout_101_port, 
                           regs(100) => DataPath_RF_bus_reg_dataout_100_port, 
                           regs(99) => DataPath_RF_bus_reg_dataout_99_port, 
                           regs(98) => DataPath_RF_bus_reg_dataout_98_port, 
                           regs(97) => DataPath_RF_bus_reg_dataout_97_port, 
                           regs(96) => DataPath_RF_bus_reg_dataout_96_port, 
                           regs(95) => DataPath_RF_bus_reg_dataout_95_port, 
                           regs(94) => DataPath_RF_bus_reg_dataout_94_port, 
                           regs(93) => DataPath_RF_bus_reg_dataout_93_port, 
                           regs(92) => DataPath_RF_bus_reg_dataout_92_port, 
                           regs(91) => DataPath_RF_bus_reg_dataout_91_port, 
                           regs(90) => DataPath_RF_bus_reg_dataout_90_port, 
                           regs(89) => DataPath_RF_bus_reg_dataout_89_port, 
                           regs(88) => DataPath_RF_bus_reg_dataout_88_port, 
                           regs(87) => DataPath_RF_bus_reg_dataout_87_port, 
                           regs(86) => DataPath_RF_bus_reg_dataout_86_port, 
                           regs(85) => DataPath_RF_bus_reg_dataout_85_port, 
                           regs(84) => DataPath_RF_bus_reg_dataout_84_port, 
                           regs(83) => DataPath_RF_bus_reg_dataout_83_port, 
                           regs(82) => DataPath_RF_bus_reg_dataout_82_port, 
                           regs(81) => DataPath_RF_bus_reg_dataout_81_port, 
                           regs(80) => DataPath_RF_bus_reg_dataout_80_port, 
                           regs(79) => DataPath_RF_bus_reg_dataout_79_port, 
                           regs(78) => DataPath_RF_bus_reg_dataout_78_port, 
                           regs(77) => DataPath_RF_bus_reg_dataout_77_port, 
                           regs(76) => DataPath_RF_bus_reg_dataout_76_port, 
                           regs(75) => DataPath_RF_bus_reg_dataout_75_port, 
                           regs(74) => DataPath_RF_bus_reg_dataout_74_port, 
                           regs(73) => DataPath_RF_bus_reg_dataout_73_port, 
                           regs(72) => DataPath_RF_bus_reg_dataout_72_port, 
                           regs(71) => DataPath_RF_bus_reg_dataout_71_port, 
                           regs(70) => DataPath_RF_bus_reg_dataout_70_port, 
                           regs(69) => DataPath_RF_bus_reg_dataout_69_port, 
                           regs(68) => DataPath_RF_bus_reg_dataout_68_port, 
                           regs(67) => DataPath_RF_bus_reg_dataout_67_port, 
                           regs(66) => DataPath_RF_bus_reg_dataout_66_port, 
                           regs(65) => DataPath_RF_bus_reg_dataout_65_port, 
                           regs(64) => DataPath_RF_bus_reg_dataout_64_port, 
                           regs(63) => DataPath_RF_bus_reg_dataout_63_port, 
                           regs(62) => DataPath_RF_bus_reg_dataout_62_port, 
                           regs(61) => DataPath_RF_bus_reg_dataout_61_port, 
                           regs(60) => DataPath_RF_bus_reg_dataout_60_port, 
                           regs(59) => DataPath_RF_bus_reg_dataout_59_port, 
                           regs(58) => DataPath_RF_bus_reg_dataout_58_port, 
                           regs(57) => DataPath_RF_bus_reg_dataout_57_port, 
                           regs(56) => DataPath_RF_bus_reg_dataout_56_port, 
                           regs(55) => DataPath_RF_bus_reg_dataout_55_port, 
                           regs(54) => DataPath_RF_bus_reg_dataout_54_port, 
                           regs(53) => DataPath_RF_bus_reg_dataout_53_port, 
                           regs(52) => DataPath_RF_bus_reg_dataout_52_port, 
                           regs(51) => DataPath_RF_bus_reg_dataout_51_port, 
                           regs(50) => DataPath_RF_bus_reg_dataout_50_port, 
                           regs(49) => DataPath_RF_bus_reg_dataout_49_port, 
                           regs(48) => DataPath_RF_bus_reg_dataout_48_port, 
                           regs(47) => DataPath_RF_bus_reg_dataout_47_port, 
                           regs(46) => DataPath_RF_bus_reg_dataout_46_port, 
                           regs(45) => DataPath_RF_bus_reg_dataout_45_port, 
                           regs(44) => DataPath_RF_bus_reg_dataout_44_port, 
                           regs(43) => DataPath_RF_bus_reg_dataout_43_port, 
                           regs(42) => DataPath_RF_bus_reg_dataout_42_port, 
                           regs(41) => DataPath_RF_bus_reg_dataout_41_port, 
                           regs(40) => DataPath_RF_bus_reg_dataout_40_port, 
                           regs(39) => DataPath_RF_bus_reg_dataout_39_port, 
                           regs(38) => DataPath_RF_bus_reg_dataout_38_port, 
                           regs(37) => DataPath_RF_bus_reg_dataout_37_port, 
                           regs(36) => DataPath_RF_bus_reg_dataout_36_port, 
                           regs(35) => DataPath_RF_bus_reg_dataout_35_port, 
                           regs(34) => DataPath_RF_bus_reg_dataout_34_port, 
                           regs(33) => DataPath_RF_bus_reg_dataout_33_port, 
                           regs(32) => DataPath_RF_bus_reg_dataout_32_port, 
                           regs(31) => DataPath_RF_bus_reg_dataout_31_port, 
                           regs(30) => DataPath_RF_bus_reg_dataout_30_port, 
                           regs(29) => DataPath_RF_bus_reg_dataout_29_port, 
                           regs(28) => DataPath_RF_bus_reg_dataout_28_port, 
                           regs(27) => DataPath_RF_bus_reg_dataout_27_port, 
                           regs(26) => DataPath_RF_bus_reg_dataout_26_port, 
                           regs(25) => DataPath_RF_bus_reg_dataout_25_port, 
                           regs(24) => DataPath_RF_bus_reg_dataout_24_port, 
                           regs(23) => DataPath_RF_bus_reg_dataout_23_port, 
                           regs(22) => DataPath_RF_bus_reg_dataout_22_port, 
                           regs(21) => DataPath_RF_bus_reg_dataout_21_port, 
                           regs(20) => DataPath_RF_bus_reg_dataout_20_port, 
                           regs(19) => DataPath_RF_bus_reg_dataout_19_port, 
                           regs(18) => DataPath_RF_bus_reg_dataout_18_port, 
                           regs(17) => DataPath_RF_bus_reg_dataout_17_port, 
                           regs(16) => DataPath_RF_bus_reg_dataout_16_port, 
                           regs(15) => DataPath_RF_bus_reg_dataout_15_port, 
                           regs(14) => DataPath_RF_bus_reg_dataout_14_port, 
                           regs(13) => DataPath_RF_bus_reg_dataout_13_port, 
                           regs(12) => DataPath_RF_bus_reg_dataout_12_port, 
                           regs(11) => DataPath_RF_bus_reg_dataout_11_port, 
                           regs(10) => DataPath_RF_bus_reg_dataout_10_port, 
                           regs(9) => DataPath_RF_bus_reg_dataout_9_port, 
                           regs(8) => DataPath_RF_bus_reg_dataout_8_port, 
                           regs(7) => DataPath_RF_bus_reg_dataout_7_port, 
                           regs(6) => DataPath_RF_bus_reg_dataout_6_port, 
                           regs(5) => DataPath_RF_bus_reg_dataout_5_port, 
                           regs(4) => DataPath_RF_bus_reg_dataout_4_port, 
                           regs(3) => DataPath_RF_bus_reg_dataout_3_port, 
                           regs(2) => DataPath_RF_bus_reg_dataout_2_port, 
                           regs(1) => DataPath_RF_bus_reg_dataout_1_port, 
                           regs(0) => DataPath_RF_bus_reg_dataout_0_port, 
                           win(4) => DataPath_RF_c_swin_4_port, win(3) => 
                           DataPath_RF_c_swin_3_port, win(2) => 
                           DataPath_RF_c_swin_2_port, win(1) => 
                           DataPath_RF_c_swin_1_port, win(0) => 
                           DataPath_RF_c_swin_0_port, curr_proc_regs(511) => 
                           DataPath_RF_bus_sel_savedwin_data_511_port, 
                           curr_proc_regs(510) => 
                           DataPath_RF_bus_sel_savedwin_data_510_port, 
                           curr_proc_regs(509) => 
                           DataPath_RF_bus_sel_savedwin_data_509_port, 
                           curr_proc_regs(508) => 
                           DataPath_RF_bus_sel_savedwin_data_508_port, 
                           curr_proc_regs(507) => 
                           DataPath_RF_bus_sel_savedwin_data_507_port, 
                           curr_proc_regs(506) => 
                           DataPath_RF_bus_sel_savedwin_data_506_port, 
                           curr_proc_regs(505) => 
                           DataPath_RF_bus_sel_savedwin_data_505_port, 
                           curr_proc_regs(504) => 
                           DataPath_RF_bus_sel_savedwin_data_504_port, 
                           curr_proc_regs(503) => 
                           DataPath_RF_bus_sel_savedwin_data_503_port, 
                           curr_proc_regs(502) => 
                           DataPath_RF_bus_sel_savedwin_data_502_port, 
                           curr_proc_regs(501) => 
                           DataPath_RF_bus_sel_savedwin_data_501_port, 
                           curr_proc_regs(500) => 
                           DataPath_RF_bus_sel_savedwin_data_500_port, 
                           curr_proc_regs(499) => 
                           DataPath_RF_bus_sel_savedwin_data_499_port, 
                           curr_proc_regs(498) => 
                           DataPath_RF_bus_sel_savedwin_data_498_port, 
                           curr_proc_regs(497) => 
                           DataPath_RF_bus_sel_savedwin_data_497_port, 
                           curr_proc_regs(496) => 
                           DataPath_RF_bus_sel_savedwin_data_496_port, 
                           curr_proc_regs(495) => 
                           DataPath_RF_bus_sel_savedwin_data_495_port, 
                           curr_proc_regs(494) => 
                           DataPath_RF_bus_sel_savedwin_data_494_port, 
                           curr_proc_regs(493) => 
                           DataPath_RF_bus_sel_savedwin_data_493_port, 
                           curr_proc_regs(492) => 
                           DataPath_RF_bus_sel_savedwin_data_492_port, 
                           curr_proc_regs(491) => 
                           DataPath_RF_bus_sel_savedwin_data_491_port, 
                           curr_proc_regs(490) => 
                           DataPath_RF_bus_sel_savedwin_data_490_port, 
                           curr_proc_regs(489) => 
                           DataPath_RF_bus_sel_savedwin_data_489_port, 
                           curr_proc_regs(488) => 
                           DataPath_RF_bus_sel_savedwin_data_488_port, 
                           curr_proc_regs(487) => 
                           DataPath_RF_bus_sel_savedwin_data_487_port, 
                           curr_proc_regs(486) => 
                           DataPath_RF_bus_sel_savedwin_data_486_port, 
                           curr_proc_regs(485) => 
                           DataPath_RF_bus_sel_savedwin_data_485_port, 
                           curr_proc_regs(484) => 
                           DataPath_RF_bus_sel_savedwin_data_484_port, 
                           curr_proc_regs(483) => 
                           DataPath_RF_bus_sel_savedwin_data_483_port, 
                           curr_proc_regs(482) => 
                           DataPath_RF_bus_sel_savedwin_data_482_port, 
                           curr_proc_regs(481) => 
                           DataPath_RF_bus_sel_savedwin_data_481_port, 
                           curr_proc_regs(480) => 
                           DataPath_RF_bus_sel_savedwin_data_480_port, 
                           curr_proc_regs(479) => 
                           DataPath_RF_bus_sel_savedwin_data_479_port, 
                           curr_proc_regs(478) => 
                           DataPath_RF_bus_sel_savedwin_data_478_port, 
                           curr_proc_regs(477) => 
                           DataPath_RF_bus_sel_savedwin_data_477_port, 
                           curr_proc_regs(476) => 
                           DataPath_RF_bus_sel_savedwin_data_476_port, 
                           curr_proc_regs(475) => 
                           DataPath_RF_bus_sel_savedwin_data_475_port, 
                           curr_proc_regs(474) => 
                           DataPath_RF_bus_sel_savedwin_data_474_port, 
                           curr_proc_regs(473) => 
                           DataPath_RF_bus_sel_savedwin_data_473_port, 
                           curr_proc_regs(472) => 
                           DataPath_RF_bus_sel_savedwin_data_472_port, 
                           curr_proc_regs(471) => 
                           DataPath_RF_bus_sel_savedwin_data_471_port, 
                           curr_proc_regs(470) => 
                           DataPath_RF_bus_sel_savedwin_data_470_port, 
                           curr_proc_regs(469) => 
                           DataPath_RF_bus_sel_savedwin_data_469_port, 
                           curr_proc_regs(468) => 
                           DataPath_RF_bus_sel_savedwin_data_468_port, 
                           curr_proc_regs(467) => 
                           DataPath_RF_bus_sel_savedwin_data_467_port, 
                           curr_proc_regs(466) => 
                           DataPath_RF_bus_sel_savedwin_data_466_port, 
                           curr_proc_regs(465) => 
                           DataPath_RF_bus_sel_savedwin_data_465_port, 
                           curr_proc_regs(464) => 
                           DataPath_RF_bus_sel_savedwin_data_464_port, 
                           curr_proc_regs(463) => 
                           DataPath_RF_bus_sel_savedwin_data_463_port, 
                           curr_proc_regs(462) => 
                           DataPath_RF_bus_sel_savedwin_data_462_port, 
                           curr_proc_regs(461) => 
                           DataPath_RF_bus_sel_savedwin_data_461_port, 
                           curr_proc_regs(460) => 
                           DataPath_RF_bus_sel_savedwin_data_460_port, 
                           curr_proc_regs(459) => 
                           DataPath_RF_bus_sel_savedwin_data_459_port, 
                           curr_proc_regs(458) => 
                           DataPath_RF_bus_sel_savedwin_data_458_port, 
                           curr_proc_regs(457) => 
                           DataPath_RF_bus_sel_savedwin_data_457_port, 
                           curr_proc_regs(456) => 
                           DataPath_RF_bus_sel_savedwin_data_456_port, 
                           curr_proc_regs(455) => 
                           DataPath_RF_bus_sel_savedwin_data_455_port, 
                           curr_proc_regs(454) => 
                           DataPath_RF_bus_sel_savedwin_data_454_port, 
                           curr_proc_regs(453) => 
                           DataPath_RF_bus_sel_savedwin_data_453_port, 
                           curr_proc_regs(452) => 
                           DataPath_RF_bus_sel_savedwin_data_452_port, 
                           curr_proc_regs(451) => 
                           DataPath_RF_bus_sel_savedwin_data_451_port, 
                           curr_proc_regs(450) => 
                           DataPath_RF_bus_sel_savedwin_data_450_port, 
                           curr_proc_regs(449) => 
                           DataPath_RF_bus_sel_savedwin_data_449_port, 
                           curr_proc_regs(448) => 
                           DataPath_RF_bus_sel_savedwin_data_448_port, 
                           curr_proc_regs(447) => 
                           DataPath_RF_bus_sel_savedwin_data_447_port, 
                           curr_proc_regs(446) => 
                           DataPath_RF_bus_sel_savedwin_data_446_port, 
                           curr_proc_regs(445) => 
                           DataPath_RF_bus_sel_savedwin_data_445_port, 
                           curr_proc_regs(444) => 
                           DataPath_RF_bus_sel_savedwin_data_444_port, 
                           curr_proc_regs(443) => 
                           DataPath_RF_bus_sel_savedwin_data_443_port, 
                           curr_proc_regs(442) => 
                           DataPath_RF_bus_sel_savedwin_data_442_port, 
                           curr_proc_regs(441) => 
                           DataPath_RF_bus_sel_savedwin_data_441_port, 
                           curr_proc_regs(440) => 
                           DataPath_RF_bus_sel_savedwin_data_440_port, 
                           curr_proc_regs(439) => 
                           DataPath_RF_bus_sel_savedwin_data_439_port, 
                           curr_proc_regs(438) => 
                           DataPath_RF_bus_sel_savedwin_data_438_port, 
                           curr_proc_regs(437) => 
                           DataPath_RF_bus_sel_savedwin_data_437_port, 
                           curr_proc_regs(436) => 
                           DataPath_RF_bus_sel_savedwin_data_436_port, 
                           curr_proc_regs(435) => 
                           DataPath_RF_bus_sel_savedwin_data_435_port, 
                           curr_proc_regs(434) => 
                           DataPath_RF_bus_sel_savedwin_data_434_port, 
                           curr_proc_regs(433) => 
                           DataPath_RF_bus_sel_savedwin_data_433_port, 
                           curr_proc_regs(432) => 
                           DataPath_RF_bus_sel_savedwin_data_432_port, 
                           curr_proc_regs(431) => 
                           DataPath_RF_bus_sel_savedwin_data_431_port, 
                           curr_proc_regs(430) => 
                           DataPath_RF_bus_sel_savedwin_data_430_port, 
                           curr_proc_regs(429) => 
                           DataPath_RF_bus_sel_savedwin_data_429_port, 
                           curr_proc_regs(428) => 
                           DataPath_RF_bus_sel_savedwin_data_428_port, 
                           curr_proc_regs(427) => 
                           DataPath_RF_bus_sel_savedwin_data_427_port, 
                           curr_proc_regs(426) => 
                           DataPath_RF_bus_sel_savedwin_data_426_port, 
                           curr_proc_regs(425) => 
                           DataPath_RF_bus_sel_savedwin_data_425_port, 
                           curr_proc_regs(424) => 
                           DataPath_RF_bus_sel_savedwin_data_424_port, 
                           curr_proc_regs(423) => 
                           DataPath_RF_bus_sel_savedwin_data_423_port, 
                           curr_proc_regs(422) => 
                           DataPath_RF_bus_sel_savedwin_data_422_port, 
                           curr_proc_regs(421) => 
                           DataPath_RF_bus_sel_savedwin_data_421_port, 
                           curr_proc_regs(420) => 
                           DataPath_RF_bus_sel_savedwin_data_420_port, 
                           curr_proc_regs(419) => 
                           DataPath_RF_bus_sel_savedwin_data_419_port, 
                           curr_proc_regs(418) => 
                           DataPath_RF_bus_sel_savedwin_data_418_port, 
                           curr_proc_regs(417) => 
                           DataPath_RF_bus_sel_savedwin_data_417_port, 
                           curr_proc_regs(416) => 
                           DataPath_RF_bus_sel_savedwin_data_416_port, 
                           curr_proc_regs(415) => 
                           DataPath_RF_bus_sel_savedwin_data_415_port, 
                           curr_proc_regs(414) => 
                           DataPath_RF_bus_sel_savedwin_data_414_port, 
                           curr_proc_regs(413) => 
                           DataPath_RF_bus_sel_savedwin_data_413_port, 
                           curr_proc_regs(412) => 
                           DataPath_RF_bus_sel_savedwin_data_412_port, 
                           curr_proc_regs(411) => 
                           DataPath_RF_bus_sel_savedwin_data_411_port, 
                           curr_proc_regs(410) => 
                           DataPath_RF_bus_sel_savedwin_data_410_port, 
                           curr_proc_regs(409) => 
                           DataPath_RF_bus_sel_savedwin_data_409_port, 
                           curr_proc_regs(408) => 
                           DataPath_RF_bus_sel_savedwin_data_408_port, 
                           curr_proc_regs(407) => 
                           DataPath_RF_bus_sel_savedwin_data_407_port, 
                           curr_proc_regs(406) => 
                           DataPath_RF_bus_sel_savedwin_data_406_port, 
                           curr_proc_regs(405) => 
                           DataPath_RF_bus_sel_savedwin_data_405_port, 
                           curr_proc_regs(404) => 
                           DataPath_RF_bus_sel_savedwin_data_404_port, 
                           curr_proc_regs(403) => 
                           DataPath_RF_bus_sel_savedwin_data_403_port, 
                           curr_proc_regs(402) => 
                           DataPath_RF_bus_sel_savedwin_data_402_port, 
                           curr_proc_regs(401) => 
                           DataPath_RF_bus_sel_savedwin_data_401_port, 
                           curr_proc_regs(400) => 
                           DataPath_RF_bus_sel_savedwin_data_400_port, 
                           curr_proc_regs(399) => 
                           DataPath_RF_bus_sel_savedwin_data_399_port, 
                           curr_proc_regs(398) => 
                           DataPath_RF_bus_sel_savedwin_data_398_port, 
                           curr_proc_regs(397) => 
                           DataPath_RF_bus_sel_savedwin_data_397_port, 
                           curr_proc_regs(396) => 
                           DataPath_RF_bus_sel_savedwin_data_396_port, 
                           curr_proc_regs(395) => 
                           DataPath_RF_bus_sel_savedwin_data_395_port, 
                           curr_proc_regs(394) => 
                           DataPath_RF_bus_sel_savedwin_data_394_port, 
                           curr_proc_regs(393) => 
                           DataPath_RF_bus_sel_savedwin_data_393_port, 
                           curr_proc_regs(392) => 
                           DataPath_RF_bus_sel_savedwin_data_392_port, 
                           curr_proc_regs(391) => 
                           DataPath_RF_bus_sel_savedwin_data_391_port, 
                           curr_proc_regs(390) => 
                           DataPath_RF_bus_sel_savedwin_data_390_port, 
                           curr_proc_regs(389) => 
                           DataPath_RF_bus_sel_savedwin_data_389_port, 
                           curr_proc_regs(388) => 
                           DataPath_RF_bus_sel_savedwin_data_388_port, 
                           curr_proc_regs(387) => 
                           DataPath_RF_bus_sel_savedwin_data_387_port, 
                           curr_proc_regs(386) => 
                           DataPath_RF_bus_sel_savedwin_data_386_port, 
                           curr_proc_regs(385) => 
                           DataPath_RF_bus_sel_savedwin_data_385_port, 
                           curr_proc_regs(384) => 
                           DataPath_RF_bus_sel_savedwin_data_384_port, 
                           curr_proc_regs(383) => 
                           DataPath_RF_bus_sel_savedwin_data_383_port, 
                           curr_proc_regs(382) => 
                           DataPath_RF_bus_sel_savedwin_data_382_port, 
                           curr_proc_regs(381) => 
                           DataPath_RF_bus_sel_savedwin_data_381_port, 
                           curr_proc_regs(380) => 
                           DataPath_RF_bus_sel_savedwin_data_380_port, 
                           curr_proc_regs(379) => 
                           DataPath_RF_bus_sel_savedwin_data_379_port, 
                           curr_proc_regs(378) => 
                           DataPath_RF_bus_sel_savedwin_data_378_port, 
                           curr_proc_regs(377) => 
                           DataPath_RF_bus_sel_savedwin_data_377_port, 
                           curr_proc_regs(376) => 
                           DataPath_RF_bus_sel_savedwin_data_376_port, 
                           curr_proc_regs(375) => 
                           DataPath_RF_bus_sel_savedwin_data_375_port, 
                           curr_proc_regs(374) => 
                           DataPath_RF_bus_sel_savedwin_data_374_port, 
                           curr_proc_regs(373) => 
                           DataPath_RF_bus_sel_savedwin_data_373_port, 
                           curr_proc_regs(372) => 
                           DataPath_RF_bus_sel_savedwin_data_372_port, 
                           curr_proc_regs(371) => 
                           DataPath_RF_bus_sel_savedwin_data_371_port, 
                           curr_proc_regs(370) => 
                           DataPath_RF_bus_sel_savedwin_data_370_port, 
                           curr_proc_regs(369) => 
                           DataPath_RF_bus_sel_savedwin_data_369_port, 
                           curr_proc_regs(368) => 
                           DataPath_RF_bus_sel_savedwin_data_368_port, 
                           curr_proc_regs(367) => 
                           DataPath_RF_bus_sel_savedwin_data_367_port, 
                           curr_proc_regs(366) => 
                           DataPath_RF_bus_sel_savedwin_data_366_port, 
                           curr_proc_regs(365) => 
                           DataPath_RF_bus_sel_savedwin_data_365_port, 
                           curr_proc_regs(364) => 
                           DataPath_RF_bus_sel_savedwin_data_364_port, 
                           curr_proc_regs(363) => 
                           DataPath_RF_bus_sel_savedwin_data_363_port, 
                           curr_proc_regs(362) => 
                           DataPath_RF_bus_sel_savedwin_data_362_port, 
                           curr_proc_regs(361) => 
                           DataPath_RF_bus_sel_savedwin_data_361_port, 
                           curr_proc_regs(360) => 
                           DataPath_RF_bus_sel_savedwin_data_360_port, 
                           curr_proc_regs(359) => 
                           DataPath_RF_bus_sel_savedwin_data_359_port, 
                           curr_proc_regs(358) => 
                           DataPath_RF_bus_sel_savedwin_data_358_port, 
                           curr_proc_regs(357) => 
                           DataPath_RF_bus_sel_savedwin_data_357_port, 
                           curr_proc_regs(356) => 
                           DataPath_RF_bus_sel_savedwin_data_356_port, 
                           curr_proc_regs(355) => 
                           DataPath_RF_bus_sel_savedwin_data_355_port, 
                           curr_proc_regs(354) => 
                           DataPath_RF_bus_sel_savedwin_data_354_port, 
                           curr_proc_regs(353) => 
                           DataPath_RF_bus_sel_savedwin_data_353_port, 
                           curr_proc_regs(352) => 
                           DataPath_RF_bus_sel_savedwin_data_352_port, 
                           curr_proc_regs(351) => 
                           DataPath_RF_bus_sel_savedwin_data_351_port, 
                           curr_proc_regs(350) => 
                           DataPath_RF_bus_sel_savedwin_data_350_port, 
                           curr_proc_regs(349) => 
                           DataPath_RF_bus_sel_savedwin_data_349_port, 
                           curr_proc_regs(348) => 
                           DataPath_RF_bus_sel_savedwin_data_348_port, 
                           curr_proc_regs(347) => 
                           DataPath_RF_bus_sel_savedwin_data_347_port, 
                           curr_proc_regs(346) => 
                           DataPath_RF_bus_sel_savedwin_data_346_port, 
                           curr_proc_regs(345) => 
                           DataPath_RF_bus_sel_savedwin_data_345_port, 
                           curr_proc_regs(344) => 
                           DataPath_RF_bus_sel_savedwin_data_344_port, 
                           curr_proc_regs(343) => 
                           DataPath_RF_bus_sel_savedwin_data_343_port, 
                           curr_proc_regs(342) => 
                           DataPath_RF_bus_sel_savedwin_data_342_port, 
                           curr_proc_regs(341) => 
                           DataPath_RF_bus_sel_savedwin_data_341_port, 
                           curr_proc_regs(340) => 
                           DataPath_RF_bus_sel_savedwin_data_340_port, 
                           curr_proc_regs(339) => 
                           DataPath_RF_bus_sel_savedwin_data_339_port, 
                           curr_proc_regs(338) => 
                           DataPath_RF_bus_sel_savedwin_data_338_port, 
                           curr_proc_regs(337) => 
                           DataPath_RF_bus_sel_savedwin_data_337_port, 
                           curr_proc_regs(336) => 
                           DataPath_RF_bus_sel_savedwin_data_336_port, 
                           curr_proc_regs(335) => 
                           DataPath_RF_bus_sel_savedwin_data_335_port, 
                           curr_proc_regs(334) => 
                           DataPath_RF_bus_sel_savedwin_data_334_port, 
                           curr_proc_regs(333) => 
                           DataPath_RF_bus_sel_savedwin_data_333_port, 
                           curr_proc_regs(332) => 
                           DataPath_RF_bus_sel_savedwin_data_332_port, 
                           curr_proc_regs(331) => 
                           DataPath_RF_bus_sel_savedwin_data_331_port, 
                           curr_proc_regs(330) => 
                           DataPath_RF_bus_sel_savedwin_data_330_port, 
                           curr_proc_regs(329) => 
                           DataPath_RF_bus_sel_savedwin_data_329_port, 
                           curr_proc_regs(328) => 
                           DataPath_RF_bus_sel_savedwin_data_328_port, 
                           curr_proc_regs(327) => 
                           DataPath_RF_bus_sel_savedwin_data_327_port, 
                           curr_proc_regs(326) => 
                           DataPath_RF_bus_sel_savedwin_data_326_port, 
                           curr_proc_regs(325) => 
                           DataPath_RF_bus_sel_savedwin_data_325_port, 
                           curr_proc_regs(324) => 
                           DataPath_RF_bus_sel_savedwin_data_324_port, 
                           curr_proc_regs(323) => 
                           DataPath_RF_bus_sel_savedwin_data_323_port, 
                           curr_proc_regs(322) => 
                           DataPath_RF_bus_sel_savedwin_data_322_port, 
                           curr_proc_regs(321) => 
                           DataPath_RF_bus_sel_savedwin_data_321_port, 
                           curr_proc_regs(320) => 
                           DataPath_RF_bus_sel_savedwin_data_320_port, 
                           curr_proc_regs(319) => 
                           DataPath_RF_bus_sel_savedwin_data_319_port, 
                           curr_proc_regs(318) => 
                           DataPath_RF_bus_sel_savedwin_data_318_port, 
                           curr_proc_regs(317) => 
                           DataPath_RF_bus_sel_savedwin_data_317_port, 
                           curr_proc_regs(316) => 
                           DataPath_RF_bus_sel_savedwin_data_316_port, 
                           curr_proc_regs(315) => 
                           DataPath_RF_bus_sel_savedwin_data_315_port, 
                           curr_proc_regs(314) => 
                           DataPath_RF_bus_sel_savedwin_data_314_port, 
                           curr_proc_regs(313) => 
                           DataPath_RF_bus_sel_savedwin_data_313_port, 
                           curr_proc_regs(312) => 
                           DataPath_RF_bus_sel_savedwin_data_312_port, 
                           curr_proc_regs(311) => 
                           DataPath_RF_bus_sel_savedwin_data_311_port, 
                           curr_proc_regs(310) => 
                           DataPath_RF_bus_sel_savedwin_data_310_port, 
                           curr_proc_regs(309) => 
                           DataPath_RF_bus_sel_savedwin_data_309_port, 
                           curr_proc_regs(308) => 
                           DataPath_RF_bus_sel_savedwin_data_308_port, 
                           curr_proc_regs(307) => 
                           DataPath_RF_bus_sel_savedwin_data_307_port, 
                           curr_proc_regs(306) => 
                           DataPath_RF_bus_sel_savedwin_data_306_port, 
                           curr_proc_regs(305) => 
                           DataPath_RF_bus_sel_savedwin_data_305_port, 
                           curr_proc_regs(304) => 
                           DataPath_RF_bus_sel_savedwin_data_304_port, 
                           curr_proc_regs(303) => 
                           DataPath_RF_bus_sel_savedwin_data_303_port, 
                           curr_proc_regs(302) => 
                           DataPath_RF_bus_sel_savedwin_data_302_port, 
                           curr_proc_regs(301) => 
                           DataPath_RF_bus_sel_savedwin_data_301_port, 
                           curr_proc_regs(300) => 
                           DataPath_RF_bus_sel_savedwin_data_300_port, 
                           curr_proc_regs(299) => 
                           DataPath_RF_bus_sel_savedwin_data_299_port, 
                           curr_proc_regs(298) => 
                           DataPath_RF_bus_sel_savedwin_data_298_port, 
                           curr_proc_regs(297) => 
                           DataPath_RF_bus_sel_savedwin_data_297_port, 
                           curr_proc_regs(296) => 
                           DataPath_RF_bus_sel_savedwin_data_296_port, 
                           curr_proc_regs(295) => 
                           DataPath_RF_bus_sel_savedwin_data_295_port, 
                           curr_proc_regs(294) => 
                           DataPath_RF_bus_sel_savedwin_data_294_port, 
                           curr_proc_regs(293) => 
                           DataPath_RF_bus_sel_savedwin_data_293_port, 
                           curr_proc_regs(292) => 
                           DataPath_RF_bus_sel_savedwin_data_292_port, 
                           curr_proc_regs(291) => 
                           DataPath_RF_bus_sel_savedwin_data_291_port, 
                           curr_proc_regs(290) => 
                           DataPath_RF_bus_sel_savedwin_data_290_port, 
                           curr_proc_regs(289) => 
                           DataPath_RF_bus_sel_savedwin_data_289_port, 
                           curr_proc_regs(288) => 
                           DataPath_RF_bus_sel_savedwin_data_288_port, 
                           curr_proc_regs(287) => 
                           DataPath_RF_bus_sel_savedwin_data_287_port, 
                           curr_proc_regs(286) => 
                           DataPath_RF_bus_sel_savedwin_data_286_port, 
                           curr_proc_regs(285) => 
                           DataPath_RF_bus_sel_savedwin_data_285_port, 
                           curr_proc_regs(284) => 
                           DataPath_RF_bus_sel_savedwin_data_284_port, 
                           curr_proc_regs(283) => 
                           DataPath_RF_bus_sel_savedwin_data_283_port, 
                           curr_proc_regs(282) => 
                           DataPath_RF_bus_sel_savedwin_data_282_port, 
                           curr_proc_regs(281) => 
                           DataPath_RF_bus_sel_savedwin_data_281_port, 
                           curr_proc_regs(280) => 
                           DataPath_RF_bus_sel_savedwin_data_280_port, 
                           curr_proc_regs(279) => 
                           DataPath_RF_bus_sel_savedwin_data_279_port, 
                           curr_proc_regs(278) => 
                           DataPath_RF_bus_sel_savedwin_data_278_port, 
                           curr_proc_regs(277) => 
                           DataPath_RF_bus_sel_savedwin_data_277_port, 
                           curr_proc_regs(276) => 
                           DataPath_RF_bus_sel_savedwin_data_276_port, 
                           curr_proc_regs(275) => 
                           DataPath_RF_bus_sel_savedwin_data_275_port, 
                           curr_proc_regs(274) => 
                           DataPath_RF_bus_sel_savedwin_data_274_port, 
                           curr_proc_regs(273) => 
                           DataPath_RF_bus_sel_savedwin_data_273_port, 
                           curr_proc_regs(272) => 
                           DataPath_RF_bus_sel_savedwin_data_272_port, 
                           curr_proc_regs(271) => 
                           DataPath_RF_bus_sel_savedwin_data_271_port, 
                           curr_proc_regs(270) => 
                           DataPath_RF_bus_sel_savedwin_data_270_port, 
                           curr_proc_regs(269) => 
                           DataPath_RF_bus_sel_savedwin_data_269_port, 
                           curr_proc_regs(268) => 
                           DataPath_RF_bus_sel_savedwin_data_268_port, 
                           curr_proc_regs(267) => 
                           DataPath_RF_bus_sel_savedwin_data_267_port, 
                           curr_proc_regs(266) => 
                           DataPath_RF_bus_sel_savedwin_data_266_port, 
                           curr_proc_regs(265) => 
                           DataPath_RF_bus_sel_savedwin_data_265_port, 
                           curr_proc_regs(264) => 
                           DataPath_RF_bus_sel_savedwin_data_264_port, 
                           curr_proc_regs(263) => 
                           DataPath_RF_bus_sel_savedwin_data_263_port, 
                           curr_proc_regs(262) => 
                           DataPath_RF_bus_sel_savedwin_data_262_port, 
                           curr_proc_regs(261) => 
                           DataPath_RF_bus_sel_savedwin_data_261_port, 
                           curr_proc_regs(260) => 
                           DataPath_RF_bus_sel_savedwin_data_260_port, 
                           curr_proc_regs(259) => 
                           DataPath_RF_bus_sel_savedwin_data_259_port, 
                           curr_proc_regs(258) => 
                           DataPath_RF_bus_sel_savedwin_data_258_port, 
                           curr_proc_regs(257) => 
                           DataPath_RF_bus_sel_savedwin_data_257_port, 
                           curr_proc_regs(256) => 
                           DataPath_RF_bus_sel_savedwin_data_256_port, 
                           curr_proc_regs(255) => 
                           DataPath_RF_bus_sel_savedwin_data_255_port, 
                           curr_proc_regs(254) => 
                           DataPath_RF_bus_sel_savedwin_data_254_port, 
                           curr_proc_regs(253) => 
                           DataPath_RF_bus_sel_savedwin_data_253_port, 
                           curr_proc_regs(252) => 
                           DataPath_RF_bus_sel_savedwin_data_252_port, 
                           curr_proc_regs(251) => 
                           DataPath_RF_bus_sel_savedwin_data_251_port, 
                           curr_proc_regs(250) => 
                           DataPath_RF_bus_sel_savedwin_data_250_port, 
                           curr_proc_regs(249) => 
                           DataPath_RF_bus_sel_savedwin_data_249_port, 
                           curr_proc_regs(248) => 
                           DataPath_RF_bus_sel_savedwin_data_248_port, 
                           curr_proc_regs(247) => 
                           DataPath_RF_bus_sel_savedwin_data_247_port, 
                           curr_proc_regs(246) => 
                           DataPath_RF_bus_sel_savedwin_data_246_port, 
                           curr_proc_regs(245) => 
                           DataPath_RF_bus_sel_savedwin_data_245_port, 
                           curr_proc_regs(244) => 
                           DataPath_RF_bus_sel_savedwin_data_244_port, 
                           curr_proc_regs(243) => 
                           DataPath_RF_bus_sel_savedwin_data_243_port, 
                           curr_proc_regs(242) => 
                           DataPath_RF_bus_sel_savedwin_data_242_port, 
                           curr_proc_regs(241) => 
                           DataPath_RF_bus_sel_savedwin_data_241_port, 
                           curr_proc_regs(240) => 
                           DataPath_RF_bus_sel_savedwin_data_240_port, 
                           curr_proc_regs(239) => 
                           DataPath_RF_bus_sel_savedwin_data_239_port, 
                           curr_proc_regs(238) => 
                           DataPath_RF_bus_sel_savedwin_data_238_port, 
                           curr_proc_regs(237) => 
                           DataPath_RF_bus_sel_savedwin_data_237_port, 
                           curr_proc_regs(236) => 
                           DataPath_RF_bus_sel_savedwin_data_236_port, 
                           curr_proc_regs(235) => 
                           DataPath_RF_bus_sel_savedwin_data_235_port, 
                           curr_proc_regs(234) => 
                           DataPath_RF_bus_sel_savedwin_data_234_port, 
                           curr_proc_regs(233) => 
                           DataPath_RF_bus_sel_savedwin_data_233_port, 
                           curr_proc_regs(232) => 
                           DataPath_RF_bus_sel_savedwin_data_232_port, 
                           curr_proc_regs(231) => 
                           DataPath_RF_bus_sel_savedwin_data_231_port, 
                           curr_proc_regs(230) => 
                           DataPath_RF_bus_sel_savedwin_data_230_port, 
                           curr_proc_regs(229) => 
                           DataPath_RF_bus_sel_savedwin_data_229_port, 
                           curr_proc_regs(228) => 
                           DataPath_RF_bus_sel_savedwin_data_228_port, 
                           curr_proc_regs(227) => 
                           DataPath_RF_bus_sel_savedwin_data_227_port, 
                           curr_proc_regs(226) => 
                           DataPath_RF_bus_sel_savedwin_data_226_port, 
                           curr_proc_regs(225) => 
                           DataPath_RF_bus_sel_savedwin_data_225_port, 
                           curr_proc_regs(224) => 
                           DataPath_RF_bus_sel_savedwin_data_224_port, 
                           curr_proc_regs(223) => 
                           DataPath_RF_bus_sel_savedwin_data_223_port, 
                           curr_proc_regs(222) => 
                           DataPath_RF_bus_sel_savedwin_data_222_port, 
                           curr_proc_regs(221) => 
                           DataPath_RF_bus_sel_savedwin_data_221_port, 
                           curr_proc_regs(220) => 
                           DataPath_RF_bus_sel_savedwin_data_220_port, 
                           curr_proc_regs(219) => 
                           DataPath_RF_bus_sel_savedwin_data_219_port, 
                           curr_proc_regs(218) => 
                           DataPath_RF_bus_sel_savedwin_data_218_port, 
                           curr_proc_regs(217) => 
                           DataPath_RF_bus_sel_savedwin_data_217_port, 
                           curr_proc_regs(216) => 
                           DataPath_RF_bus_sel_savedwin_data_216_port, 
                           curr_proc_regs(215) => 
                           DataPath_RF_bus_sel_savedwin_data_215_port, 
                           curr_proc_regs(214) => 
                           DataPath_RF_bus_sel_savedwin_data_214_port, 
                           curr_proc_regs(213) => 
                           DataPath_RF_bus_sel_savedwin_data_213_port, 
                           curr_proc_regs(212) => 
                           DataPath_RF_bus_sel_savedwin_data_212_port, 
                           curr_proc_regs(211) => 
                           DataPath_RF_bus_sel_savedwin_data_211_port, 
                           curr_proc_regs(210) => 
                           DataPath_RF_bus_sel_savedwin_data_210_port, 
                           curr_proc_regs(209) => 
                           DataPath_RF_bus_sel_savedwin_data_209_port, 
                           curr_proc_regs(208) => 
                           DataPath_RF_bus_sel_savedwin_data_208_port, 
                           curr_proc_regs(207) => 
                           DataPath_RF_bus_sel_savedwin_data_207_port, 
                           curr_proc_regs(206) => 
                           DataPath_RF_bus_sel_savedwin_data_206_port, 
                           curr_proc_regs(205) => 
                           DataPath_RF_bus_sel_savedwin_data_205_port, 
                           curr_proc_regs(204) => 
                           DataPath_RF_bus_sel_savedwin_data_204_port, 
                           curr_proc_regs(203) => 
                           DataPath_RF_bus_sel_savedwin_data_203_port, 
                           curr_proc_regs(202) => 
                           DataPath_RF_bus_sel_savedwin_data_202_port, 
                           curr_proc_regs(201) => 
                           DataPath_RF_bus_sel_savedwin_data_201_port, 
                           curr_proc_regs(200) => 
                           DataPath_RF_bus_sel_savedwin_data_200_port, 
                           curr_proc_regs(199) => 
                           DataPath_RF_bus_sel_savedwin_data_199_port, 
                           curr_proc_regs(198) => 
                           DataPath_RF_bus_sel_savedwin_data_198_port, 
                           curr_proc_regs(197) => 
                           DataPath_RF_bus_sel_savedwin_data_197_port, 
                           curr_proc_regs(196) => 
                           DataPath_RF_bus_sel_savedwin_data_196_port, 
                           curr_proc_regs(195) => 
                           DataPath_RF_bus_sel_savedwin_data_195_port, 
                           curr_proc_regs(194) => 
                           DataPath_RF_bus_sel_savedwin_data_194_port, 
                           curr_proc_regs(193) => 
                           DataPath_RF_bus_sel_savedwin_data_193_port, 
                           curr_proc_regs(192) => 
                           DataPath_RF_bus_sel_savedwin_data_192_port, 
                           curr_proc_regs(191) => 
                           DataPath_RF_bus_sel_savedwin_data_191_port, 
                           curr_proc_regs(190) => 
                           DataPath_RF_bus_sel_savedwin_data_190_port, 
                           curr_proc_regs(189) => 
                           DataPath_RF_bus_sel_savedwin_data_189_port, 
                           curr_proc_regs(188) => 
                           DataPath_RF_bus_sel_savedwin_data_188_port, 
                           curr_proc_regs(187) => 
                           DataPath_RF_bus_sel_savedwin_data_187_port, 
                           curr_proc_regs(186) => 
                           DataPath_RF_bus_sel_savedwin_data_186_port, 
                           curr_proc_regs(185) => 
                           DataPath_RF_bus_sel_savedwin_data_185_port, 
                           curr_proc_regs(184) => 
                           DataPath_RF_bus_sel_savedwin_data_184_port, 
                           curr_proc_regs(183) => 
                           DataPath_RF_bus_sel_savedwin_data_183_port, 
                           curr_proc_regs(182) => 
                           DataPath_RF_bus_sel_savedwin_data_182_port, 
                           curr_proc_regs(181) => 
                           DataPath_RF_bus_sel_savedwin_data_181_port, 
                           curr_proc_regs(180) => 
                           DataPath_RF_bus_sel_savedwin_data_180_port, 
                           curr_proc_regs(179) => 
                           DataPath_RF_bus_sel_savedwin_data_179_port, 
                           curr_proc_regs(178) => 
                           DataPath_RF_bus_sel_savedwin_data_178_port, 
                           curr_proc_regs(177) => 
                           DataPath_RF_bus_sel_savedwin_data_177_port, 
                           curr_proc_regs(176) => 
                           DataPath_RF_bus_sel_savedwin_data_176_port, 
                           curr_proc_regs(175) => 
                           DataPath_RF_bus_sel_savedwin_data_175_port, 
                           curr_proc_regs(174) => 
                           DataPath_RF_bus_sel_savedwin_data_174_port, 
                           curr_proc_regs(173) => 
                           DataPath_RF_bus_sel_savedwin_data_173_port, 
                           curr_proc_regs(172) => 
                           DataPath_RF_bus_sel_savedwin_data_172_port, 
                           curr_proc_regs(171) => 
                           DataPath_RF_bus_sel_savedwin_data_171_port, 
                           curr_proc_regs(170) => 
                           DataPath_RF_bus_sel_savedwin_data_170_port, 
                           curr_proc_regs(169) => 
                           DataPath_RF_bus_sel_savedwin_data_169_port, 
                           curr_proc_regs(168) => 
                           DataPath_RF_bus_sel_savedwin_data_168_port, 
                           curr_proc_regs(167) => 
                           DataPath_RF_bus_sel_savedwin_data_167_port, 
                           curr_proc_regs(166) => 
                           DataPath_RF_bus_sel_savedwin_data_166_port, 
                           curr_proc_regs(165) => 
                           DataPath_RF_bus_sel_savedwin_data_165_port, 
                           curr_proc_regs(164) => 
                           DataPath_RF_bus_sel_savedwin_data_164_port, 
                           curr_proc_regs(163) => 
                           DataPath_RF_bus_sel_savedwin_data_163_port, 
                           curr_proc_regs(162) => 
                           DataPath_RF_bus_sel_savedwin_data_162_port, 
                           curr_proc_regs(161) => 
                           DataPath_RF_bus_sel_savedwin_data_161_port, 
                           curr_proc_regs(160) => 
                           DataPath_RF_bus_sel_savedwin_data_160_port, 
                           curr_proc_regs(159) => 
                           DataPath_RF_bus_sel_savedwin_data_159_port, 
                           curr_proc_regs(158) => 
                           DataPath_RF_bus_sel_savedwin_data_158_port, 
                           curr_proc_regs(157) => 
                           DataPath_RF_bus_sel_savedwin_data_157_port, 
                           curr_proc_regs(156) => 
                           DataPath_RF_bus_sel_savedwin_data_156_port, 
                           curr_proc_regs(155) => 
                           DataPath_RF_bus_sel_savedwin_data_155_port, 
                           curr_proc_regs(154) => 
                           DataPath_RF_bus_sel_savedwin_data_154_port, 
                           curr_proc_regs(153) => 
                           DataPath_RF_bus_sel_savedwin_data_153_port, 
                           curr_proc_regs(152) => 
                           DataPath_RF_bus_sel_savedwin_data_152_port, 
                           curr_proc_regs(151) => 
                           DataPath_RF_bus_sel_savedwin_data_151_port, 
                           curr_proc_regs(150) => 
                           DataPath_RF_bus_sel_savedwin_data_150_port, 
                           curr_proc_regs(149) => 
                           DataPath_RF_bus_sel_savedwin_data_149_port, 
                           curr_proc_regs(148) => 
                           DataPath_RF_bus_sel_savedwin_data_148_port, 
                           curr_proc_regs(147) => 
                           DataPath_RF_bus_sel_savedwin_data_147_port, 
                           curr_proc_regs(146) => 
                           DataPath_RF_bus_sel_savedwin_data_146_port, 
                           curr_proc_regs(145) => 
                           DataPath_RF_bus_sel_savedwin_data_145_port, 
                           curr_proc_regs(144) => 
                           DataPath_RF_bus_sel_savedwin_data_144_port, 
                           curr_proc_regs(143) => 
                           DataPath_RF_bus_sel_savedwin_data_143_port, 
                           curr_proc_regs(142) => 
                           DataPath_RF_bus_sel_savedwin_data_142_port, 
                           curr_proc_regs(141) => 
                           DataPath_RF_bus_sel_savedwin_data_141_port, 
                           curr_proc_regs(140) => 
                           DataPath_RF_bus_sel_savedwin_data_140_port, 
                           curr_proc_regs(139) => 
                           DataPath_RF_bus_sel_savedwin_data_139_port, 
                           curr_proc_regs(138) => 
                           DataPath_RF_bus_sel_savedwin_data_138_port, 
                           curr_proc_regs(137) => 
                           DataPath_RF_bus_sel_savedwin_data_137_port, 
                           curr_proc_regs(136) => 
                           DataPath_RF_bus_sel_savedwin_data_136_port, 
                           curr_proc_regs(135) => 
                           DataPath_RF_bus_sel_savedwin_data_135_port, 
                           curr_proc_regs(134) => 
                           DataPath_RF_bus_sel_savedwin_data_134_port, 
                           curr_proc_regs(133) => 
                           DataPath_RF_bus_sel_savedwin_data_133_port, 
                           curr_proc_regs(132) => 
                           DataPath_RF_bus_sel_savedwin_data_132_port, 
                           curr_proc_regs(131) => 
                           DataPath_RF_bus_sel_savedwin_data_131_port, 
                           curr_proc_regs(130) => 
                           DataPath_RF_bus_sel_savedwin_data_130_port, 
                           curr_proc_regs(129) => 
                           DataPath_RF_bus_sel_savedwin_data_129_port, 
                           curr_proc_regs(128) => 
                           DataPath_RF_bus_sel_savedwin_data_128_port, 
                           curr_proc_regs(127) => 
                           DataPath_RF_bus_sel_savedwin_data_127_port, 
                           curr_proc_regs(126) => 
                           DataPath_RF_bus_sel_savedwin_data_126_port, 
                           curr_proc_regs(125) => 
                           DataPath_RF_bus_sel_savedwin_data_125_port, 
                           curr_proc_regs(124) => 
                           DataPath_RF_bus_sel_savedwin_data_124_port, 
                           curr_proc_regs(123) => 
                           DataPath_RF_bus_sel_savedwin_data_123_port, 
                           curr_proc_regs(122) => 
                           DataPath_RF_bus_sel_savedwin_data_122_port, 
                           curr_proc_regs(121) => 
                           DataPath_RF_bus_sel_savedwin_data_121_port, 
                           curr_proc_regs(120) => 
                           DataPath_RF_bus_sel_savedwin_data_120_port, 
                           curr_proc_regs(119) => 
                           DataPath_RF_bus_sel_savedwin_data_119_port, 
                           curr_proc_regs(118) => 
                           DataPath_RF_bus_sel_savedwin_data_118_port, 
                           curr_proc_regs(117) => 
                           DataPath_RF_bus_sel_savedwin_data_117_port, 
                           curr_proc_regs(116) => 
                           DataPath_RF_bus_sel_savedwin_data_116_port, 
                           curr_proc_regs(115) => 
                           DataPath_RF_bus_sel_savedwin_data_115_port, 
                           curr_proc_regs(114) => 
                           DataPath_RF_bus_sel_savedwin_data_114_port, 
                           curr_proc_regs(113) => 
                           DataPath_RF_bus_sel_savedwin_data_113_port, 
                           curr_proc_regs(112) => 
                           DataPath_RF_bus_sel_savedwin_data_112_port, 
                           curr_proc_regs(111) => 
                           DataPath_RF_bus_sel_savedwin_data_111_port, 
                           curr_proc_regs(110) => 
                           DataPath_RF_bus_sel_savedwin_data_110_port, 
                           curr_proc_regs(109) => 
                           DataPath_RF_bus_sel_savedwin_data_109_port, 
                           curr_proc_regs(108) => 
                           DataPath_RF_bus_sel_savedwin_data_108_port, 
                           curr_proc_regs(107) => 
                           DataPath_RF_bus_sel_savedwin_data_107_port, 
                           curr_proc_regs(106) => 
                           DataPath_RF_bus_sel_savedwin_data_106_port, 
                           curr_proc_regs(105) => 
                           DataPath_RF_bus_sel_savedwin_data_105_port, 
                           curr_proc_regs(104) => 
                           DataPath_RF_bus_sel_savedwin_data_104_port, 
                           curr_proc_regs(103) => 
                           DataPath_RF_bus_sel_savedwin_data_103_port, 
                           curr_proc_regs(102) => 
                           DataPath_RF_bus_sel_savedwin_data_102_port, 
                           curr_proc_regs(101) => 
                           DataPath_RF_bus_sel_savedwin_data_101_port, 
                           curr_proc_regs(100) => 
                           DataPath_RF_bus_sel_savedwin_data_100_port, 
                           curr_proc_regs(99) => 
                           DataPath_RF_bus_sel_savedwin_data_99_port, 
                           curr_proc_regs(98) => 
                           DataPath_RF_bus_sel_savedwin_data_98_port, 
                           curr_proc_regs(97) => 
                           DataPath_RF_bus_sel_savedwin_data_97_port, 
                           curr_proc_regs(96) => 
                           DataPath_RF_bus_sel_savedwin_data_96_port, 
                           curr_proc_regs(95) => 
                           DataPath_RF_bus_sel_savedwin_data_95_port, 
                           curr_proc_regs(94) => 
                           DataPath_RF_bus_sel_savedwin_data_94_port, 
                           curr_proc_regs(93) => 
                           DataPath_RF_bus_sel_savedwin_data_93_port, 
                           curr_proc_regs(92) => 
                           DataPath_RF_bus_sel_savedwin_data_92_port, 
                           curr_proc_regs(91) => 
                           DataPath_RF_bus_sel_savedwin_data_91_port, 
                           curr_proc_regs(90) => 
                           DataPath_RF_bus_sel_savedwin_data_90_port, 
                           curr_proc_regs(89) => 
                           DataPath_RF_bus_sel_savedwin_data_89_port, 
                           curr_proc_regs(88) => 
                           DataPath_RF_bus_sel_savedwin_data_88_port, 
                           curr_proc_regs(87) => 
                           DataPath_RF_bus_sel_savedwin_data_87_port, 
                           curr_proc_regs(86) => 
                           DataPath_RF_bus_sel_savedwin_data_86_port, 
                           curr_proc_regs(85) => 
                           DataPath_RF_bus_sel_savedwin_data_85_port, 
                           curr_proc_regs(84) => 
                           DataPath_RF_bus_sel_savedwin_data_84_port, 
                           curr_proc_regs(83) => 
                           DataPath_RF_bus_sel_savedwin_data_83_port, 
                           curr_proc_regs(82) => 
                           DataPath_RF_bus_sel_savedwin_data_82_port, 
                           curr_proc_regs(81) => 
                           DataPath_RF_bus_sel_savedwin_data_81_port, 
                           curr_proc_regs(80) => 
                           DataPath_RF_bus_sel_savedwin_data_80_port, 
                           curr_proc_regs(79) => 
                           DataPath_RF_bus_sel_savedwin_data_79_port, 
                           curr_proc_regs(78) => 
                           DataPath_RF_bus_sel_savedwin_data_78_port, 
                           curr_proc_regs(77) => 
                           DataPath_RF_bus_sel_savedwin_data_77_port, 
                           curr_proc_regs(76) => 
                           DataPath_RF_bus_sel_savedwin_data_76_port, 
                           curr_proc_regs(75) => 
                           DataPath_RF_bus_sel_savedwin_data_75_port, 
                           curr_proc_regs(74) => 
                           DataPath_RF_bus_sel_savedwin_data_74_port, 
                           curr_proc_regs(73) => 
                           DataPath_RF_bus_sel_savedwin_data_73_port, 
                           curr_proc_regs(72) => 
                           DataPath_RF_bus_sel_savedwin_data_72_port, 
                           curr_proc_regs(71) => 
                           DataPath_RF_bus_sel_savedwin_data_71_port, 
                           curr_proc_regs(70) => 
                           DataPath_RF_bus_sel_savedwin_data_70_port, 
                           curr_proc_regs(69) => 
                           DataPath_RF_bus_sel_savedwin_data_69_port, 
                           curr_proc_regs(68) => 
                           DataPath_RF_bus_sel_savedwin_data_68_port, 
                           curr_proc_regs(67) => 
                           DataPath_RF_bus_sel_savedwin_data_67_port, 
                           curr_proc_regs(66) => 
                           DataPath_RF_bus_sel_savedwin_data_66_port, 
                           curr_proc_regs(65) => 
                           DataPath_RF_bus_sel_savedwin_data_65_port, 
                           curr_proc_regs(64) => 
                           DataPath_RF_bus_sel_savedwin_data_64_port, 
                           curr_proc_regs(63) => 
                           DataPath_RF_bus_sel_savedwin_data_63_port, 
                           curr_proc_regs(62) => 
                           DataPath_RF_bus_sel_savedwin_data_62_port, 
                           curr_proc_regs(61) => 
                           DataPath_RF_bus_sel_savedwin_data_61_port, 
                           curr_proc_regs(60) => 
                           DataPath_RF_bus_sel_savedwin_data_60_port, 
                           curr_proc_regs(59) => 
                           DataPath_RF_bus_sel_savedwin_data_59_port, 
                           curr_proc_regs(58) => 
                           DataPath_RF_bus_sel_savedwin_data_58_port, 
                           curr_proc_regs(57) => 
                           DataPath_RF_bus_sel_savedwin_data_57_port, 
                           curr_proc_regs(56) => 
                           DataPath_RF_bus_sel_savedwin_data_56_port, 
                           curr_proc_regs(55) => 
                           DataPath_RF_bus_sel_savedwin_data_55_port, 
                           curr_proc_regs(54) => 
                           DataPath_RF_bus_sel_savedwin_data_54_port, 
                           curr_proc_regs(53) => 
                           DataPath_RF_bus_sel_savedwin_data_53_port, 
                           curr_proc_regs(52) => 
                           DataPath_RF_bus_sel_savedwin_data_52_port, 
                           curr_proc_regs(51) => 
                           DataPath_RF_bus_sel_savedwin_data_51_port, 
                           curr_proc_regs(50) => 
                           DataPath_RF_bus_sel_savedwin_data_50_port, 
                           curr_proc_regs(49) => 
                           DataPath_RF_bus_sel_savedwin_data_49_port, 
                           curr_proc_regs(48) => 
                           DataPath_RF_bus_sel_savedwin_data_48_port, 
                           curr_proc_regs(47) => 
                           DataPath_RF_bus_sel_savedwin_data_47_port, 
                           curr_proc_regs(46) => 
                           DataPath_RF_bus_sel_savedwin_data_46_port, 
                           curr_proc_regs(45) => 
                           DataPath_RF_bus_sel_savedwin_data_45_port, 
                           curr_proc_regs(44) => 
                           DataPath_RF_bus_sel_savedwin_data_44_port, 
                           curr_proc_regs(43) => 
                           DataPath_RF_bus_sel_savedwin_data_43_port, 
                           curr_proc_regs(42) => 
                           DataPath_RF_bus_sel_savedwin_data_42_port, 
                           curr_proc_regs(41) => 
                           DataPath_RF_bus_sel_savedwin_data_41_port, 
                           curr_proc_regs(40) => 
                           DataPath_RF_bus_sel_savedwin_data_40_port, 
                           curr_proc_regs(39) => 
                           DataPath_RF_bus_sel_savedwin_data_39_port, 
                           curr_proc_regs(38) => 
                           DataPath_RF_bus_sel_savedwin_data_38_port, 
                           curr_proc_regs(37) => 
                           DataPath_RF_bus_sel_savedwin_data_37_port, 
                           curr_proc_regs(36) => 
                           DataPath_RF_bus_sel_savedwin_data_36_port, 
                           curr_proc_regs(35) => 
                           DataPath_RF_bus_sel_savedwin_data_35_port, 
                           curr_proc_regs(34) => 
                           DataPath_RF_bus_sel_savedwin_data_34_port, 
                           curr_proc_regs(33) => 
                           DataPath_RF_bus_sel_savedwin_data_33_port, 
                           curr_proc_regs(32) => 
                           DataPath_RF_bus_sel_savedwin_data_32_port, 
                           curr_proc_regs(31) => 
                           DataPath_RF_bus_sel_savedwin_data_31_port, 
                           curr_proc_regs(30) => 
                           DataPath_RF_bus_sel_savedwin_data_30_port, 
                           curr_proc_regs(29) => 
                           DataPath_RF_bus_sel_savedwin_data_29_port, 
                           curr_proc_regs(28) => 
                           DataPath_RF_bus_sel_savedwin_data_28_port, 
                           curr_proc_regs(27) => 
                           DataPath_RF_bus_sel_savedwin_data_27_port, 
                           curr_proc_regs(26) => 
                           DataPath_RF_bus_sel_savedwin_data_26_port, 
                           curr_proc_regs(25) => 
                           DataPath_RF_bus_sel_savedwin_data_25_port, 
                           curr_proc_regs(24) => 
                           DataPath_RF_bus_sel_savedwin_data_24_port, 
                           curr_proc_regs(23) => 
                           DataPath_RF_bus_sel_savedwin_data_23_port, 
                           curr_proc_regs(22) => 
                           DataPath_RF_bus_sel_savedwin_data_22_port, 
                           curr_proc_regs(21) => 
                           DataPath_RF_bus_sel_savedwin_data_21_port, 
                           curr_proc_regs(20) => 
                           DataPath_RF_bus_sel_savedwin_data_20_port, 
                           curr_proc_regs(19) => 
                           DataPath_RF_bus_sel_savedwin_data_19_port, 
                           curr_proc_regs(18) => 
                           DataPath_RF_bus_sel_savedwin_data_18_port, 
                           curr_proc_regs(17) => 
                           DataPath_RF_bus_sel_savedwin_data_17_port, 
                           curr_proc_regs(16) => 
                           DataPath_RF_bus_sel_savedwin_data_16_port, 
                           curr_proc_regs(15) => 
                           DataPath_RF_bus_sel_savedwin_data_15_port, 
                           curr_proc_regs(14) => 
                           DataPath_RF_bus_sel_savedwin_data_14_port, 
                           curr_proc_regs(13) => 
                           DataPath_RF_bus_sel_savedwin_data_13_port, 
                           curr_proc_regs(12) => 
                           DataPath_RF_bus_sel_savedwin_data_12_port, 
                           curr_proc_regs(11) => 
                           DataPath_RF_bus_sel_savedwin_data_11_port, 
                           curr_proc_regs(10) => 
                           DataPath_RF_bus_sel_savedwin_data_10_port, 
                           curr_proc_regs(9) => 
                           DataPath_RF_bus_sel_savedwin_data_9_port, 
                           curr_proc_regs(8) => 
                           DataPath_RF_bus_sel_savedwin_data_8_port, 
                           curr_proc_regs(7) => 
                           DataPath_RF_bus_sel_savedwin_data_7_port, 
                           curr_proc_regs(6) => 
                           DataPath_RF_bus_sel_savedwin_data_6_port, 
                           curr_proc_regs(5) => 
                           DataPath_RF_bus_sel_savedwin_data_5_port, 
                           curr_proc_regs(4) => 
                           DataPath_RF_bus_sel_savedwin_data_4_port, 
                           curr_proc_regs(3) => 
                           DataPath_RF_bus_sel_savedwin_data_3_port, 
                           curr_proc_regs(2) => 
                           DataPath_RF_bus_sel_savedwin_data_2_port, 
                           curr_proc_regs(1) => 
                           DataPath_RF_bus_sel_savedwin_data_1_port, 
                           curr_proc_regs(0) => 
                           DataPath_RF_bus_sel_savedwin_data_0_port);
   DataPath_RF_RDPORT1 : mux_N32_M5_1 port map( S(4) => n10863, S(3) => n10864,
                           S(2) => n10865, S(1) => n10866, S(0) => n10867, 
                           Q(1023) => 
                           DataPath_RF_bus_selected_win_data_767_port, Q(1022) 
                           => DataPath_RF_bus_selected_win_data_766_port, 
                           Q(1021) => 
                           DataPath_RF_bus_selected_win_data_765_port, Q(1020) 
                           => DataPath_RF_bus_selected_win_data_764_port, 
                           Q(1019) => 
                           DataPath_RF_bus_selected_win_data_763_port, Q(1018) 
                           => DataPath_RF_bus_selected_win_data_762_port, 
                           Q(1017) => 
                           DataPath_RF_bus_selected_win_data_761_port, Q(1016) 
                           => DataPath_RF_bus_selected_win_data_760_port, 
                           Q(1015) => 
                           DataPath_RF_bus_selected_win_data_759_port, Q(1014) 
                           => DataPath_RF_bus_selected_win_data_758_port, 
                           Q(1013) => 
                           DataPath_RF_bus_selected_win_data_757_port, Q(1012) 
                           => DataPath_RF_bus_selected_win_data_756_port, 
                           Q(1011) => 
                           DataPath_RF_bus_selected_win_data_755_port, Q(1010) 
                           => DataPath_RF_bus_selected_win_data_754_port, 
                           Q(1009) => 
                           DataPath_RF_bus_selected_win_data_753_port, Q(1008) 
                           => DataPath_RF_bus_selected_win_data_752_port, 
                           Q(1007) => 
                           DataPath_RF_bus_selected_win_data_751_port, Q(1006) 
                           => DataPath_RF_bus_selected_win_data_750_port, 
                           Q(1005) => 
                           DataPath_RF_bus_selected_win_data_749_port, Q(1004) 
                           => DataPath_RF_bus_selected_win_data_748_port, 
                           Q(1003) => 
                           DataPath_RF_bus_selected_win_data_747_port, Q(1002) 
                           => DataPath_RF_bus_selected_win_data_746_port, 
                           Q(1001) => 
                           DataPath_RF_bus_selected_win_data_745_port, Q(1000) 
                           => DataPath_RF_bus_selected_win_data_744_port, 
                           Q(999) => DataPath_RF_bus_selected_win_data_743_port
                           , Q(998) => 
                           DataPath_RF_bus_selected_win_data_742_port, Q(997) 
                           => DataPath_RF_bus_selected_win_data_741_port, 
                           Q(996) => DataPath_RF_bus_selected_win_data_740_port
                           , Q(995) => 
                           DataPath_RF_bus_selected_win_data_739_port, Q(994) 
                           => DataPath_RF_bus_selected_win_data_738_port, 
                           Q(993) => DataPath_RF_bus_selected_win_data_737_port
                           , Q(992) => 
                           DataPath_RF_bus_selected_win_data_736_port, Q(991) 
                           => DataPath_RF_bus_selected_win_data_735_port, 
                           Q(990) => DataPath_RF_bus_selected_win_data_734_port
                           , Q(989) => 
                           DataPath_RF_bus_selected_win_data_733_port, Q(988) 
                           => DataPath_RF_bus_selected_win_data_732_port, 
                           Q(987) => DataPath_RF_bus_selected_win_data_731_port
                           , Q(986) => 
                           DataPath_RF_bus_selected_win_data_730_port, Q(985) 
                           => DataPath_RF_bus_selected_win_data_729_port, 
                           Q(984) => DataPath_RF_bus_selected_win_data_728_port
                           , Q(983) => 
                           DataPath_RF_bus_selected_win_data_727_port, Q(982) 
                           => DataPath_RF_bus_selected_win_data_726_port, 
                           Q(981) => DataPath_RF_bus_selected_win_data_725_port
                           , Q(980) => 
                           DataPath_RF_bus_selected_win_data_724_port, Q(979) 
                           => DataPath_RF_bus_selected_win_data_723_port, 
                           Q(978) => DataPath_RF_bus_selected_win_data_722_port
                           , Q(977) => 
                           DataPath_RF_bus_selected_win_data_721_port, Q(976) 
                           => DataPath_RF_bus_selected_win_data_720_port, 
                           Q(975) => DataPath_RF_bus_selected_win_data_719_port
                           , Q(974) => 
                           DataPath_RF_bus_selected_win_data_718_port, Q(973) 
                           => DataPath_RF_bus_selected_win_data_717_port, 
                           Q(972) => DataPath_RF_bus_selected_win_data_716_port
                           , Q(971) => 
                           DataPath_RF_bus_selected_win_data_715_port, Q(970) 
                           => DataPath_RF_bus_selected_win_data_714_port, 
                           Q(969) => DataPath_RF_bus_selected_win_data_713_port
                           , Q(968) => 
                           DataPath_RF_bus_selected_win_data_712_port, Q(967) 
                           => DataPath_RF_bus_selected_win_data_711_port, 
                           Q(966) => DataPath_RF_bus_selected_win_data_710_port
                           , Q(965) => 
                           DataPath_RF_bus_selected_win_data_709_port, Q(964) 
                           => DataPath_RF_bus_selected_win_data_708_port, 
                           Q(963) => DataPath_RF_bus_selected_win_data_707_port
                           , Q(962) => 
                           DataPath_RF_bus_selected_win_data_706_port, Q(961) 
                           => DataPath_RF_bus_selected_win_data_705_port, 
                           Q(960) => DataPath_RF_bus_selected_win_data_704_port
                           , Q(959) => 
                           DataPath_RF_bus_selected_win_data_703_port, Q(958) 
                           => DataPath_RF_bus_selected_win_data_702_port, 
                           Q(957) => DataPath_RF_bus_selected_win_data_701_port
                           , Q(956) => 
                           DataPath_RF_bus_selected_win_data_700_port, Q(955) 
                           => DataPath_RF_bus_selected_win_data_699_port, 
                           Q(954) => DataPath_RF_bus_selected_win_data_698_port
                           , Q(953) => 
                           DataPath_RF_bus_selected_win_data_697_port, Q(952) 
                           => DataPath_RF_bus_selected_win_data_696_port, 
                           Q(951) => DataPath_RF_bus_selected_win_data_695_port
                           , Q(950) => 
                           DataPath_RF_bus_selected_win_data_694_port, Q(949) 
                           => DataPath_RF_bus_selected_win_data_693_port, 
                           Q(948) => DataPath_RF_bus_selected_win_data_692_port
                           , Q(947) => 
                           DataPath_RF_bus_selected_win_data_691_port, Q(946) 
                           => DataPath_RF_bus_selected_win_data_690_port, 
                           Q(945) => DataPath_RF_bus_selected_win_data_689_port
                           , Q(944) => 
                           DataPath_RF_bus_selected_win_data_688_port, Q(943) 
                           => DataPath_RF_bus_selected_win_data_687_port, 
                           Q(942) => DataPath_RF_bus_selected_win_data_686_port
                           , Q(941) => 
                           DataPath_RF_bus_selected_win_data_685_port, Q(940) 
                           => DataPath_RF_bus_selected_win_data_684_port, 
                           Q(939) => DataPath_RF_bus_selected_win_data_683_port
                           , Q(938) => 
                           DataPath_RF_bus_selected_win_data_682_port, Q(937) 
                           => DataPath_RF_bus_selected_win_data_681_port, 
                           Q(936) => DataPath_RF_bus_selected_win_data_680_port
                           , Q(935) => 
                           DataPath_RF_bus_selected_win_data_679_port, Q(934) 
                           => DataPath_RF_bus_selected_win_data_678_port, 
                           Q(933) => DataPath_RF_bus_selected_win_data_677_port
                           , Q(932) => 
                           DataPath_RF_bus_selected_win_data_676_port, Q(931) 
                           => DataPath_RF_bus_selected_win_data_675_port, 
                           Q(930) => DataPath_RF_bus_selected_win_data_674_port
                           , Q(929) => 
                           DataPath_RF_bus_selected_win_data_673_port, Q(928) 
                           => DataPath_RF_bus_selected_win_data_672_port, 
                           Q(927) => DataPath_RF_bus_selected_win_data_671_port
                           , Q(926) => 
                           DataPath_RF_bus_selected_win_data_670_port, Q(925) 
                           => DataPath_RF_bus_selected_win_data_669_port, 
                           Q(924) => DataPath_RF_bus_selected_win_data_668_port
                           , Q(923) => 
                           DataPath_RF_bus_selected_win_data_667_port, Q(922) 
                           => DataPath_RF_bus_selected_win_data_666_port, 
                           Q(921) => DataPath_RF_bus_selected_win_data_665_port
                           , Q(920) => 
                           DataPath_RF_bus_selected_win_data_664_port, Q(919) 
                           => DataPath_RF_bus_selected_win_data_663_port, 
                           Q(918) => DataPath_RF_bus_selected_win_data_662_port
                           , Q(917) => 
                           DataPath_RF_bus_selected_win_data_661_port, Q(916) 
                           => DataPath_RF_bus_selected_win_data_660_port, 
                           Q(915) => DataPath_RF_bus_selected_win_data_659_port
                           , Q(914) => 
                           DataPath_RF_bus_selected_win_data_658_port, Q(913) 
                           => DataPath_RF_bus_selected_win_data_657_port, 
                           Q(912) => DataPath_RF_bus_selected_win_data_656_port
                           , Q(911) => 
                           DataPath_RF_bus_selected_win_data_655_port, Q(910) 
                           => DataPath_RF_bus_selected_win_data_654_port, 
                           Q(909) => DataPath_RF_bus_selected_win_data_653_port
                           , Q(908) => 
                           DataPath_RF_bus_selected_win_data_652_port, Q(907) 
                           => DataPath_RF_bus_selected_win_data_651_port, 
                           Q(906) => DataPath_RF_bus_selected_win_data_650_port
                           , Q(905) => 
                           DataPath_RF_bus_selected_win_data_649_port, Q(904) 
                           => DataPath_RF_bus_selected_win_data_648_port, 
                           Q(903) => DataPath_RF_bus_selected_win_data_647_port
                           , Q(902) => 
                           DataPath_RF_bus_selected_win_data_646_port, Q(901) 
                           => DataPath_RF_bus_selected_win_data_645_port, 
                           Q(900) => DataPath_RF_bus_selected_win_data_644_port
                           , Q(899) => 
                           DataPath_RF_bus_selected_win_data_643_port, Q(898) 
                           => DataPath_RF_bus_selected_win_data_642_port, 
                           Q(897) => DataPath_RF_bus_selected_win_data_641_port
                           , Q(896) => 
                           DataPath_RF_bus_selected_win_data_640_port, Q(895) 
                           => DataPath_RF_bus_selected_win_data_639_port, 
                           Q(894) => DataPath_RF_bus_selected_win_data_638_port
                           , Q(893) => 
                           DataPath_RF_bus_selected_win_data_637_port, Q(892) 
                           => DataPath_RF_bus_selected_win_data_636_port, 
                           Q(891) => DataPath_RF_bus_selected_win_data_635_port
                           , Q(890) => 
                           DataPath_RF_bus_selected_win_data_634_port, Q(889) 
                           => DataPath_RF_bus_selected_win_data_633_port, 
                           Q(888) => DataPath_RF_bus_selected_win_data_632_port
                           , Q(887) => 
                           DataPath_RF_bus_selected_win_data_631_port, Q(886) 
                           => DataPath_RF_bus_selected_win_data_630_port, 
                           Q(885) => DataPath_RF_bus_selected_win_data_629_port
                           , Q(884) => 
                           DataPath_RF_bus_selected_win_data_628_port, Q(883) 
                           => DataPath_RF_bus_selected_win_data_627_port, 
                           Q(882) => DataPath_RF_bus_selected_win_data_626_port
                           , Q(881) => 
                           DataPath_RF_bus_selected_win_data_625_port, Q(880) 
                           => DataPath_RF_bus_selected_win_data_624_port, 
                           Q(879) => DataPath_RF_bus_selected_win_data_623_port
                           , Q(878) => 
                           DataPath_RF_bus_selected_win_data_622_port, Q(877) 
                           => DataPath_RF_bus_selected_win_data_621_port, 
                           Q(876) => DataPath_RF_bus_selected_win_data_620_port
                           , Q(875) => 
                           DataPath_RF_bus_selected_win_data_619_port, Q(874) 
                           => DataPath_RF_bus_selected_win_data_618_port, 
                           Q(873) => DataPath_RF_bus_selected_win_data_617_port
                           , Q(872) => 
                           DataPath_RF_bus_selected_win_data_616_port, Q(871) 
                           => DataPath_RF_bus_selected_win_data_615_port, 
                           Q(870) => DataPath_RF_bus_selected_win_data_614_port
                           , Q(869) => 
                           DataPath_RF_bus_selected_win_data_613_port, Q(868) 
                           => DataPath_RF_bus_selected_win_data_612_port, 
                           Q(867) => DataPath_RF_bus_selected_win_data_611_port
                           , Q(866) => 
                           DataPath_RF_bus_selected_win_data_610_port, Q(865) 
                           => DataPath_RF_bus_selected_win_data_609_port, 
                           Q(864) => DataPath_RF_bus_selected_win_data_608_port
                           , Q(863) => 
                           DataPath_RF_bus_selected_win_data_607_port, Q(862) 
                           => DataPath_RF_bus_selected_win_data_606_port, 
                           Q(861) => DataPath_RF_bus_selected_win_data_605_port
                           , Q(860) => 
                           DataPath_RF_bus_selected_win_data_604_port, Q(859) 
                           => DataPath_RF_bus_selected_win_data_603_port, 
                           Q(858) => DataPath_RF_bus_selected_win_data_602_port
                           , Q(857) => 
                           DataPath_RF_bus_selected_win_data_601_port, Q(856) 
                           => DataPath_RF_bus_selected_win_data_600_port, 
                           Q(855) => DataPath_RF_bus_selected_win_data_599_port
                           , Q(854) => 
                           DataPath_RF_bus_selected_win_data_598_port, Q(853) 
                           => DataPath_RF_bus_selected_win_data_597_port, 
                           Q(852) => DataPath_RF_bus_selected_win_data_596_port
                           , Q(851) => 
                           DataPath_RF_bus_selected_win_data_595_port, Q(850) 
                           => DataPath_RF_bus_selected_win_data_594_port, 
                           Q(849) => DataPath_RF_bus_selected_win_data_593_port
                           , Q(848) => 
                           DataPath_RF_bus_selected_win_data_592_port, Q(847) 
                           => DataPath_RF_bus_selected_win_data_591_port, 
                           Q(846) => DataPath_RF_bus_selected_win_data_590_port
                           , Q(845) => 
                           DataPath_RF_bus_selected_win_data_589_port, Q(844) 
                           => DataPath_RF_bus_selected_win_data_588_port, 
                           Q(843) => DataPath_RF_bus_selected_win_data_587_port
                           , Q(842) => 
                           DataPath_RF_bus_selected_win_data_586_port, Q(841) 
                           => DataPath_RF_bus_selected_win_data_585_port, 
                           Q(840) => DataPath_RF_bus_selected_win_data_584_port
                           , Q(839) => 
                           DataPath_RF_bus_selected_win_data_583_port, Q(838) 
                           => DataPath_RF_bus_selected_win_data_582_port, 
                           Q(837) => DataPath_RF_bus_selected_win_data_581_port
                           , Q(836) => 
                           DataPath_RF_bus_selected_win_data_580_port, Q(835) 
                           => DataPath_RF_bus_selected_win_data_579_port, 
                           Q(834) => DataPath_RF_bus_selected_win_data_578_port
                           , Q(833) => 
                           DataPath_RF_bus_selected_win_data_577_port, Q(832) 
                           => DataPath_RF_bus_selected_win_data_576_port, 
                           Q(831) => DataPath_RF_bus_selected_win_data_575_port
                           , Q(830) => 
                           DataPath_RF_bus_selected_win_data_574_port, Q(829) 
                           => DataPath_RF_bus_selected_win_data_573_port, 
                           Q(828) => DataPath_RF_bus_selected_win_data_572_port
                           , Q(827) => 
                           DataPath_RF_bus_selected_win_data_571_port, Q(826) 
                           => DataPath_RF_bus_selected_win_data_570_port, 
                           Q(825) => DataPath_RF_bus_selected_win_data_569_port
                           , Q(824) => 
                           DataPath_RF_bus_selected_win_data_568_port, Q(823) 
                           => DataPath_RF_bus_selected_win_data_567_port, 
                           Q(822) => DataPath_RF_bus_selected_win_data_566_port
                           , Q(821) => 
                           DataPath_RF_bus_selected_win_data_565_port, Q(820) 
                           => DataPath_RF_bus_selected_win_data_564_port, 
                           Q(819) => DataPath_RF_bus_selected_win_data_563_port
                           , Q(818) => 
                           DataPath_RF_bus_selected_win_data_562_port, Q(817) 
                           => DataPath_RF_bus_selected_win_data_561_port, 
                           Q(816) => DataPath_RF_bus_selected_win_data_560_port
                           , Q(815) => 
                           DataPath_RF_bus_selected_win_data_559_port, Q(814) 
                           => DataPath_RF_bus_selected_win_data_558_port, 
                           Q(813) => DataPath_RF_bus_selected_win_data_557_port
                           , Q(812) => 
                           DataPath_RF_bus_selected_win_data_556_port, Q(811) 
                           => DataPath_RF_bus_selected_win_data_555_port, 
                           Q(810) => DataPath_RF_bus_selected_win_data_554_port
                           , Q(809) => 
                           DataPath_RF_bus_selected_win_data_553_port, Q(808) 
                           => DataPath_RF_bus_selected_win_data_552_port, 
                           Q(807) => DataPath_RF_bus_selected_win_data_551_port
                           , Q(806) => 
                           DataPath_RF_bus_selected_win_data_550_port, Q(805) 
                           => DataPath_RF_bus_selected_win_data_549_port, 
                           Q(804) => DataPath_RF_bus_selected_win_data_548_port
                           , Q(803) => 
                           DataPath_RF_bus_selected_win_data_547_port, Q(802) 
                           => DataPath_RF_bus_selected_win_data_546_port, 
                           Q(801) => DataPath_RF_bus_selected_win_data_545_port
                           , Q(800) => 
                           DataPath_RF_bus_selected_win_data_544_port, Q(799) 
                           => DataPath_RF_bus_selected_win_data_543_port, 
                           Q(798) => DataPath_RF_bus_selected_win_data_542_port
                           , Q(797) => 
                           DataPath_RF_bus_selected_win_data_541_port, Q(796) 
                           => DataPath_RF_bus_selected_win_data_540_port, 
                           Q(795) => DataPath_RF_bus_selected_win_data_539_port
                           , Q(794) => 
                           DataPath_RF_bus_selected_win_data_538_port, Q(793) 
                           => DataPath_RF_bus_selected_win_data_537_port, 
                           Q(792) => DataPath_RF_bus_selected_win_data_536_port
                           , Q(791) => 
                           DataPath_RF_bus_selected_win_data_535_port, Q(790) 
                           => DataPath_RF_bus_selected_win_data_534_port, 
                           Q(789) => DataPath_RF_bus_selected_win_data_533_port
                           , Q(788) => 
                           DataPath_RF_bus_selected_win_data_532_port, Q(787) 
                           => DataPath_RF_bus_selected_win_data_531_port, 
                           Q(786) => DataPath_RF_bus_selected_win_data_530_port
                           , Q(785) => 
                           DataPath_RF_bus_selected_win_data_529_port, Q(784) 
                           => DataPath_RF_bus_selected_win_data_528_port, 
                           Q(783) => DataPath_RF_bus_selected_win_data_527_port
                           , Q(782) => 
                           DataPath_RF_bus_selected_win_data_526_port, Q(781) 
                           => DataPath_RF_bus_selected_win_data_525_port, 
                           Q(780) => DataPath_RF_bus_selected_win_data_524_port
                           , Q(779) => 
                           DataPath_RF_bus_selected_win_data_523_port, Q(778) 
                           => DataPath_RF_bus_selected_win_data_522_port, 
                           Q(777) => DataPath_RF_bus_selected_win_data_521_port
                           , Q(776) => 
                           DataPath_RF_bus_selected_win_data_520_port, Q(775) 
                           => DataPath_RF_bus_selected_win_data_519_port, 
                           Q(774) => DataPath_RF_bus_selected_win_data_518_port
                           , Q(773) => 
                           DataPath_RF_bus_selected_win_data_517_port, Q(772) 
                           => DataPath_RF_bus_selected_win_data_516_port, 
                           Q(771) => DataPath_RF_bus_selected_win_data_515_port
                           , Q(770) => 
                           DataPath_RF_bus_selected_win_data_514_port, Q(769) 
                           => DataPath_RF_bus_selected_win_data_513_port, 
                           Q(768) => DataPath_RF_bus_selected_win_data_512_port
                           , Q(767) => 
                           DataPath_RF_bus_selected_win_data_511_port, Q(766) 
                           => DataPath_RF_bus_selected_win_data_510_port, 
                           Q(765) => DataPath_RF_bus_selected_win_data_509_port
                           , Q(764) => 
                           DataPath_RF_bus_selected_win_data_508_port, Q(763) 
                           => DataPath_RF_bus_selected_win_data_507_port, 
                           Q(762) => DataPath_RF_bus_selected_win_data_506_port
                           , Q(761) => 
                           DataPath_RF_bus_selected_win_data_505_port, Q(760) 
                           => DataPath_RF_bus_selected_win_data_504_port, 
                           Q(759) => DataPath_RF_bus_selected_win_data_503_port
                           , Q(758) => 
                           DataPath_RF_bus_selected_win_data_502_port, Q(757) 
                           => DataPath_RF_bus_selected_win_data_501_port, 
                           Q(756) => DataPath_RF_bus_selected_win_data_500_port
                           , Q(755) => 
                           DataPath_RF_bus_selected_win_data_499_port, Q(754) 
                           => DataPath_RF_bus_selected_win_data_498_port, 
                           Q(753) => DataPath_RF_bus_selected_win_data_497_port
                           , Q(752) => 
                           DataPath_RF_bus_selected_win_data_496_port, Q(751) 
                           => DataPath_RF_bus_selected_win_data_495_port, 
                           Q(750) => DataPath_RF_bus_selected_win_data_494_port
                           , Q(749) => 
                           DataPath_RF_bus_selected_win_data_493_port, Q(748) 
                           => DataPath_RF_bus_selected_win_data_492_port, 
                           Q(747) => DataPath_RF_bus_selected_win_data_491_port
                           , Q(746) => 
                           DataPath_RF_bus_selected_win_data_490_port, Q(745) 
                           => DataPath_RF_bus_selected_win_data_489_port, 
                           Q(744) => DataPath_RF_bus_selected_win_data_488_port
                           , Q(743) => 
                           DataPath_RF_bus_selected_win_data_487_port, Q(742) 
                           => DataPath_RF_bus_selected_win_data_486_port, 
                           Q(741) => DataPath_RF_bus_selected_win_data_485_port
                           , Q(740) => 
                           DataPath_RF_bus_selected_win_data_484_port, Q(739) 
                           => DataPath_RF_bus_selected_win_data_483_port, 
                           Q(738) => DataPath_RF_bus_selected_win_data_482_port
                           , Q(737) => 
                           DataPath_RF_bus_selected_win_data_481_port, Q(736) 
                           => DataPath_RF_bus_selected_win_data_480_port, 
                           Q(735) => DataPath_RF_bus_selected_win_data_479_port
                           , Q(734) => 
                           DataPath_RF_bus_selected_win_data_478_port, Q(733) 
                           => DataPath_RF_bus_selected_win_data_477_port, 
                           Q(732) => DataPath_RF_bus_selected_win_data_476_port
                           , Q(731) => 
                           DataPath_RF_bus_selected_win_data_475_port, Q(730) 
                           => DataPath_RF_bus_selected_win_data_474_port, 
                           Q(729) => DataPath_RF_bus_selected_win_data_473_port
                           , Q(728) => 
                           DataPath_RF_bus_selected_win_data_472_port, Q(727) 
                           => DataPath_RF_bus_selected_win_data_471_port, 
                           Q(726) => DataPath_RF_bus_selected_win_data_470_port
                           , Q(725) => 
                           DataPath_RF_bus_selected_win_data_469_port, Q(724) 
                           => DataPath_RF_bus_selected_win_data_468_port, 
                           Q(723) => DataPath_RF_bus_selected_win_data_467_port
                           , Q(722) => 
                           DataPath_RF_bus_selected_win_data_466_port, Q(721) 
                           => DataPath_RF_bus_selected_win_data_465_port, 
                           Q(720) => DataPath_RF_bus_selected_win_data_464_port
                           , Q(719) => 
                           DataPath_RF_bus_selected_win_data_463_port, Q(718) 
                           => DataPath_RF_bus_selected_win_data_462_port, 
                           Q(717) => DataPath_RF_bus_selected_win_data_461_port
                           , Q(716) => 
                           DataPath_RF_bus_selected_win_data_460_port, Q(715) 
                           => DataPath_RF_bus_selected_win_data_459_port, 
                           Q(714) => DataPath_RF_bus_selected_win_data_458_port
                           , Q(713) => 
                           DataPath_RF_bus_selected_win_data_457_port, Q(712) 
                           => DataPath_RF_bus_selected_win_data_456_port, 
                           Q(711) => DataPath_RF_bus_selected_win_data_455_port
                           , Q(710) => 
                           DataPath_RF_bus_selected_win_data_454_port, Q(709) 
                           => DataPath_RF_bus_selected_win_data_453_port, 
                           Q(708) => DataPath_RF_bus_selected_win_data_452_port
                           , Q(707) => 
                           DataPath_RF_bus_selected_win_data_451_port, Q(706) 
                           => DataPath_RF_bus_selected_win_data_450_port, 
                           Q(705) => DataPath_RF_bus_selected_win_data_449_port
                           , Q(704) => 
                           DataPath_RF_bus_selected_win_data_448_port, Q(703) 
                           => DataPath_RF_bus_selected_win_data_447_port, 
                           Q(702) => DataPath_RF_bus_selected_win_data_446_port
                           , Q(701) => 
                           DataPath_RF_bus_selected_win_data_445_port, Q(700) 
                           => DataPath_RF_bus_selected_win_data_444_port, 
                           Q(699) => DataPath_RF_bus_selected_win_data_443_port
                           , Q(698) => 
                           DataPath_RF_bus_selected_win_data_442_port, Q(697) 
                           => DataPath_RF_bus_selected_win_data_441_port, 
                           Q(696) => DataPath_RF_bus_selected_win_data_440_port
                           , Q(695) => 
                           DataPath_RF_bus_selected_win_data_439_port, Q(694) 
                           => DataPath_RF_bus_selected_win_data_438_port, 
                           Q(693) => DataPath_RF_bus_selected_win_data_437_port
                           , Q(692) => 
                           DataPath_RF_bus_selected_win_data_436_port, Q(691) 
                           => DataPath_RF_bus_selected_win_data_435_port, 
                           Q(690) => DataPath_RF_bus_selected_win_data_434_port
                           , Q(689) => 
                           DataPath_RF_bus_selected_win_data_433_port, Q(688) 
                           => DataPath_RF_bus_selected_win_data_432_port, 
                           Q(687) => DataPath_RF_bus_selected_win_data_431_port
                           , Q(686) => 
                           DataPath_RF_bus_selected_win_data_430_port, Q(685) 
                           => DataPath_RF_bus_selected_win_data_429_port, 
                           Q(684) => DataPath_RF_bus_selected_win_data_428_port
                           , Q(683) => 
                           DataPath_RF_bus_selected_win_data_427_port, Q(682) 
                           => DataPath_RF_bus_selected_win_data_426_port, 
                           Q(681) => DataPath_RF_bus_selected_win_data_425_port
                           , Q(680) => 
                           DataPath_RF_bus_selected_win_data_424_port, Q(679) 
                           => DataPath_RF_bus_selected_win_data_423_port, 
                           Q(678) => DataPath_RF_bus_selected_win_data_422_port
                           , Q(677) => 
                           DataPath_RF_bus_selected_win_data_421_port, Q(676) 
                           => DataPath_RF_bus_selected_win_data_420_port, 
                           Q(675) => DataPath_RF_bus_selected_win_data_419_port
                           , Q(674) => 
                           DataPath_RF_bus_selected_win_data_418_port, Q(673) 
                           => DataPath_RF_bus_selected_win_data_417_port, 
                           Q(672) => DataPath_RF_bus_selected_win_data_416_port
                           , Q(671) => 
                           DataPath_RF_bus_selected_win_data_415_port, Q(670) 
                           => DataPath_RF_bus_selected_win_data_414_port, 
                           Q(669) => DataPath_RF_bus_selected_win_data_413_port
                           , Q(668) => 
                           DataPath_RF_bus_selected_win_data_412_port, Q(667) 
                           => DataPath_RF_bus_selected_win_data_411_port, 
                           Q(666) => DataPath_RF_bus_selected_win_data_410_port
                           , Q(665) => 
                           DataPath_RF_bus_selected_win_data_409_port, Q(664) 
                           => DataPath_RF_bus_selected_win_data_408_port, 
                           Q(663) => DataPath_RF_bus_selected_win_data_407_port
                           , Q(662) => 
                           DataPath_RF_bus_selected_win_data_406_port, Q(661) 
                           => DataPath_RF_bus_selected_win_data_405_port, 
                           Q(660) => DataPath_RF_bus_selected_win_data_404_port
                           , Q(659) => 
                           DataPath_RF_bus_selected_win_data_403_port, Q(658) 
                           => DataPath_RF_bus_selected_win_data_402_port, 
                           Q(657) => DataPath_RF_bus_selected_win_data_401_port
                           , Q(656) => 
                           DataPath_RF_bus_selected_win_data_400_port, Q(655) 
                           => DataPath_RF_bus_selected_win_data_399_port, 
                           Q(654) => DataPath_RF_bus_selected_win_data_398_port
                           , Q(653) => 
                           DataPath_RF_bus_selected_win_data_397_port, Q(652) 
                           => DataPath_RF_bus_selected_win_data_396_port, 
                           Q(651) => DataPath_RF_bus_selected_win_data_395_port
                           , Q(650) => 
                           DataPath_RF_bus_selected_win_data_394_port, Q(649) 
                           => DataPath_RF_bus_selected_win_data_393_port, 
                           Q(648) => DataPath_RF_bus_selected_win_data_392_port
                           , Q(647) => 
                           DataPath_RF_bus_selected_win_data_391_port, Q(646) 
                           => DataPath_RF_bus_selected_win_data_390_port, 
                           Q(645) => DataPath_RF_bus_selected_win_data_389_port
                           , Q(644) => 
                           DataPath_RF_bus_selected_win_data_388_port, Q(643) 
                           => DataPath_RF_bus_selected_win_data_387_port, 
                           Q(642) => DataPath_RF_bus_selected_win_data_386_port
                           , Q(641) => 
                           DataPath_RF_bus_selected_win_data_385_port, Q(640) 
                           => DataPath_RF_bus_selected_win_data_384_port, 
                           Q(639) => DataPath_RF_bus_selected_win_data_383_port
                           , Q(638) => 
                           DataPath_RF_bus_selected_win_data_382_port, Q(637) 
                           => DataPath_RF_bus_selected_win_data_381_port, 
                           Q(636) => DataPath_RF_bus_selected_win_data_380_port
                           , Q(635) => 
                           DataPath_RF_bus_selected_win_data_379_port, Q(634) 
                           => DataPath_RF_bus_selected_win_data_378_port, 
                           Q(633) => DataPath_RF_bus_selected_win_data_377_port
                           , Q(632) => 
                           DataPath_RF_bus_selected_win_data_376_port, Q(631) 
                           => DataPath_RF_bus_selected_win_data_375_port, 
                           Q(630) => DataPath_RF_bus_selected_win_data_374_port
                           , Q(629) => 
                           DataPath_RF_bus_selected_win_data_373_port, Q(628) 
                           => DataPath_RF_bus_selected_win_data_372_port, 
                           Q(627) => DataPath_RF_bus_selected_win_data_371_port
                           , Q(626) => 
                           DataPath_RF_bus_selected_win_data_370_port, Q(625) 
                           => DataPath_RF_bus_selected_win_data_369_port, 
                           Q(624) => DataPath_RF_bus_selected_win_data_368_port
                           , Q(623) => 
                           DataPath_RF_bus_selected_win_data_367_port, Q(622) 
                           => DataPath_RF_bus_selected_win_data_366_port, 
                           Q(621) => DataPath_RF_bus_selected_win_data_365_port
                           , Q(620) => 
                           DataPath_RF_bus_selected_win_data_364_port, Q(619) 
                           => DataPath_RF_bus_selected_win_data_363_port, 
                           Q(618) => DataPath_RF_bus_selected_win_data_362_port
                           , Q(617) => 
                           DataPath_RF_bus_selected_win_data_361_port, Q(616) 
                           => DataPath_RF_bus_selected_win_data_360_port, 
                           Q(615) => DataPath_RF_bus_selected_win_data_359_port
                           , Q(614) => 
                           DataPath_RF_bus_selected_win_data_358_port, Q(613) 
                           => DataPath_RF_bus_selected_win_data_357_port, 
                           Q(612) => DataPath_RF_bus_selected_win_data_356_port
                           , Q(611) => 
                           DataPath_RF_bus_selected_win_data_355_port, Q(610) 
                           => DataPath_RF_bus_selected_win_data_354_port, 
                           Q(609) => DataPath_RF_bus_selected_win_data_353_port
                           , Q(608) => 
                           DataPath_RF_bus_selected_win_data_352_port, Q(607) 
                           => DataPath_RF_bus_selected_win_data_351_port, 
                           Q(606) => DataPath_RF_bus_selected_win_data_350_port
                           , Q(605) => 
                           DataPath_RF_bus_selected_win_data_349_port, Q(604) 
                           => DataPath_RF_bus_selected_win_data_348_port, 
                           Q(603) => DataPath_RF_bus_selected_win_data_347_port
                           , Q(602) => 
                           DataPath_RF_bus_selected_win_data_346_port, Q(601) 
                           => DataPath_RF_bus_selected_win_data_345_port, 
                           Q(600) => DataPath_RF_bus_selected_win_data_344_port
                           , Q(599) => 
                           DataPath_RF_bus_selected_win_data_343_port, Q(598) 
                           => DataPath_RF_bus_selected_win_data_342_port, 
                           Q(597) => DataPath_RF_bus_selected_win_data_341_port
                           , Q(596) => 
                           DataPath_RF_bus_selected_win_data_340_port, Q(595) 
                           => DataPath_RF_bus_selected_win_data_339_port, 
                           Q(594) => DataPath_RF_bus_selected_win_data_338_port
                           , Q(593) => 
                           DataPath_RF_bus_selected_win_data_337_port, Q(592) 
                           => DataPath_RF_bus_selected_win_data_336_port, 
                           Q(591) => DataPath_RF_bus_selected_win_data_335_port
                           , Q(590) => 
                           DataPath_RF_bus_selected_win_data_334_port, Q(589) 
                           => DataPath_RF_bus_selected_win_data_333_port, 
                           Q(588) => DataPath_RF_bus_selected_win_data_332_port
                           , Q(587) => 
                           DataPath_RF_bus_selected_win_data_331_port, Q(586) 
                           => DataPath_RF_bus_selected_win_data_330_port, 
                           Q(585) => DataPath_RF_bus_selected_win_data_329_port
                           , Q(584) => 
                           DataPath_RF_bus_selected_win_data_328_port, Q(583) 
                           => DataPath_RF_bus_selected_win_data_327_port, 
                           Q(582) => DataPath_RF_bus_selected_win_data_326_port
                           , Q(581) => 
                           DataPath_RF_bus_selected_win_data_325_port, Q(580) 
                           => DataPath_RF_bus_selected_win_data_324_port, 
                           Q(579) => DataPath_RF_bus_selected_win_data_323_port
                           , Q(578) => 
                           DataPath_RF_bus_selected_win_data_322_port, Q(577) 
                           => DataPath_RF_bus_selected_win_data_321_port, 
                           Q(576) => DataPath_RF_bus_selected_win_data_320_port
                           , Q(575) => 
                           DataPath_RF_bus_selected_win_data_319_port, Q(574) 
                           => DataPath_RF_bus_selected_win_data_318_port, 
                           Q(573) => DataPath_RF_bus_selected_win_data_317_port
                           , Q(572) => 
                           DataPath_RF_bus_selected_win_data_316_port, Q(571) 
                           => DataPath_RF_bus_selected_win_data_315_port, 
                           Q(570) => DataPath_RF_bus_selected_win_data_314_port
                           , Q(569) => 
                           DataPath_RF_bus_selected_win_data_313_port, Q(568) 
                           => DataPath_RF_bus_selected_win_data_312_port, 
                           Q(567) => DataPath_RF_bus_selected_win_data_311_port
                           , Q(566) => 
                           DataPath_RF_bus_selected_win_data_310_port, Q(565) 
                           => DataPath_RF_bus_selected_win_data_309_port, 
                           Q(564) => DataPath_RF_bus_selected_win_data_308_port
                           , Q(563) => 
                           DataPath_RF_bus_selected_win_data_307_port, Q(562) 
                           => DataPath_RF_bus_selected_win_data_306_port, 
                           Q(561) => DataPath_RF_bus_selected_win_data_305_port
                           , Q(560) => 
                           DataPath_RF_bus_selected_win_data_304_port, Q(559) 
                           => DataPath_RF_bus_selected_win_data_303_port, 
                           Q(558) => DataPath_RF_bus_selected_win_data_302_port
                           , Q(557) => 
                           DataPath_RF_bus_selected_win_data_301_port, Q(556) 
                           => DataPath_RF_bus_selected_win_data_300_port, 
                           Q(555) => DataPath_RF_bus_selected_win_data_299_port
                           , Q(554) => 
                           DataPath_RF_bus_selected_win_data_298_port, Q(553) 
                           => DataPath_RF_bus_selected_win_data_297_port, 
                           Q(552) => DataPath_RF_bus_selected_win_data_296_port
                           , Q(551) => 
                           DataPath_RF_bus_selected_win_data_295_port, Q(550) 
                           => DataPath_RF_bus_selected_win_data_294_port, 
                           Q(549) => DataPath_RF_bus_selected_win_data_293_port
                           , Q(548) => 
                           DataPath_RF_bus_selected_win_data_292_port, Q(547) 
                           => DataPath_RF_bus_selected_win_data_291_port, 
                           Q(546) => DataPath_RF_bus_selected_win_data_290_port
                           , Q(545) => 
                           DataPath_RF_bus_selected_win_data_289_port, Q(544) 
                           => DataPath_RF_bus_selected_win_data_288_port, 
                           Q(543) => DataPath_RF_bus_selected_win_data_287_port
                           , Q(542) => 
                           DataPath_RF_bus_selected_win_data_286_port, Q(541) 
                           => DataPath_RF_bus_selected_win_data_285_port, 
                           Q(540) => DataPath_RF_bus_selected_win_data_284_port
                           , Q(539) => 
                           DataPath_RF_bus_selected_win_data_283_port, Q(538) 
                           => DataPath_RF_bus_selected_win_data_282_port, 
                           Q(537) => DataPath_RF_bus_selected_win_data_281_port
                           , Q(536) => 
                           DataPath_RF_bus_selected_win_data_280_port, Q(535) 
                           => DataPath_RF_bus_selected_win_data_279_port, 
                           Q(534) => DataPath_RF_bus_selected_win_data_278_port
                           , Q(533) => 
                           DataPath_RF_bus_selected_win_data_277_port, Q(532) 
                           => DataPath_RF_bus_selected_win_data_276_port, 
                           Q(531) => DataPath_RF_bus_selected_win_data_275_port
                           , Q(530) => 
                           DataPath_RF_bus_selected_win_data_274_port, Q(529) 
                           => DataPath_RF_bus_selected_win_data_273_port, 
                           Q(528) => DataPath_RF_bus_selected_win_data_272_port
                           , Q(527) => 
                           DataPath_RF_bus_selected_win_data_271_port, Q(526) 
                           => DataPath_RF_bus_selected_win_data_270_port, 
                           Q(525) => DataPath_RF_bus_selected_win_data_269_port
                           , Q(524) => 
                           DataPath_RF_bus_selected_win_data_268_port, Q(523) 
                           => DataPath_RF_bus_selected_win_data_267_port, 
                           Q(522) => DataPath_RF_bus_selected_win_data_266_port
                           , Q(521) => 
                           DataPath_RF_bus_selected_win_data_265_port, Q(520) 
                           => DataPath_RF_bus_selected_win_data_264_port, 
                           Q(519) => DataPath_RF_bus_selected_win_data_263_port
                           , Q(518) => 
                           DataPath_RF_bus_selected_win_data_262_port, Q(517) 
                           => DataPath_RF_bus_selected_win_data_261_port, 
                           Q(516) => DataPath_RF_bus_selected_win_data_260_port
                           , Q(515) => 
                           DataPath_RF_bus_selected_win_data_259_port, Q(514) 
                           => DataPath_RF_bus_selected_win_data_258_port, 
                           Q(513) => DataPath_RF_bus_selected_win_data_257_port
                           , Q(512) => 
                           DataPath_RF_bus_selected_win_data_256_port, Q(511) 
                           => DataPath_RF_bus_selected_win_data_255_port, 
                           Q(510) => DataPath_RF_bus_selected_win_data_254_port
                           , Q(509) => 
                           DataPath_RF_bus_selected_win_data_253_port, Q(508) 
                           => DataPath_RF_bus_selected_win_data_252_port, 
                           Q(507) => DataPath_RF_bus_selected_win_data_251_port
                           , Q(506) => 
                           DataPath_RF_bus_selected_win_data_250_port, Q(505) 
                           => DataPath_RF_bus_selected_win_data_249_port, 
                           Q(504) => DataPath_RF_bus_selected_win_data_248_port
                           , Q(503) => 
                           DataPath_RF_bus_selected_win_data_247_port, Q(502) 
                           => DataPath_RF_bus_selected_win_data_246_port, 
                           Q(501) => DataPath_RF_bus_selected_win_data_245_port
                           , Q(500) => 
                           DataPath_RF_bus_selected_win_data_244_port, Q(499) 
                           => DataPath_RF_bus_selected_win_data_243_port, 
                           Q(498) => DataPath_RF_bus_selected_win_data_242_port
                           , Q(497) => 
                           DataPath_RF_bus_selected_win_data_241_port, Q(496) 
                           => DataPath_RF_bus_selected_win_data_240_port, 
                           Q(495) => DataPath_RF_bus_selected_win_data_239_port
                           , Q(494) => 
                           DataPath_RF_bus_selected_win_data_238_port, Q(493) 
                           => DataPath_RF_bus_selected_win_data_237_port, 
                           Q(492) => DataPath_RF_bus_selected_win_data_236_port
                           , Q(491) => 
                           DataPath_RF_bus_selected_win_data_235_port, Q(490) 
                           => DataPath_RF_bus_selected_win_data_234_port, 
                           Q(489) => DataPath_RF_bus_selected_win_data_233_port
                           , Q(488) => 
                           DataPath_RF_bus_selected_win_data_232_port, Q(487) 
                           => DataPath_RF_bus_selected_win_data_231_port, 
                           Q(486) => DataPath_RF_bus_selected_win_data_230_port
                           , Q(485) => 
                           DataPath_RF_bus_selected_win_data_229_port, Q(484) 
                           => DataPath_RF_bus_selected_win_data_228_port, 
                           Q(483) => DataPath_RF_bus_selected_win_data_227_port
                           , Q(482) => 
                           DataPath_RF_bus_selected_win_data_226_port, Q(481) 
                           => DataPath_RF_bus_selected_win_data_225_port, 
                           Q(480) => DataPath_RF_bus_selected_win_data_224_port
                           , Q(479) => 
                           DataPath_RF_bus_selected_win_data_223_port, Q(478) 
                           => DataPath_RF_bus_selected_win_data_222_port, 
                           Q(477) => DataPath_RF_bus_selected_win_data_221_port
                           , Q(476) => 
                           DataPath_RF_bus_selected_win_data_220_port, Q(475) 
                           => DataPath_RF_bus_selected_win_data_219_port, 
                           Q(474) => DataPath_RF_bus_selected_win_data_218_port
                           , Q(473) => 
                           DataPath_RF_bus_selected_win_data_217_port, Q(472) 
                           => DataPath_RF_bus_selected_win_data_216_port, 
                           Q(471) => DataPath_RF_bus_selected_win_data_215_port
                           , Q(470) => 
                           DataPath_RF_bus_selected_win_data_214_port, Q(469) 
                           => DataPath_RF_bus_selected_win_data_213_port, 
                           Q(468) => DataPath_RF_bus_selected_win_data_212_port
                           , Q(467) => 
                           DataPath_RF_bus_selected_win_data_211_port, Q(466) 
                           => DataPath_RF_bus_selected_win_data_210_port, 
                           Q(465) => DataPath_RF_bus_selected_win_data_209_port
                           , Q(464) => 
                           DataPath_RF_bus_selected_win_data_208_port, Q(463) 
                           => DataPath_RF_bus_selected_win_data_207_port, 
                           Q(462) => DataPath_RF_bus_selected_win_data_206_port
                           , Q(461) => 
                           DataPath_RF_bus_selected_win_data_205_port, Q(460) 
                           => DataPath_RF_bus_selected_win_data_204_port, 
                           Q(459) => DataPath_RF_bus_selected_win_data_203_port
                           , Q(458) => 
                           DataPath_RF_bus_selected_win_data_202_port, Q(457) 
                           => DataPath_RF_bus_selected_win_data_201_port, 
                           Q(456) => DataPath_RF_bus_selected_win_data_200_port
                           , Q(455) => 
                           DataPath_RF_bus_selected_win_data_199_port, Q(454) 
                           => DataPath_RF_bus_selected_win_data_198_port, 
                           Q(453) => DataPath_RF_bus_selected_win_data_197_port
                           , Q(452) => 
                           DataPath_RF_bus_selected_win_data_196_port, Q(451) 
                           => DataPath_RF_bus_selected_win_data_195_port, 
                           Q(450) => DataPath_RF_bus_selected_win_data_194_port
                           , Q(449) => 
                           DataPath_RF_bus_selected_win_data_193_port, Q(448) 
                           => DataPath_RF_bus_selected_win_data_192_port, 
                           Q(447) => DataPath_RF_bus_selected_win_data_191_port
                           , Q(446) => 
                           DataPath_RF_bus_selected_win_data_190_port, Q(445) 
                           => DataPath_RF_bus_selected_win_data_189_port, 
                           Q(444) => DataPath_RF_bus_selected_win_data_188_port
                           , Q(443) => 
                           DataPath_RF_bus_selected_win_data_187_port, Q(442) 
                           => DataPath_RF_bus_selected_win_data_186_port, 
                           Q(441) => DataPath_RF_bus_selected_win_data_185_port
                           , Q(440) => 
                           DataPath_RF_bus_selected_win_data_184_port, Q(439) 
                           => DataPath_RF_bus_selected_win_data_183_port, 
                           Q(438) => DataPath_RF_bus_selected_win_data_182_port
                           , Q(437) => 
                           DataPath_RF_bus_selected_win_data_181_port, Q(436) 
                           => DataPath_RF_bus_selected_win_data_180_port, 
                           Q(435) => DataPath_RF_bus_selected_win_data_179_port
                           , Q(434) => 
                           DataPath_RF_bus_selected_win_data_178_port, Q(433) 
                           => DataPath_RF_bus_selected_win_data_177_port, 
                           Q(432) => DataPath_RF_bus_selected_win_data_176_port
                           , Q(431) => 
                           DataPath_RF_bus_selected_win_data_175_port, Q(430) 
                           => DataPath_RF_bus_selected_win_data_174_port, 
                           Q(429) => DataPath_RF_bus_selected_win_data_173_port
                           , Q(428) => 
                           DataPath_RF_bus_selected_win_data_172_port, Q(427) 
                           => DataPath_RF_bus_selected_win_data_171_port, 
                           Q(426) => DataPath_RF_bus_selected_win_data_170_port
                           , Q(425) => 
                           DataPath_RF_bus_selected_win_data_169_port, Q(424) 
                           => DataPath_RF_bus_selected_win_data_168_port, 
                           Q(423) => DataPath_RF_bus_selected_win_data_167_port
                           , Q(422) => 
                           DataPath_RF_bus_selected_win_data_166_port, Q(421) 
                           => DataPath_RF_bus_selected_win_data_165_port, 
                           Q(420) => DataPath_RF_bus_selected_win_data_164_port
                           , Q(419) => 
                           DataPath_RF_bus_selected_win_data_163_port, Q(418) 
                           => DataPath_RF_bus_selected_win_data_162_port, 
                           Q(417) => DataPath_RF_bus_selected_win_data_161_port
                           , Q(416) => 
                           DataPath_RF_bus_selected_win_data_160_port, Q(415) 
                           => DataPath_RF_bus_selected_win_data_159_port, 
                           Q(414) => DataPath_RF_bus_selected_win_data_158_port
                           , Q(413) => 
                           DataPath_RF_bus_selected_win_data_157_port, Q(412) 
                           => DataPath_RF_bus_selected_win_data_156_port, 
                           Q(411) => DataPath_RF_bus_selected_win_data_155_port
                           , Q(410) => 
                           DataPath_RF_bus_selected_win_data_154_port, Q(409) 
                           => DataPath_RF_bus_selected_win_data_153_port, 
                           Q(408) => DataPath_RF_bus_selected_win_data_152_port
                           , Q(407) => 
                           DataPath_RF_bus_selected_win_data_151_port, Q(406) 
                           => DataPath_RF_bus_selected_win_data_150_port, 
                           Q(405) => DataPath_RF_bus_selected_win_data_149_port
                           , Q(404) => 
                           DataPath_RF_bus_selected_win_data_148_port, Q(403) 
                           => DataPath_RF_bus_selected_win_data_147_port, 
                           Q(402) => DataPath_RF_bus_selected_win_data_146_port
                           , Q(401) => 
                           DataPath_RF_bus_selected_win_data_145_port, Q(400) 
                           => DataPath_RF_bus_selected_win_data_144_port, 
                           Q(399) => DataPath_RF_bus_selected_win_data_143_port
                           , Q(398) => 
                           DataPath_RF_bus_selected_win_data_142_port, Q(397) 
                           => DataPath_RF_bus_selected_win_data_141_port, 
                           Q(396) => DataPath_RF_bus_selected_win_data_140_port
                           , Q(395) => 
                           DataPath_RF_bus_selected_win_data_139_port, Q(394) 
                           => DataPath_RF_bus_selected_win_data_138_port, 
                           Q(393) => DataPath_RF_bus_selected_win_data_137_port
                           , Q(392) => 
                           DataPath_RF_bus_selected_win_data_136_port, Q(391) 
                           => DataPath_RF_bus_selected_win_data_135_port, 
                           Q(390) => DataPath_RF_bus_selected_win_data_134_port
                           , Q(389) => 
                           DataPath_RF_bus_selected_win_data_133_port, Q(388) 
                           => DataPath_RF_bus_selected_win_data_132_port, 
                           Q(387) => DataPath_RF_bus_selected_win_data_131_port
                           , Q(386) => 
                           DataPath_RF_bus_selected_win_data_130_port, Q(385) 
                           => DataPath_RF_bus_selected_win_data_129_port, 
                           Q(384) => DataPath_RF_bus_selected_win_data_128_port
                           , Q(383) => 
                           DataPath_RF_bus_selected_win_data_127_port, Q(382) 
                           => DataPath_RF_bus_selected_win_data_126_port, 
                           Q(381) => DataPath_RF_bus_selected_win_data_125_port
                           , Q(380) => 
                           DataPath_RF_bus_selected_win_data_124_port, Q(379) 
                           => DataPath_RF_bus_selected_win_data_123_port, 
                           Q(378) => DataPath_RF_bus_selected_win_data_122_port
                           , Q(377) => 
                           DataPath_RF_bus_selected_win_data_121_port, Q(376) 
                           => DataPath_RF_bus_selected_win_data_120_port, 
                           Q(375) => DataPath_RF_bus_selected_win_data_119_port
                           , Q(374) => 
                           DataPath_RF_bus_selected_win_data_118_port, Q(373) 
                           => DataPath_RF_bus_selected_win_data_117_port, 
                           Q(372) => DataPath_RF_bus_selected_win_data_116_port
                           , Q(371) => 
                           DataPath_RF_bus_selected_win_data_115_port, Q(370) 
                           => DataPath_RF_bus_selected_win_data_114_port, 
                           Q(369) => DataPath_RF_bus_selected_win_data_113_port
                           , Q(368) => 
                           DataPath_RF_bus_selected_win_data_112_port, Q(367) 
                           => DataPath_RF_bus_selected_win_data_111_port, 
                           Q(366) => DataPath_RF_bus_selected_win_data_110_port
                           , Q(365) => 
                           DataPath_RF_bus_selected_win_data_109_port, Q(364) 
                           => DataPath_RF_bus_selected_win_data_108_port, 
                           Q(363) => DataPath_RF_bus_selected_win_data_107_port
                           , Q(362) => 
                           DataPath_RF_bus_selected_win_data_106_port, Q(361) 
                           => DataPath_RF_bus_selected_win_data_105_port, 
                           Q(360) => DataPath_RF_bus_selected_win_data_104_port
                           , Q(359) => 
                           DataPath_RF_bus_selected_win_data_103_port, Q(358) 
                           => DataPath_RF_bus_selected_win_data_102_port, 
                           Q(357) => DataPath_RF_bus_selected_win_data_101_port
                           , Q(356) => 
                           DataPath_RF_bus_selected_win_data_100_port, Q(355) 
                           => DataPath_RF_bus_selected_win_data_99_port, Q(354)
                           => DataPath_RF_bus_selected_win_data_98_port, Q(353)
                           => DataPath_RF_bus_selected_win_data_97_port, Q(352)
                           => DataPath_RF_bus_selected_win_data_96_port, Q(351)
                           => DataPath_RF_bus_selected_win_data_95_port, Q(350)
                           => DataPath_RF_bus_selected_win_data_94_port, Q(349)
                           => DataPath_RF_bus_selected_win_data_93_port, Q(348)
                           => DataPath_RF_bus_selected_win_data_92_port, Q(347)
                           => DataPath_RF_bus_selected_win_data_91_port, Q(346)
                           => DataPath_RF_bus_selected_win_data_90_port, Q(345)
                           => DataPath_RF_bus_selected_win_data_89_port, Q(344)
                           => DataPath_RF_bus_selected_win_data_88_port, Q(343)
                           => DataPath_RF_bus_selected_win_data_87_port, Q(342)
                           => DataPath_RF_bus_selected_win_data_86_port, Q(341)
                           => DataPath_RF_bus_selected_win_data_85_port, Q(340)
                           => DataPath_RF_bus_selected_win_data_84_port, Q(339)
                           => DataPath_RF_bus_selected_win_data_83_port, Q(338)
                           => DataPath_RF_bus_selected_win_data_82_port, Q(337)
                           => DataPath_RF_bus_selected_win_data_81_port, Q(336)
                           => DataPath_RF_bus_selected_win_data_80_port, Q(335)
                           => DataPath_RF_bus_selected_win_data_79_port, Q(334)
                           => DataPath_RF_bus_selected_win_data_78_port, Q(333)
                           => DataPath_RF_bus_selected_win_data_77_port, Q(332)
                           => DataPath_RF_bus_selected_win_data_76_port, Q(331)
                           => DataPath_RF_bus_selected_win_data_75_port, Q(330)
                           => DataPath_RF_bus_selected_win_data_74_port, Q(329)
                           => DataPath_RF_bus_selected_win_data_73_port, Q(328)
                           => DataPath_RF_bus_selected_win_data_72_port, Q(327)
                           => DataPath_RF_bus_selected_win_data_71_port, Q(326)
                           => DataPath_RF_bus_selected_win_data_70_port, Q(325)
                           => DataPath_RF_bus_selected_win_data_69_port, Q(324)
                           => DataPath_RF_bus_selected_win_data_68_port, Q(323)
                           => DataPath_RF_bus_selected_win_data_67_port, Q(322)
                           => DataPath_RF_bus_selected_win_data_66_port, Q(321)
                           => DataPath_RF_bus_selected_win_data_65_port, Q(320)
                           => DataPath_RF_bus_selected_win_data_64_port, Q(319)
                           => DataPath_RF_bus_selected_win_data_63_port, Q(318)
                           => DataPath_RF_bus_selected_win_data_62_port, Q(317)
                           => DataPath_RF_bus_selected_win_data_61_port, Q(316)
                           => DataPath_RF_bus_selected_win_data_60_port, Q(315)
                           => DataPath_RF_bus_selected_win_data_59_port, Q(314)
                           => DataPath_RF_bus_selected_win_data_58_port, Q(313)
                           => DataPath_RF_bus_selected_win_data_57_port, Q(312)
                           => DataPath_RF_bus_selected_win_data_56_port, Q(311)
                           => DataPath_RF_bus_selected_win_data_55_port, Q(310)
                           => DataPath_RF_bus_selected_win_data_54_port, Q(309)
                           => DataPath_RF_bus_selected_win_data_53_port, Q(308)
                           => DataPath_RF_bus_selected_win_data_52_port, Q(307)
                           => DataPath_RF_bus_selected_win_data_51_port, Q(306)
                           => DataPath_RF_bus_selected_win_data_50_port, Q(305)
                           => DataPath_RF_bus_selected_win_data_49_port, Q(304)
                           => DataPath_RF_bus_selected_win_data_48_port, Q(303)
                           => DataPath_RF_bus_selected_win_data_47_port, Q(302)
                           => DataPath_RF_bus_selected_win_data_46_port, Q(301)
                           => DataPath_RF_bus_selected_win_data_45_port, Q(300)
                           => DataPath_RF_bus_selected_win_data_44_port, Q(299)
                           => DataPath_RF_bus_selected_win_data_43_port, Q(298)
                           => DataPath_RF_bus_selected_win_data_42_port, Q(297)
                           => DataPath_RF_bus_selected_win_data_41_port, Q(296)
                           => DataPath_RF_bus_selected_win_data_40_port, Q(295)
                           => DataPath_RF_bus_selected_win_data_39_port, Q(294)
                           => DataPath_RF_bus_selected_win_data_38_port, Q(293)
                           => DataPath_RF_bus_selected_win_data_37_port, Q(292)
                           => DataPath_RF_bus_selected_win_data_36_port, Q(291)
                           => DataPath_RF_bus_selected_win_data_35_port, Q(290)
                           => DataPath_RF_bus_selected_win_data_34_port, Q(289)
                           => DataPath_RF_bus_selected_win_data_33_port, Q(288)
                           => DataPath_RF_bus_selected_win_data_32_port, Q(287)
                           => DataPath_RF_bus_selected_win_data_31_port, Q(286)
                           => DataPath_RF_bus_selected_win_data_30_port, Q(285)
                           => DataPath_RF_bus_selected_win_data_29_port, Q(284)
                           => DataPath_RF_bus_selected_win_data_28_port, Q(283)
                           => DataPath_RF_bus_selected_win_data_27_port, Q(282)
                           => DataPath_RF_bus_selected_win_data_26_port, Q(281)
                           => DataPath_RF_bus_selected_win_data_25_port, Q(280)
                           => DataPath_RF_bus_selected_win_data_24_port, Q(279)
                           => DataPath_RF_bus_selected_win_data_23_port, Q(278)
                           => DataPath_RF_bus_selected_win_data_22_port, Q(277)
                           => DataPath_RF_bus_selected_win_data_21_port, Q(276)
                           => DataPath_RF_bus_selected_win_data_20_port, Q(275)
                           => DataPath_RF_bus_selected_win_data_19_port, Q(274)
                           => DataPath_RF_bus_selected_win_data_18_port, Q(273)
                           => DataPath_RF_bus_selected_win_data_17_port, Q(272)
                           => DataPath_RF_bus_selected_win_data_16_port, Q(271)
                           => DataPath_RF_bus_selected_win_data_15_port, Q(270)
                           => DataPath_RF_bus_selected_win_data_14_port, Q(269)
                           => DataPath_RF_bus_selected_win_data_13_port, Q(268)
                           => DataPath_RF_bus_selected_win_data_12_port, Q(267)
                           => DataPath_RF_bus_selected_win_data_11_port, Q(266)
                           => DataPath_RF_bus_selected_win_data_10_port, Q(265)
                           => DataPath_RF_bus_selected_win_data_9_port, Q(264) 
                           => DataPath_RF_bus_selected_win_data_8_port, Q(263) 
                           => DataPath_RF_bus_selected_win_data_7_port, Q(262) 
                           => DataPath_RF_bus_selected_win_data_6_port, Q(261) 
                           => DataPath_RF_bus_selected_win_data_5_port, Q(260) 
                           => DataPath_RF_bus_selected_win_data_4_port, Q(259) 
                           => DataPath_RF_bus_selected_win_data_3_port, Q(258) 
                           => DataPath_RF_bus_selected_win_data_2_port, Q(257) 
                           => DataPath_RF_bus_selected_win_data_1_port, Q(256) 
                           => DataPath_RF_bus_selected_win_data_0_port, Q(255) 
                           => DataPath_RF_bus_complete_win_data_255_port, 
                           Q(254) => DataPath_RF_bus_complete_win_data_254_port
                           , Q(253) => 
                           DataPath_RF_bus_complete_win_data_253_port, Q(252) 
                           => DataPath_RF_bus_complete_win_data_252_port, 
                           Q(251) => DataPath_RF_bus_complete_win_data_251_port
                           , Q(250) => 
                           DataPath_RF_bus_complete_win_data_250_port, Q(249) 
                           => DataPath_RF_bus_complete_win_data_249_port, 
                           Q(248) => DataPath_RF_bus_complete_win_data_248_port
                           , Q(247) => 
                           DataPath_RF_bus_complete_win_data_247_port, Q(246) 
                           => DataPath_RF_bus_complete_win_data_246_port, 
                           Q(245) => DataPath_RF_bus_complete_win_data_245_port
                           , Q(244) => 
                           DataPath_RF_bus_complete_win_data_244_port, Q(243) 
                           => DataPath_RF_bus_complete_win_data_243_port, 
                           Q(242) => DataPath_RF_bus_complete_win_data_242_port
                           , Q(241) => 
                           DataPath_RF_bus_complete_win_data_241_port, Q(240) 
                           => DataPath_RF_bus_complete_win_data_240_port, 
                           Q(239) => DataPath_RF_bus_complete_win_data_239_port
                           , Q(238) => 
                           DataPath_RF_bus_complete_win_data_238_port, Q(237) 
                           => DataPath_RF_bus_complete_win_data_237_port, 
                           Q(236) => DataPath_RF_bus_complete_win_data_236_port
                           , Q(235) => 
                           DataPath_RF_bus_complete_win_data_235_port, Q(234) 
                           => DataPath_RF_bus_complete_win_data_234_port, 
                           Q(233) => DataPath_RF_bus_complete_win_data_233_port
                           , Q(232) => 
                           DataPath_RF_bus_complete_win_data_232_port, Q(231) 
                           => DataPath_RF_bus_complete_win_data_231_port, 
                           Q(230) => DataPath_RF_bus_complete_win_data_230_port
                           , Q(229) => 
                           DataPath_RF_bus_complete_win_data_229_port, Q(228) 
                           => DataPath_RF_bus_complete_win_data_228_port, 
                           Q(227) => DataPath_RF_bus_complete_win_data_227_port
                           , Q(226) => 
                           DataPath_RF_bus_complete_win_data_226_port, Q(225) 
                           => DataPath_RF_bus_complete_win_data_225_port, 
                           Q(224) => DataPath_RF_bus_complete_win_data_224_port
                           , Q(223) => 
                           DataPath_RF_bus_complete_win_data_223_port, Q(222) 
                           => DataPath_RF_bus_complete_win_data_222_port, 
                           Q(221) => DataPath_RF_bus_complete_win_data_221_port
                           , Q(220) => 
                           DataPath_RF_bus_complete_win_data_220_port, Q(219) 
                           => DataPath_RF_bus_complete_win_data_219_port, 
                           Q(218) => DataPath_RF_bus_complete_win_data_218_port
                           , Q(217) => 
                           DataPath_RF_bus_complete_win_data_217_port, Q(216) 
                           => DataPath_RF_bus_complete_win_data_216_port, 
                           Q(215) => DataPath_RF_bus_complete_win_data_215_port
                           , Q(214) => 
                           DataPath_RF_bus_complete_win_data_214_port, Q(213) 
                           => DataPath_RF_bus_complete_win_data_213_port, 
                           Q(212) => DataPath_RF_bus_complete_win_data_212_port
                           , Q(211) => 
                           DataPath_RF_bus_complete_win_data_211_port, Q(210) 
                           => DataPath_RF_bus_complete_win_data_210_port, 
                           Q(209) => DataPath_RF_bus_complete_win_data_209_port
                           , Q(208) => 
                           DataPath_RF_bus_complete_win_data_208_port, Q(207) 
                           => DataPath_RF_bus_complete_win_data_207_port, 
                           Q(206) => DataPath_RF_bus_complete_win_data_206_port
                           , Q(205) => 
                           DataPath_RF_bus_complete_win_data_205_port, Q(204) 
                           => DataPath_RF_bus_complete_win_data_204_port, 
                           Q(203) => DataPath_RF_bus_complete_win_data_203_port
                           , Q(202) => 
                           DataPath_RF_bus_complete_win_data_202_port, Q(201) 
                           => DataPath_RF_bus_complete_win_data_201_port, 
                           Q(200) => DataPath_RF_bus_complete_win_data_200_port
                           , Q(199) => 
                           DataPath_RF_bus_complete_win_data_199_port, Q(198) 
                           => DataPath_RF_bus_complete_win_data_198_port, 
                           Q(197) => DataPath_RF_bus_complete_win_data_197_port
                           , Q(196) => 
                           DataPath_RF_bus_complete_win_data_196_port, Q(195) 
                           => DataPath_RF_bus_complete_win_data_195_port, 
                           Q(194) => DataPath_RF_bus_complete_win_data_194_port
                           , Q(193) => 
                           DataPath_RF_bus_complete_win_data_193_port, Q(192) 
                           => DataPath_RF_bus_complete_win_data_192_port, 
                           Q(191) => DataPath_RF_bus_complete_win_data_191_port
                           , Q(190) => 
                           DataPath_RF_bus_complete_win_data_190_port, Q(189) 
                           => DataPath_RF_bus_complete_win_data_189_port, 
                           Q(188) => DataPath_RF_bus_complete_win_data_188_port
                           , Q(187) => 
                           DataPath_RF_bus_complete_win_data_187_port, Q(186) 
                           => DataPath_RF_bus_complete_win_data_186_port, 
                           Q(185) => DataPath_RF_bus_complete_win_data_185_port
                           , Q(184) => 
                           DataPath_RF_bus_complete_win_data_184_port, Q(183) 
                           => DataPath_RF_bus_complete_win_data_183_port, 
                           Q(182) => DataPath_RF_bus_complete_win_data_182_port
                           , Q(181) => 
                           DataPath_RF_bus_complete_win_data_181_port, Q(180) 
                           => DataPath_RF_bus_complete_win_data_180_port, 
                           Q(179) => DataPath_RF_bus_complete_win_data_179_port
                           , Q(178) => 
                           DataPath_RF_bus_complete_win_data_178_port, Q(177) 
                           => DataPath_RF_bus_complete_win_data_177_port, 
                           Q(176) => DataPath_RF_bus_complete_win_data_176_port
                           , Q(175) => 
                           DataPath_RF_bus_complete_win_data_175_port, Q(174) 
                           => DataPath_RF_bus_complete_win_data_174_port, 
                           Q(173) => DataPath_RF_bus_complete_win_data_173_port
                           , Q(172) => 
                           DataPath_RF_bus_complete_win_data_172_port, Q(171) 
                           => DataPath_RF_bus_complete_win_data_171_port, 
                           Q(170) => DataPath_RF_bus_complete_win_data_170_port
                           , Q(169) => 
                           DataPath_RF_bus_complete_win_data_169_port, Q(168) 
                           => DataPath_RF_bus_complete_win_data_168_port, 
                           Q(167) => DataPath_RF_bus_complete_win_data_167_port
                           , Q(166) => 
                           DataPath_RF_bus_complete_win_data_166_port, Q(165) 
                           => DataPath_RF_bus_complete_win_data_165_port, 
                           Q(164) => DataPath_RF_bus_complete_win_data_164_port
                           , Q(163) => 
                           DataPath_RF_bus_complete_win_data_163_port, Q(162) 
                           => DataPath_RF_bus_complete_win_data_162_port, 
                           Q(161) => DataPath_RF_bus_complete_win_data_161_port
                           , Q(160) => 
                           DataPath_RF_bus_complete_win_data_160_port, Q(159) 
                           => DataPath_RF_bus_complete_win_data_159_port, 
                           Q(158) => DataPath_RF_bus_complete_win_data_158_port
                           , Q(157) => 
                           DataPath_RF_bus_complete_win_data_157_port, Q(156) 
                           => DataPath_RF_bus_complete_win_data_156_port, 
                           Q(155) => DataPath_RF_bus_complete_win_data_155_port
                           , Q(154) => 
                           DataPath_RF_bus_complete_win_data_154_port, Q(153) 
                           => DataPath_RF_bus_complete_win_data_153_port, 
                           Q(152) => DataPath_RF_bus_complete_win_data_152_port
                           , Q(151) => 
                           DataPath_RF_bus_complete_win_data_151_port, Q(150) 
                           => DataPath_RF_bus_complete_win_data_150_port, 
                           Q(149) => DataPath_RF_bus_complete_win_data_149_port
                           , Q(148) => 
                           DataPath_RF_bus_complete_win_data_148_port, Q(147) 
                           => DataPath_RF_bus_complete_win_data_147_port, 
                           Q(146) => DataPath_RF_bus_complete_win_data_146_port
                           , Q(145) => 
                           DataPath_RF_bus_complete_win_data_145_port, Q(144) 
                           => DataPath_RF_bus_complete_win_data_144_port, 
                           Q(143) => DataPath_RF_bus_complete_win_data_143_port
                           , Q(142) => 
                           DataPath_RF_bus_complete_win_data_142_port, Q(141) 
                           => DataPath_RF_bus_complete_win_data_141_port, 
                           Q(140) => DataPath_RF_bus_complete_win_data_140_port
                           , Q(139) => 
                           DataPath_RF_bus_complete_win_data_139_port, Q(138) 
                           => DataPath_RF_bus_complete_win_data_138_port, 
                           Q(137) => DataPath_RF_bus_complete_win_data_137_port
                           , Q(136) => 
                           DataPath_RF_bus_complete_win_data_136_port, Q(135) 
                           => DataPath_RF_bus_complete_win_data_135_port, 
                           Q(134) => DataPath_RF_bus_complete_win_data_134_port
                           , Q(133) => 
                           DataPath_RF_bus_complete_win_data_133_port, Q(132) 
                           => DataPath_RF_bus_complete_win_data_132_port, 
                           Q(131) => DataPath_RF_bus_complete_win_data_131_port
                           , Q(130) => 
                           DataPath_RF_bus_complete_win_data_130_port, Q(129) 
                           => DataPath_RF_bus_complete_win_data_129_port, 
                           Q(128) => DataPath_RF_bus_complete_win_data_128_port
                           , Q(127) => 
                           DataPath_RF_bus_complete_win_data_127_port, Q(126) 
                           => DataPath_RF_bus_complete_win_data_126_port, 
                           Q(125) => DataPath_RF_bus_complete_win_data_125_port
                           , Q(124) => 
                           DataPath_RF_bus_complete_win_data_124_port, Q(123) 
                           => DataPath_RF_bus_complete_win_data_123_port, 
                           Q(122) => DataPath_RF_bus_complete_win_data_122_port
                           , Q(121) => 
                           DataPath_RF_bus_complete_win_data_121_port, Q(120) 
                           => DataPath_RF_bus_complete_win_data_120_port, 
                           Q(119) => DataPath_RF_bus_complete_win_data_119_port
                           , Q(118) => 
                           DataPath_RF_bus_complete_win_data_118_port, Q(117) 
                           => DataPath_RF_bus_complete_win_data_117_port, 
                           Q(116) => DataPath_RF_bus_complete_win_data_116_port
                           , Q(115) => 
                           DataPath_RF_bus_complete_win_data_115_port, Q(114) 
                           => DataPath_RF_bus_complete_win_data_114_port, 
                           Q(113) => DataPath_RF_bus_complete_win_data_113_port
                           , Q(112) => 
                           DataPath_RF_bus_complete_win_data_112_port, Q(111) 
                           => DataPath_RF_bus_complete_win_data_111_port, 
                           Q(110) => DataPath_RF_bus_complete_win_data_110_port
                           , Q(109) => 
                           DataPath_RF_bus_complete_win_data_109_port, Q(108) 
                           => DataPath_RF_bus_complete_win_data_108_port, 
                           Q(107) => DataPath_RF_bus_complete_win_data_107_port
                           , Q(106) => 
                           DataPath_RF_bus_complete_win_data_106_port, Q(105) 
                           => DataPath_RF_bus_complete_win_data_105_port, 
                           Q(104) => DataPath_RF_bus_complete_win_data_104_port
                           , Q(103) => 
                           DataPath_RF_bus_complete_win_data_103_port, Q(102) 
                           => DataPath_RF_bus_complete_win_data_102_port, 
                           Q(101) => DataPath_RF_bus_complete_win_data_101_port
                           , Q(100) => 
                           DataPath_RF_bus_complete_win_data_100_port, Q(99) =>
                           DataPath_RF_bus_complete_win_data_99_port, Q(98) => 
                           DataPath_RF_bus_complete_win_data_98_port, Q(97) => 
                           DataPath_RF_bus_complete_win_data_97_port, Q(96) => 
                           DataPath_RF_bus_complete_win_data_96_port, Q(95) => 
                           DataPath_RF_bus_complete_win_data_95_port, Q(94) => 
                           DataPath_RF_bus_complete_win_data_94_port, Q(93) => 
                           DataPath_RF_bus_complete_win_data_93_port, Q(92) => 
                           DataPath_RF_bus_complete_win_data_92_port, Q(91) => 
                           DataPath_RF_bus_complete_win_data_91_port, Q(90) => 
                           DataPath_RF_bus_complete_win_data_90_port, Q(89) => 
                           DataPath_RF_bus_complete_win_data_89_port, Q(88) => 
                           DataPath_RF_bus_complete_win_data_88_port, Q(87) => 
                           DataPath_RF_bus_complete_win_data_87_port, Q(86) => 
                           DataPath_RF_bus_complete_win_data_86_port, Q(85) => 
                           DataPath_RF_bus_complete_win_data_85_port, Q(84) => 
                           DataPath_RF_bus_complete_win_data_84_port, Q(83) => 
                           DataPath_RF_bus_complete_win_data_83_port, Q(82) => 
                           DataPath_RF_bus_complete_win_data_82_port, Q(81) => 
                           DataPath_RF_bus_complete_win_data_81_port, Q(80) => 
                           DataPath_RF_bus_complete_win_data_80_port, Q(79) => 
                           DataPath_RF_bus_complete_win_data_79_port, Q(78) => 
                           DataPath_RF_bus_complete_win_data_78_port, Q(77) => 
                           DataPath_RF_bus_complete_win_data_77_port, Q(76) => 
                           DataPath_RF_bus_complete_win_data_76_port, Q(75) => 
                           DataPath_RF_bus_complete_win_data_75_port, Q(74) => 
                           DataPath_RF_bus_complete_win_data_74_port, Q(73) => 
                           DataPath_RF_bus_complete_win_data_73_port, Q(72) => 
                           DataPath_RF_bus_complete_win_data_72_port, Q(71) => 
                           DataPath_RF_bus_complete_win_data_71_port, Q(70) => 
                           DataPath_RF_bus_complete_win_data_70_port, Q(69) => 
                           DataPath_RF_bus_complete_win_data_69_port, Q(68) => 
                           DataPath_RF_bus_complete_win_data_68_port, Q(67) => 
                           DataPath_RF_bus_complete_win_data_67_port, Q(66) => 
                           DataPath_RF_bus_complete_win_data_66_port, Q(65) => 
                           DataPath_RF_bus_complete_win_data_65_port, Q(64) => 
                           DataPath_RF_bus_complete_win_data_64_port, Q(63) => 
                           DataPath_RF_bus_complete_win_data_63_port, Q(62) => 
                           DataPath_RF_bus_complete_win_data_62_port, Q(61) => 
                           DataPath_RF_bus_complete_win_data_61_port, Q(60) => 
                           DataPath_RF_bus_complete_win_data_60_port, Q(59) => 
                           DataPath_RF_bus_complete_win_data_59_port, Q(58) => 
                           DataPath_RF_bus_complete_win_data_58_port, Q(57) => 
                           DataPath_RF_bus_complete_win_data_57_port, Q(56) => 
                           DataPath_RF_bus_complete_win_data_56_port, Q(55) => 
                           DataPath_RF_bus_complete_win_data_55_port, Q(54) => 
                           DataPath_RF_bus_complete_win_data_54_port, Q(53) => 
                           DataPath_RF_bus_complete_win_data_53_port, Q(52) => 
                           DataPath_RF_bus_complete_win_data_52_port, Q(51) => 
                           DataPath_RF_bus_complete_win_data_51_port, Q(50) => 
                           DataPath_RF_bus_complete_win_data_50_port, Q(49) => 
                           DataPath_RF_bus_complete_win_data_49_port, Q(48) => 
                           DataPath_RF_bus_complete_win_data_48_port, Q(47) => 
                           DataPath_RF_bus_complete_win_data_47_port, Q(46) => 
                           DataPath_RF_bus_complete_win_data_46_port, Q(45) => 
                           DataPath_RF_bus_complete_win_data_45_port, Q(44) => 
                           DataPath_RF_bus_complete_win_data_44_port, Q(43) => 
                           DataPath_RF_bus_complete_win_data_43_port, Q(42) => 
                           DataPath_RF_bus_complete_win_data_42_port, Q(41) => 
                           DataPath_RF_bus_complete_win_data_41_port, Q(40) => 
                           DataPath_RF_bus_complete_win_data_40_port, Q(39) => 
                           DataPath_RF_bus_complete_win_data_39_port, Q(38) => 
                           DataPath_RF_bus_complete_win_data_38_port, Q(37) => 
                           DataPath_RF_bus_complete_win_data_37_port, Q(36) => 
                           DataPath_RF_bus_complete_win_data_36_port, Q(35) => 
                           DataPath_RF_bus_complete_win_data_35_port, Q(34) => 
                           DataPath_RF_bus_complete_win_data_34_port, Q(33) => 
                           DataPath_RF_bus_complete_win_data_33_port, Q(32) => 
                           DataPath_RF_bus_complete_win_data_32_port, Q(31) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(30) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(29) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(28) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(27) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(26) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(25) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(24) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(23) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(22) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(21) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(20) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(19) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(18) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(17) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(16) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(15) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(14) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(13) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(12) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(11) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(10) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(9) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(8) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(7) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(6) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(5) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(4) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(3) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(2) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(1) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(0) => 
                           DataPath_RF_bus_complete_win_data_0_port, Y(31) => 
                           DataPath_RF_internal_out2_31_port, Y(30) => 
                           DataPath_RF_internal_out2_30_port, Y(29) => 
                           DataPath_RF_internal_out2_29_port, Y(28) => 
                           DataPath_RF_internal_out2_28_port, Y(27) => 
                           DataPath_RF_internal_out2_27_port, Y(26) => 
                           DataPath_RF_internal_out2_26_port, Y(25) => 
                           DataPath_RF_internal_out2_25_port, Y(24) => 
                           DataPath_RF_internal_out2_24_port, Y(23) => 
                           DataPath_RF_internal_out2_23_port, Y(22) => 
                           DataPath_RF_internal_out2_22_port, Y(21) => 
                           DataPath_RF_internal_out2_21_port, Y(20) => 
                           DataPath_RF_internal_out2_20_port, Y(19) => 
                           DataPath_RF_internal_out2_19_port, Y(18) => 
                           DataPath_RF_internal_out2_18_port, Y(17) => 
                           DataPath_RF_internal_out2_17_port, Y(16) => 
                           DataPath_RF_internal_out2_16_port, Y(15) => 
                           DataPath_RF_internal_out2_15_port, Y(14) => 
                           DataPath_RF_internal_out2_14_port, Y(13) => 
                           DataPath_RF_internal_out2_13_port, Y(12) => 
                           DataPath_RF_internal_out2_12_port, Y(11) => 
                           DataPath_RF_internal_out2_11_port, Y(10) => 
                           DataPath_RF_internal_out2_10_port, Y(9) => 
                           DataPath_RF_internal_out2_9_port, Y(8) => 
                           DataPath_RF_internal_out2_8_port, Y(7) => 
                           DataPath_RF_internal_out2_7_port, Y(6) => 
                           DataPath_RF_internal_out2_6_port, Y(5) => 
                           DataPath_RF_internal_out2_5_port, Y(4) => 
                           DataPath_RF_internal_out2_4_port, Y(3) => 
                           DataPath_RF_internal_out2_3_port, Y(2) => 
                           DataPath_RF_internal_out2_2_port, Y(1) => 
                           DataPath_RF_internal_out2_1_port, Y(0) => 
                           DataPath_RF_internal_out2_0_port);
   DataPath_RF_RDPORT0 : mux_N32_M5_0 port map( S(4) => n10858, S(3) => n10859,
                           S(2) => n10860, S(1) => n10861, S(0) => n10862, 
                           Q(1023) => 
                           DataPath_RF_bus_selected_win_data_767_port, Q(1022) 
                           => DataPath_RF_bus_selected_win_data_766_port, 
                           Q(1021) => 
                           DataPath_RF_bus_selected_win_data_765_port, Q(1020) 
                           => DataPath_RF_bus_selected_win_data_764_port, 
                           Q(1019) => 
                           DataPath_RF_bus_selected_win_data_763_port, Q(1018) 
                           => DataPath_RF_bus_selected_win_data_762_port, 
                           Q(1017) => 
                           DataPath_RF_bus_selected_win_data_761_port, Q(1016) 
                           => DataPath_RF_bus_selected_win_data_760_port, 
                           Q(1015) => 
                           DataPath_RF_bus_selected_win_data_759_port, Q(1014) 
                           => DataPath_RF_bus_selected_win_data_758_port, 
                           Q(1013) => 
                           DataPath_RF_bus_selected_win_data_757_port, Q(1012) 
                           => DataPath_RF_bus_selected_win_data_756_port, 
                           Q(1011) => 
                           DataPath_RF_bus_selected_win_data_755_port, Q(1010) 
                           => DataPath_RF_bus_selected_win_data_754_port, 
                           Q(1009) => 
                           DataPath_RF_bus_selected_win_data_753_port, Q(1008) 
                           => DataPath_RF_bus_selected_win_data_752_port, 
                           Q(1007) => 
                           DataPath_RF_bus_selected_win_data_751_port, Q(1006) 
                           => DataPath_RF_bus_selected_win_data_750_port, 
                           Q(1005) => 
                           DataPath_RF_bus_selected_win_data_749_port, Q(1004) 
                           => DataPath_RF_bus_selected_win_data_748_port, 
                           Q(1003) => 
                           DataPath_RF_bus_selected_win_data_747_port, Q(1002) 
                           => DataPath_RF_bus_selected_win_data_746_port, 
                           Q(1001) => 
                           DataPath_RF_bus_selected_win_data_745_port, Q(1000) 
                           => DataPath_RF_bus_selected_win_data_744_port, 
                           Q(999) => DataPath_RF_bus_selected_win_data_743_port
                           , Q(998) => 
                           DataPath_RF_bus_selected_win_data_742_port, Q(997) 
                           => DataPath_RF_bus_selected_win_data_741_port, 
                           Q(996) => DataPath_RF_bus_selected_win_data_740_port
                           , Q(995) => 
                           DataPath_RF_bus_selected_win_data_739_port, Q(994) 
                           => DataPath_RF_bus_selected_win_data_738_port, 
                           Q(993) => DataPath_RF_bus_selected_win_data_737_port
                           , Q(992) => 
                           DataPath_RF_bus_selected_win_data_736_port, Q(991) 
                           => DataPath_RF_bus_selected_win_data_735_port, 
                           Q(990) => DataPath_RF_bus_selected_win_data_734_port
                           , Q(989) => 
                           DataPath_RF_bus_selected_win_data_733_port, Q(988) 
                           => DataPath_RF_bus_selected_win_data_732_port, 
                           Q(987) => DataPath_RF_bus_selected_win_data_731_port
                           , Q(986) => 
                           DataPath_RF_bus_selected_win_data_730_port, Q(985) 
                           => DataPath_RF_bus_selected_win_data_729_port, 
                           Q(984) => DataPath_RF_bus_selected_win_data_728_port
                           , Q(983) => 
                           DataPath_RF_bus_selected_win_data_727_port, Q(982) 
                           => DataPath_RF_bus_selected_win_data_726_port, 
                           Q(981) => DataPath_RF_bus_selected_win_data_725_port
                           , Q(980) => 
                           DataPath_RF_bus_selected_win_data_724_port, Q(979) 
                           => DataPath_RF_bus_selected_win_data_723_port, 
                           Q(978) => DataPath_RF_bus_selected_win_data_722_port
                           , Q(977) => 
                           DataPath_RF_bus_selected_win_data_721_port, Q(976) 
                           => DataPath_RF_bus_selected_win_data_720_port, 
                           Q(975) => DataPath_RF_bus_selected_win_data_719_port
                           , Q(974) => 
                           DataPath_RF_bus_selected_win_data_718_port, Q(973) 
                           => DataPath_RF_bus_selected_win_data_717_port, 
                           Q(972) => DataPath_RF_bus_selected_win_data_716_port
                           , Q(971) => 
                           DataPath_RF_bus_selected_win_data_715_port, Q(970) 
                           => DataPath_RF_bus_selected_win_data_714_port, 
                           Q(969) => DataPath_RF_bus_selected_win_data_713_port
                           , Q(968) => 
                           DataPath_RF_bus_selected_win_data_712_port, Q(967) 
                           => DataPath_RF_bus_selected_win_data_711_port, 
                           Q(966) => DataPath_RF_bus_selected_win_data_710_port
                           , Q(965) => 
                           DataPath_RF_bus_selected_win_data_709_port, Q(964) 
                           => DataPath_RF_bus_selected_win_data_708_port, 
                           Q(963) => DataPath_RF_bus_selected_win_data_707_port
                           , Q(962) => 
                           DataPath_RF_bus_selected_win_data_706_port, Q(961) 
                           => DataPath_RF_bus_selected_win_data_705_port, 
                           Q(960) => DataPath_RF_bus_selected_win_data_704_port
                           , Q(959) => 
                           DataPath_RF_bus_selected_win_data_703_port, Q(958) 
                           => DataPath_RF_bus_selected_win_data_702_port, 
                           Q(957) => DataPath_RF_bus_selected_win_data_701_port
                           , Q(956) => 
                           DataPath_RF_bus_selected_win_data_700_port, Q(955) 
                           => DataPath_RF_bus_selected_win_data_699_port, 
                           Q(954) => DataPath_RF_bus_selected_win_data_698_port
                           , Q(953) => 
                           DataPath_RF_bus_selected_win_data_697_port, Q(952) 
                           => DataPath_RF_bus_selected_win_data_696_port, 
                           Q(951) => DataPath_RF_bus_selected_win_data_695_port
                           , Q(950) => 
                           DataPath_RF_bus_selected_win_data_694_port, Q(949) 
                           => DataPath_RF_bus_selected_win_data_693_port, 
                           Q(948) => DataPath_RF_bus_selected_win_data_692_port
                           , Q(947) => 
                           DataPath_RF_bus_selected_win_data_691_port, Q(946) 
                           => DataPath_RF_bus_selected_win_data_690_port, 
                           Q(945) => DataPath_RF_bus_selected_win_data_689_port
                           , Q(944) => 
                           DataPath_RF_bus_selected_win_data_688_port, Q(943) 
                           => DataPath_RF_bus_selected_win_data_687_port, 
                           Q(942) => DataPath_RF_bus_selected_win_data_686_port
                           , Q(941) => 
                           DataPath_RF_bus_selected_win_data_685_port, Q(940) 
                           => DataPath_RF_bus_selected_win_data_684_port, 
                           Q(939) => DataPath_RF_bus_selected_win_data_683_port
                           , Q(938) => 
                           DataPath_RF_bus_selected_win_data_682_port, Q(937) 
                           => DataPath_RF_bus_selected_win_data_681_port, 
                           Q(936) => DataPath_RF_bus_selected_win_data_680_port
                           , Q(935) => 
                           DataPath_RF_bus_selected_win_data_679_port, Q(934) 
                           => DataPath_RF_bus_selected_win_data_678_port, 
                           Q(933) => DataPath_RF_bus_selected_win_data_677_port
                           , Q(932) => 
                           DataPath_RF_bus_selected_win_data_676_port, Q(931) 
                           => DataPath_RF_bus_selected_win_data_675_port, 
                           Q(930) => DataPath_RF_bus_selected_win_data_674_port
                           , Q(929) => 
                           DataPath_RF_bus_selected_win_data_673_port, Q(928) 
                           => DataPath_RF_bus_selected_win_data_672_port, 
                           Q(927) => DataPath_RF_bus_selected_win_data_671_port
                           , Q(926) => 
                           DataPath_RF_bus_selected_win_data_670_port, Q(925) 
                           => DataPath_RF_bus_selected_win_data_669_port, 
                           Q(924) => DataPath_RF_bus_selected_win_data_668_port
                           , Q(923) => 
                           DataPath_RF_bus_selected_win_data_667_port, Q(922) 
                           => DataPath_RF_bus_selected_win_data_666_port, 
                           Q(921) => DataPath_RF_bus_selected_win_data_665_port
                           , Q(920) => 
                           DataPath_RF_bus_selected_win_data_664_port, Q(919) 
                           => DataPath_RF_bus_selected_win_data_663_port, 
                           Q(918) => DataPath_RF_bus_selected_win_data_662_port
                           , Q(917) => 
                           DataPath_RF_bus_selected_win_data_661_port, Q(916) 
                           => DataPath_RF_bus_selected_win_data_660_port, 
                           Q(915) => DataPath_RF_bus_selected_win_data_659_port
                           , Q(914) => 
                           DataPath_RF_bus_selected_win_data_658_port, Q(913) 
                           => DataPath_RF_bus_selected_win_data_657_port, 
                           Q(912) => DataPath_RF_bus_selected_win_data_656_port
                           , Q(911) => 
                           DataPath_RF_bus_selected_win_data_655_port, Q(910) 
                           => DataPath_RF_bus_selected_win_data_654_port, 
                           Q(909) => DataPath_RF_bus_selected_win_data_653_port
                           , Q(908) => 
                           DataPath_RF_bus_selected_win_data_652_port, Q(907) 
                           => DataPath_RF_bus_selected_win_data_651_port, 
                           Q(906) => DataPath_RF_bus_selected_win_data_650_port
                           , Q(905) => 
                           DataPath_RF_bus_selected_win_data_649_port, Q(904) 
                           => DataPath_RF_bus_selected_win_data_648_port, 
                           Q(903) => DataPath_RF_bus_selected_win_data_647_port
                           , Q(902) => 
                           DataPath_RF_bus_selected_win_data_646_port, Q(901) 
                           => DataPath_RF_bus_selected_win_data_645_port, 
                           Q(900) => DataPath_RF_bus_selected_win_data_644_port
                           , Q(899) => 
                           DataPath_RF_bus_selected_win_data_643_port, Q(898) 
                           => DataPath_RF_bus_selected_win_data_642_port, 
                           Q(897) => DataPath_RF_bus_selected_win_data_641_port
                           , Q(896) => 
                           DataPath_RF_bus_selected_win_data_640_port, Q(895) 
                           => DataPath_RF_bus_selected_win_data_639_port, 
                           Q(894) => DataPath_RF_bus_selected_win_data_638_port
                           , Q(893) => 
                           DataPath_RF_bus_selected_win_data_637_port, Q(892) 
                           => DataPath_RF_bus_selected_win_data_636_port, 
                           Q(891) => DataPath_RF_bus_selected_win_data_635_port
                           , Q(890) => 
                           DataPath_RF_bus_selected_win_data_634_port, Q(889) 
                           => DataPath_RF_bus_selected_win_data_633_port, 
                           Q(888) => DataPath_RF_bus_selected_win_data_632_port
                           , Q(887) => 
                           DataPath_RF_bus_selected_win_data_631_port, Q(886) 
                           => DataPath_RF_bus_selected_win_data_630_port, 
                           Q(885) => DataPath_RF_bus_selected_win_data_629_port
                           , Q(884) => 
                           DataPath_RF_bus_selected_win_data_628_port, Q(883) 
                           => DataPath_RF_bus_selected_win_data_627_port, 
                           Q(882) => DataPath_RF_bus_selected_win_data_626_port
                           , Q(881) => 
                           DataPath_RF_bus_selected_win_data_625_port, Q(880) 
                           => DataPath_RF_bus_selected_win_data_624_port, 
                           Q(879) => DataPath_RF_bus_selected_win_data_623_port
                           , Q(878) => 
                           DataPath_RF_bus_selected_win_data_622_port, Q(877) 
                           => DataPath_RF_bus_selected_win_data_621_port, 
                           Q(876) => DataPath_RF_bus_selected_win_data_620_port
                           , Q(875) => 
                           DataPath_RF_bus_selected_win_data_619_port, Q(874) 
                           => DataPath_RF_bus_selected_win_data_618_port, 
                           Q(873) => DataPath_RF_bus_selected_win_data_617_port
                           , Q(872) => 
                           DataPath_RF_bus_selected_win_data_616_port, Q(871) 
                           => DataPath_RF_bus_selected_win_data_615_port, 
                           Q(870) => DataPath_RF_bus_selected_win_data_614_port
                           , Q(869) => 
                           DataPath_RF_bus_selected_win_data_613_port, Q(868) 
                           => DataPath_RF_bus_selected_win_data_612_port, 
                           Q(867) => DataPath_RF_bus_selected_win_data_611_port
                           , Q(866) => 
                           DataPath_RF_bus_selected_win_data_610_port, Q(865) 
                           => DataPath_RF_bus_selected_win_data_609_port, 
                           Q(864) => DataPath_RF_bus_selected_win_data_608_port
                           , Q(863) => 
                           DataPath_RF_bus_selected_win_data_607_port, Q(862) 
                           => DataPath_RF_bus_selected_win_data_606_port, 
                           Q(861) => DataPath_RF_bus_selected_win_data_605_port
                           , Q(860) => 
                           DataPath_RF_bus_selected_win_data_604_port, Q(859) 
                           => DataPath_RF_bus_selected_win_data_603_port, 
                           Q(858) => DataPath_RF_bus_selected_win_data_602_port
                           , Q(857) => 
                           DataPath_RF_bus_selected_win_data_601_port, Q(856) 
                           => DataPath_RF_bus_selected_win_data_600_port, 
                           Q(855) => DataPath_RF_bus_selected_win_data_599_port
                           , Q(854) => 
                           DataPath_RF_bus_selected_win_data_598_port, Q(853) 
                           => DataPath_RF_bus_selected_win_data_597_port, 
                           Q(852) => DataPath_RF_bus_selected_win_data_596_port
                           , Q(851) => 
                           DataPath_RF_bus_selected_win_data_595_port, Q(850) 
                           => DataPath_RF_bus_selected_win_data_594_port, 
                           Q(849) => DataPath_RF_bus_selected_win_data_593_port
                           , Q(848) => 
                           DataPath_RF_bus_selected_win_data_592_port, Q(847) 
                           => DataPath_RF_bus_selected_win_data_591_port, 
                           Q(846) => DataPath_RF_bus_selected_win_data_590_port
                           , Q(845) => 
                           DataPath_RF_bus_selected_win_data_589_port, Q(844) 
                           => DataPath_RF_bus_selected_win_data_588_port, 
                           Q(843) => DataPath_RF_bus_selected_win_data_587_port
                           , Q(842) => 
                           DataPath_RF_bus_selected_win_data_586_port, Q(841) 
                           => DataPath_RF_bus_selected_win_data_585_port, 
                           Q(840) => DataPath_RF_bus_selected_win_data_584_port
                           , Q(839) => 
                           DataPath_RF_bus_selected_win_data_583_port, Q(838) 
                           => DataPath_RF_bus_selected_win_data_582_port, 
                           Q(837) => DataPath_RF_bus_selected_win_data_581_port
                           , Q(836) => 
                           DataPath_RF_bus_selected_win_data_580_port, Q(835) 
                           => DataPath_RF_bus_selected_win_data_579_port, 
                           Q(834) => DataPath_RF_bus_selected_win_data_578_port
                           , Q(833) => 
                           DataPath_RF_bus_selected_win_data_577_port, Q(832) 
                           => DataPath_RF_bus_selected_win_data_576_port, 
                           Q(831) => DataPath_RF_bus_selected_win_data_575_port
                           , Q(830) => 
                           DataPath_RF_bus_selected_win_data_574_port, Q(829) 
                           => DataPath_RF_bus_selected_win_data_573_port, 
                           Q(828) => DataPath_RF_bus_selected_win_data_572_port
                           , Q(827) => 
                           DataPath_RF_bus_selected_win_data_571_port, Q(826) 
                           => DataPath_RF_bus_selected_win_data_570_port, 
                           Q(825) => DataPath_RF_bus_selected_win_data_569_port
                           , Q(824) => 
                           DataPath_RF_bus_selected_win_data_568_port, Q(823) 
                           => DataPath_RF_bus_selected_win_data_567_port, 
                           Q(822) => DataPath_RF_bus_selected_win_data_566_port
                           , Q(821) => 
                           DataPath_RF_bus_selected_win_data_565_port, Q(820) 
                           => DataPath_RF_bus_selected_win_data_564_port, 
                           Q(819) => DataPath_RF_bus_selected_win_data_563_port
                           , Q(818) => 
                           DataPath_RF_bus_selected_win_data_562_port, Q(817) 
                           => DataPath_RF_bus_selected_win_data_561_port, 
                           Q(816) => DataPath_RF_bus_selected_win_data_560_port
                           , Q(815) => 
                           DataPath_RF_bus_selected_win_data_559_port, Q(814) 
                           => DataPath_RF_bus_selected_win_data_558_port, 
                           Q(813) => DataPath_RF_bus_selected_win_data_557_port
                           , Q(812) => 
                           DataPath_RF_bus_selected_win_data_556_port, Q(811) 
                           => DataPath_RF_bus_selected_win_data_555_port, 
                           Q(810) => DataPath_RF_bus_selected_win_data_554_port
                           , Q(809) => 
                           DataPath_RF_bus_selected_win_data_553_port, Q(808) 
                           => DataPath_RF_bus_selected_win_data_552_port, 
                           Q(807) => DataPath_RF_bus_selected_win_data_551_port
                           , Q(806) => 
                           DataPath_RF_bus_selected_win_data_550_port, Q(805) 
                           => DataPath_RF_bus_selected_win_data_549_port, 
                           Q(804) => DataPath_RF_bus_selected_win_data_548_port
                           , Q(803) => 
                           DataPath_RF_bus_selected_win_data_547_port, Q(802) 
                           => DataPath_RF_bus_selected_win_data_546_port, 
                           Q(801) => DataPath_RF_bus_selected_win_data_545_port
                           , Q(800) => 
                           DataPath_RF_bus_selected_win_data_544_port, Q(799) 
                           => DataPath_RF_bus_selected_win_data_543_port, 
                           Q(798) => DataPath_RF_bus_selected_win_data_542_port
                           , Q(797) => 
                           DataPath_RF_bus_selected_win_data_541_port, Q(796) 
                           => DataPath_RF_bus_selected_win_data_540_port, 
                           Q(795) => DataPath_RF_bus_selected_win_data_539_port
                           , Q(794) => 
                           DataPath_RF_bus_selected_win_data_538_port, Q(793) 
                           => DataPath_RF_bus_selected_win_data_537_port, 
                           Q(792) => DataPath_RF_bus_selected_win_data_536_port
                           , Q(791) => 
                           DataPath_RF_bus_selected_win_data_535_port, Q(790) 
                           => DataPath_RF_bus_selected_win_data_534_port, 
                           Q(789) => DataPath_RF_bus_selected_win_data_533_port
                           , Q(788) => 
                           DataPath_RF_bus_selected_win_data_532_port, Q(787) 
                           => DataPath_RF_bus_selected_win_data_531_port, 
                           Q(786) => DataPath_RF_bus_selected_win_data_530_port
                           , Q(785) => 
                           DataPath_RF_bus_selected_win_data_529_port, Q(784) 
                           => DataPath_RF_bus_selected_win_data_528_port, 
                           Q(783) => DataPath_RF_bus_selected_win_data_527_port
                           , Q(782) => 
                           DataPath_RF_bus_selected_win_data_526_port, Q(781) 
                           => DataPath_RF_bus_selected_win_data_525_port, 
                           Q(780) => DataPath_RF_bus_selected_win_data_524_port
                           , Q(779) => 
                           DataPath_RF_bus_selected_win_data_523_port, Q(778) 
                           => DataPath_RF_bus_selected_win_data_522_port, 
                           Q(777) => DataPath_RF_bus_selected_win_data_521_port
                           , Q(776) => 
                           DataPath_RF_bus_selected_win_data_520_port, Q(775) 
                           => DataPath_RF_bus_selected_win_data_519_port, 
                           Q(774) => DataPath_RF_bus_selected_win_data_518_port
                           , Q(773) => 
                           DataPath_RF_bus_selected_win_data_517_port, Q(772) 
                           => DataPath_RF_bus_selected_win_data_516_port, 
                           Q(771) => DataPath_RF_bus_selected_win_data_515_port
                           , Q(770) => 
                           DataPath_RF_bus_selected_win_data_514_port, Q(769) 
                           => DataPath_RF_bus_selected_win_data_513_port, 
                           Q(768) => DataPath_RF_bus_selected_win_data_512_port
                           , Q(767) => 
                           DataPath_RF_bus_selected_win_data_511_port, Q(766) 
                           => DataPath_RF_bus_selected_win_data_510_port, 
                           Q(765) => DataPath_RF_bus_selected_win_data_509_port
                           , Q(764) => 
                           DataPath_RF_bus_selected_win_data_508_port, Q(763) 
                           => DataPath_RF_bus_selected_win_data_507_port, 
                           Q(762) => DataPath_RF_bus_selected_win_data_506_port
                           , Q(761) => 
                           DataPath_RF_bus_selected_win_data_505_port, Q(760) 
                           => DataPath_RF_bus_selected_win_data_504_port, 
                           Q(759) => DataPath_RF_bus_selected_win_data_503_port
                           , Q(758) => 
                           DataPath_RF_bus_selected_win_data_502_port, Q(757) 
                           => DataPath_RF_bus_selected_win_data_501_port, 
                           Q(756) => DataPath_RF_bus_selected_win_data_500_port
                           , Q(755) => 
                           DataPath_RF_bus_selected_win_data_499_port, Q(754) 
                           => DataPath_RF_bus_selected_win_data_498_port, 
                           Q(753) => DataPath_RF_bus_selected_win_data_497_port
                           , Q(752) => 
                           DataPath_RF_bus_selected_win_data_496_port, Q(751) 
                           => DataPath_RF_bus_selected_win_data_495_port, 
                           Q(750) => DataPath_RF_bus_selected_win_data_494_port
                           , Q(749) => 
                           DataPath_RF_bus_selected_win_data_493_port, Q(748) 
                           => DataPath_RF_bus_selected_win_data_492_port, 
                           Q(747) => DataPath_RF_bus_selected_win_data_491_port
                           , Q(746) => 
                           DataPath_RF_bus_selected_win_data_490_port, Q(745) 
                           => DataPath_RF_bus_selected_win_data_489_port, 
                           Q(744) => DataPath_RF_bus_selected_win_data_488_port
                           , Q(743) => 
                           DataPath_RF_bus_selected_win_data_487_port, Q(742) 
                           => DataPath_RF_bus_selected_win_data_486_port, 
                           Q(741) => DataPath_RF_bus_selected_win_data_485_port
                           , Q(740) => 
                           DataPath_RF_bus_selected_win_data_484_port, Q(739) 
                           => DataPath_RF_bus_selected_win_data_483_port, 
                           Q(738) => DataPath_RF_bus_selected_win_data_482_port
                           , Q(737) => 
                           DataPath_RF_bus_selected_win_data_481_port, Q(736) 
                           => DataPath_RF_bus_selected_win_data_480_port, 
                           Q(735) => DataPath_RF_bus_selected_win_data_479_port
                           , Q(734) => 
                           DataPath_RF_bus_selected_win_data_478_port, Q(733) 
                           => DataPath_RF_bus_selected_win_data_477_port, 
                           Q(732) => DataPath_RF_bus_selected_win_data_476_port
                           , Q(731) => 
                           DataPath_RF_bus_selected_win_data_475_port, Q(730) 
                           => DataPath_RF_bus_selected_win_data_474_port, 
                           Q(729) => DataPath_RF_bus_selected_win_data_473_port
                           , Q(728) => 
                           DataPath_RF_bus_selected_win_data_472_port, Q(727) 
                           => DataPath_RF_bus_selected_win_data_471_port, 
                           Q(726) => DataPath_RF_bus_selected_win_data_470_port
                           , Q(725) => 
                           DataPath_RF_bus_selected_win_data_469_port, Q(724) 
                           => DataPath_RF_bus_selected_win_data_468_port, 
                           Q(723) => DataPath_RF_bus_selected_win_data_467_port
                           , Q(722) => 
                           DataPath_RF_bus_selected_win_data_466_port, Q(721) 
                           => DataPath_RF_bus_selected_win_data_465_port, 
                           Q(720) => DataPath_RF_bus_selected_win_data_464_port
                           , Q(719) => 
                           DataPath_RF_bus_selected_win_data_463_port, Q(718) 
                           => DataPath_RF_bus_selected_win_data_462_port, 
                           Q(717) => DataPath_RF_bus_selected_win_data_461_port
                           , Q(716) => 
                           DataPath_RF_bus_selected_win_data_460_port, Q(715) 
                           => DataPath_RF_bus_selected_win_data_459_port, 
                           Q(714) => DataPath_RF_bus_selected_win_data_458_port
                           , Q(713) => 
                           DataPath_RF_bus_selected_win_data_457_port, Q(712) 
                           => DataPath_RF_bus_selected_win_data_456_port, 
                           Q(711) => DataPath_RF_bus_selected_win_data_455_port
                           , Q(710) => 
                           DataPath_RF_bus_selected_win_data_454_port, Q(709) 
                           => DataPath_RF_bus_selected_win_data_453_port, 
                           Q(708) => DataPath_RF_bus_selected_win_data_452_port
                           , Q(707) => 
                           DataPath_RF_bus_selected_win_data_451_port, Q(706) 
                           => DataPath_RF_bus_selected_win_data_450_port, 
                           Q(705) => DataPath_RF_bus_selected_win_data_449_port
                           , Q(704) => 
                           DataPath_RF_bus_selected_win_data_448_port, Q(703) 
                           => DataPath_RF_bus_selected_win_data_447_port, 
                           Q(702) => DataPath_RF_bus_selected_win_data_446_port
                           , Q(701) => 
                           DataPath_RF_bus_selected_win_data_445_port, Q(700) 
                           => DataPath_RF_bus_selected_win_data_444_port, 
                           Q(699) => DataPath_RF_bus_selected_win_data_443_port
                           , Q(698) => 
                           DataPath_RF_bus_selected_win_data_442_port, Q(697) 
                           => DataPath_RF_bus_selected_win_data_441_port, 
                           Q(696) => DataPath_RF_bus_selected_win_data_440_port
                           , Q(695) => 
                           DataPath_RF_bus_selected_win_data_439_port, Q(694) 
                           => DataPath_RF_bus_selected_win_data_438_port, 
                           Q(693) => DataPath_RF_bus_selected_win_data_437_port
                           , Q(692) => 
                           DataPath_RF_bus_selected_win_data_436_port, Q(691) 
                           => DataPath_RF_bus_selected_win_data_435_port, 
                           Q(690) => DataPath_RF_bus_selected_win_data_434_port
                           , Q(689) => 
                           DataPath_RF_bus_selected_win_data_433_port, Q(688) 
                           => DataPath_RF_bus_selected_win_data_432_port, 
                           Q(687) => DataPath_RF_bus_selected_win_data_431_port
                           , Q(686) => 
                           DataPath_RF_bus_selected_win_data_430_port, Q(685) 
                           => DataPath_RF_bus_selected_win_data_429_port, 
                           Q(684) => DataPath_RF_bus_selected_win_data_428_port
                           , Q(683) => 
                           DataPath_RF_bus_selected_win_data_427_port, Q(682) 
                           => DataPath_RF_bus_selected_win_data_426_port, 
                           Q(681) => DataPath_RF_bus_selected_win_data_425_port
                           , Q(680) => 
                           DataPath_RF_bus_selected_win_data_424_port, Q(679) 
                           => DataPath_RF_bus_selected_win_data_423_port, 
                           Q(678) => DataPath_RF_bus_selected_win_data_422_port
                           , Q(677) => 
                           DataPath_RF_bus_selected_win_data_421_port, Q(676) 
                           => DataPath_RF_bus_selected_win_data_420_port, 
                           Q(675) => DataPath_RF_bus_selected_win_data_419_port
                           , Q(674) => 
                           DataPath_RF_bus_selected_win_data_418_port, Q(673) 
                           => DataPath_RF_bus_selected_win_data_417_port, 
                           Q(672) => DataPath_RF_bus_selected_win_data_416_port
                           , Q(671) => 
                           DataPath_RF_bus_selected_win_data_415_port, Q(670) 
                           => DataPath_RF_bus_selected_win_data_414_port, 
                           Q(669) => DataPath_RF_bus_selected_win_data_413_port
                           , Q(668) => 
                           DataPath_RF_bus_selected_win_data_412_port, Q(667) 
                           => DataPath_RF_bus_selected_win_data_411_port, 
                           Q(666) => DataPath_RF_bus_selected_win_data_410_port
                           , Q(665) => 
                           DataPath_RF_bus_selected_win_data_409_port, Q(664) 
                           => DataPath_RF_bus_selected_win_data_408_port, 
                           Q(663) => DataPath_RF_bus_selected_win_data_407_port
                           , Q(662) => 
                           DataPath_RF_bus_selected_win_data_406_port, Q(661) 
                           => DataPath_RF_bus_selected_win_data_405_port, 
                           Q(660) => DataPath_RF_bus_selected_win_data_404_port
                           , Q(659) => 
                           DataPath_RF_bus_selected_win_data_403_port, Q(658) 
                           => DataPath_RF_bus_selected_win_data_402_port, 
                           Q(657) => DataPath_RF_bus_selected_win_data_401_port
                           , Q(656) => 
                           DataPath_RF_bus_selected_win_data_400_port, Q(655) 
                           => DataPath_RF_bus_selected_win_data_399_port, 
                           Q(654) => DataPath_RF_bus_selected_win_data_398_port
                           , Q(653) => 
                           DataPath_RF_bus_selected_win_data_397_port, Q(652) 
                           => DataPath_RF_bus_selected_win_data_396_port, 
                           Q(651) => DataPath_RF_bus_selected_win_data_395_port
                           , Q(650) => 
                           DataPath_RF_bus_selected_win_data_394_port, Q(649) 
                           => DataPath_RF_bus_selected_win_data_393_port, 
                           Q(648) => DataPath_RF_bus_selected_win_data_392_port
                           , Q(647) => 
                           DataPath_RF_bus_selected_win_data_391_port, Q(646) 
                           => DataPath_RF_bus_selected_win_data_390_port, 
                           Q(645) => DataPath_RF_bus_selected_win_data_389_port
                           , Q(644) => 
                           DataPath_RF_bus_selected_win_data_388_port, Q(643) 
                           => DataPath_RF_bus_selected_win_data_387_port, 
                           Q(642) => DataPath_RF_bus_selected_win_data_386_port
                           , Q(641) => 
                           DataPath_RF_bus_selected_win_data_385_port, Q(640) 
                           => DataPath_RF_bus_selected_win_data_384_port, 
                           Q(639) => DataPath_RF_bus_selected_win_data_383_port
                           , Q(638) => 
                           DataPath_RF_bus_selected_win_data_382_port, Q(637) 
                           => DataPath_RF_bus_selected_win_data_381_port, 
                           Q(636) => DataPath_RF_bus_selected_win_data_380_port
                           , Q(635) => 
                           DataPath_RF_bus_selected_win_data_379_port, Q(634) 
                           => DataPath_RF_bus_selected_win_data_378_port, 
                           Q(633) => DataPath_RF_bus_selected_win_data_377_port
                           , Q(632) => 
                           DataPath_RF_bus_selected_win_data_376_port, Q(631) 
                           => DataPath_RF_bus_selected_win_data_375_port, 
                           Q(630) => DataPath_RF_bus_selected_win_data_374_port
                           , Q(629) => 
                           DataPath_RF_bus_selected_win_data_373_port, Q(628) 
                           => DataPath_RF_bus_selected_win_data_372_port, 
                           Q(627) => DataPath_RF_bus_selected_win_data_371_port
                           , Q(626) => 
                           DataPath_RF_bus_selected_win_data_370_port, Q(625) 
                           => DataPath_RF_bus_selected_win_data_369_port, 
                           Q(624) => DataPath_RF_bus_selected_win_data_368_port
                           , Q(623) => 
                           DataPath_RF_bus_selected_win_data_367_port, Q(622) 
                           => DataPath_RF_bus_selected_win_data_366_port, 
                           Q(621) => DataPath_RF_bus_selected_win_data_365_port
                           , Q(620) => 
                           DataPath_RF_bus_selected_win_data_364_port, Q(619) 
                           => DataPath_RF_bus_selected_win_data_363_port, 
                           Q(618) => DataPath_RF_bus_selected_win_data_362_port
                           , Q(617) => 
                           DataPath_RF_bus_selected_win_data_361_port, Q(616) 
                           => DataPath_RF_bus_selected_win_data_360_port, 
                           Q(615) => DataPath_RF_bus_selected_win_data_359_port
                           , Q(614) => 
                           DataPath_RF_bus_selected_win_data_358_port, Q(613) 
                           => DataPath_RF_bus_selected_win_data_357_port, 
                           Q(612) => DataPath_RF_bus_selected_win_data_356_port
                           , Q(611) => 
                           DataPath_RF_bus_selected_win_data_355_port, Q(610) 
                           => DataPath_RF_bus_selected_win_data_354_port, 
                           Q(609) => DataPath_RF_bus_selected_win_data_353_port
                           , Q(608) => 
                           DataPath_RF_bus_selected_win_data_352_port, Q(607) 
                           => DataPath_RF_bus_selected_win_data_351_port, 
                           Q(606) => DataPath_RF_bus_selected_win_data_350_port
                           , Q(605) => 
                           DataPath_RF_bus_selected_win_data_349_port, Q(604) 
                           => DataPath_RF_bus_selected_win_data_348_port, 
                           Q(603) => DataPath_RF_bus_selected_win_data_347_port
                           , Q(602) => 
                           DataPath_RF_bus_selected_win_data_346_port, Q(601) 
                           => DataPath_RF_bus_selected_win_data_345_port, 
                           Q(600) => DataPath_RF_bus_selected_win_data_344_port
                           , Q(599) => 
                           DataPath_RF_bus_selected_win_data_343_port, Q(598) 
                           => DataPath_RF_bus_selected_win_data_342_port, 
                           Q(597) => DataPath_RF_bus_selected_win_data_341_port
                           , Q(596) => 
                           DataPath_RF_bus_selected_win_data_340_port, Q(595) 
                           => DataPath_RF_bus_selected_win_data_339_port, 
                           Q(594) => DataPath_RF_bus_selected_win_data_338_port
                           , Q(593) => 
                           DataPath_RF_bus_selected_win_data_337_port, Q(592) 
                           => DataPath_RF_bus_selected_win_data_336_port, 
                           Q(591) => DataPath_RF_bus_selected_win_data_335_port
                           , Q(590) => 
                           DataPath_RF_bus_selected_win_data_334_port, Q(589) 
                           => DataPath_RF_bus_selected_win_data_333_port, 
                           Q(588) => DataPath_RF_bus_selected_win_data_332_port
                           , Q(587) => 
                           DataPath_RF_bus_selected_win_data_331_port, Q(586) 
                           => DataPath_RF_bus_selected_win_data_330_port, 
                           Q(585) => DataPath_RF_bus_selected_win_data_329_port
                           , Q(584) => 
                           DataPath_RF_bus_selected_win_data_328_port, Q(583) 
                           => DataPath_RF_bus_selected_win_data_327_port, 
                           Q(582) => DataPath_RF_bus_selected_win_data_326_port
                           , Q(581) => 
                           DataPath_RF_bus_selected_win_data_325_port, Q(580) 
                           => DataPath_RF_bus_selected_win_data_324_port, 
                           Q(579) => DataPath_RF_bus_selected_win_data_323_port
                           , Q(578) => 
                           DataPath_RF_bus_selected_win_data_322_port, Q(577) 
                           => DataPath_RF_bus_selected_win_data_321_port, 
                           Q(576) => DataPath_RF_bus_selected_win_data_320_port
                           , Q(575) => 
                           DataPath_RF_bus_selected_win_data_319_port, Q(574) 
                           => DataPath_RF_bus_selected_win_data_318_port, 
                           Q(573) => DataPath_RF_bus_selected_win_data_317_port
                           , Q(572) => 
                           DataPath_RF_bus_selected_win_data_316_port, Q(571) 
                           => DataPath_RF_bus_selected_win_data_315_port, 
                           Q(570) => DataPath_RF_bus_selected_win_data_314_port
                           , Q(569) => 
                           DataPath_RF_bus_selected_win_data_313_port, Q(568) 
                           => DataPath_RF_bus_selected_win_data_312_port, 
                           Q(567) => DataPath_RF_bus_selected_win_data_311_port
                           , Q(566) => 
                           DataPath_RF_bus_selected_win_data_310_port, Q(565) 
                           => DataPath_RF_bus_selected_win_data_309_port, 
                           Q(564) => DataPath_RF_bus_selected_win_data_308_port
                           , Q(563) => 
                           DataPath_RF_bus_selected_win_data_307_port, Q(562) 
                           => DataPath_RF_bus_selected_win_data_306_port, 
                           Q(561) => DataPath_RF_bus_selected_win_data_305_port
                           , Q(560) => 
                           DataPath_RF_bus_selected_win_data_304_port, Q(559) 
                           => DataPath_RF_bus_selected_win_data_303_port, 
                           Q(558) => DataPath_RF_bus_selected_win_data_302_port
                           , Q(557) => 
                           DataPath_RF_bus_selected_win_data_301_port, Q(556) 
                           => DataPath_RF_bus_selected_win_data_300_port, 
                           Q(555) => DataPath_RF_bus_selected_win_data_299_port
                           , Q(554) => 
                           DataPath_RF_bus_selected_win_data_298_port, Q(553) 
                           => DataPath_RF_bus_selected_win_data_297_port, 
                           Q(552) => DataPath_RF_bus_selected_win_data_296_port
                           , Q(551) => 
                           DataPath_RF_bus_selected_win_data_295_port, Q(550) 
                           => DataPath_RF_bus_selected_win_data_294_port, 
                           Q(549) => DataPath_RF_bus_selected_win_data_293_port
                           , Q(548) => 
                           DataPath_RF_bus_selected_win_data_292_port, Q(547) 
                           => DataPath_RF_bus_selected_win_data_291_port, 
                           Q(546) => DataPath_RF_bus_selected_win_data_290_port
                           , Q(545) => 
                           DataPath_RF_bus_selected_win_data_289_port, Q(544) 
                           => DataPath_RF_bus_selected_win_data_288_port, 
                           Q(543) => DataPath_RF_bus_selected_win_data_287_port
                           , Q(542) => 
                           DataPath_RF_bus_selected_win_data_286_port, Q(541) 
                           => DataPath_RF_bus_selected_win_data_285_port, 
                           Q(540) => DataPath_RF_bus_selected_win_data_284_port
                           , Q(539) => 
                           DataPath_RF_bus_selected_win_data_283_port, Q(538) 
                           => DataPath_RF_bus_selected_win_data_282_port, 
                           Q(537) => DataPath_RF_bus_selected_win_data_281_port
                           , Q(536) => 
                           DataPath_RF_bus_selected_win_data_280_port, Q(535) 
                           => DataPath_RF_bus_selected_win_data_279_port, 
                           Q(534) => DataPath_RF_bus_selected_win_data_278_port
                           , Q(533) => 
                           DataPath_RF_bus_selected_win_data_277_port, Q(532) 
                           => DataPath_RF_bus_selected_win_data_276_port, 
                           Q(531) => DataPath_RF_bus_selected_win_data_275_port
                           , Q(530) => 
                           DataPath_RF_bus_selected_win_data_274_port, Q(529) 
                           => DataPath_RF_bus_selected_win_data_273_port, 
                           Q(528) => DataPath_RF_bus_selected_win_data_272_port
                           , Q(527) => 
                           DataPath_RF_bus_selected_win_data_271_port, Q(526) 
                           => DataPath_RF_bus_selected_win_data_270_port, 
                           Q(525) => DataPath_RF_bus_selected_win_data_269_port
                           , Q(524) => 
                           DataPath_RF_bus_selected_win_data_268_port, Q(523) 
                           => DataPath_RF_bus_selected_win_data_267_port, 
                           Q(522) => DataPath_RF_bus_selected_win_data_266_port
                           , Q(521) => 
                           DataPath_RF_bus_selected_win_data_265_port, Q(520) 
                           => DataPath_RF_bus_selected_win_data_264_port, 
                           Q(519) => DataPath_RF_bus_selected_win_data_263_port
                           , Q(518) => 
                           DataPath_RF_bus_selected_win_data_262_port, Q(517) 
                           => DataPath_RF_bus_selected_win_data_261_port, 
                           Q(516) => DataPath_RF_bus_selected_win_data_260_port
                           , Q(515) => 
                           DataPath_RF_bus_selected_win_data_259_port, Q(514) 
                           => DataPath_RF_bus_selected_win_data_258_port, 
                           Q(513) => DataPath_RF_bus_selected_win_data_257_port
                           , Q(512) => 
                           DataPath_RF_bus_selected_win_data_256_port, Q(511) 
                           => DataPath_RF_bus_selected_win_data_255_port, 
                           Q(510) => DataPath_RF_bus_selected_win_data_254_port
                           , Q(509) => 
                           DataPath_RF_bus_selected_win_data_253_port, Q(508) 
                           => DataPath_RF_bus_selected_win_data_252_port, 
                           Q(507) => DataPath_RF_bus_selected_win_data_251_port
                           , Q(506) => 
                           DataPath_RF_bus_selected_win_data_250_port, Q(505) 
                           => DataPath_RF_bus_selected_win_data_249_port, 
                           Q(504) => DataPath_RF_bus_selected_win_data_248_port
                           , Q(503) => 
                           DataPath_RF_bus_selected_win_data_247_port, Q(502) 
                           => DataPath_RF_bus_selected_win_data_246_port, 
                           Q(501) => DataPath_RF_bus_selected_win_data_245_port
                           , Q(500) => 
                           DataPath_RF_bus_selected_win_data_244_port, Q(499) 
                           => DataPath_RF_bus_selected_win_data_243_port, 
                           Q(498) => DataPath_RF_bus_selected_win_data_242_port
                           , Q(497) => 
                           DataPath_RF_bus_selected_win_data_241_port, Q(496) 
                           => DataPath_RF_bus_selected_win_data_240_port, 
                           Q(495) => DataPath_RF_bus_selected_win_data_239_port
                           , Q(494) => 
                           DataPath_RF_bus_selected_win_data_238_port, Q(493) 
                           => DataPath_RF_bus_selected_win_data_237_port, 
                           Q(492) => DataPath_RF_bus_selected_win_data_236_port
                           , Q(491) => 
                           DataPath_RF_bus_selected_win_data_235_port, Q(490) 
                           => DataPath_RF_bus_selected_win_data_234_port, 
                           Q(489) => DataPath_RF_bus_selected_win_data_233_port
                           , Q(488) => 
                           DataPath_RF_bus_selected_win_data_232_port, Q(487) 
                           => DataPath_RF_bus_selected_win_data_231_port, 
                           Q(486) => DataPath_RF_bus_selected_win_data_230_port
                           , Q(485) => 
                           DataPath_RF_bus_selected_win_data_229_port, Q(484) 
                           => DataPath_RF_bus_selected_win_data_228_port, 
                           Q(483) => DataPath_RF_bus_selected_win_data_227_port
                           , Q(482) => 
                           DataPath_RF_bus_selected_win_data_226_port, Q(481) 
                           => DataPath_RF_bus_selected_win_data_225_port, 
                           Q(480) => DataPath_RF_bus_selected_win_data_224_port
                           , Q(479) => 
                           DataPath_RF_bus_selected_win_data_223_port, Q(478) 
                           => DataPath_RF_bus_selected_win_data_222_port, 
                           Q(477) => DataPath_RF_bus_selected_win_data_221_port
                           , Q(476) => 
                           DataPath_RF_bus_selected_win_data_220_port, Q(475) 
                           => DataPath_RF_bus_selected_win_data_219_port, 
                           Q(474) => DataPath_RF_bus_selected_win_data_218_port
                           , Q(473) => 
                           DataPath_RF_bus_selected_win_data_217_port, Q(472) 
                           => DataPath_RF_bus_selected_win_data_216_port, 
                           Q(471) => DataPath_RF_bus_selected_win_data_215_port
                           , Q(470) => 
                           DataPath_RF_bus_selected_win_data_214_port, Q(469) 
                           => DataPath_RF_bus_selected_win_data_213_port, 
                           Q(468) => DataPath_RF_bus_selected_win_data_212_port
                           , Q(467) => 
                           DataPath_RF_bus_selected_win_data_211_port, Q(466) 
                           => DataPath_RF_bus_selected_win_data_210_port, 
                           Q(465) => DataPath_RF_bus_selected_win_data_209_port
                           , Q(464) => 
                           DataPath_RF_bus_selected_win_data_208_port, Q(463) 
                           => DataPath_RF_bus_selected_win_data_207_port, 
                           Q(462) => DataPath_RF_bus_selected_win_data_206_port
                           , Q(461) => 
                           DataPath_RF_bus_selected_win_data_205_port, Q(460) 
                           => DataPath_RF_bus_selected_win_data_204_port, 
                           Q(459) => DataPath_RF_bus_selected_win_data_203_port
                           , Q(458) => 
                           DataPath_RF_bus_selected_win_data_202_port, Q(457) 
                           => DataPath_RF_bus_selected_win_data_201_port, 
                           Q(456) => DataPath_RF_bus_selected_win_data_200_port
                           , Q(455) => 
                           DataPath_RF_bus_selected_win_data_199_port, Q(454) 
                           => DataPath_RF_bus_selected_win_data_198_port, 
                           Q(453) => DataPath_RF_bus_selected_win_data_197_port
                           , Q(452) => 
                           DataPath_RF_bus_selected_win_data_196_port, Q(451) 
                           => DataPath_RF_bus_selected_win_data_195_port, 
                           Q(450) => DataPath_RF_bus_selected_win_data_194_port
                           , Q(449) => 
                           DataPath_RF_bus_selected_win_data_193_port, Q(448) 
                           => DataPath_RF_bus_selected_win_data_192_port, 
                           Q(447) => DataPath_RF_bus_selected_win_data_191_port
                           , Q(446) => 
                           DataPath_RF_bus_selected_win_data_190_port, Q(445) 
                           => DataPath_RF_bus_selected_win_data_189_port, 
                           Q(444) => DataPath_RF_bus_selected_win_data_188_port
                           , Q(443) => 
                           DataPath_RF_bus_selected_win_data_187_port, Q(442) 
                           => DataPath_RF_bus_selected_win_data_186_port, 
                           Q(441) => DataPath_RF_bus_selected_win_data_185_port
                           , Q(440) => 
                           DataPath_RF_bus_selected_win_data_184_port, Q(439) 
                           => DataPath_RF_bus_selected_win_data_183_port, 
                           Q(438) => DataPath_RF_bus_selected_win_data_182_port
                           , Q(437) => 
                           DataPath_RF_bus_selected_win_data_181_port, Q(436) 
                           => DataPath_RF_bus_selected_win_data_180_port, 
                           Q(435) => DataPath_RF_bus_selected_win_data_179_port
                           , Q(434) => 
                           DataPath_RF_bus_selected_win_data_178_port, Q(433) 
                           => DataPath_RF_bus_selected_win_data_177_port, 
                           Q(432) => DataPath_RF_bus_selected_win_data_176_port
                           , Q(431) => 
                           DataPath_RF_bus_selected_win_data_175_port, Q(430) 
                           => DataPath_RF_bus_selected_win_data_174_port, 
                           Q(429) => DataPath_RF_bus_selected_win_data_173_port
                           , Q(428) => 
                           DataPath_RF_bus_selected_win_data_172_port, Q(427) 
                           => DataPath_RF_bus_selected_win_data_171_port, 
                           Q(426) => DataPath_RF_bus_selected_win_data_170_port
                           , Q(425) => 
                           DataPath_RF_bus_selected_win_data_169_port, Q(424) 
                           => DataPath_RF_bus_selected_win_data_168_port, 
                           Q(423) => DataPath_RF_bus_selected_win_data_167_port
                           , Q(422) => 
                           DataPath_RF_bus_selected_win_data_166_port, Q(421) 
                           => DataPath_RF_bus_selected_win_data_165_port, 
                           Q(420) => DataPath_RF_bus_selected_win_data_164_port
                           , Q(419) => 
                           DataPath_RF_bus_selected_win_data_163_port, Q(418) 
                           => DataPath_RF_bus_selected_win_data_162_port, 
                           Q(417) => DataPath_RF_bus_selected_win_data_161_port
                           , Q(416) => 
                           DataPath_RF_bus_selected_win_data_160_port, Q(415) 
                           => DataPath_RF_bus_selected_win_data_159_port, 
                           Q(414) => DataPath_RF_bus_selected_win_data_158_port
                           , Q(413) => 
                           DataPath_RF_bus_selected_win_data_157_port, Q(412) 
                           => DataPath_RF_bus_selected_win_data_156_port, 
                           Q(411) => DataPath_RF_bus_selected_win_data_155_port
                           , Q(410) => 
                           DataPath_RF_bus_selected_win_data_154_port, Q(409) 
                           => DataPath_RF_bus_selected_win_data_153_port, 
                           Q(408) => DataPath_RF_bus_selected_win_data_152_port
                           , Q(407) => 
                           DataPath_RF_bus_selected_win_data_151_port, Q(406) 
                           => DataPath_RF_bus_selected_win_data_150_port, 
                           Q(405) => DataPath_RF_bus_selected_win_data_149_port
                           , Q(404) => 
                           DataPath_RF_bus_selected_win_data_148_port, Q(403) 
                           => DataPath_RF_bus_selected_win_data_147_port, 
                           Q(402) => DataPath_RF_bus_selected_win_data_146_port
                           , Q(401) => 
                           DataPath_RF_bus_selected_win_data_145_port, Q(400) 
                           => DataPath_RF_bus_selected_win_data_144_port, 
                           Q(399) => DataPath_RF_bus_selected_win_data_143_port
                           , Q(398) => 
                           DataPath_RF_bus_selected_win_data_142_port, Q(397) 
                           => DataPath_RF_bus_selected_win_data_141_port, 
                           Q(396) => DataPath_RF_bus_selected_win_data_140_port
                           , Q(395) => 
                           DataPath_RF_bus_selected_win_data_139_port, Q(394) 
                           => DataPath_RF_bus_selected_win_data_138_port, 
                           Q(393) => DataPath_RF_bus_selected_win_data_137_port
                           , Q(392) => 
                           DataPath_RF_bus_selected_win_data_136_port, Q(391) 
                           => DataPath_RF_bus_selected_win_data_135_port, 
                           Q(390) => DataPath_RF_bus_selected_win_data_134_port
                           , Q(389) => 
                           DataPath_RF_bus_selected_win_data_133_port, Q(388) 
                           => DataPath_RF_bus_selected_win_data_132_port, 
                           Q(387) => DataPath_RF_bus_selected_win_data_131_port
                           , Q(386) => 
                           DataPath_RF_bus_selected_win_data_130_port, Q(385) 
                           => DataPath_RF_bus_selected_win_data_129_port, 
                           Q(384) => DataPath_RF_bus_selected_win_data_128_port
                           , Q(383) => 
                           DataPath_RF_bus_selected_win_data_127_port, Q(382) 
                           => DataPath_RF_bus_selected_win_data_126_port, 
                           Q(381) => DataPath_RF_bus_selected_win_data_125_port
                           , Q(380) => 
                           DataPath_RF_bus_selected_win_data_124_port, Q(379) 
                           => DataPath_RF_bus_selected_win_data_123_port, 
                           Q(378) => DataPath_RF_bus_selected_win_data_122_port
                           , Q(377) => 
                           DataPath_RF_bus_selected_win_data_121_port, Q(376) 
                           => DataPath_RF_bus_selected_win_data_120_port, 
                           Q(375) => DataPath_RF_bus_selected_win_data_119_port
                           , Q(374) => 
                           DataPath_RF_bus_selected_win_data_118_port, Q(373) 
                           => DataPath_RF_bus_selected_win_data_117_port, 
                           Q(372) => DataPath_RF_bus_selected_win_data_116_port
                           , Q(371) => 
                           DataPath_RF_bus_selected_win_data_115_port, Q(370) 
                           => DataPath_RF_bus_selected_win_data_114_port, 
                           Q(369) => DataPath_RF_bus_selected_win_data_113_port
                           , Q(368) => 
                           DataPath_RF_bus_selected_win_data_112_port, Q(367) 
                           => DataPath_RF_bus_selected_win_data_111_port, 
                           Q(366) => DataPath_RF_bus_selected_win_data_110_port
                           , Q(365) => 
                           DataPath_RF_bus_selected_win_data_109_port, Q(364) 
                           => DataPath_RF_bus_selected_win_data_108_port, 
                           Q(363) => DataPath_RF_bus_selected_win_data_107_port
                           , Q(362) => 
                           DataPath_RF_bus_selected_win_data_106_port, Q(361) 
                           => DataPath_RF_bus_selected_win_data_105_port, 
                           Q(360) => DataPath_RF_bus_selected_win_data_104_port
                           , Q(359) => 
                           DataPath_RF_bus_selected_win_data_103_port, Q(358) 
                           => DataPath_RF_bus_selected_win_data_102_port, 
                           Q(357) => DataPath_RF_bus_selected_win_data_101_port
                           , Q(356) => 
                           DataPath_RF_bus_selected_win_data_100_port, Q(355) 
                           => DataPath_RF_bus_selected_win_data_99_port, Q(354)
                           => DataPath_RF_bus_selected_win_data_98_port, Q(353)
                           => DataPath_RF_bus_selected_win_data_97_port, Q(352)
                           => DataPath_RF_bus_selected_win_data_96_port, Q(351)
                           => DataPath_RF_bus_selected_win_data_95_port, Q(350)
                           => DataPath_RF_bus_selected_win_data_94_port, Q(349)
                           => DataPath_RF_bus_selected_win_data_93_port, Q(348)
                           => DataPath_RF_bus_selected_win_data_92_port, Q(347)
                           => DataPath_RF_bus_selected_win_data_91_port, Q(346)
                           => DataPath_RF_bus_selected_win_data_90_port, Q(345)
                           => DataPath_RF_bus_selected_win_data_89_port, Q(344)
                           => DataPath_RF_bus_selected_win_data_88_port, Q(343)
                           => DataPath_RF_bus_selected_win_data_87_port, Q(342)
                           => DataPath_RF_bus_selected_win_data_86_port, Q(341)
                           => DataPath_RF_bus_selected_win_data_85_port, Q(340)
                           => DataPath_RF_bus_selected_win_data_84_port, Q(339)
                           => DataPath_RF_bus_selected_win_data_83_port, Q(338)
                           => DataPath_RF_bus_selected_win_data_82_port, Q(337)
                           => DataPath_RF_bus_selected_win_data_81_port, Q(336)
                           => DataPath_RF_bus_selected_win_data_80_port, Q(335)
                           => DataPath_RF_bus_selected_win_data_79_port, Q(334)
                           => DataPath_RF_bus_selected_win_data_78_port, Q(333)
                           => DataPath_RF_bus_selected_win_data_77_port, Q(332)
                           => DataPath_RF_bus_selected_win_data_76_port, Q(331)
                           => DataPath_RF_bus_selected_win_data_75_port, Q(330)
                           => DataPath_RF_bus_selected_win_data_74_port, Q(329)
                           => DataPath_RF_bus_selected_win_data_73_port, Q(328)
                           => DataPath_RF_bus_selected_win_data_72_port, Q(327)
                           => DataPath_RF_bus_selected_win_data_71_port, Q(326)
                           => DataPath_RF_bus_selected_win_data_70_port, Q(325)
                           => DataPath_RF_bus_selected_win_data_69_port, Q(324)
                           => DataPath_RF_bus_selected_win_data_68_port, Q(323)
                           => DataPath_RF_bus_selected_win_data_67_port, Q(322)
                           => DataPath_RF_bus_selected_win_data_66_port, Q(321)
                           => DataPath_RF_bus_selected_win_data_65_port, Q(320)
                           => DataPath_RF_bus_selected_win_data_64_port, Q(319)
                           => DataPath_RF_bus_selected_win_data_63_port, Q(318)
                           => DataPath_RF_bus_selected_win_data_62_port, Q(317)
                           => DataPath_RF_bus_selected_win_data_61_port, Q(316)
                           => DataPath_RF_bus_selected_win_data_60_port, Q(315)
                           => DataPath_RF_bus_selected_win_data_59_port, Q(314)
                           => DataPath_RF_bus_selected_win_data_58_port, Q(313)
                           => DataPath_RF_bus_selected_win_data_57_port, Q(312)
                           => DataPath_RF_bus_selected_win_data_56_port, Q(311)
                           => DataPath_RF_bus_selected_win_data_55_port, Q(310)
                           => DataPath_RF_bus_selected_win_data_54_port, Q(309)
                           => DataPath_RF_bus_selected_win_data_53_port, Q(308)
                           => DataPath_RF_bus_selected_win_data_52_port, Q(307)
                           => DataPath_RF_bus_selected_win_data_51_port, Q(306)
                           => DataPath_RF_bus_selected_win_data_50_port, Q(305)
                           => DataPath_RF_bus_selected_win_data_49_port, Q(304)
                           => DataPath_RF_bus_selected_win_data_48_port, Q(303)
                           => DataPath_RF_bus_selected_win_data_47_port, Q(302)
                           => DataPath_RF_bus_selected_win_data_46_port, Q(301)
                           => DataPath_RF_bus_selected_win_data_45_port, Q(300)
                           => DataPath_RF_bus_selected_win_data_44_port, Q(299)
                           => DataPath_RF_bus_selected_win_data_43_port, Q(298)
                           => DataPath_RF_bus_selected_win_data_42_port, Q(297)
                           => DataPath_RF_bus_selected_win_data_41_port, Q(296)
                           => DataPath_RF_bus_selected_win_data_40_port, Q(295)
                           => DataPath_RF_bus_selected_win_data_39_port, Q(294)
                           => DataPath_RF_bus_selected_win_data_38_port, Q(293)
                           => DataPath_RF_bus_selected_win_data_37_port, Q(292)
                           => DataPath_RF_bus_selected_win_data_36_port, Q(291)
                           => DataPath_RF_bus_selected_win_data_35_port, Q(290)
                           => DataPath_RF_bus_selected_win_data_34_port, Q(289)
                           => DataPath_RF_bus_selected_win_data_33_port, Q(288)
                           => DataPath_RF_bus_selected_win_data_32_port, Q(287)
                           => DataPath_RF_bus_selected_win_data_31_port, Q(286)
                           => DataPath_RF_bus_selected_win_data_30_port, Q(285)
                           => DataPath_RF_bus_selected_win_data_29_port, Q(284)
                           => DataPath_RF_bus_selected_win_data_28_port, Q(283)
                           => DataPath_RF_bus_selected_win_data_27_port, Q(282)
                           => DataPath_RF_bus_selected_win_data_26_port, Q(281)
                           => DataPath_RF_bus_selected_win_data_25_port, Q(280)
                           => DataPath_RF_bus_selected_win_data_24_port, Q(279)
                           => DataPath_RF_bus_selected_win_data_23_port, Q(278)
                           => DataPath_RF_bus_selected_win_data_22_port, Q(277)
                           => DataPath_RF_bus_selected_win_data_21_port, Q(276)
                           => DataPath_RF_bus_selected_win_data_20_port, Q(275)
                           => DataPath_RF_bus_selected_win_data_19_port, Q(274)
                           => DataPath_RF_bus_selected_win_data_18_port, Q(273)
                           => DataPath_RF_bus_selected_win_data_17_port, Q(272)
                           => DataPath_RF_bus_selected_win_data_16_port, Q(271)
                           => DataPath_RF_bus_selected_win_data_15_port, Q(270)
                           => DataPath_RF_bus_selected_win_data_14_port, Q(269)
                           => DataPath_RF_bus_selected_win_data_13_port, Q(268)
                           => DataPath_RF_bus_selected_win_data_12_port, Q(267)
                           => DataPath_RF_bus_selected_win_data_11_port, Q(266)
                           => DataPath_RF_bus_selected_win_data_10_port, Q(265)
                           => DataPath_RF_bus_selected_win_data_9_port, Q(264) 
                           => DataPath_RF_bus_selected_win_data_8_port, Q(263) 
                           => DataPath_RF_bus_selected_win_data_7_port, Q(262) 
                           => DataPath_RF_bus_selected_win_data_6_port, Q(261) 
                           => DataPath_RF_bus_selected_win_data_5_port, Q(260) 
                           => DataPath_RF_bus_selected_win_data_4_port, Q(259) 
                           => DataPath_RF_bus_selected_win_data_3_port, Q(258) 
                           => DataPath_RF_bus_selected_win_data_2_port, Q(257) 
                           => DataPath_RF_bus_selected_win_data_1_port, Q(256) 
                           => DataPath_RF_bus_selected_win_data_0_port, Q(255) 
                           => DataPath_RF_bus_complete_win_data_255_port, 
                           Q(254) => DataPath_RF_bus_complete_win_data_254_port
                           , Q(253) => 
                           DataPath_RF_bus_complete_win_data_253_port, Q(252) 
                           => DataPath_RF_bus_complete_win_data_252_port, 
                           Q(251) => DataPath_RF_bus_complete_win_data_251_port
                           , Q(250) => 
                           DataPath_RF_bus_complete_win_data_250_port, Q(249) 
                           => DataPath_RF_bus_complete_win_data_249_port, 
                           Q(248) => DataPath_RF_bus_complete_win_data_248_port
                           , Q(247) => 
                           DataPath_RF_bus_complete_win_data_247_port, Q(246) 
                           => DataPath_RF_bus_complete_win_data_246_port, 
                           Q(245) => DataPath_RF_bus_complete_win_data_245_port
                           , Q(244) => 
                           DataPath_RF_bus_complete_win_data_244_port, Q(243) 
                           => DataPath_RF_bus_complete_win_data_243_port, 
                           Q(242) => DataPath_RF_bus_complete_win_data_242_port
                           , Q(241) => 
                           DataPath_RF_bus_complete_win_data_241_port, Q(240) 
                           => DataPath_RF_bus_complete_win_data_240_port, 
                           Q(239) => DataPath_RF_bus_complete_win_data_239_port
                           , Q(238) => 
                           DataPath_RF_bus_complete_win_data_238_port, Q(237) 
                           => DataPath_RF_bus_complete_win_data_237_port, 
                           Q(236) => DataPath_RF_bus_complete_win_data_236_port
                           , Q(235) => 
                           DataPath_RF_bus_complete_win_data_235_port, Q(234) 
                           => DataPath_RF_bus_complete_win_data_234_port, 
                           Q(233) => DataPath_RF_bus_complete_win_data_233_port
                           , Q(232) => 
                           DataPath_RF_bus_complete_win_data_232_port, Q(231) 
                           => DataPath_RF_bus_complete_win_data_231_port, 
                           Q(230) => DataPath_RF_bus_complete_win_data_230_port
                           , Q(229) => 
                           DataPath_RF_bus_complete_win_data_229_port, Q(228) 
                           => DataPath_RF_bus_complete_win_data_228_port, 
                           Q(227) => DataPath_RF_bus_complete_win_data_227_port
                           , Q(226) => 
                           DataPath_RF_bus_complete_win_data_226_port, Q(225) 
                           => DataPath_RF_bus_complete_win_data_225_port, 
                           Q(224) => DataPath_RF_bus_complete_win_data_224_port
                           , Q(223) => 
                           DataPath_RF_bus_complete_win_data_223_port, Q(222) 
                           => DataPath_RF_bus_complete_win_data_222_port, 
                           Q(221) => DataPath_RF_bus_complete_win_data_221_port
                           , Q(220) => 
                           DataPath_RF_bus_complete_win_data_220_port, Q(219) 
                           => DataPath_RF_bus_complete_win_data_219_port, 
                           Q(218) => DataPath_RF_bus_complete_win_data_218_port
                           , Q(217) => 
                           DataPath_RF_bus_complete_win_data_217_port, Q(216) 
                           => DataPath_RF_bus_complete_win_data_216_port, 
                           Q(215) => DataPath_RF_bus_complete_win_data_215_port
                           , Q(214) => 
                           DataPath_RF_bus_complete_win_data_214_port, Q(213) 
                           => DataPath_RF_bus_complete_win_data_213_port, 
                           Q(212) => DataPath_RF_bus_complete_win_data_212_port
                           , Q(211) => 
                           DataPath_RF_bus_complete_win_data_211_port, Q(210) 
                           => DataPath_RF_bus_complete_win_data_210_port, 
                           Q(209) => DataPath_RF_bus_complete_win_data_209_port
                           , Q(208) => 
                           DataPath_RF_bus_complete_win_data_208_port, Q(207) 
                           => DataPath_RF_bus_complete_win_data_207_port, 
                           Q(206) => DataPath_RF_bus_complete_win_data_206_port
                           , Q(205) => 
                           DataPath_RF_bus_complete_win_data_205_port, Q(204) 
                           => DataPath_RF_bus_complete_win_data_204_port, 
                           Q(203) => DataPath_RF_bus_complete_win_data_203_port
                           , Q(202) => 
                           DataPath_RF_bus_complete_win_data_202_port, Q(201) 
                           => DataPath_RF_bus_complete_win_data_201_port, 
                           Q(200) => DataPath_RF_bus_complete_win_data_200_port
                           , Q(199) => 
                           DataPath_RF_bus_complete_win_data_199_port, Q(198) 
                           => DataPath_RF_bus_complete_win_data_198_port, 
                           Q(197) => DataPath_RF_bus_complete_win_data_197_port
                           , Q(196) => 
                           DataPath_RF_bus_complete_win_data_196_port, Q(195) 
                           => DataPath_RF_bus_complete_win_data_195_port, 
                           Q(194) => DataPath_RF_bus_complete_win_data_194_port
                           , Q(193) => 
                           DataPath_RF_bus_complete_win_data_193_port, Q(192) 
                           => DataPath_RF_bus_complete_win_data_192_port, 
                           Q(191) => DataPath_RF_bus_complete_win_data_191_port
                           , Q(190) => 
                           DataPath_RF_bus_complete_win_data_190_port, Q(189) 
                           => DataPath_RF_bus_complete_win_data_189_port, 
                           Q(188) => DataPath_RF_bus_complete_win_data_188_port
                           , Q(187) => 
                           DataPath_RF_bus_complete_win_data_187_port, Q(186) 
                           => DataPath_RF_bus_complete_win_data_186_port, 
                           Q(185) => DataPath_RF_bus_complete_win_data_185_port
                           , Q(184) => 
                           DataPath_RF_bus_complete_win_data_184_port, Q(183) 
                           => DataPath_RF_bus_complete_win_data_183_port, 
                           Q(182) => DataPath_RF_bus_complete_win_data_182_port
                           , Q(181) => 
                           DataPath_RF_bus_complete_win_data_181_port, Q(180) 
                           => DataPath_RF_bus_complete_win_data_180_port, 
                           Q(179) => DataPath_RF_bus_complete_win_data_179_port
                           , Q(178) => 
                           DataPath_RF_bus_complete_win_data_178_port, Q(177) 
                           => DataPath_RF_bus_complete_win_data_177_port, 
                           Q(176) => DataPath_RF_bus_complete_win_data_176_port
                           , Q(175) => 
                           DataPath_RF_bus_complete_win_data_175_port, Q(174) 
                           => DataPath_RF_bus_complete_win_data_174_port, 
                           Q(173) => DataPath_RF_bus_complete_win_data_173_port
                           , Q(172) => 
                           DataPath_RF_bus_complete_win_data_172_port, Q(171) 
                           => DataPath_RF_bus_complete_win_data_171_port, 
                           Q(170) => DataPath_RF_bus_complete_win_data_170_port
                           , Q(169) => 
                           DataPath_RF_bus_complete_win_data_169_port, Q(168) 
                           => DataPath_RF_bus_complete_win_data_168_port, 
                           Q(167) => DataPath_RF_bus_complete_win_data_167_port
                           , Q(166) => 
                           DataPath_RF_bus_complete_win_data_166_port, Q(165) 
                           => DataPath_RF_bus_complete_win_data_165_port, 
                           Q(164) => DataPath_RF_bus_complete_win_data_164_port
                           , Q(163) => 
                           DataPath_RF_bus_complete_win_data_163_port, Q(162) 
                           => DataPath_RF_bus_complete_win_data_162_port, 
                           Q(161) => DataPath_RF_bus_complete_win_data_161_port
                           , Q(160) => 
                           DataPath_RF_bus_complete_win_data_160_port, Q(159) 
                           => DataPath_RF_bus_complete_win_data_159_port, 
                           Q(158) => DataPath_RF_bus_complete_win_data_158_port
                           , Q(157) => 
                           DataPath_RF_bus_complete_win_data_157_port, Q(156) 
                           => DataPath_RF_bus_complete_win_data_156_port, 
                           Q(155) => DataPath_RF_bus_complete_win_data_155_port
                           , Q(154) => 
                           DataPath_RF_bus_complete_win_data_154_port, Q(153) 
                           => DataPath_RF_bus_complete_win_data_153_port, 
                           Q(152) => DataPath_RF_bus_complete_win_data_152_port
                           , Q(151) => 
                           DataPath_RF_bus_complete_win_data_151_port, Q(150) 
                           => DataPath_RF_bus_complete_win_data_150_port, 
                           Q(149) => DataPath_RF_bus_complete_win_data_149_port
                           , Q(148) => 
                           DataPath_RF_bus_complete_win_data_148_port, Q(147) 
                           => DataPath_RF_bus_complete_win_data_147_port, 
                           Q(146) => DataPath_RF_bus_complete_win_data_146_port
                           , Q(145) => 
                           DataPath_RF_bus_complete_win_data_145_port, Q(144) 
                           => DataPath_RF_bus_complete_win_data_144_port, 
                           Q(143) => DataPath_RF_bus_complete_win_data_143_port
                           , Q(142) => 
                           DataPath_RF_bus_complete_win_data_142_port, Q(141) 
                           => DataPath_RF_bus_complete_win_data_141_port, 
                           Q(140) => DataPath_RF_bus_complete_win_data_140_port
                           , Q(139) => 
                           DataPath_RF_bus_complete_win_data_139_port, Q(138) 
                           => DataPath_RF_bus_complete_win_data_138_port, 
                           Q(137) => DataPath_RF_bus_complete_win_data_137_port
                           , Q(136) => 
                           DataPath_RF_bus_complete_win_data_136_port, Q(135) 
                           => DataPath_RF_bus_complete_win_data_135_port, 
                           Q(134) => DataPath_RF_bus_complete_win_data_134_port
                           , Q(133) => 
                           DataPath_RF_bus_complete_win_data_133_port, Q(132) 
                           => DataPath_RF_bus_complete_win_data_132_port, 
                           Q(131) => DataPath_RF_bus_complete_win_data_131_port
                           , Q(130) => 
                           DataPath_RF_bus_complete_win_data_130_port, Q(129) 
                           => DataPath_RF_bus_complete_win_data_129_port, 
                           Q(128) => DataPath_RF_bus_complete_win_data_128_port
                           , Q(127) => 
                           DataPath_RF_bus_complete_win_data_127_port, Q(126) 
                           => DataPath_RF_bus_complete_win_data_126_port, 
                           Q(125) => DataPath_RF_bus_complete_win_data_125_port
                           , Q(124) => 
                           DataPath_RF_bus_complete_win_data_124_port, Q(123) 
                           => DataPath_RF_bus_complete_win_data_123_port, 
                           Q(122) => DataPath_RF_bus_complete_win_data_122_port
                           , Q(121) => 
                           DataPath_RF_bus_complete_win_data_121_port, Q(120) 
                           => DataPath_RF_bus_complete_win_data_120_port, 
                           Q(119) => DataPath_RF_bus_complete_win_data_119_port
                           , Q(118) => 
                           DataPath_RF_bus_complete_win_data_118_port, Q(117) 
                           => DataPath_RF_bus_complete_win_data_117_port, 
                           Q(116) => DataPath_RF_bus_complete_win_data_116_port
                           , Q(115) => 
                           DataPath_RF_bus_complete_win_data_115_port, Q(114) 
                           => DataPath_RF_bus_complete_win_data_114_port, 
                           Q(113) => DataPath_RF_bus_complete_win_data_113_port
                           , Q(112) => 
                           DataPath_RF_bus_complete_win_data_112_port, Q(111) 
                           => DataPath_RF_bus_complete_win_data_111_port, 
                           Q(110) => DataPath_RF_bus_complete_win_data_110_port
                           , Q(109) => 
                           DataPath_RF_bus_complete_win_data_109_port, Q(108) 
                           => DataPath_RF_bus_complete_win_data_108_port, 
                           Q(107) => DataPath_RF_bus_complete_win_data_107_port
                           , Q(106) => 
                           DataPath_RF_bus_complete_win_data_106_port, Q(105) 
                           => DataPath_RF_bus_complete_win_data_105_port, 
                           Q(104) => DataPath_RF_bus_complete_win_data_104_port
                           , Q(103) => 
                           DataPath_RF_bus_complete_win_data_103_port, Q(102) 
                           => DataPath_RF_bus_complete_win_data_102_port, 
                           Q(101) => DataPath_RF_bus_complete_win_data_101_port
                           , Q(100) => 
                           DataPath_RF_bus_complete_win_data_100_port, Q(99) =>
                           DataPath_RF_bus_complete_win_data_99_port, Q(98) => 
                           DataPath_RF_bus_complete_win_data_98_port, Q(97) => 
                           DataPath_RF_bus_complete_win_data_97_port, Q(96) => 
                           DataPath_RF_bus_complete_win_data_96_port, Q(95) => 
                           DataPath_RF_bus_complete_win_data_95_port, Q(94) => 
                           DataPath_RF_bus_complete_win_data_94_port, Q(93) => 
                           DataPath_RF_bus_complete_win_data_93_port, Q(92) => 
                           DataPath_RF_bus_complete_win_data_92_port, Q(91) => 
                           DataPath_RF_bus_complete_win_data_91_port, Q(90) => 
                           DataPath_RF_bus_complete_win_data_90_port, Q(89) => 
                           DataPath_RF_bus_complete_win_data_89_port, Q(88) => 
                           DataPath_RF_bus_complete_win_data_88_port, Q(87) => 
                           DataPath_RF_bus_complete_win_data_87_port, Q(86) => 
                           DataPath_RF_bus_complete_win_data_86_port, Q(85) => 
                           DataPath_RF_bus_complete_win_data_85_port, Q(84) => 
                           DataPath_RF_bus_complete_win_data_84_port, Q(83) => 
                           DataPath_RF_bus_complete_win_data_83_port, Q(82) => 
                           DataPath_RF_bus_complete_win_data_82_port, Q(81) => 
                           DataPath_RF_bus_complete_win_data_81_port, Q(80) => 
                           DataPath_RF_bus_complete_win_data_80_port, Q(79) => 
                           DataPath_RF_bus_complete_win_data_79_port, Q(78) => 
                           DataPath_RF_bus_complete_win_data_78_port, Q(77) => 
                           DataPath_RF_bus_complete_win_data_77_port, Q(76) => 
                           DataPath_RF_bus_complete_win_data_76_port, Q(75) => 
                           DataPath_RF_bus_complete_win_data_75_port, Q(74) => 
                           DataPath_RF_bus_complete_win_data_74_port, Q(73) => 
                           DataPath_RF_bus_complete_win_data_73_port, Q(72) => 
                           DataPath_RF_bus_complete_win_data_72_port, Q(71) => 
                           DataPath_RF_bus_complete_win_data_71_port, Q(70) => 
                           DataPath_RF_bus_complete_win_data_70_port, Q(69) => 
                           DataPath_RF_bus_complete_win_data_69_port, Q(68) => 
                           DataPath_RF_bus_complete_win_data_68_port, Q(67) => 
                           DataPath_RF_bus_complete_win_data_67_port, Q(66) => 
                           DataPath_RF_bus_complete_win_data_66_port, Q(65) => 
                           DataPath_RF_bus_complete_win_data_65_port, Q(64) => 
                           DataPath_RF_bus_complete_win_data_64_port, Q(63) => 
                           DataPath_RF_bus_complete_win_data_63_port, Q(62) => 
                           DataPath_RF_bus_complete_win_data_62_port, Q(61) => 
                           DataPath_RF_bus_complete_win_data_61_port, Q(60) => 
                           DataPath_RF_bus_complete_win_data_60_port, Q(59) => 
                           DataPath_RF_bus_complete_win_data_59_port, Q(58) => 
                           DataPath_RF_bus_complete_win_data_58_port, Q(57) => 
                           DataPath_RF_bus_complete_win_data_57_port, Q(56) => 
                           DataPath_RF_bus_complete_win_data_56_port, Q(55) => 
                           DataPath_RF_bus_complete_win_data_55_port, Q(54) => 
                           DataPath_RF_bus_complete_win_data_54_port, Q(53) => 
                           DataPath_RF_bus_complete_win_data_53_port, Q(52) => 
                           DataPath_RF_bus_complete_win_data_52_port, Q(51) => 
                           DataPath_RF_bus_complete_win_data_51_port, Q(50) => 
                           DataPath_RF_bus_complete_win_data_50_port, Q(49) => 
                           DataPath_RF_bus_complete_win_data_49_port, Q(48) => 
                           DataPath_RF_bus_complete_win_data_48_port, Q(47) => 
                           DataPath_RF_bus_complete_win_data_47_port, Q(46) => 
                           DataPath_RF_bus_complete_win_data_46_port, Q(45) => 
                           DataPath_RF_bus_complete_win_data_45_port, Q(44) => 
                           DataPath_RF_bus_complete_win_data_44_port, Q(43) => 
                           DataPath_RF_bus_complete_win_data_43_port, Q(42) => 
                           DataPath_RF_bus_complete_win_data_42_port, Q(41) => 
                           DataPath_RF_bus_complete_win_data_41_port, Q(40) => 
                           DataPath_RF_bus_complete_win_data_40_port, Q(39) => 
                           DataPath_RF_bus_complete_win_data_39_port, Q(38) => 
                           DataPath_RF_bus_complete_win_data_38_port, Q(37) => 
                           DataPath_RF_bus_complete_win_data_37_port, Q(36) => 
                           DataPath_RF_bus_complete_win_data_36_port, Q(35) => 
                           DataPath_RF_bus_complete_win_data_35_port, Q(34) => 
                           DataPath_RF_bus_complete_win_data_34_port, Q(33) => 
                           DataPath_RF_bus_complete_win_data_33_port, Q(32) => 
                           DataPath_RF_bus_complete_win_data_32_port, Q(31) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(30) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(29) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(28) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(27) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(26) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(25) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(24) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(23) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(22) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(21) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(20) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(19) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(18) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(17) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(16) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(15) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(14) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(13) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(12) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(11) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(10) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(9) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(8) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(7) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(6) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(5) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(4) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(3) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(2) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(1) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(0) => 
                           DataPath_RF_bus_complete_win_data_0_port, Y(31) => 
                           DataPath_RF_internal_out1_31_port, Y(30) => 
                           DataPath_RF_internal_out1_30_port, Y(29) => 
                           DataPath_RF_internal_out1_29_port, Y(28) => 
                           DataPath_RF_internal_out1_28_port, Y(27) => 
                           DataPath_RF_internal_out1_27_port, Y(26) => 
                           DataPath_RF_internal_out1_26_port, Y(25) => 
                           DataPath_RF_internal_out1_25_port, Y(24) => 
                           DataPath_RF_internal_out1_24_port, Y(23) => 
                           DataPath_RF_internal_out1_23_port, Y(22) => 
                           DataPath_RF_internal_out1_22_port, Y(21) => 
                           DataPath_RF_internal_out1_21_port, Y(20) => 
                           DataPath_RF_internal_out1_20_port, Y(19) => 
                           DataPath_RF_internal_out1_19_port, Y(18) => 
                           DataPath_RF_internal_out1_18_port, Y(17) => 
                           DataPath_RF_internal_out1_17_port, Y(16) => 
                           DataPath_RF_internal_out1_16_port, Y(15) => 
                           DataPath_RF_internal_out1_15_port, Y(14) => 
                           DataPath_RF_internal_out1_14_port, Y(13) => 
                           DataPath_RF_internal_out1_13_port, Y(12) => 
                           DataPath_RF_internal_out1_12_port, Y(11) => 
                           DataPath_RF_internal_out1_11_port, Y(10) => 
                           DataPath_RF_internal_out1_10_port, Y(9) => 
                           DataPath_RF_internal_out1_9_port, Y(8) => 
                           DataPath_RF_internal_out1_8_port, Y(7) => 
                           DataPath_RF_internal_out1_7_port, Y(6) => 
                           DataPath_RF_internal_out1_6_port, Y(5) => 
                           DataPath_RF_internal_out1_5_port, Y(4) => 
                           DataPath_RF_internal_out1_4_port, Y(3) => 
                           DataPath_RF_internal_out1_3_port, Y(2) => 
                           DataPath_RF_internal_out1_2_port, Y(1) => 
                           DataPath_RF_internal_out1_1_port, Y(0) => 
                           DataPath_RF_internal_out1_0_port);
   DataPath_RF_SEL_BLK : select_block_NBIT_DATA32_N8_F5 port map( regs(2559) =>
                           DataPath_RF_bus_reg_dataout_2559_port, regs(2558) =>
                           DataPath_RF_bus_reg_dataout_2558_port, regs(2557) =>
                           DataPath_RF_bus_reg_dataout_2557_port, regs(2556) =>
                           DataPath_RF_bus_reg_dataout_2556_port, regs(2555) =>
                           DataPath_RF_bus_reg_dataout_2555_port, regs(2554) =>
                           DataPath_RF_bus_reg_dataout_2554_port, regs(2553) =>
                           DataPath_RF_bus_reg_dataout_2553_port, regs(2552) =>
                           DataPath_RF_bus_reg_dataout_2552_port, regs(2551) =>
                           DataPath_RF_bus_reg_dataout_2551_port, regs(2550) =>
                           DataPath_RF_bus_reg_dataout_2550_port, regs(2549) =>
                           DataPath_RF_bus_reg_dataout_2549_port, regs(2548) =>
                           DataPath_RF_bus_reg_dataout_2548_port, regs(2547) =>
                           DataPath_RF_bus_reg_dataout_2547_port, regs(2546) =>
                           DataPath_RF_bus_reg_dataout_2546_port, regs(2545) =>
                           DataPath_RF_bus_reg_dataout_2545_port, regs(2544) =>
                           DataPath_RF_bus_reg_dataout_2544_port, regs(2543) =>
                           DataPath_RF_bus_reg_dataout_2543_port, regs(2542) =>
                           DataPath_RF_bus_reg_dataout_2542_port, regs(2541) =>
                           DataPath_RF_bus_reg_dataout_2541_port, regs(2540) =>
                           DataPath_RF_bus_reg_dataout_2540_port, regs(2539) =>
                           DataPath_RF_bus_reg_dataout_2539_port, regs(2538) =>
                           DataPath_RF_bus_reg_dataout_2538_port, regs(2537) =>
                           DataPath_RF_bus_reg_dataout_2537_port, regs(2536) =>
                           DataPath_RF_bus_reg_dataout_2536_port, regs(2535) =>
                           DataPath_RF_bus_reg_dataout_2535_port, regs(2534) =>
                           DataPath_RF_bus_reg_dataout_2534_port, regs(2533) =>
                           DataPath_RF_bus_reg_dataout_2533_port, regs(2532) =>
                           DataPath_RF_bus_reg_dataout_2532_port, regs(2531) =>
                           DataPath_RF_bus_reg_dataout_2531_port, regs(2530) =>
                           DataPath_RF_bus_reg_dataout_2530_port, regs(2529) =>
                           DataPath_RF_bus_reg_dataout_2529_port, regs(2528) =>
                           DataPath_RF_bus_reg_dataout_2528_port, regs(2527) =>
                           DataPath_RF_bus_reg_dataout_2527_port, regs(2526) =>
                           DataPath_RF_bus_reg_dataout_2526_port, regs(2525) =>
                           DataPath_RF_bus_reg_dataout_2525_port, regs(2524) =>
                           DataPath_RF_bus_reg_dataout_2524_port, regs(2523) =>
                           DataPath_RF_bus_reg_dataout_2523_port, regs(2522) =>
                           DataPath_RF_bus_reg_dataout_2522_port, regs(2521) =>
                           DataPath_RF_bus_reg_dataout_2521_port, regs(2520) =>
                           DataPath_RF_bus_reg_dataout_2520_port, regs(2519) =>
                           DataPath_RF_bus_reg_dataout_2519_port, regs(2518) =>
                           DataPath_RF_bus_reg_dataout_2518_port, regs(2517) =>
                           DataPath_RF_bus_reg_dataout_2517_port, regs(2516) =>
                           DataPath_RF_bus_reg_dataout_2516_port, regs(2515) =>
                           DataPath_RF_bus_reg_dataout_2515_port, regs(2514) =>
                           DataPath_RF_bus_reg_dataout_2514_port, regs(2513) =>
                           DataPath_RF_bus_reg_dataout_2513_port, regs(2512) =>
                           DataPath_RF_bus_reg_dataout_2512_port, regs(2511) =>
                           DataPath_RF_bus_reg_dataout_2511_port, regs(2510) =>
                           DataPath_RF_bus_reg_dataout_2510_port, regs(2509) =>
                           DataPath_RF_bus_reg_dataout_2509_port, regs(2508) =>
                           DataPath_RF_bus_reg_dataout_2508_port, regs(2507) =>
                           DataPath_RF_bus_reg_dataout_2507_port, regs(2506) =>
                           DataPath_RF_bus_reg_dataout_2506_port, regs(2505) =>
                           DataPath_RF_bus_reg_dataout_2505_port, regs(2504) =>
                           DataPath_RF_bus_reg_dataout_2504_port, regs(2503) =>
                           DataPath_RF_bus_reg_dataout_2503_port, regs(2502) =>
                           DataPath_RF_bus_reg_dataout_2502_port, regs(2501) =>
                           DataPath_RF_bus_reg_dataout_2501_port, regs(2500) =>
                           DataPath_RF_bus_reg_dataout_2500_port, regs(2499) =>
                           DataPath_RF_bus_reg_dataout_2499_port, regs(2498) =>
                           DataPath_RF_bus_reg_dataout_2498_port, regs(2497) =>
                           DataPath_RF_bus_reg_dataout_2497_port, regs(2496) =>
                           DataPath_RF_bus_reg_dataout_2496_port, regs(2495) =>
                           DataPath_RF_bus_reg_dataout_2495_port, regs(2494) =>
                           DataPath_RF_bus_reg_dataout_2494_port, regs(2493) =>
                           DataPath_RF_bus_reg_dataout_2493_port, regs(2492) =>
                           DataPath_RF_bus_reg_dataout_2492_port, regs(2491) =>
                           DataPath_RF_bus_reg_dataout_2491_port, regs(2490) =>
                           DataPath_RF_bus_reg_dataout_2490_port, regs(2489) =>
                           DataPath_RF_bus_reg_dataout_2489_port, regs(2488) =>
                           DataPath_RF_bus_reg_dataout_2488_port, regs(2487) =>
                           DataPath_RF_bus_reg_dataout_2487_port, regs(2486) =>
                           DataPath_RF_bus_reg_dataout_2486_port, regs(2485) =>
                           DataPath_RF_bus_reg_dataout_2485_port, regs(2484) =>
                           DataPath_RF_bus_reg_dataout_2484_port, regs(2483) =>
                           DataPath_RF_bus_reg_dataout_2483_port, regs(2482) =>
                           DataPath_RF_bus_reg_dataout_2482_port, regs(2481) =>
                           DataPath_RF_bus_reg_dataout_2481_port, regs(2480) =>
                           DataPath_RF_bus_reg_dataout_2480_port, regs(2479) =>
                           DataPath_RF_bus_reg_dataout_2479_port, regs(2478) =>
                           DataPath_RF_bus_reg_dataout_2478_port, regs(2477) =>
                           DataPath_RF_bus_reg_dataout_2477_port, regs(2476) =>
                           DataPath_RF_bus_reg_dataout_2476_port, regs(2475) =>
                           DataPath_RF_bus_reg_dataout_2475_port, regs(2474) =>
                           DataPath_RF_bus_reg_dataout_2474_port, regs(2473) =>
                           DataPath_RF_bus_reg_dataout_2473_port, regs(2472) =>
                           DataPath_RF_bus_reg_dataout_2472_port, regs(2471) =>
                           DataPath_RF_bus_reg_dataout_2471_port, regs(2470) =>
                           DataPath_RF_bus_reg_dataout_2470_port, regs(2469) =>
                           DataPath_RF_bus_reg_dataout_2469_port, regs(2468) =>
                           DataPath_RF_bus_reg_dataout_2468_port, regs(2467) =>
                           DataPath_RF_bus_reg_dataout_2467_port, regs(2466) =>
                           DataPath_RF_bus_reg_dataout_2466_port, regs(2465) =>
                           DataPath_RF_bus_reg_dataout_2465_port, regs(2464) =>
                           DataPath_RF_bus_reg_dataout_2464_port, regs(2463) =>
                           DataPath_RF_bus_reg_dataout_2463_port, regs(2462) =>
                           DataPath_RF_bus_reg_dataout_2462_port, regs(2461) =>
                           DataPath_RF_bus_reg_dataout_2461_port, regs(2460) =>
                           DataPath_RF_bus_reg_dataout_2460_port, regs(2459) =>
                           DataPath_RF_bus_reg_dataout_2459_port, regs(2458) =>
                           DataPath_RF_bus_reg_dataout_2458_port, regs(2457) =>
                           DataPath_RF_bus_reg_dataout_2457_port, regs(2456) =>
                           DataPath_RF_bus_reg_dataout_2456_port, regs(2455) =>
                           DataPath_RF_bus_reg_dataout_2455_port, regs(2454) =>
                           DataPath_RF_bus_reg_dataout_2454_port, regs(2453) =>
                           DataPath_RF_bus_reg_dataout_2453_port, regs(2452) =>
                           DataPath_RF_bus_reg_dataout_2452_port, regs(2451) =>
                           DataPath_RF_bus_reg_dataout_2451_port, regs(2450) =>
                           DataPath_RF_bus_reg_dataout_2450_port, regs(2449) =>
                           DataPath_RF_bus_reg_dataout_2449_port, regs(2448) =>
                           DataPath_RF_bus_reg_dataout_2448_port, regs(2447) =>
                           DataPath_RF_bus_reg_dataout_2447_port, regs(2446) =>
                           DataPath_RF_bus_reg_dataout_2446_port, regs(2445) =>
                           DataPath_RF_bus_reg_dataout_2445_port, regs(2444) =>
                           DataPath_RF_bus_reg_dataout_2444_port, regs(2443) =>
                           DataPath_RF_bus_reg_dataout_2443_port, regs(2442) =>
                           DataPath_RF_bus_reg_dataout_2442_port, regs(2441) =>
                           DataPath_RF_bus_reg_dataout_2441_port, regs(2440) =>
                           DataPath_RF_bus_reg_dataout_2440_port, regs(2439) =>
                           DataPath_RF_bus_reg_dataout_2439_port, regs(2438) =>
                           DataPath_RF_bus_reg_dataout_2438_port, regs(2437) =>
                           DataPath_RF_bus_reg_dataout_2437_port, regs(2436) =>
                           DataPath_RF_bus_reg_dataout_2436_port, regs(2435) =>
                           DataPath_RF_bus_reg_dataout_2435_port, regs(2434) =>
                           DataPath_RF_bus_reg_dataout_2434_port, regs(2433) =>
                           DataPath_RF_bus_reg_dataout_2433_port, regs(2432) =>
                           DataPath_RF_bus_reg_dataout_2432_port, regs(2431) =>
                           DataPath_RF_bus_reg_dataout_2431_port, regs(2430) =>
                           DataPath_RF_bus_reg_dataout_2430_port, regs(2429) =>
                           DataPath_RF_bus_reg_dataout_2429_port, regs(2428) =>
                           DataPath_RF_bus_reg_dataout_2428_port, regs(2427) =>
                           DataPath_RF_bus_reg_dataout_2427_port, regs(2426) =>
                           DataPath_RF_bus_reg_dataout_2426_port, regs(2425) =>
                           DataPath_RF_bus_reg_dataout_2425_port, regs(2424) =>
                           DataPath_RF_bus_reg_dataout_2424_port, regs(2423) =>
                           DataPath_RF_bus_reg_dataout_2423_port, regs(2422) =>
                           DataPath_RF_bus_reg_dataout_2422_port, regs(2421) =>
                           DataPath_RF_bus_reg_dataout_2421_port, regs(2420) =>
                           DataPath_RF_bus_reg_dataout_2420_port, regs(2419) =>
                           DataPath_RF_bus_reg_dataout_2419_port, regs(2418) =>
                           DataPath_RF_bus_reg_dataout_2418_port, regs(2417) =>
                           DataPath_RF_bus_reg_dataout_2417_port, regs(2416) =>
                           DataPath_RF_bus_reg_dataout_2416_port, regs(2415) =>
                           DataPath_RF_bus_reg_dataout_2415_port, regs(2414) =>
                           DataPath_RF_bus_reg_dataout_2414_port, regs(2413) =>
                           DataPath_RF_bus_reg_dataout_2413_port, regs(2412) =>
                           DataPath_RF_bus_reg_dataout_2412_port, regs(2411) =>
                           DataPath_RF_bus_reg_dataout_2411_port, regs(2410) =>
                           DataPath_RF_bus_reg_dataout_2410_port, regs(2409) =>
                           DataPath_RF_bus_reg_dataout_2409_port, regs(2408) =>
                           DataPath_RF_bus_reg_dataout_2408_port, regs(2407) =>
                           DataPath_RF_bus_reg_dataout_2407_port, regs(2406) =>
                           DataPath_RF_bus_reg_dataout_2406_port, regs(2405) =>
                           DataPath_RF_bus_reg_dataout_2405_port, regs(2404) =>
                           DataPath_RF_bus_reg_dataout_2404_port, regs(2403) =>
                           DataPath_RF_bus_reg_dataout_2403_port, regs(2402) =>
                           DataPath_RF_bus_reg_dataout_2402_port, regs(2401) =>
                           DataPath_RF_bus_reg_dataout_2401_port, regs(2400) =>
                           DataPath_RF_bus_reg_dataout_2400_port, regs(2399) =>
                           DataPath_RF_bus_reg_dataout_2399_port, regs(2398) =>
                           DataPath_RF_bus_reg_dataout_2398_port, regs(2397) =>
                           DataPath_RF_bus_reg_dataout_2397_port, regs(2396) =>
                           DataPath_RF_bus_reg_dataout_2396_port, regs(2395) =>
                           DataPath_RF_bus_reg_dataout_2395_port, regs(2394) =>
                           DataPath_RF_bus_reg_dataout_2394_port, regs(2393) =>
                           DataPath_RF_bus_reg_dataout_2393_port, regs(2392) =>
                           DataPath_RF_bus_reg_dataout_2392_port, regs(2391) =>
                           DataPath_RF_bus_reg_dataout_2391_port, regs(2390) =>
                           DataPath_RF_bus_reg_dataout_2390_port, regs(2389) =>
                           DataPath_RF_bus_reg_dataout_2389_port, regs(2388) =>
                           DataPath_RF_bus_reg_dataout_2388_port, regs(2387) =>
                           DataPath_RF_bus_reg_dataout_2387_port, regs(2386) =>
                           DataPath_RF_bus_reg_dataout_2386_port, regs(2385) =>
                           DataPath_RF_bus_reg_dataout_2385_port, regs(2384) =>
                           DataPath_RF_bus_reg_dataout_2384_port, regs(2383) =>
                           DataPath_RF_bus_reg_dataout_2383_port, regs(2382) =>
                           DataPath_RF_bus_reg_dataout_2382_port, regs(2381) =>
                           DataPath_RF_bus_reg_dataout_2381_port, regs(2380) =>
                           DataPath_RF_bus_reg_dataout_2380_port, regs(2379) =>
                           DataPath_RF_bus_reg_dataout_2379_port, regs(2378) =>
                           DataPath_RF_bus_reg_dataout_2378_port, regs(2377) =>
                           DataPath_RF_bus_reg_dataout_2377_port, regs(2376) =>
                           DataPath_RF_bus_reg_dataout_2376_port, regs(2375) =>
                           DataPath_RF_bus_reg_dataout_2375_port, regs(2374) =>
                           DataPath_RF_bus_reg_dataout_2374_port, regs(2373) =>
                           DataPath_RF_bus_reg_dataout_2373_port, regs(2372) =>
                           DataPath_RF_bus_reg_dataout_2372_port, regs(2371) =>
                           DataPath_RF_bus_reg_dataout_2371_port, regs(2370) =>
                           DataPath_RF_bus_reg_dataout_2370_port, regs(2369) =>
                           DataPath_RF_bus_reg_dataout_2369_port, regs(2368) =>
                           DataPath_RF_bus_reg_dataout_2368_port, regs(2367) =>
                           DataPath_RF_bus_reg_dataout_2367_port, regs(2366) =>
                           DataPath_RF_bus_reg_dataout_2366_port, regs(2365) =>
                           DataPath_RF_bus_reg_dataout_2365_port, regs(2364) =>
                           DataPath_RF_bus_reg_dataout_2364_port, regs(2363) =>
                           DataPath_RF_bus_reg_dataout_2363_port, regs(2362) =>
                           DataPath_RF_bus_reg_dataout_2362_port, regs(2361) =>
                           DataPath_RF_bus_reg_dataout_2361_port, regs(2360) =>
                           DataPath_RF_bus_reg_dataout_2360_port, regs(2359) =>
                           DataPath_RF_bus_reg_dataout_2359_port, regs(2358) =>
                           DataPath_RF_bus_reg_dataout_2358_port, regs(2357) =>
                           DataPath_RF_bus_reg_dataout_2357_port, regs(2356) =>
                           DataPath_RF_bus_reg_dataout_2356_port, regs(2355) =>
                           DataPath_RF_bus_reg_dataout_2355_port, regs(2354) =>
                           DataPath_RF_bus_reg_dataout_2354_port, regs(2353) =>
                           DataPath_RF_bus_reg_dataout_2353_port, regs(2352) =>
                           DataPath_RF_bus_reg_dataout_2352_port, regs(2351) =>
                           DataPath_RF_bus_reg_dataout_2351_port, regs(2350) =>
                           DataPath_RF_bus_reg_dataout_2350_port, regs(2349) =>
                           DataPath_RF_bus_reg_dataout_2349_port, regs(2348) =>
                           DataPath_RF_bus_reg_dataout_2348_port, regs(2347) =>
                           DataPath_RF_bus_reg_dataout_2347_port, regs(2346) =>
                           DataPath_RF_bus_reg_dataout_2346_port, regs(2345) =>
                           DataPath_RF_bus_reg_dataout_2345_port, regs(2344) =>
                           DataPath_RF_bus_reg_dataout_2344_port, regs(2343) =>
                           DataPath_RF_bus_reg_dataout_2343_port, regs(2342) =>
                           DataPath_RF_bus_reg_dataout_2342_port, regs(2341) =>
                           DataPath_RF_bus_reg_dataout_2341_port, regs(2340) =>
                           DataPath_RF_bus_reg_dataout_2340_port, regs(2339) =>
                           DataPath_RF_bus_reg_dataout_2339_port, regs(2338) =>
                           DataPath_RF_bus_reg_dataout_2338_port, regs(2337) =>
                           DataPath_RF_bus_reg_dataout_2337_port, regs(2336) =>
                           DataPath_RF_bus_reg_dataout_2336_port, regs(2335) =>
                           DataPath_RF_bus_reg_dataout_2335_port, regs(2334) =>
                           DataPath_RF_bus_reg_dataout_2334_port, regs(2333) =>
                           DataPath_RF_bus_reg_dataout_2333_port, regs(2332) =>
                           DataPath_RF_bus_reg_dataout_2332_port, regs(2331) =>
                           DataPath_RF_bus_reg_dataout_2331_port, regs(2330) =>
                           DataPath_RF_bus_reg_dataout_2330_port, regs(2329) =>
                           DataPath_RF_bus_reg_dataout_2329_port, regs(2328) =>
                           DataPath_RF_bus_reg_dataout_2328_port, regs(2327) =>
                           DataPath_RF_bus_reg_dataout_2327_port, regs(2326) =>
                           DataPath_RF_bus_reg_dataout_2326_port, regs(2325) =>
                           DataPath_RF_bus_reg_dataout_2325_port, regs(2324) =>
                           DataPath_RF_bus_reg_dataout_2324_port, regs(2323) =>
                           DataPath_RF_bus_reg_dataout_2323_port, regs(2322) =>
                           DataPath_RF_bus_reg_dataout_2322_port, regs(2321) =>
                           DataPath_RF_bus_reg_dataout_2321_port, regs(2320) =>
                           DataPath_RF_bus_reg_dataout_2320_port, regs(2319) =>
                           DataPath_RF_bus_reg_dataout_2319_port, regs(2318) =>
                           DataPath_RF_bus_reg_dataout_2318_port, regs(2317) =>
                           DataPath_RF_bus_reg_dataout_2317_port, regs(2316) =>
                           DataPath_RF_bus_reg_dataout_2316_port, regs(2315) =>
                           DataPath_RF_bus_reg_dataout_2315_port, regs(2314) =>
                           DataPath_RF_bus_reg_dataout_2314_port, regs(2313) =>
                           DataPath_RF_bus_reg_dataout_2313_port, regs(2312) =>
                           DataPath_RF_bus_reg_dataout_2312_port, regs(2311) =>
                           DataPath_RF_bus_reg_dataout_2311_port, regs(2310) =>
                           DataPath_RF_bus_reg_dataout_2310_port, regs(2309) =>
                           DataPath_RF_bus_reg_dataout_2309_port, regs(2308) =>
                           DataPath_RF_bus_reg_dataout_2308_port, regs(2307) =>
                           DataPath_RF_bus_reg_dataout_2307_port, regs(2306) =>
                           DataPath_RF_bus_reg_dataout_2306_port, regs(2305) =>
                           DataPath_RF_bus_reg_dataout_2305_port, regs(2304) =>
                           DataPath_RF_bus_reg_dataout_2304_port, regs(2303) =>
                           DataPath_RF_bus_reg_dataout_2303_port, regs(2302) =>
                           DataPath_RF_bus_reg_dataout_2302_port, regs(2301) =>
                           DataPath_RF_bus_reg_dataout_2301_port, regs(2300) =>
                           DataPath_RF_bus_reg_dataout_2300_port, regs(2299) =>
                           DataPath_RF_bus_reg_dataout_2299_port, regs(2298) =>
                           DataPath_RF_bus_reg_dataout_2298_port, regs(2297) =>
                           DataPath_RF_bus_reg_dataout_2297_port, regs(2296) =>
                           DataPath_RF_bus_reg_dataout_2296_port, regs(2295) =>
                           DataPath_RF_bus_reg_dataout_2295_port, regs(2294) =>
                           DataPath_RF_bus_reg_dataout_2294_port, regs(2293) =>
                           DataPath_RF_bus_reg_dataout_2293_port, regs(2292) =>
                           DataPath_RF_bus_reg_dataout_2292_port, regs(2291) =>
                           DataPath_RF_bus_reg_dataout_2291_port, regs(2290) =>
                           DataPath_RF_bus_reg_dataout_2290_port, regs(2289) =>
                           DataPath_RF_bus_reg_dataout_2289_port, regs(2288) =>
                           DataPath_RF_bus_reg_dataout_2288_port, regs(2287) =>
                           DataPath_RF_bus_reg_dataout_2287_port, regs(2286) =>
                           DataPath_RF_bus_reg_dataout_2286_port, regs(2285) =>
                           DataPath_RF_bus_reg_dataout_2285_port, regs(2284) =>
                           DataPath_RF_bus_reg_dataout_2284_port, regs(2283) =>
                           DataPath_RF_bus_reg_dataout_2283_port, regs(2282) =>
                           DataPath_RF_bus_reg_dataout_2282_port, regs(2281) =>
                           DataPath_RF_bus_reg_dataout_2281_port, regs(2280) =>
                           DataPath_RF_bus_reg_dataout_2280_port, regs(2279) =>
                           DataPath_RF_bus_reg_dataout_2279_port, regs(2278) =>
                           DataPath_RF_bus_reg_dataout_2278_port, regs(2277) =>
                           DataPath_RF_bus_reg_dataout_2277_port, regs(2276) =>
                           DataPath_RF_bus_reg_dataout_2276_port, regs(2275) =>
                           DataPath_RF_bus_reg_dataout_2275_port, regs(2274) =>
                           DataPath_RF_bus_reg_dataout_2274_port, regs(2273) =>
                           DataPath_RF_bus_reg_dataout_2273_port, regs(2272) =>
                           DataPath_RF_bus_reg_dataout_2272_port, regs(2271) =>
                           DataPath_RF_bus_reg_dataout_2271_port, regs(2270) =>
                           DataPath_RF_bus_reg_dataout_2270_port, regs(2269) =>
                           DataPath_RF_bus_reg_dataout_2269_port, regs(2268) =>
                           DataPath_RF_bus_reg_dataout_2268_port, regs(2267) =>
                           DataPath_RF_bus_reg_dataout_2267_port, regs(2266) =>
                           DataPath_RF_bus_reg_dataout_2266_port, regs(2265) =>
                           DataPath_RF_bus_reg_dataout_2265_port, regs(2264) =>
                           DataPath_RF_bus_reg_dataout_2264_port, regs(2263) =>
                           DataPath_RF_bus_reg_dataout_2263_port, regs(2262) =>
                           DataPath_RF_bus_reg_dataout_2262_port, regs(2261) =>
                           DataPath_RF_bus_reg_dataout_2261_port, regs(2260) =>
                           DataPath_RF_bus_reg_dataout_2260_port, regs(2259) =>
                           DataPath_RF_bus_reg_dataout_2259_port, regs(2258) =>
                           DataPath_RF_bus_reg_dataout_2258_port, regs(2257) =>
                           DataPath_RF_bus_reg_dataout_2257_port, regs(2256) =>
                           DataPath_RF_bus_reg_dataout_2256_port, regs(2255) =>
                           DataPath_RF_bus_reg_dataout_2255_port, regs(2254) =>
                           DataPath_RF_bus_reg_dataout_2254_port, regs(2253) =>
                           DataPath_RF_bus_reg_dataout_2253_port, regs(2252) =>
                           DataPath_RF_bus_reg_dataout_2252_port, regs(2251) =>
                           DataPath_RF_bus_reg_dataout_2251_port, regs(2250) =>
                           DataPath_RF_bus_reg_dataout_2250_port, regs(2249) =>
                           DataPath_RF_bus_reg_dataout_2249_port, regs(2248) =>
                           DataPath_RF_bus_reg_dataout_2248_port, regs(2247) =>
                           DataPath_RF_bus_reg_dataout_2247_port, regs(2246) =>
                           DataPath_RF_bus_reg_dataout_2246_port, regs(2245) =>
                           DataPath_RF_bus_reg_dataout_2245_port, regs(2244) =>
                           DataPath_RF_bus_reg_dataout_2244_port, regs(2243) =>
                           DataPath_RF_bus_reg_dataout_2243_port, regs(2242) =>
                           DataPath_RF_bus_reg_dataout_2242_port, regs(2241) =>
                           DataPath_RF_bus_reg_dataout_2241_port, regs(2240) =>
                           DataPath_RF_bus_reg_dataout_2240_port, regs(2239) =>
                           DataPath_RF_bus_reg_dataout_2239_port, regs(2238) =>
                           DataPath_RF_bus_reg_dataout_2238_port, regs(2237) =>
                           DataPath_RF_bus_reg_dataout_2237_port, regs(2236) =>
                           DataPath_RF_bus_reg_dataout_2236_port, regs(2235) =>
                           DataPath_RF_bus_reg_dataout_2235_port, regs(2234) =>
                           DataPath_RF_bus_reg_dataout_2234_port, regs(2233) =>
                           DataPath_RF_bus_reg_dataout_2233_port, regs(2232) =>
                           DataPath_RF_bus_reg_dataout_2232_port, regs(2231) =>
                           DataPath_RF_bus_reg_dataout_2231_port, regs(2230) =>
                           DataPath_RF_bus_reg_dataout_2230_port, regs(2229) =>
                           DataPath_RF_bus_reg_dataout_2229_port, regs(2228) =>
                           DataPath_RF_bus_reg_dataout_2228_port, regs(2227) =>
                           DataPath_RF_bus_reg_dataout_2227_port, regs(2226) =>
                           DataPath_RF_bus_reg_dataout_2226_port, regs(2225) =>
                           DataPath_RF_bus_reg_dataout_2225_port, regs(2224) =>
                           DataPath_RF_bus_reg_dataout_2224_port, regs(2223) =>
                           DataPath_RF_bus_reg_dataout_2223_port, regs(2222) =>
                           DataPath_RF_bus_reg_dataout_2222_port, regs(2221) =>
                           DataPath_RF_bus_reg_dataout_2221_port, regs(2220) =>
                           DataPath_RF_bus_reg_dataout_2220_port, regs(2219) =>
                           DataPath_RF_bus_reg_dataout_2219_port, regs(2218) =>
                           DataPath_RF_bus_reg_dataout_2218_port, regs(2217) =>
                           DataPath_RF_bus_reg_dataout_2217_port, regs(2216) =>
                           DataPath_RF_bus_reg_dataout_2216_port, regs(2215) =>
                           DataPath_RF_bus_reg_dataout_2215_port, regs(2214) =>
                           DataPath_RF_bus_reg_dataout_2214_port, regs(2213) =>
                           DataPath_RF_bus_reg_dataout_2213_port, regs(2212) =>
                           DataPath_RF_bus_reg_dataout_2212_port, regs(2211) =>
                           DataPath_RF_bus_reg_dataout_2211_port, regs(2210) =>
                           DataPath_RF_bus_reg_dataout_2210_port, regs(2209) =>
                           DataPath_RF_bus_reg_dataout_2209_port, regs(2208) =>
                           DataPath_RF_bus_reg_dataout_2208_port, regs(2207) =>
                           DataPath_RF_bus_reg_dataout_2207_port, regs(2206) =>
                           DataPath_RF_bus_reg_dataout_2206_port, regs(2205) =>
                           DataPath_RF_bus_reg_dataout_2205_port, regs(2204) =>
                           DataPath_RF_bus_reg_dataout_2204_port, regs(2203) =>
                           DataPath_RF_bus_reg_dataout_2203_port, regs(2202) =>
                           DataPath_RF_bus_reg_dataout_2202_port, regs(2201) =>
                           DataPath_RF_bus_reg_dataout_2201_port, regs(2200) =>
                           DataPath_RF_bus_reg_dataout_2200_port, regs(2199) =>
                           DataPath_RF_bus_reg_dataout_2199_port, regs(2198) =>
                           DataPath_RF_bus_reg_dataout_2198_port, regs(2197) =>
                           DataPath_RF_bus_reg_dataout_2197_port, regs(2196) =>
                           DataPath_RF_bus_reg_dataout_2196_port, regs(2195) =>
                           DataPath_RF_bus_reg_dataout_2195_port, regs(2194) =>
                           DataPath_RF_bus_reg_dataout_2194_port, regs(2193) =>
                           DataPath_RF_bus_reg_dataout_2193_port, regs(2192) =>
                           DataPath_RF_bus_reg_dataout_2192_port, regs(2191) =>
                           DataPath_RF_bus_reg_dataout_2191_port, regs(2190) =>
                           DataPath_RF_bus_reg_dataout_2190_port, regs(2189) =>
                           DataPath_RF_bus_reg_dataout_2189_port, regs(2188) =>
                           DataPath_RF_bus_reg_dataout_2188_port, regs(2187) =>
                           DataPath_RF_bus_reg_dataout_2187_port, regs(2186) =>
                           DataPath_RF_bus_reg_dataout_2186_port, regs(2185) =>
                           DataPath_RF_bus_reg_dataout_2185_port, regs(2184) =>
                           DataPath_RF_bus_reg_dataout_2184_port, regs(2183) =>
                           DataPath_RF_bus_reg_dataout_2183_port, regs(2182) =>
                           DataPath_RF_bus_reg_dataout_2182_port, regs(2181) =>
                           DataPath_RF_bus_reg_dataout_2181_port, regs(2180) =>
                           DataPath_RF_bus_reg_dataout_2180_port, regs(2179) =>
                           DataPath_RF_bus_reg_dataout_2179_port, regs(2178) =>
                           DataPath_RF_bus_reg_dataout_2178_port, regs(2177) =>
                           DataPath_RF_bus_reg_dataout_2177_port, regs(2176) =>
                           DataPath_RF_bus_reg_dataout_2176_port, regs(2175) =>
                           DataPath_RF_bus_reg_dataout_2175_port, regs(2174) =>
                           DataPath_RF_bus_reg_dataout_2174_port, regs(2173) =>
                           DataPath_RF_bus_reg_dataout_2173_port, regs(2172) =>
                           DataPath_RF_bus_reg_dataout_2172_port, regs(2171) =>
                           DataPath_RF_bus_reg_dataout_2171_port, regs(2170) =>
                           DataPath_RF_bus_reg_dataout_2170_port, regs(2169) =>
                           DataPath_RF_bus_reg_dataout_2169_port, regs(2168) =>
                           DataPath_RF_bus_reg_dataout_2168_port, regs(2167) =>
                           DataPath_RF_bus_reg_dataout_2167_port, regs(2166) =>
                           DataPath_RF_bus_reg_dataout_2166_port, regs(2165) =>
                           DataPath_RF_bus_reg_dataout_2165_port, regs(2164) =>
                           DataPath_RF_bus_reg_dataout_2164_port, regs(2163) =>
                           DataPath_RF_bus_reg_dataout_2163_port, regs(2162) =>
                           DataPath_RF_bus_reg_dataout_2162_port, regs(2161) =>
                           DataPath_RF_bus_reg_dataout_2161_port, regs(2160) =>
                           DataPath_RF_bus_reg_dataout_2160_port, regs(2159) =>
                           DataPath_RF_bus_reg_dataout_2159_port, regs(2158) =>
                           DataPath_RF_bus_reg_dataout_2158_port, regs(2157) =>
                           DataPath_RF_bus_reg_dataout_2157_port, regs(2156) =>
                           DataPath_RF_bus_reg_dataout_2156_port, regs(2155) =>
                           DataPath_RF_bus_reg_dataout_2155_port, regs(2154) =>
                           DataPath_RF_bus_reg_dataout_2154_port, regs(2153) =>
                           DataPath_RF_bus_reg_dataout_2153_port, regs(2152) =>
                           DataPath_RF_bus_reg_dataout_2152_port, regs(2151) =>
                           DataPath_RF_bus_reg_dataout_2151_port, regs(2150) =>
                           DataPath_RF_bus_reg_dataout_2150_port, regs(2149) =>
                           DataPath_RF_bus_reg_dataout_2149_port, regs(2148) =>
                           DataPath_RF_bus_reg_dataout_2148_port, regs(2147) =>
                           DataPath_RF_bus_reg_dataout_2147_port, regs(2146) =>
                           DataPath_RF_bus_reg_dataout_2146_port, regs(2145) =>
                           DataPath_RF_bus_reg_dataout_2145_port, regs(2144) =>
                           DataPath_RF_bus_reg_dataout_2144_port, regs(2143) =>
                           DataPath_RF_bus_reg_dataout_2143_port, regs(2142) =>
                           DataPath_RF_bus_reg_dataout_2142_port, regs(2141) =>
                           DataPath_RF_bus_reg_dataout_2141_port, regs(2140) =>
                           DataPath_RF_bus_reg_dataout_2140_port, regs(2139) =>
                           DataPath_RF_bus_reg_dataout_2139_port, regs(2138) =>
                           DataPath_RF_bus_reg_dataout_2138_port, regs(2137) =>
                           DataPath_RF_bus_reg_dataout_2137_port, regs(2136) =>
                           DataPath_RF_bus_reg_dataout_2136_port, regs(2135) =>
                           DataPath_RF_bus_reg_dataout_2135_port, regs(2134) =>
                           DataPath_RF_bus_reg_dataout_2134_port, regs(2133) =>
                           DataPath_RF_bus_reg_dataout_2133_port, regs(2132) =>
                           DataPath_RF_bus_reg_dataout_2132_port, regs(2131) =>
                           DataPath_RF_bus_reg_dataout_2131_port, regs(2130) =>
                           DataPath_RF_bus_reg_dataout_2130_port, regs(2129) =>
                           DataPath_RF_bus_reg_dataout_2129_port, regs(2128) =>
                           DataPath_RF_bus_reg_dataout_2128_port, regs(2127) =>
                           DataPath_RF_bus_reg_dataout_2127_port, regs(2126) =>
                           DataPath_RF_bus_reg_dataout_2126_port, regs(2125) =>
                           DataPath_RF_bus_reg_dataout_2125_port, regs(2124) =>
                           DataPath_RF_bus_reg_dataout_2124_port, regs(2123) =>
                           DataPath_RF_bus_reg_dataout_2123_port, regs(2122) =>
                           DataPath_RF_bus_reg_dataout_2122_port, regs(2121) =>
                           DataPath_RF_bus_reg_dataout_2121_port, regs(2120) =>
                           DataPath_RF_bus_reg_dataout_2120_port, regs(2119) =>
                           DataPath_RF_bus_reg_dataout_2119_port, regs(2118) =>
                           DataPath_RF_bus_reg_dataout_2118_port, regs(2117) =>
                           DataPath_RF_bus_reg_dataout_2117_port, regs(2116) =>
                           DataPath_RF_bus_reg_dataout_2116_port, regs(2115) =>
                           DataPath_RF_bus_reg_dataout_2115_port, regs(2114) =>
                           DataPath_RF_bus_reg_dataout_2114_port, regs(2113) =>
                           DataPath_RF_bus_reg_dataout_2113_port, regs(2112) =>
                           DataPath_RF_bus_reg_dataout_2112_port, regs(2111) =>
                           DataPath_RF_bus_reg_dataout_2111_port, regs(2110) =>
                           DataPath_RF_bus_reg_dataout_2110_port, regs(2109) =>
                           DataPath_RF_bus_reg_dataout_2109_port, regs(2108) =>
                           DataPath_RF_bus_reg_dataout_2108_port, regs(2107) =>
                           DataPath_RF_bus_reg_dataout_2107_port, regs(2106) =>
                           DataPath_RF_bus_reg_dataout_2106_port, regs(2105) =>
                           DataPath_RF_bus_reg_dataout_2105_port, regs(2104) =>
                           DataPath_RF_bus_reg_dataout_2104_port, regs(2103) =>
                           DataPath_RF_bus_reg_dataout_2103_port, regs(2102) =>
                           DataPath_RF_bus_reg_dataout_2102_port, regs(2101) =>
                           DataPath_RF_bus_reg_dataout_2101_port, regs(2100) =>
                           DataPath_RF_bus_reg_dataout_2100_port, regs(2099) =>
                           DataPath_RF_bus_reg_dataout_2099_port, regs(2098) =>
                           DataPath_RF_bus_reg_dataout_2098_port, regs(2097) =>
                           DataPath_RF_bus_reg_dataout_2097_port, regs(2096) =>
                           DataPath_RF_bus_reg_dataout_2096_port, regs(2095) =>
                           DataPath_RF_bus_reg_dataout_2095_port, regs(2094) =>
                           DataPath_RF_bus_reg_dataout_2094_port, regs(2093) =>
                           DataPath_RF_bus_reg_dataout_2093_port, regs(2092) =>
                           DataPath_RF_bus_reg_dataout_2092_port, regs(2091) =>
                           DataPath_RF_bus_reg_dataout_2091_port, regs(2090) =>
                           DataPath_RF_bus_reg_dataout_2090_port, regs(2089) =>
                           DataPath_RF_bus_reg_dataout_2089_port, regs(2088) =>
                           DataPath_RF_bus_reg_dataout_2088_port, regs(2087) =>
                           DataPath_RF_bus_reg_dataout_2087_port, regs(2086) =>
                           DataPath_RF_bus_reg_dataout_2086_port, regs(2085) =>
                           DataPath_RF_bus_reg_dataout_2085_port, regs(2084) =>
                           DataPath_RF_bus_reg_dataout_2084_port, regs(2083) =>
                           DataPath_RF_bus_reg_dataout_2083_port, regs(2082) =>
                           DataPath_RF_bus_reg_dataout_2082_port, regs(2081) =>
                           DataPath_RF_bus_reg_dataout_2081_port, regs(2080) =>
                           DataPath_RF_bus_reg_dataout_2080_port, regs(2079) =>
                           DataPath_RF_bus_reg_dataout_2079_port, regs(2078) =>
                           DataPath_RF_bus_reg_dataout_2078_port, regs(2077) =>
                           DataPath_RF_bus_reg_dataout_2077_port, regs(2076) =>
                           DataPath_RF_bus_reg_dataout_2076_port, regs(2075) =>
                           DataPath_RF_bus_reg_dataout_2075_port, regs(2074) =>
                           DataPath_RF_bus_reg_dataout_2074_port, regs(2073) =>
                           DataPath_RF_bus_reg_dataout_2073_port, regs(2072) =>
                           DataPath_RF_bus_reg_dataout_2072_port, regs(2071) =>
                           DataPath_RF_bus_reg_dataout_2071_port, regs(2070) =>
                           DataPath_RF_bus_reg_dataout_2070_port, regs(2069) =>
                           DataPath_RF_bus_reg_dataout_2069_port, regs(2068) =>
                           DataPath_RF_bus_reg_dataout_2068_port, regs(2067) =>
                           DataPath_RF_bus_reg_dataout_2067_port, regs(2066) =>
                           DataPath_RF_bus_reg_dataout_2066_port, regs(2065) =>
                           DataPath_RF_bus_reg_dataout_2065_port, regs(2064) =>
                           DataPath_RF_bus_reg_dataout_2064_port, regs(2063) =>
                           DataPath_RF_bus_reg_dataout_2063_port, regs(2062) =>
                           DataPath_RF_bus_reg_dataout_2062_port, regs(2061) =>
                           DataPath_RF_bus_reg_dataout_2061_port, regs(2060) =>
                           DataPath_RF_bus_reg_dataout_2060_port, regs(2059) =>
                           DataPath_RF_bus_reg_dataout_2059_port, regs(2058) =>
                           DataPath_RF_bus_reg_dataout_2058_port, regs(2057) =>
                           DataPath_RF_bus_reg_dataout_2057_port, regs(2056) =>
                           DataPath_RF_bus_reg_dataout_2056_port, regs(2055) =>
                           DataPath_RF_bus_reg_dataout_2055_port, regs(2054) =>
                           DataPath_RF_bus_reg_dataout_2054_port, regs(2053) =>
                           DataPath_RF_bus_reg_dataout_2053_port, regs(2052) =>
                           DataPath_RF_bus_reg_dataout_2052_port, regs(2051) =>
                           DataPath_RF_bus_reg_dataout_2051_port, regs(2050) =>
                           DataPath_RF_bus_reg_dataout_2050_port, regs(2049) =>
                           DataPath_RF_bus_reg_dataout_2049_port, regs(2048) =>
                           DataPath_RF_bus_reg_dataout_2048_port, regs(2047) =>
                           DataPath_RF_bus_reg_dataout_2047_port, regs(2046) =>
                           DataPath_RF_bus_reg_dataout_2046_port, regs(2045) =>
                           DataPath_RF_bus_reg_dataout_2045_port, regs(2044) =>
                           DataPath_RF_bus_reg_dataout_2044_port, regs(2043) =>
                           DataPath_RF_bus_reg_dataout_2043_port, regs(2042) =>
                           DataPath_RF_bus_reg_dataout_2042_port, regs(2041) =>
                           DataPath_RF_bus_reg_dataout_2041_port, regs(2040) =>
                           DataPath_RF_bus_reg_dataout_2040_port, regs(2039) =>
                           DataPath_RF_bus_reg_dataout_2039_port, regs(2038) =>
                           DataPath_RF_bus_reg_dataout_2038_port, regs(2037) =>
                           DataPath_RF_bus_reg_dataout_2037_port, regs(2036) =>
                           DataPath_RF_bus_reg_dataout_2036_port, regs(2035) =>
                           DataPath_RF_bus_reg_dataout_2035_port, regs(2034) =>
                           DataPath_RF_bus_reg_dataout_2034_port, regs(2033) =>
                           DataPath_RF_bus_reg_dataout_2033_port, regs(2032) =>
                           DataPath_RF_bus_reg_dataout_2032_port, regs(2031) =>
                           DataPath_RF_bus_reg_dataout_2031_port, regs(2030) =>
                           DataPath_RF_bus_reg_dataout_2030_port, regs(2029) =>
                           DataPath_RF_bus_reg_dataout_2029_port, regs(2028) =>
                           DataPath_RF_bus_reg_dataout_2028_port, regs(2027) =>
                           DataPath_RF_bus_reg_dataout_2027_port, regs(2026) =>
                           DataPath_RF_bus_reg_dataout_2026_port, regs(2025) =>
                           DataPath_RF_bus_reg_dataout_2025_port, regs(2024) =>
                           DataPath_RF_bus_reg_dataout_2024_port, regs(2023) =>
                           DataPath_RF_bus_reg_dataout_2023_port, regs(2022) =>
                           DataPath_RF_bus_reg_dataout_2022_port, regs(2021) =>
                           DataPath_RF_bus_reg_dataout_2021_port, regs(2020) =>
                           DataPath_RF_bus_reg_dataout_2020_port, regs(2019) =>
                           DataPath_RF_bus_reg_dataout_2019_port, regs(2018) =>
                           DataPath_RF_bus_reg_dataout_2018_port, regs(2017) =>
                           DataPath_RF_bus_reg_dataout_2017_port, regs(2016) =>
                           DataPath_RF_bus_reg_dataout_2016_port, regs(2015) =>
                           DataPath_RF_bus_reg_dataout_2015_port, regs(2014) =>
                           DataPath_RF_bus_reg_dataout_2014_port, regs(2013) =>
                           DataPath_RF_bus_reg_dataout_2013_port, regs(2012) =>
                           DataPath_RF_bus_reg_dataout_2012_port, regs(2011) =>
                           DataPath_RF_bus_reg_dataout_2011_port, regs(2010) =>
                           DataPath_RF_bus_reg_dataout_2010_port, regs(2009) =>
                           DataPath_RF_bus_reg_dataout_2009_port, regs(2008) =>
                           DataPath_RF_bus_reg_dataout_2008_port, regs(2007) =>
                           DataPath_RF_bus_reg_dataout_2007_port, regs(2006) =>
                           DataPath_RF_bus_reg_dataout_2006_port, regs(2005) =>
                           DataPath_RF_bus_reg_dataout_2005_port, regs(2004) =>
                           DataPath_RF_bus_reg_dataout_2004_port, regs(2003) =>
                           DataPath_RF_bus_reg_dataout_2003_port, regs(2002) =>
                           DataPath_RF_bus_reg_dataout_2002_port, regs(2001) =>
                           DataPath_RF_bus_reg_dataout_2001_port, regs(2000) =>
                           DataPath_RF_bus_reg_dataout_2000_port, regs(1999) =>
                           DataPath_RF_bus_reg_dataout_1999_port, regs(1998) =>
                           DataPath_RF_bus_reg_dataout_1998_port, regs(1997) =>
                           DataPath_RF_bus_reg_dataout_1997_port, regs(1996) =>
                           DataPath_RF_bus_reg_dataout_1996_port, regs(1995) =>
                           DataPath_RF_bus_reg_dataout_1995_port, regs(1994) =>
                           DataPath_RF_bus_reg_dataout_1994_port, regs(1993) =>
                           DataPath_RF_bus_reg_dataout_1993_port, regs(1992) =>
                           DataPath_RF_bus_reg_dataout_1992_port, regs(1991) =>
                           DataPath_RF_bus_reg_dataout_1991_port, regs(1990) =>
                           DataPath_RF_bus_reg_dataout_1990_port, regs(1989) =>
                           DataPath_RF_bus_reg_dataout_1989_port, regs(1988) =>
                           DataPath_RF_bus_reg_dataout_1988_port, regs(1987) =>
                           DataPath_RF_bus_reg_dataout_1987_port, regs(1986) =>
                           DataPath_RF_bus_reg_dataout_1986_port, regs(1985) =>
                           DataPath_RF_bus_reg_dataout_1985_port, regs(1984) =>
                           DataPath_RF_bus_reg_dataout_1984_port, regs(1983) =>
                           DataPath_RF_bus_reg_dataout_1983_port, regs(1982) =>
                           DataPath_RF_bus_reg_dataout_1982_port, regs(1981) =>
                           DataPath_RF_bus_reg_dataout_1981_port, regs(1980) =>
                           DataPath_RF_bus_reg_dataout_1980_port, regs(1979) =>
                           DataPath_RF_bus_reg_dataout_1979_port, regs(1978) =>
                           DataPath_RF_bus_reg_dataout_1978_port, regs(1977) =>
                           DataPath_RF_bus_reg_dataout_1977_port, regs(1976) =>
                           DataPath_RF_bus_reg_dataout_1976_port, regs(1975) =>
                           DataPath_RF_bus_reg_dataout_1975_port, regs(1974) =>
                           DataPath_RF_bus_reg_dataout_1974_port, regs(1973) =>
                           DataPath_RF_bus_reg_dataout_1973_port, regs(1972) =>
                           DataPath_RF_bus_reg_dataout_1972_port, regs(1971) =>
                           DataPath_RF_bus_reg_dataout_1971_port, regs(1970) =>
                           DataPath_RF_bus_reg_dataout_1970_port, regs(1969) =>
                           DataPath_RF_bus_reg_dataout_1969_port, regs(1968) =>
                           DataPath_RF_bus_reg_dataout_1968_port, regs(1967) =>
                           DataPath_RF_bus_reg_dataout_1967_port, regs(1966) =>
                           DataPath_RF_bus_reg_dataout_1966_port, regs(1965) =>
                           DataPath_RF_bus_reg_dataout_1965_port, regs(1964) =>
                           DataPath_RF_bus_reg_dataout_1964_port, regs(1963) =>
                           DataPath_RF_bus_reg_dataout_1963_port, regs(1962) =>
                           DataPath_RF_bus_reg_dataout_1962_port, regs(1961) =>
                           DataPath_RF_bus_reg_dataout_1961_port, regs(1960) =>
                           DataPath_RF_bus_reg_dataout_1960_port, regs(1959) =>
                           DataPath_RF_bus_reg_dataout_1959_port, regs(1958) =>
                           DataPath_RF_bus_reg_dataout_1958_port, regs(1957) =>
                           DataPath_RF_bus_reg_dataout_1957_port, regs(1956) =>
                           DataPath_RF_bus_reg_dataout_1956_port, regs(1955) =>
                           DataPath_RF_bus_reg_dataout_1955_port, regs(1954) =>
                           DataPath_RF_bus_reg_dataout_1954_port, regs(1953) =>
                           DataPath_RF_bus_reg_dataout_1953_port, regs(1952) =>
                           DataPath_RF_bus_reg_dataout_1952_port, regs(1951) =>
                           DataPath_RF_bus_reg_dataout_1951_port, regs(1950) =>
                           DataPath_RF_bus_reg_dataout_1950_port, regs(1949) =>
                           DataPath_RF_bus_reg_dataout_1949_port, regs(1948) =>
                           DataPath_RF_bus_reg_dataout_1948_port, regs(1947) =>
                           DataPath_RF_bus_reg_dataout_1947_port, regs(1946) =>
                           DataPath_RF_bus_reg_dataout_1946_port, regs(1945) =>
                           DataPath_RF_bus_reg_dataout_1945_port, regs(1944) =>
                           DataPath_RF_bus_reg_dataout_1944_port, regs(1943) =>
                           DataPath_RF_bus_reg_dataout_1943_port, regs(1942) =>
                           DataPath_RF_bus_reg_dataout_1942_port, regs(1941) =>
                           DataPath_RF_bus_reg_dataout_1941_port, regs(1940) =>
                           DataPath_RF_bus_reg_dataout_1940_port, regs(1939) =>
                           DataPath_RF_bus_reg_dataout_1939_port, regs(1938) =>
                           DataPath_RF_bus_reg_dataout_1938_port, regs(1937) =>
                           DataPath_RF_bus_reg_dataout_1937_port, regs(1936) =>
                           DataPath_RF_bus_reg_dataout_1936_port, regs(1935) =>
                           DataPath_RF_bus_reg_dataout_1935_port, regs(1934) =>
                           DataPath_RF_bus_reg_dataout_1934_port, regs(1933) =>
                           DataPath_RF_bus_reg_dataout_1933_port, regs(1932) =>
                           DataPath_RF_bus_reg_dataout_1932_port, regs(1931) =>
                           DataPath_RF_bus_reg_dataout_1931_port, regs(1930) =>
                           DataPath_RF_bus_reg_dataout_1930_port, regs(1929) =>
                           DataPath_RF_bus_reg_dataout_1929_port, regs(1928) =>
                           DataPath_RF_bus_reg_dataout_1928_port, regs(1927) =>
                           DataPath_RF_bus_reg_dataout_1927_port, regs(1926) =>
                           DataPath_RF_bus_reg_dataout_1926_port, regs(1925) =>
                           DataPath_RF_bus_reg_dataout_1925_port, regs(1924) =>
                           DataPath_RF_bus_reg_dataout_1924_port, regs(1923) =>
                           DataPath_RF_bus_reg_dataout_1923_port, regs(1922) =>
                           DataPath_RF_bus_reg_dataout_1922_port, regs(1921) =>
                           DataPath_RF_bus_reg_dataout_1921_port, regs(1920) =>
                           DataPath_RF_bus_reg_dataout_1920_port, regs(1919) =>
                           DataPath_RF_bus_reg_dataout_1919_port, regs(1918) =>
                           DataPath_RF_bus_reg_dataout_1918_port, regs(1917) =>
                           DataPath_RF_bus_reg_dataout_1917_port, regs(1916) =>
                           DataPath_RF_bus_reg_dataout_1916_port, regs(1915) =>
                           DataPath_RF_bus_reg_dataout_1915_port, regs(1914) =>
                           DataPath_RF_bus_reg_dataout_1914_port, regs(1913) =>
                           DataPath_RF_bus_reg_dataout_1913_port, regs(1912) =>
                           DataPath_RF_bus_reg_dataout_1912_port, regs(1911) =>
                           DataPath_RF_bus_reg_dataout_1911_port, regs(1910) =>
                           DataPath_RF_bus_reg_dataout_1910_port, regs(1909) =>
                           DataPath_RF_bus_reg_dataout_1909_port, regs(1908) =>
                           DataPath_RF_bus_reg_dataout_1908_port, regs(1907) =>
                           DataPath_RF_bus_reg_dataout_1907_port, regs(1906) =>
                           DataPath_RF_bus_reg_dataout_1906_port, regs(1905) =>
                           DataPath_RF_bus_reg_dataout_1905_port, regs(1904) =>
                           DataPath_RF_bus_reg_dataout_1904_port, regs(1903) =>
                           DataPath_RF_bus_reg_dataout_1903_port, regs(1902) =>
                           DataPath_RF_bus_reg_dataout_1902_port, regs(1901) =>
                           DataPath_RF_bus_reg_dataout_1901_port, regs(1900) =>
                           DataPath_RF_bus_reg_dataout_1900_port, regs(1899) =>
                           DataPath_RF_bus_reg_dataout_1899_port, regs(1898) =>
                           DataPath_RF_bus_reg_dataout_1898_port, regs(1897) =>
                           DataPath_RF_bus_reg_dataout_1897_port, regs(1896) =>
                           DataPath_RF_bus_reg_dataout_1896_port, regs(1895) =>
                           DataPath_RF_bus_reg_dataout_1895_port, regs(1894) =>
                           DataPath_RF_bus_reg_dataout_1894_port, regs(1893) =>
                           DataPath_RF_bus_reg_dataout_1893_port, regs(1892) =>
                           DataPath_RF_bus_reg_dataout_1892_port, regs(1891) =>
                           DataPath_RF_bus_reg_dataout_1891_port, regs(1890) =>
                           DataPath_RF_bus_reg_dataout_1890_port, regs(1889) =>
                           DataPath_RF_bus_reg_dataout_1889_port, regs(1888) =>
                           DataPath_RF_bus_reg_dataout_1888_port, regs(1887) =>
                           DataPath_RF_bus_reg_dataout_1887_port, regs(1886) =>
                           DataPath_RF_bus_reg_dataout_1886_port, regs(1885) =>
                           DataPath_RF_bus_reg_dataout_1885_port, regs(1884) =>
                           DataPath_RF_bus_reg_dataout_1884_port, regs(1883) =>
                           DataPath_RF_bus_reg_dataout_1883_port, regs(1882) =>
                           DataPath_RF_bus_reg_dataout_1882_port, regs(1881) =>
                           DataPath_RF_bus_reg_dataout_1881_port, regs(1880) =>
                           DataPath_RF_bus_reg_dataout_1880_port, regs(1879) =>
                           DataPath_RF_bus_reg_dataout_1879_port, regs(1878) =>
                           DataPath_RF_bus_reg_dataout_1878_port, regs(1877) =>
                           DataPath_RF_bus_reg_dataout_1877_port, regs(1876) =>
                           DataPath_RF_bus_reg_dataout_1876_port, regs(1875) =>
                           DataPath_RF_bus_reg_dataout_1875_port, regs(1874) =>
                           DataPath_RF_bus_reg_dataout_1874_port, regs(1873) =>
                           DataPath_RF_bus_reg_dataout_1873_port, regs(1872) =>
                           DataPath_RF_bus_reg_dataout_1872_port, regs(1871) =>
                           DataPath_RF_bus_reg_dataout_1871_port, regs(1870) =>
                           DataPath_RF_bus_reg_dataout_1870_port, regs(1869) =>
                           DataPath_RF_bus_reg_dataout_1869_port, regs(1868) =>
                           DataPath_RF_bus_reg_dataout_1868_port, regs(1867) =>
                           DataPath_RF_bus_reg_dataout_1867_port, regs(1866) =>
                           DataPath_RF_bus_reg_dataout_1866_port, regs(1865) =>
                           DataPath_RF_bus_reg_dataout_1865_port, regs(1864) =>
                           DataPath_RF_bus_reg_dataout_1864_port, regs(1863) =>
                           DataPath_RF_bus_reg_dataout_1863_port, regs(1862) =>
                           DataPath_RF_bus_reg_dataout_1862_port, regs(1861) =>
                           DataPath_RF_bus_reg_dataout_1861_port, regs(1860) =>
                           DataPath_RF_bus_reg_dataout_1860_port, regs(1859) =>
                           DataPath_RF_bus_reg_dataout_1859_port, regs(1858) =>
                           DataPath_RF_bus_reg_dataout_1858_port, regs(1857) =>
                           DataPath_RF_bus_reg_dataout_1857_port, regs(1856) =>
                           DataPath_RF_bus_reg_dataout_1856_port, regs(1855) =>
                           DataPath_RF_bus_reg_dataout_1855_port, regs(1854) =>
                           DataPath_RF_bus_reg_dataout_1854_port, regs(1853) =>
                           DataPath_RF_bus_reg_dataout_1853_port, regs(1852) =>
                           DataPath_RF_bus_reg_dataout_1852_port, regs(1851) =>
                           DataPath_RF_bus_reg_dataout_1851_port, regs(1850) =>
                           DataPath_RF_bus_reg_dataout_1850_port, regs(1849) =>
                           DataPath_RF_bus_reg_dataout_1849_port, regs(1848) =>
                           DataPath_RF_bus_reg_dataout_1848_port, regs(1847) =>
                           DataPath_RF_bus_reg_dataout_1847_port, regs(1846) =>
                           DataPath_RF_bus_reg_dataout_1846_port, regs(1845) =>
                           DataPath_RF_bus_reg_dataout_1845_port, regs(1844) =>
                           DataPath_RF_bus_reg_dataout_1844_port, regs(1843) =>
                           DataPath_RF_bus_reg_dataout_1843_port, regs(1842) =>
                           DataPath_RF_bus_reg_dataout_1842_port, regs(1841) =>
                           DataPath_RF_bus_reg_dataout_1841_port, regs(1840) =>
                           DataPath_RF_bus_reg_dataout_1840_port, regs(1839) =>
                           DataPath_RF_bus_reg_dataout_1839_port, regs(1838) =>
                           DataPath_RF_bus_reg_dataout_1838_port, regs(1837) =>
                           DataPath_RF_bus_reg_dataout_1837_port, regs(1836) =>
                           DataPath_RF_bus_reg_dataout_1836_port, regs(1835) =>
                           DataPath_RF_bus_reg_dataout_1835_port, regs(1834) =>
                           DataPath_RF_bus_reg_dataout_1834_port, regs(1833) =>
                           DataPath_RF_bus_reg_dataout_1833_port, regs(1832) =>
                           DataPath_RF_bus_reg_dataout_1832_port, regs(1831) =>
                           DataPath_RF_bus_reg_dataout_1831_port, regs(1830) =>
                           DataPath_RF_bus_reg_dataout_1830_port, regs(1829) =>
                           DataPath_RF_bus_reg_dataout_1829_port, regs(1828) =>
                           DataPath_RF_bus_reg_dataout_1828_port, regs(1827) =>
                           DataPath_RF_bus_reg_dataout_1827_port, regs(1826) =>
                           DataPath_RF_bus_reg_dataout_1826_port, regs(1825) =>
                           DataPath_RF_bus_reg_dataout_1825_port, regs(1824) =>
                           DataPath_RF_bus_reg_dataout_1824_port, regs(1823) =>
                           DataPath_RF_bus_reg_dataout_1823_port, regs(1822) =>
                           DataPath_RF_bus_reg_dataout_1822_port, regs(1821) =>
                           DataPath_RF_bus_reg_dataout_1821_port, regs(1820) =>
                           DataPath_RF_bus_reg_dataout_1820_port, regs(1819) =>
                           DataPath_RF_bus_reg_dataout_1819_port, regs(1818) =>
                           DataPath_RF_bus_reg_dataout_1818_port, regs(1817) =>
                           DataPath_RF_bus_reg_dataout_1817_port, regs(1816) =>
                           DataPath_RF_bus_reg_dataout_1816_port, regs(1815) =>
                           DataPath_RF_bus_reg_dataout_1815_port, regs(1814) =>
                           DataPath_RF_bus_reg_dataout_1814_port, regs(1813) =>
                           DataPath_RF_bus_reg_dataout_1813_port, regs(1812) =>
                           DataPath_RF_bus_reg_dataout_1812_port, regs(1811) =>
                           DataPath_RF_bus_reg_dataout_1811_port, regs(1810) =>
                           DataPath_RF_bus_reg_dataout_1810_port, regs(1809) =>
                           DataPath_RF_bus_reg_dataout_1809_port, regs(1808) =>
                           DataPath_RF_bus_reg_dataout_1808_port, regs(1807) =>
                           DataPath_RF_bus_reg_dataout_1807_port, regs(1806) =>
                           DataPath_RF_bus_reg_dataout_1806_port, regs(1805) =>
                           DataPath_RF_bus_reg_dataout_1805_port, regs(1804) =>
                           DataPath_RF_bus_reg_dataout_1804_port, regs(1803) =>
                           DataPath_RF_bus_reg_dataout_1803_port, regs(1802) =>
                           DataPath_RF_bus_reg_dataout_1802_port, regs(1801) =>
                           DataPath_RF_bus_reg_dataout_1801_port, regs(1800) =>
                           DataPath_RF_bus_reg_dataout_1800_port, regs(1799) =>
                           DataPath_RF_bus_reg_dataout_1799_port, regs(1798) =>
                           DataPath_RF_bus_reg_dataout_1798_port, regs(1797) =>
                           DataPath_RF_bus_reg_dataout_1797_port, regs(1796) =>
                           DataPath_RF_bus_reg_dataout_1796_port, regs(1795) =>
                           DataPath_RF_bus_reg_dataout_1795_port, regs(1794) =>
                           DataPath_RF_bus_reg_dataout_1794_port, regs(1793) =>
                           DataPath_RF_bus_reg_dataout_1793_port, regs(1792) =>
                           DataPath_RF_bus_reg_dataout_1792_port, regs(1791) =>
                           DataPath_RF_bus_reg_dataout_1791_port, regs(1790) =>
                           DataPath_RF_bus_reg_dataout_1790_port, regs(1789) =>
                           DataPath_RF_bus_reg_dataout_1789_port, regs(1788) =>
                           DataPath_RF_bus_reg_dataout_1788_port, regs(1787) =>
                           DataPath_RF_bus_reg_dataout_1787_port, regs(1786) =>
                           DataPath_RF_bus_reg_dataout_1786_port, regs(1785) =>
                           DataPath_RF_bus_reg_dataout_1785_port, regs(1784) =>
                           DataPath_RF_bus_reg_dataout_1784_port, regs(1783) =>
                           DataPath_RF_bus_reg_dataout_1783_port, regs(1782) =>
                           DataPath_RF_bus_reg_dataout_1782_port, regs(1781) =>
                           DataPath_RF_bus_reg_dataout_1781_port, regs(1780) =>
                           DataPath_RF_bus_reg_dataout_1780_port, regs(1779) =>
                           DataPath_RF_bus_reg_dataout_1779_port, regs(1778) =>
                           DataPath_RF_bus_reg_dataout_1778_port, regs(1777) =>
                           DataPath_RF_bus_reg_dataout_1777_port, regs(1776) =>
                           DataPath_RF_bus_reg_dataout_1776_port, regs(1775) =>
                           DataPath_RF_bus_reg_dataout_1775_port, regs(1774) =>
                           DataPath_RF_bus_reg_dataout_1774_port, regs(1773) =>
                           DataPath_RF_bus_reg_dataout_1773_port, regs(1772) =>
                           DataPath_RF_bus_reg_dataout_1772_port, regs(1771) =>
                           DataPath_RF_bus_reg_dataout_1771_port, regs(1770) =>
                           DataPath_RF_bus_reg_dataout_1770_port, regs(1769) =>
                           DataPath_RF_bus_reg_dataout_1769_port, regs(1768) =>
                           DataPath_RF_bus_reg_dataout_1768_port, regs(1767) =>
                           DataPath_RF_bus_reg_dataout_1767_port, regs(1766) =>
                           DataPath_RF_bus_reg_dataout_1766_port, regs(1765) =>
                           DataPath_RF_bus_reg_dataout_1765_port, regs(1764) =>
                           DataPath_RF_bus_reg_dataout_1764_port, regs(1763) =>
                           DataPath_RF_bus_reg_dataout_1763_port, regs(1762) =>
                           DataPath_RF_bus_reg_dataout_1762_port, regs(1761) =>
                           DataPath_RF_bus_reg_dataout_1761_port, regs(1760) =>
                           DataPath_RF_bus_reg_dataout_1760_port, regs(1759) =>
                           DataPath_RF_bus_reg_dataout_1759_port, regs(1758) =>
                           DataPath_RF_bus_reg_dataout_1758_port, regs(1757) =>
                           DataPath_RF_bus_reg_dataout_1757_port, regs(1756) =>
                           DataPath_RF_bus_reg_dataout_1756_port, regs(1755) =>
                           DataPath_RF_bus_reg_dataout_1755_port, regs(1754) =>
                           DataPath_RF_bus_reg_dataout_1754_port, regs(1753) =>
                           DataPath_RF_bus_reg_dataout_1753_port, regs(1752) =>
                           DataPath_RF_bus_reg_dataout_1752_port, regs(1751) =>
                           DataPath_RF_bus_reg_dataout_1751_port, regs(1750) =>
                           DataPath_RF_bus_reg_dataout_1750_port, regs(1749) =>
                           DataPath_RF_bus_reg_dataout_1749_port, regs(1748) =>
                           DataPath_RF_bus_reg_dataout_1748_port, regs(1747) =>
                           DataPath_RF_bus_reg_dataout_1747_port, regs(1746) =>
                           DataPath_RF_bus_reg_dataout_1746_port, regs(1745) =>
                           DataPath_RF_bus_reg_dataout_1745_port, regs(1744) =>
                           DataPath_RF_bus_reg_dataout_1744_port, regs(1743) =>
                           DataPath_RF_bus_reg_dataout_1743_port, regs(1742) =>
                           DataPath_RF_bus_reg_dataout_1742_port, regs(1741) =>
                           DataPath_RF_bus_reg_dataout_1741_port, regs(1740) =>
                           DataPath_RF_bus_reg_dataout_1740_port, regs(1739) =>
                           DataPath_RF_bus_reg_dataout_1739_port, regs(1738) =>
                           DataPath_RF_bus_reg_dataout_1738_port, regs(1737) =>
                           DataPath_RF_bus_reg_dataout_1737_port, regs(1736) =>
                           DataPath_RF_bus_reg_dataout_1736_port, regs(1735) =>
                           DataPath_RF_bus_reg_dataout_1735_port, regs(1734) =>
                           DataPath_RF_bus_reg_dataout_1734_port, regs(1733) =>
                           DataPath_RF_bus_reg_dataout_1733_port, regs(1732) =>
                           DataPath_RF_bus_reg_dataout_1732_port, regs(1731) =>
                           DataPath_RF_bus_reg_dataout_1731_port, regs(1730) =>
                           DataPath_RF_bus_reg_dataout_1730_port, regs(1729) =>
                           DataPath_RF_bus_reg_dataout_1729_port, regs(1728) =>
                           DataPath_RF_bus_reg_dataout_1728_port, regs(1727) =>
                           DataPath_RF_bus_reg_dataout_1727_port, regs(1726) =>
                           DataPath_RF_bus_reg_dataout_1726_port, regs(1725) =>
                           DataPath_RF_bus_reg_dataout_1725_port, regs(1724) =>
                           DataPath_RF_bus_reg_dataout_1724_port, regs(1723) =>
                           DataPath_RF_bus_reg_dataout_1723_port, regs(1722) =>
                           DataPath_RF_bus_reg_dataout_1722_port, regs(1721) =>
                           DataPath_RF_bus_reg_dataout_1721_port, regs(1720) =>
                           DataPath_RF_bus_reg_dataout_1720_port, regs(1719) =>
                           DataPath_RF_bus_reg_dataout_1719_port, regs(1718) =>
                           DataPath_RF_bus_reg_dataout_1718_port, regs(1717) =>
                           DataPath_RF_bus_reg_dataout_1717_port, regs(1716) =>
                           DataPath_RF_bus_reg_dataout_1716_port, regs(1715) =>
                           DataPath_RF_bus_reg_dataout_1715_port, regs(1714) =>
                           DataPath_RF_bus_reg_dataout_1714_port, regs(1713) =>
                           DataPath_RF_bus_reg_dataout_1713_port, regs(1712) =>
                           DataPath_RF_bus_reg_dataout_1712_port, regs(1711) =>
                           DataPath_RF_bus_reg_dataout_1711_port, regs(1710) =>
                           DataPath_RF_bus_reg_dataout_1710_port, regs(1709) =>
                           DataPath_RF_bus_reg_dataout_1709_port, regs(1708) =>
                           DataPath_RF_bus_reg_dataout_1708_port, regs(1707) =>
                           DataPath_RF_bus_reg_dataout_1707_port, regs(1706) =>
                           DataPath_RF_bus_reg_dataout_1706_port, regs(1705) =>
                           DataPath_RF_bus_reg_dataout_1705_port, regs(1704) =>
                           DataPath_RF_bus_reg_dataout_1704_port, regs(1703) =>
                           DataPath_RF_bus_reg_dataout_1703_port, regs(1702) =>
                           DataPath_RF_bus_reg_dataout_1702_port, regs(1701) =>
                           DataPath_RF_bus_reg_dataout_1701_port, regs(1700) =>
                           DataPath_RF_bus_reg_dataout_1700_port, regs(1699) =>
                           DataPath_RF_bus_reg_dataout_1699_port, regs(1698) =>
                           DataPath_RF_bus_reg_dataout_1698_port, regs(1697) =>
                           DataPath_RF_bus_reg_dataout_1697_port, regs(1696) =>
                           DataPath_RF_bus_reg_dataout_1696_port, regs(1695) =>
                           DataPath_RF_bus_reg_dataout_1695_port, regs(1694) =>
                           DataPath_RF_bus_reg_dataout_1694_port, regs(1693) =>
                           DataPath_RF_bus_reg_dataout_1693_port, regs(1692) =>
                           DataPath_RF_bus_reg_dataout_1692_port, regs(1691) =>
                           DataPath_RF_bus_reg_dataout_1691_port, regs(1690) =>
                           DataPath_RF_bus_reg_dataout_1690_port, regs(1689) =>
                           DataPath_RF_bus_reg_dataout_1689_port, regs(1688) =>
                           DataPath_RF_bus_reg_dataout_1688_port, regs(1687) =>
                           DataPath_RF_bus_reg_dataout_1687_port, regs(1686) =>
                           DataPath_RF_bus_reg_dataout_1686_port, regs(1685) =>
                           DataPath_RF_bus_reg_dataout_1685_port, regs(1684) =>
                           DataPath_RF_bus_reg_dataout_1684_port, regs(1683) =>
                           DataPath_RF_bus_reg_dataout_1683_port, regs(1682) =>
                           DataPath_RF_bus_reg_dataout_1682_port, regs(1681) =>
                           DataPath_RF_bus_reg_dataout_1681_port, regs(1680) =>
                           DataPath_RF_bus_reg_dataout_1680_port, regs(1679) =>
                           DataPath_RF_bus_reg_dataout_1679_port, regs(1678) =>
                           DataPath_RF_bus_reg_dataout_1678_port, regs(1677) =>
                           DataPath_RF_bus_reg_dataout_1677_port, regs(1676) =>
                           DataPath_RF_bus_reg_dataout_1676_port, regs(1675) =>
                           DataPath_RF_bus_reg_dataout_1675_port, regs(1674) =>
                           DataPath_RF_bus_reg_dataout_1674_port, regs(1673) =>
                           DataPath_RF_bus_reg_dataout_1673_port, regs(1672) =>
                           DataPath_RF_bus_reg_dataout_1672_port, regs(1671) =>
                           DataPath_RF_bus_reg_dataout_1671_port, regs(1670) =>
                           DataPath_RF_bus_reg_dataout_1670_port, regs(1669) =>
                           DataPath_RF_bus_reg_dataout_1669_port, regs(1668) =>
                           DataPath_RF_bus_reg_dataout_1668_port, regs(1667) =>
                           DataPath_RF_bus_reg_dataout_1667_port, regs(1666) =>
                           DataPath_RF_bus_reg_dataout_1666_port, regs(1665) =>
                           DataPath_RF_bus_reg_dataout_1665_port, regs(1664) =>
                           DataPath_RF_bus_reg_dataout_1664_port, regs(1663) =>
                           DataPath_RF_bus_reg_dataout_1663_port, regs(1662) =>
                           DataPath_RF_bus_reg_dataout_1662_port, regs(1661) =>
                           DataPath_RF_bus_reg_dataout_1661_port, regs(1660) =>
                           DataPath_RF_bus_reg_dataout_1660_port, regs(1659) =>
                           DataPath_RF_bus_reg_dataout_1659_port, regs(1658) =>
                           DataPath_RF_bus_reg_dataout_1658_port, regs(1657) =>
                           DataPath_RF_bus_reg_dataout_1657_port, regs(1656) =>
                           DataPath_RF_bus_reg_dataout_1656_port, regs(1655) =>
                           DataPath_RF_bus_reg_dataout_1655_port, regs(1654) =>
                           DataPath_RF_bus_reg_dataout_1654_port, regs(1653) =>
                           DataPath_RF_bus_reg_dataout_1653_port, regs(1652) =>
                           DataPath_RF_bus_reg_dataout_1652_port, regs(1651) =>
                           DataPath_RF_bus_reg_dataout_1651_port, regs(1650) =>
                           DataPath_RF_bus_reg_dataout_1650_port, regs(1649) =>
                           DataPath_RF_bus_reg_dataout_1649_port, regs(1648) =>
                           DataPath_RF_bus_reg_dataout_1648_port, regs(1647) =>
                           DataPath_RF_bus_reg_dataout_1647_port, regs(1646) =>
                           DataPath_RF_bus_reg_dataout_1646_port, regs(1645) =>
                           DataPath_RF_bus_reg_dataout_1645_port, regs(1644) =>
                           DataPath_RF_bus_reg_dataout_1644_port, regs(1643) =>
                           DataPath_RF_bus_reg_dataout_1643_port, regs(1642) =>
                           DataPath_RF_bus_reg_dataout_1642_port, regs(1641) =>
                           DataPath_RF_bus_reg_dataout_1641_port, regs(1640) =>
                           DataPath_RF_bus_reg_dataout_1640_port, regs(1639) =>
                           DataPath_RF_bus_reg_dataout_1639_port, regs(1638) =>
                           DataPath_RF_bus_reg_dataout_1638_port, regs(1637) =>
                           DataPath_RF_bus_reg_dataout_1637_port, regs(1636) =>
                           DataPath_RF_bus_reg_dataout_1636_port, regs(1635) =>
                           DataPath_RF_bus_reg_dataout_1635_port, regs(1634) =>
                           DataPath_RF_bus_reg_dataout_1634_port, regs(1633) =>
                           DataPath_RF_bus_reg_dataout_1633_port, regs(1632) =>
                           DataPath_RF_bus_reg_dataout_1632_port, regs(1631) =>
                           DataPath_RF_bus_reg_dataout_1631_port, regs(1630) =>
                           DataPath_RF_bus_reg_dataout_1630_port, regs(1629) =>
                           DataPath_RF_bus_reg_dataout_1629_port, regs(1628) =>
                           DataPath_RF_bus_reg_dataout_1628_port, regs(1627) =>
                           DataPath_RF_bus_reg_dataout_1627_port, regs(1626) =>
                           DataPath_RF_bus_reg_dataout_1626_port, regs(1625) =>
                           DataPath_RF_bus_reg_dataout_1625_port, regs(1624) =>
                           DataPath_RF_bus_reg_dataout_1624_port, regs(1623) =>
                           DataPath_RF_bus_reg_dataout_1623_port, regs(1622) =>
                           DataPath_RF_bus_reg_dataout_1622_port, regs(1621) =>
                           DataPath_RF_bus_reg_dataout_1621_port, regs(1620) =>
                           DataPath_RF_bus_reg_dataout_1620_port, regs(1619) =>
                           DataPath_RF_bus_reg_dataout_1619_port, regs(1618) =>
                           DataPath_RF_bus_reg_dataout_1618_port, regs(1617) =>
                           DataPath_RF_bus_reg_dataout_1617_port, regs(1616) =>
                           DataPath_RF_bus_reg_dataout_1616_port, regs(1615) =>
                           DataPath_RF_bus_reg_dataout_1615_port, regs(1614) =>
                           DataPath_RF_bus_reg_dataout_1614_port, regs(1613) =>
                           DataPath_RF_bus_reg_dataout_1613_port, regs(1612) =>
                           DataPath_RF_bus_reg_dataout_1612_port, regs(1611) =>
                           DataPath_RF_bus_reg_dataout_1611_port, regs(1610) =>
                           DataPath_RF_bus_reg_dataout_1610_port, regs(1609) =>
                           DataPath_RF_bus_reg_dataout_1609_port, regs(1608) =>
                           DataPath_RF_bus_reg_dataout_1608_port, regs(1607) =>
                           DataPath_RF_bus_reg_dataout_1607_port, regs(1606) =>
                           DataPath_RF_bus_reg_dataout_1606_port, regs(1605) =>
                           DataPath_RF_bus_reg_dataout_1605_port, regs(1604) =>
                           DataPath_RF_bus_reg_dataout_1604_port, regs(1603) =>
                           DataPath_RF_bus_reg_dataout_1603_port, regs(1602) =>
                           DataPath_RF_bus_reg_dataout_1602_port, regs(1601) =>
                           DataPath_RF_bus_reg_dataout_1601_port, regs(1600) =>
                           DataPath_RF_bus_reg_dataout_1600_port, regs(1599) =>
                           DataPath_RF_bus_reg_dataout_1599_port, regs(1598) =>
                           DataPath_RF_bus_reg_dataout_1598_port, regs(1597) =>
                           DataPath_RF_bus_reg_dataout_1597_port, regs(1596) =>
                           DataPath_RF_bus_reg_dataout_1596_port, regs(1595) =>
                           DataPath_RF_bus_reg_dataout_1595_port, regs(1594) =>
                           DataPath_RF_bus_reg_dataout_1594_port, regs(1593) =>
                           DataPath_RF_bus_reg_dataout_1593_port, regs(1592) =>
                           DataPath_RF_bus_reg_dataout_1592_port, regs(1591) =>
                           DataPath_RF_bus_reg_dataout_1591_port, regs(1590) =>
                           DataPath_RF_bus_reg_dataout_1590_port, regs(1589) =>
                           DataPath_RF_bus_reg_dataout_1589_port, regs(1588) =>
                           DataPath_RF_bus_reg_dataout_1588_port, regs(1587) =>
                           DataPath_RF_bus_reg_dataout_1587_port, regs(1586) =>
                           DataPath_RF_bus_reg_dataout_1586_port, regs(1585) =>
                           DataPath_RF_bus_reg_dataout_1585_port, regs(1584) =>
                           DataPath_RF_bus_reg_dataout_1584_port, regs(1583) =>
                           DataPath_RF_bus_reg_dataout_1583_port, regs(1582) =>
                           DataPath_RF_bus_reg_dataout_1582_port, regs(1581) =>
                           DataPath_RF_bus_reg_dataout_1581_port, regs(1580) =>
                           DataPath_RF_bus_reg_dataout_1580_port, regs(1579) =>
                           DataPath_RF_bus_reg_dataout_1579_port, regs(1578) =>
                           DataPath_RF_bus_reg_dataout_1578_port, regs(1577) =>
                           DataPath_RF_bus_reg_dataout_1577_port, regs(1576) =>
                           DataPath_RF_bus_reg_dataout_1576_port, regs(1575) =>
                           DataPath_RF_bus_reg_dataout_1575_port, regs(1574) =>
                           DataPath_RF_bus_reg_dataout_1574_port, regs(1573) =>
                           DataPath_RF_bus_reg_dataout_1573_port, regs(1572) =>
                           DataPath_RF_bus_reg_dataout_1572_port, regs(1571) =>
                           DataPath_RF_bus_reg_dataout_1571_port, regs(1570) =>
                           DataPath_RF_bus_reg_dataout_1570_port, regs(1569) =>
                           DataPath_RF_bus_reg_dataout_1569_port, regs(1568) =>
                           DataPath_RF_bus_reg_dataout_1568_port, regs(1567) =>
                           DataPath_RF_bus_reg_dataout_1567_port, regs(1566) =>
                           DataPath_RF_bus_reg_dataout_1566_port, regs(1565) =>
                           DataPath_RF_bus_reg_dataout_1565_port, regs(1564) =>
                           DataPath_RF_bus_reg_dataout_1564_port, regs(1563) =>
                           DataPath_RF_bus_reg_dataout_1563_port, regs(1562) =>
                           DataPath_RF_bus_reg_dataout_1562_port, regs(1561) =>
                           DataPath_RF_bus_reg_dataout_1561_port, regs(1560) =>
                           DataPath_RF_bus_reg_dataout_1560_port, regs(1559) =>
                           DataPath_RF_bus_reg_dataout_1559_port, regs(1558) =>
                           DataPath_RF_bus_reg_dataout_1558_port, regs(1557) =>
                           DataPath_RF_bus_reg_dataout_1557_port, regs(1556) =>
                           DataPath_RF_bus_reg_dataout_1556_port, regs(1555) =>
                           DataPath_RF_bus_reg_dataout_1555_port, regs(1554) =>
                           DataPath_RF_bus_reg_dataout_1554_port, regs(1553) =>
                           DataPath_RF_bus_reg_dataout_1553_port, regs(1552) =>
                           DataPath_RF_bus_reg_dataout_1552_port, regs(1551) =>
                           DataPath_RF_bus_reg_dataout_1551_port, regs(1550) =>
                           DataPath_RF_bus_reg_dataout_1550_port, regs(1549) =>
                           DataPath_RF_bus_reg_dataout_1549_port, regs(1548) =>
                           DataPath_RF_bus_reg_dataout_1548_port, regs(1547) =>
                           DataPath_RF_bus_reg_dataout_1547_port, regs(1546) =>
                           DataPath_RF_bus_reg_dataout_1546_port, regs(1545) =>
                           DataPath_RF_bus_reg_dataout_1545_port, regs(1544) =>
                           DataPath_RF_bus_reg_dataout_1544_port, regs(1543) =>
                           DataPath_RF_bus_reg_dataout_1543_port, regs(1542) =>
                           DataPath_RF_bus_reg_dataout_1542_port, regs(1541) =>
                           DataPath_RF_bus_reg_dataout_1541_port, regs(1540) =>
                           DataPath_RF_bus_reg_dataout_1540_port, regs(1539) =>
                           DataPath_RF_bus_reg_dataout_1539_port, regs(1538) =>
                           DataPath_RF_bus_reg_dataout_1538_port, regs(1537) =>
                           DataPath_RF_bus_reg_dataout_1537_port, regs(1536) =>
                           DataPath_RF_bus_reg_dataout_1536_port, regs(1535) =>
                           DataPath_RF_bus_reg_dataout_1535_port, regs(1534) =>
                           DataPath_RF_bus_reg_dataout_1534_port, regs(1533) =>
                           DataPath_RF_bus_reg_dataout_1533_port, regs(1532) =>
                           DataPath_RF_bus_reg_dataout_1532_port, regs(1531) =>
                           DataPath_RF_bus_reg_dataout_1531_port, regs(1530) =>
                           DataPath_RF_bus_reg_dataout_1530_port, regs(1529) =>
                           DataPath_RF_bus_reg_dataout_1529_port, regs(1528) =>
                           DataPath_RF_bus_reg_dataout_1528_port, regs(1527) =>
                           DataPath_RF_bus_reg_dataout_1527_port, regs(1526) =>
                           DataPath_RF_bus_reg_dataout_1526_port, regs(1525) =>
                           DataPath_RF_bus_reg_dataout_1525_port, regs(1524) =>
                           DataPath_RF_bus_reg_dataout_1524_port, regs(1523) =>
                           DataPath_RF_bus_reg_dataout_1523_port, regs(1522) =>
                           DataPath_RF_bus_reg_dataout_1522_port, regs(1521) =>
                           DataPath_RF_bus_reg_dataout_1521_port, regs(1520) =>
                           DataPath_RF_bus_reg_dataout_1520_port, regs(1519) =>
                           DataPath_RF_bus_reg_dataout_1519_port, regs(1518) =>
                           DataPath_RF_bus_reg_dataout_1518_port, regs(1517) =>
                           DataPath_RF_bus_reg_dataout_1517_port, regs(1516) =>
                           DataPath_RF_bus_reg_dataout_1516_port, regs(1515) =>
                           DataPath_RF_bus_reg_dataout_1515_port, regs(1514) =>
                           DataPath_RF_bus_reg_dataout_1514_port, regs(1513) =>
                           DataPath_RF_bus_reg_dataout_1513_port, regs(1512) =>
                           DataPath_RF_bus_reg_dataout_1512_port, regs(1511) =>
                           DataPath_RF_bus_reg_dataout_1511_port, regs(1510) =>
                           DataPath_RF_bus_reg_dataout_1510_port, regs(1509) =>
                           DataPath_RF_bus_reg_dataout_1509_port, regs(1508) =>
                           DataPath_RF_bus_reg_dataout_1508_port, regs(1507) =>
                           DataPath_RF_bus_reg_dataout_1507_port, regs(1506) =>
                           DataPath_RF_bus_reg_dataout_1506_port, regs(1505) =>
                           DataPath_RF_bus_reg_dataout_1505_port, regs(1504) =>
                           DataPath_RF_bus_reg_dataout_1504_port, regs(1503) =>
                           DataPath_RF_bus_reg_dataout_1503_port, regs(1502) =>
                           DataPath_RF_bus_reg_dataout_1502_port, regs(1501) =>
                           DataPath_RF_bus_reg_dataout_1501_port, regs(1500) =>
                           DataPath_RF_bus_reg_dataout_1500_port, regs(1499) =>
                           DataPath_RF_bus_reg_dataout_1499_port, regs(1498) =>
                           DataPath_RF_bus_reg_dataout_1498_port, regs(1497) =>
                           DataPath_RF_bus_reg_dataout_1497_port, regs(1496) =>
                           DataPath_RF_bus_reg_dataout_1496_port, regs(1495) =>
                           DataPath_RF_bus_reg_dataout_1495_port, regs(1494) =>
                           DataPath_RF_bus_reg_dataout_1494_port, regs(1493) =>
                           DataPath_RF_bus_reg_dataout_1493_port, regs(1492) =>
                           DataPath_RF_bus_reg_dataout_1492_port, regs(1491) =>
                           DataPath_RF_bus_reg_dataout_1491_port, regs(1490) =>
                           DataPath_RF_bus_reg_dataout_1490_port, regs(1489) =>
                           DataPath_RF_bus_reg_dataout_1489_port, regs(1488) =>
                           DataPath_RF_bus_reg_dataout_1488_port, regs(1487) =>
                           DataPath_RF_bus_reg_dataout_1487_port, regs(1486) =>
                           DataPath_RF_bus_reg_dataout_1486_port, regs(1485) =>
                           DataPath_RF_bus_reg_dataout_1485_port, regs(1484) =>
                           DataPath_RF_bus_reg_dataout_1484_port, regs(1483) =>
                           DataPath_RF_bus_reg_dataout_1483_port, regs(1482) =>
                           DataPath_RF_bus_reg_dataout_1482_port, regs(1481) =>
                           DataPath_RF_bus_reg_dataout_1481_port, regs(1480) =>
                           DataPath_RF_bus_reg_dataout_1480_port, regs(1479) =>
                           DataPath_RF_bus_reg_dataout_1479_port, regs(1478) =>
                           DataPath_RF_bus_reg_dataout_1478_port, regs(1477) =>
                           DataPath_RF_bus_reg_dataout_1477_port, regs(1476) =>
                           DataPath_RF_bus_reg_dataout_1476_port, regs(1475) =>
                           DataPath_RF_bus_reg_dataout_1475_port, regs(1474) =>
                           DataPath_RF_bus_reg_dataout_1474_port, regs(1473) =>
                           DataPath_RF_bus_reg_dataout_1473_port, regs(1472) =>
                           DataPath_RF_bus_reg_dataout_1472_port, regs(1471) =>
                           DataPath_RF_bus_reg_dataout_1471_port, regs(1470) =>
                           DataPath_RF_bus_reg_dataout_1470_port, regs(1469) =>
                           DataPath_RF_bus_reg_dataout_1469_port, regs(1468) =>
                           DataPath_RF_bus_reg_dataout_1468_port, regs(1467) =>
                           DataPath_RF_bus_reg_dataout_1467_port, regs(1466) =>
                           DataPath_RF_bus_reg_dataout_1466_port, regs(1465) =>
                           DataPath_RF_bus_reg_dataout_1465_port, regs(1464) =>
                           DataPath_RF_bus_reg_dataout_1464_port, regs(1463) =>
                           DataPath_RF_bus_reg_dataout_1463_port, regs(1462) =>
                           DataPath_RF_bus_reg_dataout_1462_port, regs(1461) =>
                           DataPath_RF_bus_reg_dataout_1461_port, regs(1460) =>
                           DataPath_RF_bus_reg_dataout_1460_port, regs(1459) =>
                           DataPath_RF_bus_reg_dataout_1459_port, regs(1458) =>
                           DataPath_RF_bus_reg_dataout_1458_port, regs(1457) =>
                           DataPath_RF_bus_reg_dataout_1457_port, regs(1456) =>
                           DataPath_RF_bus_reg_dataout_1456_port, regs(1455) =>
                           DataPath_RF_bus_reg_dataout_1455_port, regs(1454) =>
                           DataPath_RF_bus_reg_dataout_1454_port, regs(1453) =>
                           DataPath_RF_bus_reg_dataout_1453_port, regs(1452) =>
                           DataPath_RF_bus_reg_dataout_1452_port, regs(1451) =>
                           DataPath_RF_bus_reg_dataout_1451_port, regs(1450) =>
                           DataPath_RF_bus_reg_dataout_1450_port, regs(1449) =>
                           DataPath_RF_bus_reg_dataout_1449_port, regs(1448) =>
                           DataPath_RF_bus_reg_dataout_1448_port, regs(1447) =>
                           DataPath_RF_bus_reg_dataout_1447_port, regs(1446) =>
                           DataPath_RF_bus_reg_dataout_1446_port, regs(1445) =>
                           DataPath_RF_bus_reg_dataout_1445_port, regs(1444) =>
                           DataPath_RF_bus_reg_dataout_1444_port, regs(1443) =>
                           DataPath_RF_bus_reg_dataout_1443_port, regs(1442) =>
                           DataPath_RF_bus_reg_dataout_1442_port, regs(1441) =>
                           DataPath_RF_bus_reg_dataout_1441_port, regs(1440) =>
                           DataPath_RF_bus_reg_dataout_1440_port, regs(1439) =>
                           DataPath_RF_bus_reg_dataout_1439_port, regs(1438) =>
                           DataPath_RF_bus_reg_dataout_1438_port, regs(1437) =>
                           DataPath_RF_bus_reg_dataout_1437_port, regs(1436) =>
                           DataPath_RF_bus_reg_dataout_1436_port, regs(1435) =>
                           DataPath_RF_bus_reg_dataout_1435_port, regs(1434) =>
                           DataPath_RF_bus_reg_dataout_1434_port, regs(1433) =>
                           DataPath_RF_bus_reg_dataout_1433_port, regs(1432) =>
                           DataPath_RF_bus_reg_dataout_1432_port, regs(1431) =>
                           DataPath_RF_bus_reg_dataout_1431_port, regs(1430) =>
                           DataPath_RF_bus_reg_dataout_1430_port, regs(1429) =>
                           DataPath_RF_bus_reg_dataout_1429_port, regs(1428) =>
                           DataPath_RF_bus_reg_dataout_1428_port, regs(1427) =>
                           DataPath_RF_bus_reg_dataout_1427_port, regs(1426) =>
                           DataPath_RF_bus_reg_dataout_1426_port, regs(1425) =>
                           DataPath_RF_bus_reg_dataout_1425_port, regs(1424) =>
                           DataPath_RF_bus_reg_dataout_1424_port, regs(1423) =>
                           DataPath_RF_bus_reg_dataout_1423_port, regs(1422) =>
                           DataPath_RF_bus_reg_dataout_1422_port, regs(1421) =>
                           DataPath_RF_bus_reg_dataout_1421_port, regs(1420) =>
                           DataPath_RF_bus_reg_dataout_1420_port, regs(1419) =>
                           DataPath_RF_bus_reg_dataout_1419_port, regs(1418) =>
                           DataPath_RF_bus_reg_dataout_1418_port, regs(1417) =>
                           DataPath_RF_bus_reg_dataout_1417_port, regs(1416) =>
                           DataPath_RF_bus_reg_dataout_1416_port, regs(1415) =>
                           DataPath_RF_bus_reg_dataout_1415_port, regs(1414) =>
                           DataPath_RF_bus_reg_dataout_1414_port, regs(1413) =>
                           DataPath_RF_bus_reg_dataout_1413_port, regs(1412) =>
                           DataPath_RF_bus_reg_dataout_1412_port, regs(1411) =>
                           DataPath_RF_bus_reg_dataout_1411_port, regs(1410) =>
                           DataPath_RF_bus_reg_dataout_1410_port, regs(1409) =>
                           DataPath_RF_bus_reg_dataout_1409_port, regs(1408) =>
                           DataPath_RF_bus_reg_dataout_1408_port, regs(1407) =>
                           DataPath_RF_bus_reg_dataout_1407_port, regs(1406) =>
                           DataPath_RF_bus_reg_dataout_1406_port, regs(1405) =>
                           DataPath_RF_bus_reg_dataout_1405_port, regs(1404) =>
                           DataPath_RF_bus_reg_dataout_1404_port, regs(1403) =>
                           DataPath_RF_bus_reg_dataout_1403_port, regs(1402) =>
                           DataPath_RF_bus_reg_dataout_1402_port, regs(1401) =>
                           DataPath_RF_bus_reg_dataout_1401_port, regs(1400) =>
                           DataPath_RF_bus_reg_dataout_1400_port, regs(1399) =>
                           DataPath_RF_bus_reg_dataout_1399_port, regs(1398) =>
                           DataPath_RF_bus_reg_dataout_1398_port, regs(1397) =>
                           DataPath_RF_bus_reg_dataout_1397_port, regs(1396) =>
                           DataPath_RF_bus_reg_dataout_1396_port, regs(1395) =>
                           DataPath_RF_bus_reg_dataout_1395_port, regs(1394) =>
                           DataPath_RF_bus_reg_dataout_1394_port, regs(1393) =>
                           DataPath_RF_bus_reg_dataout_1393_port, regs(1392) =>
                           DataPath_RF_bus_reg_dataout_1392_port, regs(1391) =>
                           DataPath_RF_bus_reg_dataout_1391_port, regs(1390) =>
                           DataPath_RF_bus_reg_dataout_1390_port, regs(1389) =>
                           DataPath_RF_bus_reg_dataout_1389_port, regs(1388) =>
                           DataPath_RF_bus_reg_dataout_1388_port, regs(1387) =>
                           DataPath_RF_bus_reg_dataout_1387_port, regs(1386) =>
                           DataPath_RF_bus_reg_dataout_1386_port, regs(1385) =>
                           DataPath_RF_bus_reg_dataout_1385_port, regs(1384) =>
                           DataPath_RF_bus_reg_dataout_1384_port, regs(1383) =>
                           DataPath_RF_bus_reg_dataout_1383_port, regs(1382) =>
                           DataPath_RF_bus_reg_dataout_1382_port, regs(1381) =>
                           DataPath_RF_bus_reg_dataout_1381_port, regs(1380) =>
                           DataPath_RF_bus_reg_dataout_1380_port, regs(1379) =>
                           DataPath_RF_bus_reg_dataout_1379_port, regs(1378) =>
                           DataPath_RF_bus_reg_dataout_1378_port, regs(1377) =>
                           DataPath_RF_bus_reg_dataout_1377_port, regs(1376) =>
                           DataPath_RF_bus_reg_dataout_1376_port, regs(1375) =>
                           DataPath_RF_bus_reg_dataout_1375_port, regs(1374) =>
                           DataPath_RF_bus_reg_dataout_1374_port, regs(1373) =>
                           DataPath_RF_bus_reg_dataout_1373_port, regs(1372) =>
                           DataPath_RF_bus_reg_dataout_1372_port, regs(1371) =>
                           DataPath_RF_bus_reg_dataout_1371_port, regs(1370) =>
                           DataPath_RF_bus_reg_dataout_1370_port, regs(1369) =>
                           DataPath_RF_bus_reg_dataout_1369_port, regs(1368) =>
                           DataPath_RF_bus_reg_dataout_1368_port, regs(1367) =>
                           DataPath_RF_bus_reg_dataout_1367_port, regs(1366) =>
                           DataPath_RF_bus_reg_dataout_1366_port, regs(1365) =>
                           DataPath_RF_bus_reg_dataout_1365_port, regs(1364) =>
                           DataPath_RF_bus_reg_dataout_1364_port, regs(1363) =>
                           DataPath_RF_bus_reg_dataout_1363_port, regs(1362) =>
                           DataPath_RF_bus_reg_dataout_1362_port, regs(1361) =>
                           DataPath_RF_bus_reg_dataout_1361_port, regs(1360) =>
                           DataPath_RF_bus_reg_dataout_1360_port, regs(1359) =>
                           DataPath_RF_bus_reg_dataout_1359_port, regs(1358) =>
                           DataPath_RF_bus_reg_dataout_1358_port, regs(1357) =>
                           DataPath_RF_bus_reg_dataout_1357_port, regs(1356) =>
                           DataPath_RF_bus_reg_dataout_1356_port, regs(1355) =>
                           DataPath_RF_bus_reg_dataout_1355_port, regs(1354) =>
                           DataPath_RF_bus_reg_dataout_1354_port, regs(1353) =>
                           DataPath_RF_bus_reg_dataout_1353_port, regs(1352) =>
                           DataPath_RF_bus_reg_dataout_1352_port, regs(1351) =>
                           DataPath_RF_bus_reg_dataout_1351_port, regs(1350) =>
                           DataPath_RF_bus_reg_dataout_1350_port, regs(1349) =>
                           DataPath_RF_bus_reg_dataout_1349_port, regs(1348) =>
                           DataPath_RF_bus_reg_dataout_1348_port, regs(1347) =>
                           DataPath_RF_bus_reg_dataout_1347_port, regs(1346) =>
                           DataPath_RF_bus_reg_dataout_1346_port, regs(1345) =>
                           DataPath_RF_bus_reg_dataout_1345_port, regs(1344) =>
                           DataPath_RF_bus_reg_dataout_1344_port, regs(1343) =>
                           DataPath_RF_bus_reg_dataout_1343_port, regs(1342) =>
                           DataPath_RF_bus_reg_dataout_1342_port, regs(1341) =>
                           DataPath_RF_bus_reg_dataout_1341_port, regs(1340) =>
                           DataPath_RF_bus_reg_dataout_1340_port, regs(1339) =>
                           DataPath_RF_bus_reg_dataout_1339_port, regs(1338) =>
                           DataPath_RF_bus_reg_dataout_1338_port, regs(1337) =>
                           DataPath_RF_bus_reg_dataout_1337_port, regs(1336) =>
                           DataPath_RF_bus_reg_dataout_1336_port, regs(1335) =>
                           DataPath_RF_bus_reg_dataout_1335_port, regs(1334) =>
                           DataPath_RF_bus_reg_dataout_1334_port, regs(1333) =>
                           DataPath_RF_bus_reg_dataout_1333_port, regs(1332) =>
                           DataPath_RF_bus_reg_dataout_1332_port, regs(1331) =>
                           DataPath_RF_bus_reg_dataout_1331_port, regs(1330) =>
                           DataPath_RF_bus_reg_dataout_1330_port, regs(1329) =>
                           DataPath_RF_bus_reg_dataout_1329_port, regs(1328) =>
                           DataPath_RF_bus_reg_dataout_1328_port, regs(1327) =>
                           DataPath_RF_bus_reg_dataout_1327_port, regs(1326) =>
                           DataPath_RF_bus_reg_dataout_1326_port, regs(1325) =>
                           DataPath_RF_bus_reg_dataout_1325_port, regs(1324) =>
                           DataPath_RF_bus_reg_dataout_1324_port, regs(1323) =>
                           DataPath_RF_bus_reg_dataout_1323_port, regs(1322) =>
                           DataPath_RF_bus_reg_dataout_1322_port, regs(1321) =>
                           DataPath_RF_bus_reg_dataout_1321_port, regs(1320) =>
                           DataPath_RF_bus_reg_dataout_1320_port, regs(1319) =>
                           DataPath_RF_bus_reg_dataout_1319_port, regs(1318) =>
                           DataPath_RF_bus_reg_dataout_1318_port, regs(1317) =>
                           DataPath_RF_bus_reg_dataout_1317_port, regs(1316) =>
                           DataPath_RF_bus_reg_dataout_1316_port, regs(1315) =>
                           DataPath_RF_bus_reg_dataout_1315_port, regs(1314) =>
                           DataPath_RF_bus_reg_dataout_1314_port, regs(1313) =>
                           DataPath_RF_bus_reg_dataout_1313_port, regs(1312) =>
                           DataPath_RF_bus_reg_dataout_1312_port, regs(1311) =>
                           DataPath_RF_bus_reg_dataout_1311_port, regs(1310) =>
                           DataPath_RF_bus_reg_dataout_1310_port, regs(1309) =>
                           DataPath_RF_bus_reg_dataout_1309_port, regs(1308) =>
                           DataPath_RF_bus_reg_dataout_1308_port, regs(1307) =>
                           DataPath_RF_bus_reg_dataout_1307_port, regs(1306) =>
                           DataPath_RF_bus_reg_dataout_1306_port, regs(1305) =>
                           DataPath_RF_bus_reg_dataout_1305_port, regs(1304) =>
                           DataPath_RF_bus_reg_dataout_1304_port, regs(1303) =>
                           DataPath_RF_bus_reg_dataout_1303_port, regs(1302) =>
                           DataPath_RF_bus_reg_dataout_1302_port, regs(1301) =>
                           DataPath_RF_bus_reg_dataout_1301_port, regs(1300) =>
                           DataPath_RF_bus_reg_dataout_1300_port, regs(1299) =>
                           DataPath_RF_bus_reg_dataout_1299_port, regs(1298) =>
                           DataPath_RF_bus_reg_dataout_1298_port, regs(1297) =>
                           DataPath_RF_bus_reg_dataout_1297_port, regs(1296) =>
                           DataPath_RF_bus_reg_dataout_1296_port, regs(1295) =>
                           DataPath_RF_bus_reg_dataout_1295_port, regs(1294) =>
                           DataPath_RF_bus_reg_dataout_1294_port, regs(1293) =>
                           DataPath_RF_bus_reg_dataout_1293_port, regs(1292) =>
                           DataPath_RF_bus_reg_dataout_1292_port, regs(1291) =>
                           DataPath_RF_bus_reg_dataout_1291_port, regs(1290) =>
                           DataPath_RF_bus_reg_dataout_1290_port, regs(1289) =>
                           DataPath_RF_bus_reg_dataout_1289_port, regs(1288) =>
                           DataPath_RF_bus_reg_dataout_1288_port, regs(1287) =>
                           DataPath_RF_bus_reg_dataout_1287_port, regs(1286) =>
                           DataPath_RF_bus_reg_dataout_1286_port, regs(1285) =>
                           DataPath_RF_bus_reg_dataout_1285_port, regs(1284) =>
                           DataPath_RF_bus_reg_dataout_1284_port, regs(1283) =>
                           DataPath_RF_bus_reg_dataout_1283_port, regs(1282) =>
                           DataPath_RF_bus_reg_dataout_1282_port, regs(1281) =>
                           DataPath_RF_bus_reg_dataout_1281_port, regs(1280) =>
                           DataPath_RF_bus_reg_dataout_1280_port, regs(1279) =>
                           DataPath_RF_bus_reg_dataout_1279_port, regs(1278) =>
                           DataPath_RF_bus_reg_dataout_1278_port, regs(1277) =>
                           DataPath_RF_bus_reg_dataout_1277_port, regs(1276) =>
                           DataPath_RF_bus_reg_dataout_1276_port, regs(1275) =>
                           DataPath_RF_bus_reg_dataout_1275_port, regs(1274) =>
                           DataPath_RF_bus_reg_dataout_1274_port, regs(1273) =>
                           DataPath_RF_bus_reg_dataout_1273_port, regs(1272) =>
                           DataPath_RF_bus_reg_dataout_1272_port, regs(1271) =>
                           DataPath_RF_bus_reg_dataout_1271_port, regs(1270) =>
                           DataPath_RF_bus_reg_dataout_1270_port, regs(1269) =>
                           DataPath_RF_bus_reg_dataout_1269_port, regs(1268) =>
                           DataPath_RF_bus_reg_dataout_1268_port, regs(1267) =>
                           DataPath_RF_bus_reg_dataout_1267_port, regs(1266) =>
                           DataPath_RF_bus_reg_dataout_1266_port, regs(1265) =>
                           DataPath_RF_bus_reg_dataout_1265_port, regs(1264) =>
                           DataPath_RF_bus_reg_dataout_1264_port, regs(1263) =>
                           DataPath_RF_bus_reg_dataout_1263_port, regs(1262) =>
                           DataPath_RF_bus_reg_dataout_1262_port, regs(1261) =>
                           DataPath_RF_bus_reg_dataout_1261_port, regs(1260) =>
                           DataPath_RF_bus_reg_dataout_1260_port, regs(1259) =>
                           DataPath_RF_bus_reg_dataout_1259_port, regs(1258) =>
                           DataPath_RF_bus_reg_dataout_1258_port, regs(1257) =>
                           DataPath_RF_bus_reg_dataout_1257_port, regs(1256) =>
                           DataPath_RF_bus_reg_dataout_1256_port, regs(1255) =>
                           DataPath_RF_bus_reg_dataout_1255_port, regs(1254) =>
                           DataPath_RF_bus_reg_dataout_1254_port, regs(1253) =>
                           DataPath_RF_bus_reg_dataout_1253_port, regs(1252) =>
                           DataPath_RF_bus_reg_dataout_1252_port, regs(1251) =>
                           DataPath_RF_bus_reg_dataout_1251_port, regs(1250) =>
                           DataPath_RF_bus_reg_dataout_1250_port, regs(1249) =>
                           DataPath_RF_bus_reg_dataout_1249_port, regs(1248) =>
                           DataPath_RF_bus_reg_dataout_1248_port, regs(1247) =>
                           DataPath_RF_bus_reg_dataout_1247_port, regs(1246) =>
                           DataPath_RF_bus_reg_dataout_1246_port, regs(1245) =>
                           DataPath_RF_bus_reg_dataout_1245_port, regs(1244) =>
                           DataPath_RF_bus_reg_dataout_1244_port, regs(1243) =>
                           DataPath_RF_bus_reg_dataout_1243_port, regs(1242) =>
                           DataPath_RF_bus_reg_dataout_1242_port, regs(1241) =>
                           DataPath_RF_bus_reg_dataout_1241_port, regs(1240) =>
                           DataPath_RF_bus_reg_dataout_1240_port, regs(1239) =>
                           DataPath_RF_bus_reg_dataout_1239_port, regs(1238) =>
                           DataPath_RF_bus_reg_dataout_1238_port, regs(1237) =>
                           DataPath_RF_bus_reg_dataout_1237_port, regs(1236) =>
                           DataPath_RF_bus_reg_dataout_1236_port, regs(1235) =>
                           DataPath_RF_bus_reg_dataout_1235_port, regs(1234) =>
                           DataPath_RF_bus_reg_dataout_1234_port, regs(1233) =>
                           DataPath_RF_bus_reg_dataout_1233_port, regs(1232) =>
                           DataPath_RF_bus_reg_dataout_1232_port, regs(1231) =>
                           DataPath_RF_bus_reg_dataout_1231_port, regs(1230) =>
                           DataPath_RF_bus_reg_dataout_1230_port, regs(1229) =>
                           DataPath_RF_bus_reg_dataout_1229_port, regs(1228) =>
                           DataPath_RF_bus_reg_dataout_1228_port, regs(1227) =>
                           DataPath_RF_bus_reg_dataout_1227_port, regs(1226) =>
                           DataPath_RF_bus_reg_dataout_1226_port, regs(1225) =>
                           DataPath_RF_bus_reg_dataout_1225_port, regs(1224) =>
                           DataPath_RF_bus_reg_dataout_1224_port, regs(1223) =>
                           DataPath_RF_bus_reg_dataout_1223_port, regs(1222) =>
                           DataPath_RF_bus_reg_dataout_1222_port, regs(1221) =>
                           DataPath_RF_bus_reg_dataout_1221_port, regs(1220) =>
                           DataPath_RF_bus_reg_dataout_1220_port, regs(1219) =>
                           DataPath_RF_bus_reg_dataout_1219_port, regs(1218) =>
                           DataPath_RF_bus_reg_dataout_1218_port, regs(1217) =>
                           DataPath_RF_bus_reg_dataout_1217_port, regs(1216) =>
                           DataPath_RF_bus_reg_dataout_1216_port, regs(1215) =>
                           DataPath_RF_bus_reg_dataout_1215_port, regs(1214) =>
                           DataPath_RF_bus_reg_dataout_1214_port, regs(1213) =>
                           DataPath_RF_bus_reg_dataout_1213_port, regs(1212) =>
                           DataPath_RF_bus_reg_dataout_1212_port, regs(1211) =>
                           DataPath_RF_bus_reg_dataout_1211_port, regs(1210) =>
                           DataPath_RF_bus_reg_dataout_1210_port, regs(1209) =>
                           DataPath_RF_bus_reg_dataout_1209_port, regs(1208) =>
                           DataPath_RF_bus_reg_dataout_1208_port, regs(1207) =>
                           DataPath_RF_bus_reg_dataout_1207_port, regs(1206) =>
                           DataPath_RF_bus_reg_dataout_1206_port, regs(1205) =>
                           DataPath_RF_bus_reg_dataout_1205_port, regs(1204) =>
                           DataPath_RF_bus_reg_dataout_1204_port, regs(1203) =>
                           DataPath_RF_bus_reg_dataout_1203_port, regs(1202) =>
                           DataPath_RF_bus_reg_dataout_1202_port, regs(1201) =>
                           DataPath_RF_bus_reg_dataout_1201_port, regs(1200) =>
                           DataPath_RF_bus_reg_dataout_1200_port, regs(1199) =>
                           DataPath_RF_bus_reg_dataout_1199_port, regs(1198) =>
                           DataPath_RF_bus_reg_dataout_1198_port, regs(1197) =>
                           DataPath_RF_bus_reg_dataout_1197_port, regs(1196) =>
                           DataPath_RF_bus_reg_dataout_1196_port, regs(1195) =>
                           DataPath_RF_bus_reg_dataout_1195_port, regs(1194) =>
                           DataPath_RF_bus_reg_dataout_1194_port, regs(1193) =>
                           DataPath_RF_bus_reg_dataout_1193_port, regs(1192) =>
                           DataPath_RF_bus_reg_dataout_1192_port, regs(1191) =>
                           DataPath_RF_bus_reg_dataout_1191_port, regs(1190) =>
                           DataPath_RF_bus_reg_dataout_1190_port, regs(1189) =>
                           DataPath_RF_bus_reg_dataout_1189_port, regs(1188) =>
                           DataPath_RF_bus_reg_dataout_1188_port, regs(1187) =>
                           DataPath_RF_bus_reg_dataout_1187_port, regs(1186) =>
                           DataPath_RF_bus_reg_dataout_1186_port, regs(1185) =>
                           DataPath_RF_bus_reg_dataout_1185_port, regs(1184) =>
                           DataPath_RF_bus_reg_dataout_1184_port, regs(1183) =>
                           DataPath_RF_bus_reg_dataout_1183_port, regs(1182) =>
                           DataPath_RF_bus_reg_dataout_1182_port, regs(1181) =>
                           DataPath_RF_bus_reg_dataout_1181_port, regs(1180) =>
                           DataPath_RF_bus_reg_dataout_1180_port, regs(1179) =>
                           DataPath_RF_bus_reg_dataout_1179_port, regs(1178) =>
                           DataPath_RF_bus_reg_dataout_1178_port, regs(1177) =>
                           DataPath_RF_bus_reg_dataout_1177_port, regs(1176) =>
                           DataPath_RF_bus_reg_dataout_1176_port, regs(1175) =>
                           DataPath_RF_bus_reg_dataout_1175_port, regs(1174) =>
                           DataPath_RF_bus_reg_dataout_1174_port, regs(1173) =>
                           DataPath_RF_bus_reg_dataout_1173_port, regs(1172) =>
                           DataPath_RF_bus_reg_dataout_1172_port, regs(1171) =>
                           DataPath_RF_bus_reg_dataout_1171_port, regs(1170) =>
                           DataPath_RF_bus_reg_dataout_1170_port, regs(1169) =>
                           DataPath_RF_bus_reg_dataout_1169_port, regs(1168) =>
                           DataPath_RF_bus_reg_dataout_1168_port, regs(1167) =>
                           DataPath_RF_bus_reg_dataout_1167_port, regs(1166) =>
                           DataPath_RF_bus_reg_dataout_1166_port, regs(1165) =>
                           DataPath_RF_bus_reg_dataout_1165_port, regs(1164) =>
                           DataPath_RF_bus_reg_dataout_1164_port, regs(1163) =>
                           DataPath_RF_bus_reg_dataout_1163_port, regs(1162) =>
                           DataPath_RF_bus_reg_dataout_1162_port, regs(1161) =>
                           DataPath_RF_bus_reg_dataout_1161_port, regs(1160) =>
                           DataPath_RF_bus_reg_dataout_1160_port, regs(1159) =>
                           DataPath_RF_bus_reg_dataout_1159_port, regs(1158) =>
                           DataPath_RF_bus_reg_dataout_1158_port, regs(1157) =>
                           DataPath_RF_bus_reg_dataout_1157_port, regs(1156) =>
                           DataPath_RF_bus_reg_dataout_1156_port, regs(1155) =>
                           DataPath_RF_bus_reg_dataout_1155_port, regs(1154) =>
                           DataPath_RF_bus_reg_dataout_1154_port, regs(1153) =>
                           DataPath_RF_bus_reg_dataout_1153_port, regs(1152) =>
                           DataPath_RF_bus_reg_dataout_1152_port, regs(1151) =>
                           DataPath_RF_bus_reg_dataout_1151_port, regs(1150) =>
                           DataPath_RF_bus_reg_dataout_1150_port, regs(1149) =>
                           DataPath_RF_bus_reg_dataout_1149_port, regs(1148) =>
                           DataPath_RF_bus_reg_dataout_1148_port, regs(1147) =>
                           DataPath_RF_bus_reg_dataout_1147_port, regs(1146) =>
                           DataPath_RF_bus_reg_dataout_1146_port, regs(1145) =>
                           DataPath_RF_bus_reg_dataout_1145_port, regs(1144) =>
                           DataPath_RF_bus_reg_dataout_1144_port, regs(1143) =>
                           DataPath_RF_bus_reg_dataout_1143_port, regs(1142) =>
                           DataPath_RF_bus_reg_dataout_1142_port, regs(1141) =>
                           DataPath_RF_bus_reg_dataout_1141_port, regs(1140) =>
                           DataPath_RF_bus_reg_dataout_1140_port, regs(1139) =>
                           DataPath_RF_bus_reg_dataout_1139_port, regs(1138) =>
                           DataPath_RF_bus_reg_dataout_1138_port, regs(1137) =>
                           DataPath_RF_bus_reg_dataout_1137_port, regs(1136) =>
                           DataPath_RF_bus_reg_dataout_1136_port, regs(1135) =>
                           DataPath_RF_bus_reg_dataout_1135_port, regs(1134) =>
                           DataPath_RF_bus_reg_dataout_1134_port, regs(1133) =>
                           DataPath_RF_bus_reg_dataout_1133_port, regs(1132) =>
                           DataPath_RF_bus_reg_dataout_1132_port, regs(1131) =>
                           DataPath_RF_bus_reg_dataout_1131_port, regs(1130) =>
                           DataPath_RF_bus_reg_dataout_1130_port, regs(1129) =>
                           DataPath_RF_bus_reg_dataout_1129_port, regs(1128) =>
                           DataPath_RF_bus_reg_dataout_1128_port, regs(1127) =>
                           DataPath_RF_bus_reg_dataout_1127_port, regs(1126) =>
                           DataPath_RF_bus_reg_dataout_1126_port, regs(1125) =>
                           DataPath_RF_bus_reg_dataout_1125_port, regs(1124) =>
                           DataPath_RF_bus_reg_dataout_1124_port, regs(1123) =>
                           DataPath_RF_bus_reg_dataout_1123_port, regs(1122) =>
                           DataPath_RF_bus_reg_dataout_1122_port, regs(1121) =>
                           DataPath_RF_bus_reg_dataout_1121_port, regs(1120) =>
                           DataPath_RF_bus_reg_dataout_1120_port, regs(1119) =>
                           DataPath_RF_bus_reg_dataout_1119_port, regs(1118) =>
                           DataPath_RF_bus_reg_dataout_1118_port, regs(1117) =>
                           DataPath_RF_bus_reg_dataout_1117_port, regs(1116) =>
                           DataPath_RF_bus_reg_dataout_1116_port, regs(1115) =>
                           DataPath_RF_bus_reg_dataout_1115_port, regs(1114) =>
                           DataPath_RF_bus_reg_dataout_1114_port, regs(1113) =>
                           DataPath_RF_bus_reg_dataout_1113_port, regs(1112) =>
                           DataPath_RF_bus_reg_dataout_1112_port, regs(1111) =>
                           DataPath_RF_bus_reg_dataout_1111_port, regs(1110) =>
                           DataPath_RF_bus_reg_dataout_1110_port, regs(1109) =>
                           DataPath_RF_bus_reg_dataout_1109_port, regs(1108) =>
                           DataPath_RF_bus_reg_dataout_1108_port, regs(1107) =>
                           DataPath_RF_bus_reg_dataout_1107_port, regs(1106) =>
                           DataPath_RF_bus_reg_dataout_1106_port, regs(1105) =>
                           DataPath_RF_bus_reg_dataout_1105_port, regs(1104) =>
                           DataPath_RF_bus_reg_dataout_1104_port, regs(1103) =>
                           DataPath_RF_bus_reg_dataout_1103_port, regs(1102) =>
                           DataPath_RF_bus_reg_dataout_1102_port, regs(1101) =>
                           DataPath_RF_bus_reg_dataout_1101_port, regs(1100) =>
                           DataPath_RF_bus_reg_dataout_1100_port, regs(1099) =>
                           DataPath_RF_bus_reg_dataout_1099_port, regs(1098) =>
                           DataPath_RF_bus_reg_dataout_1098_port, regs(1097) =>
                           DataPath_RF_bus_reg_dataout_1097_port, regs(1096) =>
                           DataPath_RF_bus_reg_dataout_1096_port, regs(1095) =>
                           DataPath_RF_bus_reg_dataout_1095_port, regs(1094) =>
                           DataPath_RF_bus_reg_dataout_1094_port, regs(1093) =>
                           DataPath_RF_bus_reg_dataout_1093_port, regs(1092) =>
                           DataPath_RF_bus_reg_dataout_1092_port, regs(1091) =>
                           DataPath_RF_bus_reg_dataout_1091_port, regs(1090) =>
                           DataPath_RF_bus_reg_dataout_1090_port, regs(1089) =>
                           DataPath_RF_bus_reg_dataout_1089_port, regs(1088) =>
                           DataPath_RF_bus_reg_dataout_1088_port, regs(1087) =>
                           DataPath_RF_bus_reg_dataout_1087_port, regs(1086) =>
                           DataPath_RF_bus_reg_dataout_1086_port, regs(1085) =>
                           DataPath_RF_bus_reg_dataout_1085_port, regs(1084) =>
                           DataPath_RF_bus_reg_dataout_1084_port, regs(1083) =>
                           DataPath_RF_bus_reg_dataout_1083_port, regs(1082) =>
                           DataPath_RF_bus_reg_dataout_1082_port, regs(1081) =>
                           DataPath_RF_bus_reg_dataout_1081_port, regs(1080) =>
                           DataPath_RF_bus_reg_dataout_1080_port, regs(1079) =>
                           DataPath_RF_bus_reg_dataout_1079_port, regs(1078) =>
                           DataPath_RF_bus_reg_dataout_1078_port, regs(1077) =>
                           DataPath_RF_bus_reg_dataout_1077_port, regs(1076) =>
                           DataPath_RF_bus_reg_dataout_1076_port, regs(1075) =>
                           DataPath_RF_bus_reg_dataout_1075_port, regs(1074) =>
                           DataPath_RF_bus_reg_dataout_1074_port, regs(1073) =>
                           DataPath_RF_bus_reg_dataout_1073_port, regs(1072) =>
                           DataPath_RF_bus_reg_dataout_1072_port, regs(1071) =>
                           DataPath_RF_bus_reg_dataout_1071_port, regs(1070) =>
                           DataPath_RF_bus_reg_dataout_1070_port, regs(1069) =>
                           DataPath_RF_bus_reg_dataout_1069_port, regs(1068) =>
                           DataPath_RF_bus_reg_dataout_1068_port, regs(1067) =>
                           DataPath_RF_bus_reg_dataout_1067_port, regs(1066) =>
                           DataPath_RF_bus_reg_dataout_1066_port, regs(1065) =>
                           DataPath_RF_bus_reg_dataout_1065_port, regs(1064) =>
                           DataPath_RF_bus_reg_dataout_1064_port, regs(1063) =>
                           DataPath_RF_bus_reg_dataout_1063_port, regs(1062) =>
                           DataPath_RF_bus_reg_dataout_1062_port, regs(1061) =>
                           DataPath_RF_bus_reg_dataout_1061_port, regs(1060) =>
                           DataPath_RF_bus_reg_dataout_1060_port, regs(1059) =>
                           DataPath_RF_bus_reg_dataout_1059_port, regs(1058) =>
                           DataPath_RF_bus_reg_dataout_1058_port, regs(1057) =>
                           DataPath_RF_bus_reg_dataout_1057_port, regs(1056) =>
                           DataPath_RF_bus_reg_dataout_1056_port, regs(1055) =>
                           DataPath_RF_bus_reg_dataout_1055_port, regs(1054) =>
                           DataPath_RF_bus_reg_dataout_1054_port, regs(1053) =>
                           DataPath_RF_bus_reg_dataout_1053_port, regs(1052) =>
                           DataPath_RF_bus_reg_dataout_1052_port, regs(1051) =>
                           DataPath_RF_bus_reg_dataout_1051_port, regs(1050) =>
                           DataPath_RF_bus_reg_dataout_1050_port, regs(1049) =>
                           DataPath_RF_bus_reg_dataout_1049_port, regs(1048) =>
                           DataPath_RF_bus_reg_dataout_1048_port, regs(1047) =>
                           DataPath_RF_bus_reg_dataout_1047_port, regs(1046) =>
                           DataPath_RF_bus_reg_dataout_1046_port, regs(1045) =>
                           DataPath_RF_bus_reg_dataout_1045_port, regs(1044) =>
                           DataPath_RF_bus_reg_dataout_1044_port, regs(1043) =>
                           DataPath_RF_bus_reg_dataout_1043_port, regs(1042) =>
                           DataPath_RF_bus_reg_dataout_1042_port, regs(1041) =>
                           DataPath_RF_bus_reg_dataout_1041_port, regs(1040) =>
                           DataPath_RF_bus_reg_dataout_1040_port, regs(1039) =>
                           DataPath_RF_bus_reg_dataout_1039_port, regs(1038) =>
                           DataPath_RF_bus_reg_dataout_1038_port, regs(1037) =>
                           DataPath_RF_bus_reg_dataout_1037_port, regs(1036) =>
                           DataPath_RF_bus_reg_dataout_1036_port, regs(1035) =>
                           DataPath_RF_bus_reg_dataout_1035_port, regs(1034) =>
                           DataPath_RF_bus_reg_dataout_1034_port, regs(1033) =>
                           DataPath_RF_bus_reg_dataout_1033_port, regs(1032) =>
                           DataPath_RF_bus_reg_dataout_1032_port, regs(1031) =>
                           DataPath_RF_bus_reg_dataout_1031_port, regs(1030) =>
                           DataPath_RF_bus_reg_dataout_1030_port, regs(1029) =>
                           DataPath_RF_bus_reg_dataout_1029_port, regs(1028) =>
                           DataPath_RF_bus_reg_dataout_1028_port, regs(1027) =>
                           DataPath_RF_bus_reg_dataout_1027_port, regs(1026) =>
                           DataPath_RF_bus_reg_dataout_1026_port, regs(1025) =>
                           DataPath_RF_bus_reg_dataout_1025_port, regs(1024) =>
                           DataPath_RF_bus_reg_dataout_1024_port, regs(1023) =>
                           DataPath_RF_bus_reg_dataout_1023_port, regs(1022) =>
                           DataPath_RF_bus_reg_dataout_1022_port, regs(1021) =>
                           DataPath_RF_bus_reg_dataout_1021_port, regs(1020) =>
                           DataPath_RF_bus_reg_dataout_1020_port, regs(1019) =>
                           DataPath_RF_bus_reg_dataout_1019_port, regs(1018) =>
                           DataPath_RF_bus_reg_dataout_1018_port, regs(1017) =>
                           DataPath_RF_bus_reg_dataout_1017_port, regs(1016) =>
                           DataPath_RF_bus_reg_dataout_1016_port, regs(1015) =>
                           DataPath_RF_bus_reg_dataout_1015_port, regs(1014) =>
                           DataPath_RF_bus_reg_dataout_1014_port, regs(1013) =>
                           DataPath_RF_bus_reg_dataout_1013_port, regs(1012) =>
                           DataPath_RF_bus_reg_dataout_1012_port, regs(1011) =>
                           DataPath_RF_bus_reg_dataout_1011_port, regs(1010) =>
                           DataPath_RF_bus_reg_dataout_1010_port, regs(1009) =>
                           DataPath_RF_bus_reg_dataout_1009_port, regs(1008) =>
                           DataPath_RF_bus_reg_dataout_1008_port, regs(1007) =>
                           DataPath_RF_bus_reg_dataout_1007_port, regs(1006) =>
                           DataPath_RF_bus_reg_dataout_1006_port, regs(1005) =>
                           DataPath_RF_bus_reg_dataout_1005_port, regs(1004) =>
                           DataPath_RF_bus_reg_dataout_1004_port, regs(1003) =>
                           DataPath_RF_bus_reg_dataout_1003_port, regs(1002) =>
                           DataPath_RF_bus_reg_dataout_1002_port, regs(1001) =>
                           DataPath_RF_bus_reg_dataout_1001_port, regs(1000) =>
                           DataPath_RF_bus_reg_dataout_1000_port, regs(999) => 
                           DataPath_RF_bus_reg_dataout_999_port, regs(998) => 
                           DataPath_RF_bus_reg_dataout_998_port, regs(997) => 
                           DataPath_RF_bus_reg_dataout_997_port, regs(996) => 
                           DataPath_RF_bus_reg_dataout_996_port, regs(995) => 
                           DataPath_RF_bus_reg_dataout_995_port, regs(994) => 
                           DataPath_RF_bus_reg_dataout_994_port, regs(993) => 
                           DataPath_RF_bus_reg_dataout_993_port, regs(992) => 
                           DataPath_RF_bus_reg_dataout_992_port, regs(991) => 
                           DataPath_RF_bus_reg_dataout_991_port, regs(990) => 
                           DataPath_RF_bus_reg_dataout_990_port, regs(989) => 
                           DataPath_RF_bus_reg_dataout_989_port, regs(988) => 
                           DataPath_RF_bus_reg_dataout_988_port, regs(987) => 
                           DataPath_RF_bus_reg_dataout_987_port, regs(986) => 
                           DataPath_RF_bus_reg_dataout_986_port, regs(985) => 
                           DataPath_RF_bus_reg_dataout_985_port, regs(984) => 
                           DataPath_RF_bus_reg_dataout_984_port, regs(983) => 
                           DataPath_RF_bus_reg_dataout_983_port, regs(982) => 
                           DataPath_RF_bus_reg_dataout_982_port, regs(981) => 
                           DataPath_RF_bus_reg_dataout_981_port, regs(980) => 
                           DataPath_RF_bus_reg_dataout_980_port, regs(979) => 
                           DataPath_RF_bus_reg_dataout_979_port, regs(978) => 
                           DataPath_RF_bus_reg_dataout_978_port, regs(977) => 
                           DataPath_RF_bus_reg_dataout_977_port, regs(976) => 
                           DataPath_RF_bus_reg_dataout_976_port, regs(975) => 
                           DataPath_RF_bus_reg_dataout_975_port, regs(974) => 
                           DataPath_RF_bus_reg_dataout_974_port, regs(973) => 
                           DataPath_RF_bus_reg_dataout_973_port, regs(972) => 
                           DataPath_RF_bus_reg_dataout_972_port, regs(971) => 
                           DataPath_RF_bus_reg_dataout_971_port, regs(970) => 
                           DataPath_RF_bus_reg_dataout_970_port, regs(969) => 
                           DataPath_RF_bus_reg_dataout_969_port, regs(968) => 
                           DataPath_RF_bus_reg_dataout_968_port, regs(967) => 
                           DataPath_RF_bus_reg_dataout_967_port, regs(966) => 
                           DataPath_RF_bus_reg_dataout_966_port, regs(965) => 
                           DataPath_RF_bus_reg_dataout_965_port, regs(964) => 
                           DataPath_RF_bus_reg_dataout_964_port, regs(963) => 
                           DataPath_RF_bus_reg_dataout_963_port, regs(962) => 
                           DataPath_RF_bus_reg_dataout_962_port, regs(961) => 
                           DataPath_RF_bus_reg_dataout_961_port, regs(960) => 
                           DataPath_RF_bus_reg_dataout_960_port, regs(959) => 
                           DataPath_RF_bus_reg_dataout_959_port, regs(958) => 
                           DataPath_RF_bus_reg_dataout_958_port, regs(957) => 
                           DataPath_RF_bus_reg_dataout_957_port, regs(956) => 
                           DataPath_RF_bus_reg_dataout_956_port, regs(955) => 
                           DataPath_RF_bus_reg_dataout_955_port, regs(954) => 
                           DataPath_RF_bus_reg_dataout_954_port, regs(953) => 
                           DataPath_RF_bus_reg_dataout_953_port, regs(952) => 
                           DataPath_RF_bus_reg_dataout_952_port, regs(951) => 
                           DataPath_RF_bus_reg_dataout_951_port, regs(950) => 
                           DataPath_RF_bus_reg_dataout_950_port, regs(949) => 
                           DataPath_RF_bus_reg_dataout_949_port, regs(948) => 
                           DataPath_RF_bus_reg_dataout_948_port, regs(947) => 
                           DataPath_RF_bus_reg_dataout_947_port, regs(946) => 
                           DataPath_RF_bus_reg_dataout_946_port, regs(945) => 
                           DataPath_RF_bus_reg_dataout_945_port, regs(944) => 
                           DataPath_RF_bus_reg_dataout_944_port, regs(943) => 
                           DataPath_RF_bus_reg_dataout_943_port, regs(942) => 
                           DataPath_RF_bus_reg_dataout_942_port, regs(941) => 
                           DataPath_RF_bus_reg_dataout_941_port, regs(940) => 
                           DataPath_RF_bus_reg_dataout_940_port, regs(939) => 
                           DataPath_RF_bus_reg_dataout_939_port, regs(938) => 
                           DataPath_RF_bus_reg_dataout_938_port, regs(937) => 
                           DataPath_RF_bus_reg_dataout_937_port, regs(936) => 
                           DataPath_RF_bus_reg_dataout_936_port, regs(935) => 
                           DataPath_RF_bus_reg_dataout_935_port, regs(934) => 
                           DataPath_RF_bus_reg_dataout_934_port, regs(933) => 
                           DataPath_RF_bus_reg_dataout_933_port, regs(932) => 
                           DataPath_RF_bus_reg_dataout_932_port, regs(931) => 
                           DataPath_RF_bus_reg_dataout_931_port, regs(930) => 
                           DataPath_RF_bus_reg_dataout_930_port, regs(929) => 
                           DataPath_RF_bus_reg_dataout_929_port, regs(928) => 
                           DataPath_RF_bus_reg_dataout_928_port, regs(927) => 
                           DataPath_RF_bus_reg_dataout_927_port, regs(926) => 
                           DataPath_RF_bus_reg_dataout_926_port, regs(925) => 
                           DataPath_RF_bus_reg_dataout_925_port, regs(924) => 
                           DataPath_RF_bus_reg_dataout_924_port, regs(923) => 
                           DataPath_RF_bus_reg_dataout_923_port, regs(922) => 
                           DataPath_RF_bus_reg_dataout_922_port, regs(921) => 
                           DataPath_RF_bus_reg_dataout_921_port, regs(920) => 
                           DataPath_RF_bus_reg_dataout_920_port, regs(919) => 
                           DataPath_RF_bus_reg_dataout_919_port, regs(918) => 
                           DataPath_RF_bus_reg_dataout_918_port, regs(917) => 
                           DataPath_RF_bus_reg_dataout_917_port, regs(916) => 
                           DataPath_RF_bus_reg_dataout_916_port, regs(915) => 
                           DataPath_RF_bus_reg_dataout_915_port, regs(914) => 
                           DataPath_RF_bus_reg_dataout_914_port, regs(913) => 
                           DataPath_RF_bus_reg_dataout_913_port, regs(912) => 
                           DataPath_RF_bus_reg_dataout_912_port, regs(911) => 
                           DataPath_RF_bus_reg_dataout_911_port, regs(910) => 
                           DataPath_RF_bus_reg_dataout_910_port, regs(909) => 
                           DataPath_RF_bus_reg_dataout_909_port, regs(908) => 
                           DataPath_RF_bus_reg_dataout_908_port, regs(907) => 
                           DataPath_RF_bus_reg_dataout_907_port, regs(906) => 
                           DataPath_RF_bus_reg_dataout_906_port, regs(905) => 
                           DataPath_RF_bus_reg_dataout_905_port, regs(904) => 
                           DataPath_RF_bus_reg_dataout_904_port, regs(903) => 
                           DataPath_RF_bus_reg_dataout_903_port, regs(902) => 
                           DataPath_RF_bus_reg_dataout_902_port, regs(901) => 
                           DataPath_RF_bus_reg_dataout_901_port, regs(900) => 
                           DataPath_RF_bus_reg_dataout_900_port, regs(899) => 
                           DataPath_RF_bus_reg_dataout_899_port, regs(898) => 
                           DataPath_RF_bus_reg_dataout_898_port, regs(897) => 
                           DataPath_RF_bus_reg_dataout_897_port, regs(896) => 
                           DataPath_RF_bus_reg_dataout_896_port, regs(895) => 
                           DataPath_RF_bus_reg_dataout_895_port, regs(894) => 
                           DataPath_RF_bus_reg_dataout_894_port, regs(893) => 
                           DataPath_RF_bus_reg_dataout_893_port, regs(892) => 
                           DataPath_RF_bus_reg_dataout_892_port, regs(891) => 
                           DataPath_RF_bus_reg_dataout_891_port, regs(890) => 
                           DataPath_RF_bus_reg_dataout_890_port, regs(889) => 
                           DataPath_RF_bus_reg_dataout_889_port, regs(888) => 
                           DataPath_RF_bus_reg_dataout_888_port, regs(887) => 
                           DataPath_RF_bus_reg_dataout_887_port, regs(886) => 
                           DataPath_RF_bus_reg_dataout_886_port, regs(885) => 
                           DataPath_RF_bus_reg_dataout_885_port, regs(884) => 
                           DataPath_RF_bus_reg_dataout_884_port, regs(883) => 
                           DataPath_RF_bus_reg_dataout_883_port, regs(882) => 
                           DataPath_RF_bus_reg_dataout_882_port, regs(881) => 
                           DataPath_RF_bus_reg_dataout_881_port, regs(880) => 
                           DataPath_RF_bus_reg_dataout_880_port, regs(879) => 
                           DataPath_RF_bus_reg_dataout_879_port, regs(878) => 
                           DataPath_RF_bus_reg_dataout_878_port, regs(877) => 
                           DataPath_RF_bus_reg_dataout_877_port, regs(876) => 
                           DataPath_RF_bus_reg_dataout_876_port, regs(875) => 
                           DataPath_RF_bus_reg_dataout_875_port, regs(874) => 
                           DataPath_RF_bus_reg_dataout_874_port, regs(873) => 
                           DataPath_RF_bus_reg_dataout_873_port, regs(872) => 
                           DataPath_RF_bus_reg_dataout_872_port, regs(871) => 
                           DataPath_RF_bus_reg_dataout_871_port, regs(870) => 
                           DataPath_RF_bus_reg_dataout_870_port, regs(869) => 
                           DataPath_RF_bus_reg_dataout_869_port, regs(868) => 
                           DataPath_RF_bus_reg_dataout_868_port, regs(867) => 
                           DataPath_RF_bus_reg_dataout_867_port, regs(866) => 
                           DataPath_RF_bus_reg_dataout_866_port, regs(865) => 
                           DataPath_RF_bus_reg_dataout_865_port, regs(864) => 
                           DataPath_RF_bus_reg_dataout_864_port, regs(863) => 
                           DataPath_RF_bus_reg_dataout_863_port, regs(862) => 
                           DataPath_RF_bus_reg_dataout_862_port, regs(861) => 
                           DataPath_RF_bus_reg_dataout_861_port, regs(860) => 
                           DataPath_RF_bus_reg_dataout_860_port, regs(859) => 
                           DataPath_RF_bus_reg_dataout_859_port, regs(858) => 
                           DataPath_RF_bus_reg_dataout_858_port, regs(857) => 
                           DataPath_RF_bus_reg_dataout_857_port, regs(856) => 
                           DataPath_RF_bus_reg_dataout_856_port, regs(855) => 
                           DataPath_RF_bus_reg_dataout_855_port, regs(854) => 
                           DataPath_RF_bus_reg_dataout_854_port, regs(853) => 
                           DataPath_RF_bus_reg_dataout_853_port, regs(852) => 
                           DataPath_RF_bus_reg_dataout_852_port, regs(851) => 
                           DataPath_RF_bus_reg_dataout_851_port, regs(850) => 
                           DataPath_RF_bus_reg_dataout_850_port, regs(849) => 
                           DataPath_RF_bus_reg_dataout_849_port, regs(848) => 
                           DataPath_RF_bus_reg_dataout_848_port, regs(847) => 
                           DataPath_RF_bus_reg_dataout_847_port, regs(846) => 
                           DataPath_RF_bus_reg_dataout_846_port, regs(845) => 
                           DataPath_RF_bus_reg_dataout_845_port, regs(844) => 
                           DataPath_RF_bus_reg_dataout_844_port, regs(843) => 
                           DataPath_RF_bus_reg_dataout_843_port, regs(842) => 
                           DataPath_RF_bus_reg_dataout_842_port, regs(841) => 
                           DataPath_RF_bus_reg_dataout_841_port, regs(840) => 
                           DataPath_RF_bus_reg_dataout_840_port, regs(839) => 
                           DataPath_RF_bus_reg_dataout_839_port, regs(838) => 
                           DataPath_RF_bus_reg_dataout_838_port, regs(837) => 
                           DataPath_RF_bus_reg_dataout_837_port, regs(836) => 
                           DataPath_RF_bus_reg_dataout_836_port, regs(835) => 
                           DataPath_RF_bus_reg_dataout_835_port, regs(834) => 
                           DataPath_RF_bus_reg_dataout_834_port, regs(833) => 
                           DataPath_RF_bus_reg_dataout_833_port, regs(832) => 
                           DataPath_RF_bus_reg_dataout_832_port, regs(831) => 
                           DataPath_RF_bus_reg_dataout_831_port, regs(830) => 
                           DataPath_RF_bus_reg_dataout_830_port, regs(829) => 
                           DataPath_RF_bus_reg_dataout_829_port, regs(828) => 
                           DataPath_RF_bus_reg_dataout_828_port, regs(827) => 
                           DataPath_RF_bus_reg_dataout_827_port, regs(826) => 
                           DataPath_RF_bus_reg_dataout_826_port, regs(825) => 
                           DataPath_RF_bus_reg_dataout_825_port, regs(824) => 
                           DataPath_RF_bus_reg_dataout_824_port, regs(823) => 
                           DataPath_RF_bus_reg_dataout_823_port, regs(822) => 
                           DataPath_RF_bus_reg_dataout_822_port, regs(821) => 
                           DataPath_RF_bus_reg_dataout_821_port, regs(820) => 
                           DataPath_RF_bus_reg_dataout_820_port, regs(819) => 
                           DataPath_RF_bus_reg_dataout_819_port, regs(818) => 
                           DataPath_RF_bus_reg_dataout_818_port, regs(817) => 
                           DataPath_RF_bus_reg_dataout_817_port, regs(816) => 
                           DataPath_RF_bus_reg_dataout_816_port, regs(815) => 
                           DataPath_RF_bus_reg_dataout_815_port, regs(814) => 
                           DataPath_RF_bus_reg_dataout_814_port, regs(813) => 
                           DataPath_RF_bus_reg_dataout_813_port, regs(812) => 
                           DataPath_RF_bus_reg_dataout_812_port, regs(811) => 
                           DataPath_RF_bus_reg_dataout_811_port, regs(810) => 
                           DataPath_RF_bus_reg_dataout_810_port, regs(809) => 
                           DataPath_RF_bus_reg_dataout_809_port, regs(808) => 
                           DataPath_RF_bus_reg_dataout_808_port, regs(807) => 
                           DataPath_RF_bus_reg_dataout_807_port, regs(806) => 
                           DataPath_RF_bus_reg_dataout_806_port, regs(805) => 
                           DataPath_RF_bus_reg_dataout_805_port, regs(804) => 
                           DataPath_RF_bus_reg_dataout_804_port, regs(803) => 
                           DataPath_RF_bus_reg_dataout_803_port, regs(802) => 
                           DataPath_RF_bus_reg_dataout_802_port, regs(801) => 
                           DataPath_RF_bus_reg_dataout_801_port, regs(800) => 
                           DataPath_RF_bus_reg_dataout_800_port, regs(799) => 
                           DataPath_RF_bus_reg_dataout_799_port, regs(798) => 
                           DataPath_RF_bus_reg_dataout_798_port, regs(797) => 
                           DataPath_RF_bus_reg_dataout_797_port, regs(796) => 
                           DataPath_RF_bus_reg_dataout_796_port, regs(795) => 
                           DataPath_RF_bus_reg_dataout_795_port, regs(794) => 
                           DataPath_RF_bus_reg_dataout_794_port, regs(793) => 
                           DataPath_RF_bus_reg_dataout_793_port, regs(792) => 
                           DataPath_RF_bus_reg_dataout_792_port, regs(791) => 
                           DataPath_RF_bus_reg_dataout_791_port, regs(790) => 
                           DataPath_RF_bus_reg_dataout_790_port, regs(789) => 
                           DataPath_RF_bus_reg_dataout_789_port, regs(788) => 
                           DataPath_RF_bus_reg_dataout_788_port, regs(787) => 
                           DataPath_RF_bus_reg_dataout_787_port, regs(786) => 
                           DataPath_RF_bus_reg_dataout_786_port, regs(785) => 
                           DataPath_RF_bus_reg_dataout_785_port, regs(784) => 
                           DataPath_RF_bus_reg_dataout_784_port, regs(783) => 
                           DataPath_RF_bus_reg_dataout_783_port, regs(782) => 
                           DataPath_RF_bus_reg_dataout_782_port, regs(781) => 
                           DataPath_RF_bus_reg_dataout_781_port, regs(780) => 
                           DataPath_RF_bus_reg_dataout_780_port, regs(779) => 
                           DataPath_RF_bus_reg_dataout_779_port, regs(778) => 
                           DataPath_RF_bus_reg_dataout_778_port, regs(777) => 
                           DataPath_RF_bus_reg_dataout_777_port, regs(776) => 
                           DataPath_RF_bus_reg_dataout_776_port, regs(775) => 
                           DataPath_RF_bus_reg_dataout_775_port, regs(774) => 
                           DataPath_RF_bus_reg_dataout_774_port, regs(773) => 
                           DataPath_RF_bus_reg_dataout_773_port, regs(772) => 
                           DataPath_RF_bus_reg_dataout_772_port, regs(771) => 
                           DataPath_RF_bus_reg_dataout_771_port, regs(770) => 
                           DataPath_RF_bus_reg_dataout_770_port, regs(769) => 
                           DataPath_RF_bus_reg_dataout_769_port, regs(768) => 
                           DataPath_RF_bus_reg_dataout_768_port, regs(767) => 
                           DataPath_RF_bus_reg_dataout_767_port, regs(766) => 
                           DataPath_RF_bus_reg_dataout_766_port, regs(765) => 
                           DataPath_RF_bus_reg_dataout_765_port, regs(764) => 
                           DataPath_RF_bus_reg_dataout_764_port, regs(763) => 
                           DataPath_RF_bus_reg_dataout_763_port, regs(762) => 
                           DataPath_RF_bus_reg_dataout_762_port, regs(761) => 
                           DataPath_RF_bus_reg_dataout_761_port, regs(760) => 
                           DataPath_RF_bus_reg_dataout_760_port, regs(759) => 
                           DataPath_RF_bus_reg_dataout_759_port, regs(758) => 
                           DataPath_RF_bus_reg_dataout_758_port, regs(757) => 
                           DataPath_RF_bus_reg_dataout_757_port, regs(756) => 
                           DataPath_RF_bus_reg_dataout_756_port, regs(755) => 
                           DataPath_RF_bus_reg_dataout_755_port, regs(754) => 
                           DataPath_RF_bus_reg_dataout_754_port, regs(753) => 
                           DataPath_RF_bus_reg_dataout_753_port, regs(752) => 
                           DataPath_RF_bus_reg_dataout_752_port, regs(751) => 
                           DataPath_RF_bus_reg_dataout_751_port, regs(750) => 
                           DataPath_RF_bus_reg_dataout_750_port, regs(749) => 
                           DataPath_RF_bus_reg_dataout_749_port, regs(748) => 
                           DataPath_RF_bus_reg_dataout_748_port, regs(747) => 
                           DataPath_RF_bus_reg_dataout_747_port, regs(746) => 
                           DataPath_RF_bus_reg_dataout_746_port, regs(745) => 
                           DataPath_RF_bus_reg_dataout_745_port, regs(744) => 
                           DataPath_RF_bus_reg_dataout_744_port, regs(743) => 
                           DataPath_RF_bus_reg_dataout_743_port, regs(742) => 
                           DataPath_RF_bus_reg_dataout_742_port, regs(741) => 
                           DataPath_RF_bus_reg_dataout_741_port, regs(740) => 
                           DataPath_RF_bus_reg_dataout_740_port, regs(739) => 
                           DataPath_RF_bus_reg_dataout_739_port, regs(738) => 
                           DataPath_RF_bus_reg_dataout_738_port, regs(737) => 
                           DataPath_RF_bus_reg_dataout_737_port, regs(736) => 
                           DataPath_RF_bus_reg_dataout_736_port, regs(735) => 
                           DataPath_RF_bus_reg_dataout_735_port, regs(734) => 
                           DataPath_RF_bus_reg_dataout_734_port, regs(733) => 
                           DataPath_RF_bus_reg_dataout_733_port, regs(732) => 
                           DataPath_RF_bus_reg_dataout_732_port, regs(731) => 
                           DataPath_RF_bus_reg_dataout_731_port, regs(730) => 
                           DataPath_RF_bus_reg_dataout_730_port, regs(729) => 
                           DataPath_RF_bus_reg_dataout_729_port, regs(728) => 
                           DataPath_RF_bus_reg_dataout_728_port, regs(727) => 
                           DataPath_RF_bus_reg_dataout_727_port, regs(726) => 
                           DataPath_RF_bus_reg_dataout_726_port, regs(725) => 
                           DataPath_RF_bus_reg_dataout_725_port, regs(724) => 
                           DataPath_RF_bus_reg_dataout_724_port, regs(723) => 
                           DataPath_RF_bus_reg_dataout_723_port, regs(722) => 
                           DataPath_RF_bus_reg_dataout_722_port, regs(721) => 
                           DataPath_RF_bus_reg_dataout_721_port, regs(720) => 
                           DataPath_RF_bus_reg_dataout_720_port, regs(719) => 
                           DataPath_RF_bus_reg_dataout_719_port, regs(718) => 
                           DataPath_RF_bus_reg_dataout_718_port, regs(717) => 
                           DataPath_RF_bus_reg_dataout_717_port, regs(716) => 
                           DataPath_RF_bus_reg_dataout_716_port, regs(715) => 
                           DataPath_RF_bus_reg_dataout_715_port, regs(714) => 
                           DataPath_RF_bus_reg_dataout_714_port, regs(713) => 
                           DataPath_RF_bus_reg_dataout_713_port, regs(712) => 
                           DataPath_RF_bus_reg_dataout_712_port, regs(711) => 
                           DataPath_RF_bus_reg_dataout_711_port, regs(710) => 
                           DataPath_RF_bus_reg_dataout_710_port, regs(709) => 
                           DataPath_RF_bus_reg_dataout_709_port, regs(708) => 
                           DataPath_RF_bus_reg_dataout_708_port, regs(707) => 
                           DataPath_RF_bus_reg_dataout_707_port, regs(706) => 
                           DataPath_RF_bus_reg_dataout_706_port, regs(705) => 
                           DataPath_RF_bus_reg_dataout_705_port, regs(704) => 
                           DataPath_RF_bus_reg_dataout_704_port, regs(703) => 
                           DataPath_RF_bus_reg_dataout_703_port, regs(702) => 
                           DataPath_RF_bus_reg_dataout_702_port, regs(701) => 
                           DataPath_RF_bus_reg_dataout_701_port, regs(700) => 
                           DataPath_RF_bus_reg_dataout_700_port, regs(699) => 
                           DataPath_RF_bus_reg_dataout_699_port, regs(698) => 
                           DataPath_RF_bus_reg_dataout_698_port, regs(697) => 
                           DataPath_RF_bus_reg_dataout_697_port, regs(696) => 
                           DataPath_RF_bus_reg_dataout_696_port, regs(695) => 
                           DataPath_RF_bus_reg_dataout_695_port, regs(694) => 
                           DataPath_RF_bus_reg_dataout_694_port, regs(693) => 
                           DataPath_RF_bus_reg_dataout_693_port, regs(692) => 
                           DataPath_RF_bus_reg_dataout_692_port, regs(691) => 
                           DataPath_RF_bus_reg_dataout_691_port, regs(690) => 
                           DataPath_RF_bus_reg_dataout_690_port, regs(689) => 
                           DataPath_RF_bus_reg_dataout_689_port, regs(688) => 
                           DataPath_RF_bus_reg_dataout_688_port, regs(687) => 
                           DataPath_RF_bus_reg_dataout_687_port, regs(686) => 
                           DataPath_RF_bus_reg_dataout_686_port, regs(685) => 
                           DataPath_RF_bus_reg_dataout_685_port, regs(684) => 
                           DataPath_RF_bus_reg_dataout_684_port, regs(683) => 
                           DataPath_RF_bus_reg_dataout_683_port, regs(682) => 
                           DataPath_RF_bus_reg_dataout_682_port, regs(681) => 
                           DataPath_RF_bus_reg_dataout_681_port, regs(680) => 
                           DataPath_RF_bus_reg_dataout_680_port, regs(679) => 
                           DataPath_RF_bus_reg_dataout_679_port, regs(678) => 
                           DataPath_RF_bus_reg_dataout_678_port, regs(677) => 
                           DataPath_RF_bus_reg_dataout_677_port, regs(676) => 
                           DataPath_RF_bus_reg_dataout_676_port, regs(675) => 
                           DataPath_RF_bus_reg_dataout_675_port, regs(674) => 
                           DataPath_RF_bus_reg_dataout_674_port, regs(673) => 
                           DataPath_RF_bus_reg_dataout_673_port, regs(672) => 
                           DataPath_RF_bus_reg_dataout_672_port, regs(671) => 
                           DataPath_RF_bus_reg_dataout_671_port, regs(670) => 
                           DataPath_RF_bus_reg_dataout_670_port, regs(669) => 
                           DataPath_RF_bus_reg_dataout_669_port, regs(668) => 
                           DataPath_RF_bus_reg_dataout_668_port, regs(667) => 
                           DataPath_RF_bus_reg_dataout_667_port, regs(666) => 
                           DataPath_RF_bus_reg_dataout_666_port, regs(665) => 
                           DataPath_RF_bus_reg_dataout_665_port, regs(664) => 
                           DataPath_RF_bus_reg_dataout_664_port, regs(663) => 
                           DataPath_RF_bus_reg_dataout_663_port, regs(662) => 
                           DataPath_RF_bus_reg_dataout_662_port, regs(661) => 
                           DataPath_RF_bus_reg_dataout_661_port, regs(660) => 
                           DataPath_RF_bus_reg_dataout_660_port, regs(659) => 
                           DataPath_RF_bus_reg_dataout_659_port, regs(658) => 
                           DataPath_RF_bus_reg_dataout_658_port, regs(657) => 
                           DataPath_RF_bus_reg_dataout_657_port, regs(656) => 
                           DataPath_RF_bus_reg_dataout_656_port, regs(655) => 
                           DataPath_RF_bus_reg_dataout_655_port, regs(654) => 
                           DataPath_RF_bus_reg_dataout_654_port, regs(653) => 
                           DataPath_RF_bus_reg_dataout_653_port, regs(652) => 
                           DataPath_RF_bus_reg_dataout_652_port, regs(651) => 
                           DataPath_RF_bus_reg_dataout_651_port, regs(650) => 
                           DataPath_RF_bus_reg_dataout_650_port, regs(649) => 
                           DataPath_RF_bus_reg_dataout_649_port, regs(648) => 
                           DataPath_RF_bus_reg_dataout_648_port, regs(647) => 
                           DataPath_RF_bus_reg_dataout_647_port, regs(646) => 
                           DataPath_RF_bus_reg_dataout_646_port, regs(645) => 
                           DataPath_RF_bus_reg_dataout_645_port, regs(644) => 
                           DataPath_RF_bus_reg_dataout_644_port, regs(643) => 
                           DataPath_RF_bus_reg_dataout_643_port, regs(642) => 
                           DataPath_RF_bus_reg_dataout_642_port, regs(641) => 
                           DataPath_RF_bus_reg_dataout_641_port, regs(640) => 
                           DataPath_RF_bus_reg_dataout_640_port, regs(639) => 
                           DataPath_RF_bus_reg_dataout_639_port, regs(638) => 
                           DataPath_RF_bus_reg_dataout_638_port, regs(637) => 
                           DataPath_RF_bus_reg_dataout_637_port, regs(636) => 
                           DataPath_RF_bus_reg_dataout_636_port, regs(635) => 
                           DataPath_RF_bus_reg_dataout_635_port, regs(634) => 
                           DataPath_RF_bus_reg_dataout_634_port, regs(633) => 
                           DataPath_RF_bus_reg_dataout_633_port, regs(632) => 
                           DataPath_RF_bus_reg_dataout_632_port, regs(631) => 
                           DataPath_RF_bus_reg_dataout_631_port, regs(630) => 
                           DataPath_RF_bus_reg_dataout_630_port, regs(629) => 
                           DataPath_RF_bus_reg_dataout_629_port, regs(628) => 
                           DataPath_RF_bus_reg_dataout_628_port, regs(627) => 
                           DataPath_RF_bus_reg_dataout_627_port, regs(626) => 
                           DataPath_RF_bus_reg_dataout_626_port, regs(625) => 
                           DataPath_RF_bus_reg_dataout_625_port, regs(624) => 
                           DataPath_RF_bus_reg_dataout_624_port, regs(623) => 
                           DataPath_RF_bus_reg_dataout_623_port, regs(622) => 
                           DataPath_RF_bus_reg_dataout_622_port, regs(621) => 
                           DataPath_RF_bus_reg_dataout_621_port, regs(620) => 
                           DataPath_RF_bus_reg_dataout_620_port, regs(619) => 
                           DataPath_RF_bus_reg_dataout_619_port, regs(618) => 
                           DataPath_RF_bus_reg_dataout_618_port, regs(617) => 
                           DataPath_RF_bus_reg_dataout_617_port, regs(616) => 
                           DataPath_RF_bus_reg_dataout_616_port, regs(615) => 
                           DataPath_RF_bus_reg_dataout_615_port, regs(614) => 
                           DataPath_RF_bus_reg_dataout_614_port, regs(613) => 
                           DataPath_RF_bus_reg_dataout_613_port, regs(612) => 
                           DataPath_RF_bus_reg_dataout_612_port, regs(611) => 
                           DataPath_RF_bus_reg_dataout_611_port, regs(610) => 
                           DataPath_RF_bus_reg_dataout_610_port, regs(609) => 
                           DataPath_RF_bus_reg_dataout_609_port, regs(608) => 
                           DataPath_RF_bus_reg_dataout_608_port, regs(607) => 
                           DataPath_RF_bus_reg_dataout_607_port, regs(606) => 
                           DataPath_RF_bus_reg_dataout_606_port, regs(605) => 
                           DataPath_RF_bus_reg_dataout_605_port, regs(604) => 
                           DataPath_RF_bus_reg_dataout_604_port, regs(603) => 
                           DataPath_RF_bus_reg_dataout_603_port, regs(602) => 
                           DataPath_RF_bus_reg_dataout_602_port, regs(601) => 
                           DataPath_RF_bus_reg_dataout_601_port, regs(600) => 
                           DataPath_RF_bus_reg_dataout_600_port, regs(599) => 
                           DataPath_RF_bus_reg_dataout_599_port, regs(598) => 
                           DataPath_RF_bus_reg_dataout_598_port, regs(597) => 
                           DataPath_RF_bus_reg_dataout_597_port, regs(596) => 
                           DataPath_RF_bus_reg_dataout_596_port, regs(595) => 
                           DataPath_RF_bus_reg_dataout_595_port, regs(594) => 
                           DataPath_RF_bus_reg_dataout_594_port, regs(593) => 
                           DataPath_RF_bus_reg_dataout_593_port, regs(592) => 
                           DataPath_RF_bus_reg_dataout_592_port, regs(591) => 
                           DataPath_RF_bus_reg_dataout_591_port, regs(590) => 
                           DataPath_RF_bus_reg_dataout_590_port, regs(589) => 
                           DataPath_RF_bus_reg_dataout_589_port, regs(588) => 
                           DataPath_RF_bus_reg_dataout_588_port, regs(587) => 
                           DataPath_RF_bus_reg_dataout_587_port, regs(586) => 
                           DataPath_RF_bus_reg_dataout_586_port, regs(585) => 
                           DataPath_RF_bus_reg_dataout_585_port, regs(584) => 
                           DataPath_RF_bus_reg_dataout_584_port, regs(583) => 
                           DataPath_RF_bus_reg_dataout_583_port, regs(582) => 
                           DataPath_RF_bus_reg_dataout_582_port, regs(581) => 
                           DataPath_RF_bus_reg_dataout_581_port, regs(580) => 
                           DataPath_RF_bus_reg_dataout_580_port, regs(579) => 
                           DataPath_RF_bus_reg_dataout_579_port, regs(578) => 
                           DataPath_RF_bus_reg_dataout_578_port, regs(577) => 
                           DataPath_RF_bus_reg_dataout_577_port, regs(576) => 
                           DataPath_RF_bus_reg_dataout_576_port, regs(575) => 
                           DataPath_RF_bus_reg_dataout_575_port, regs(574) => 
                           DataPath_RF_bus_reg_dataout_574_port, regs(573) => 
                           DataPath_RF_bus_reg_dataout_573_port, regs(572) => 
                           DataPath_RF_bus_reg_dataout_572_port, regs(571) => 
                           DataPath_RF_bus_reg_dataout_571_port, regs(570) => 
                           DataPath_RF_bus_reg_dataout_570_port, regs(569) => 
                           DataPath_RF_bus_reg_dataout_569_port, regs(568) => 
                           DataPath_RF_bus_reg_dataout_568_port, regs(567) => 
                           DataPath_RF_bus_reg_dataout_567_port, regs(566) => 
                           DataPath_RF_bus_reg_dataout_566_port, regs(565) => 
                           DataPath_RF_bus_reg_dataout_565_port, regs(564) => 
                           DataPath_RF_bus_reg_dataout_564_port, regs(563) => 
                           DataPath_RF_bus_reg_dataout_563_port, regs(562) => 
                           DataPath_RF_bus_reg_dataout_562_port, regs(561) => 
                           DataPath_RF_bus_reg_dataout_561_port, regs(560) => 
                           DataPath_RF_bus_reg_dataout_560_port, regs(559) => 
                           DataPath_RF_bus_reg_dataout_559_port, regs(558) => 
                           DataPath_RF_bus_reg_dataout_558_port, regs(557) => 
                           DataPath_RF_bus_reg_dataout_557_port, regs(556) => 
                           DataPath_RF_bus_reg_dataout_556_port, regs(555) => 
                           DataPath_RF_bus_reg_dataout_555_port, regs(554) => 
                           DataPath_RF_bus_reg_dataout_554_port, regs(553) => 
                           DataPath_RF_bus_reg_dataout_553_port, regs(552) => 
                           DataPath_RF_bus_reg_dataout_552_port, regs(551) => 
                           DataPath_RF_bus_reg_dataout_551_port, regs(550) => 
                           DataPath_RF_bus_reg_dataout_550_port, regs(549) => 
                           DataPath_RF_bus_reg_dataout_549_port, regs(548) => 
                           DataPath_RF_bus_reg_dataout_548_port, regs(547) => 
                           DataPath_RF_bus_reg_dataout_547_port, regs(546) => 
                           DataPath_RF_bus_reg_dataout_546_port, regs(545) => 
                           DataPath_RF_bus_reg_dataout_545_port, regs(544) => 
                           DataPath_RF_bus_reg_dataout_544_port, regs(543) => 
                           DataPath_RF_bus_reg_dataout_543_port, regs(542) => 
                           DataPath_RF_bus_reg_dataout_542_port, regs(541) => 
                           DataPath_RF_bus_reg_dataout_541_port, regs(540) => 
                           DataPath_RF_bus_reg_dataout_540_port, regs(539) => 
                           DataPath_RF_bus_reg_dataout_539_port, regs(538) => 
                           DataPath_RF_bus_reg_dataout_538_port, regs(537) => 
                           DataPath_RF_bus_reg_dataout_537_port, regs(536) => 
                           DataPath_RF_bus_reg_dataout_536_port, regs(535) => 
                           DataPath_RF_bus_reg_dataout_535_port, regs(534) => 
                           DataPath_RF_bus_reg_dataout_534_port, regs(533) => 
                           DataPath_RF_bus_reg_dataout_533_port, regs(532) => 
                           DataPath_RF_bus_reg_dataout_532_port, regs(531) => 
                           DataPath_RF_bus_reg_dataout_531_port, regs(530) => 
                           DataPath_RF_bus_reg_dataout_530_port, regs(529) => 
                           DataPath_RF_bus_reg_dataout_529_port, regs(528) => 
                           DataPath_RF_bus_reg_dataout_528_port, regs(527) => 
                           DataPath_RF_bus_reg_dataout_527_port, regs(526) => 
                           DataPath_RF_bus_reg_dataout_526_port, regs(525) => 
                           DataPath_RF_bus_reg_dataout_525_port, regs(524) => 
                           DataPath_RF_bus_reg_dataout_524_port, regs(523) => 
                           DataPath_RF_bus_reg_dataout_523_port, regs(522) => 
                           DataPath_RF_bus_reg_dataout_522_port, regs(521) => 
                           DataPath_RF_bus_reg_dataout_521_port, regs(520) => 
                           DataPath_RF_bus_reg_dataout_520_port, regs(519) => 
                           DataPath_RF_bus_reg_dataout_519_port, regs(518) => 
                           DataPath_RF_bus_reg_dataout_518_port, regs(517) => 
                           DataPath_RF_bus_reg_dataout_517_port, regs(516) => 
                           DataPath_RF_bus_reg_dataout_516_port, regs(515) => 
                           DataPath_RF_bus_reg_dataout_515_port, regs(514) => 
                           DataPath_RF_bus_reg_dataout_514_port, regs(513) => 
                           DataPath_RF_bus_reg_dataout_513_port, regs(512) => 
                           DataPath_RF_bus_reg_dataout_512_port, regs(511) => 
                           DataPath_RF_bus_reg_dataout_511_port, regs(510) => 
                           DataPath_RF_bus_reg_dataout_510_port, regs(509) => 
                           DataPath_RF_bus_reg_dataout_509_port, regs(508) => 
                           DataPath_RF_bus_reg_dataout_508_port, regs(507) => 
                           DataPath_RF_bus_reg_dataout_507_port, regs(506) => 
                           DataPath_RF_bus_reg_dataout_506_port, regs(505) => 
                           DataPath_RF_bus_reg_dataout_505_port, regs(504) => 
                           DataPath_RF_bus_reg_dataout_504_port, regs(503) => 
                           DataPath_RF_bus_reg_dataout_503_port, regs(502) => 
                           DataPath_RF_bus_reg_dataout_502_port, regs(501) => 
                           DataPath_RF_bus_reg_dataout_501_port, regs(500) => 
                           DataPath_RF_bus_reg_dataout_500_port, regs(499) => 
                           DataPath_RF_bus_reg_dataout_499_port, regs(498) => 
                           DataPath_RF_bus_reg_dataout_498_port, regs(497) => 
                           DataPath_RF_bus_reg_dataout_497_port, regs(496) => 
                           DataPath_RF_bus_reg_dataout_496_port, regs(495) => 
                           DataPath_RF_bus_reg_dataout_495_port, regs(494) => 
                           DataPath_RF_bus_reg_dataout_494_port, regs(493) => 
                           DataPath_RF_bus_reg_dataout_493_port, regs(492) => 
                           DataPath_RF_bus_reg_dataout_492_port, regs(491) => 
                           DataPath_RF_bus_reg_dataout_491_port, regs(490) => 
                           DataPath_RF_bus_reg_dataout_490_port, regs(489) => 
                           DataPath_RF_bus_reg_dataout_489_port, regs(488) => 
                           DataPath_RF_bus_reg_dataout_488_port, regs(487) => 
                           DataPath_RF_bus_reg_dataout_487_port, regs(486) => 
                           DataPath_RF_bus_reg_dataout_486_port, regs(485) => 
                           DataPath_RF_bus_reg_dataout_485_port, regs(484) => 
                           DataPath_RF_bus_reg_dataout_484_port, regs(483) => 
                           DataPath_RF_bus_reg_dataout_483_port, regs(482) => 
                           DataPath_RF_bus_reg_dataout_482_port, regs(481) => 
                           DataPath_RF_bus_reg_dataout_481_port, regs(480) => 
                           DataPath_RF_bus_reg_dataout_480_port, regs(479) => 
                           DataPath_RF_bus_reg_dataout_479_port, regs(478) => 
                           DataPath_RF_bus_reg_dataout_478_port, regs(477) => 
                           DataPath_RF_bus_reg_dataout_477_port, regs(476) => 
                           DataPath_RF_bus_reg_dataout_476_port, regs(475) => 
                           DataPath_RF_bus_reg_dataout_475_port, regs(474) => 
                           DataPath_RF_bus_reg_dataout_474_port, regs(473) => 
                           DataPath_RF_bus_reg_dataout_473_port, regs(472) => 
                           DataPath_RF_bus_reg_dataout_472_port, regs(471) => 
                           DataPath_RF_bus_reg_dataout_471_port, regs(470) => 
                           DataPath_RF_bus_reg_dataout_470_port, regs(469) => 
                           DataPath_RF_bus_reg_dataout_469_port, regs(468) => 
                           DataPath_RF_bus_reg_dataout_468_port, regs(467) => 
                           DataPath_RF_bus_reg_dataout_467_port, regs(466) => 
                           DataPath_RF_bus_reg_dataout_466_port, regs(465) => 
                           DataPath_RF_bus_reg_dataout_465_port, regs(464) => 
                           DataPath_RF_bus_reg_dataout_464_port, regs(463) => 
                           DataPath_RF_bus_reg_dataout_463_port, regs(462) => 
                           DataPath_RF_bus_reg_dataout_462_port, regs(461) => 
                           DataPath_RF_bus_reg_dataout_461_port, regs(460) => 
                           DataPath_RF_bus_reg_dataout_460_port, regs(459) => 
                           DataPath_RF_bus_reg_dataout_459_port, regs(458) => 
                           DataPath_RF_bus_reg_dataout_458_port, regs(457) => 
                           DataPath_RF_bus_reg_dataout_457_port, regs(456) => 
                           DataPath_RF_bus_reg_dataout_456_port, regs(455) => 
                           DataPath_RF_bus_reg_dataout_455_port, regs(454) => 
                           DataPath_RF_bus_reg_dataout_454_port, regs(453) => 
                           DataPath_RF_bus_reg_dataout_453_port, regs(452) => 
                           DataPath_RF_bus_reg_dataout_452_port, regs(451) => 
                           DataPath_RF_bus_reg_dataout_451_port, regs(450) => 
                           DataPath_RF_bus_reg_dataout_450_port, regs(449) => 
                           DataPath_RF_bus_reg_dataout_449_port, regs(448) => 
                           DataPath_RF_bus_reg_dataout_448_port, regs(447) => 
                           DataPath_RF_bus_reg_dataout_447_port, regs(446) => 
                           DataPath_RF_bus_reg_dataout_446_port, regs(445) => 
                           DataPath_RF_bus_reg_dataout_445_port, regs(444) => 
                           DataPath_RF_bus_reg_dataout_444_port, regs(443) => 
                           DataPath_RF_bus_reg_dataout_443_port, regs(442) => 
                           DataPath_RF_bus_reg_dataout_442_port, regs(441) => 
                           DataPath_RF_bus_reg_dataout_441_port, regs(440) => 
                           DataPath_RF_bus_reg_dataout_440_port, regs(439) => 
                           DataPath_RF_bus_reg_dataout_439_port, regs(438) => 
                           DataPath_RF_bus_reg_dataout_438_port, regs(437) => 
                           DataPath_RF_bus_reg_dataout_437_port, regs(436) => 
                           DataPath_RF_bus_reg_dataout_436_port, regs(435) => 
                           DataPath_RF_bus_reg_dataout_435_port, regs(434) => 
                           DataPath_RF_bus_reg_dataout_434_port, regs(433) => 
                           DataPath_RF_bus_reg_dataout_433_port, regs(432) => 
                           DataPath_RF_bus_reg_dataout_432_port, regs(431) => 
                           DataPath_RF_bus_reg_dataout_431_port, regs(430) => 
                           DataPath_RF_bus_reg_dataout_430_port, regs(429) => 
                           DataPath_RF_bus_reg_dataout_429_port, regs(428) => 
                           DataPath_RF_bus_reg_dataout_428_port, regs(427) => 
                           DataPath_RF_bus_reg_dataout_427_port, regs(426) => 
                           DataPath_RF_bus_reg_dataout_426_port, regs(425) => 
                           DataPath_RF_bus_reg_dataout_425_port, regs(424) => 
                           DataPath_RF_bus_reg_dataout_424_port, regs(423) => 
                           DataPath_RF_bus_reg_dataout_423_port, regs(422) => 
                           DataPath_RF_bus_reg_dataout_422_port, regs(421) => 
                           DataPath_RF_bus_reg_dataout_421_port, regs(420) => 
                           DataPath_RF_bus_reg_dataout_420_port, regs(419) => 
                           DataPath_RF_bus_reg_dataout_419_port, regs(418) => 
                           DataPath_RF_bus_reg_dataout_418_port, regs(417) => 
                           DataPath_RF_bus_reg_dataout_417_port, regs(416) => 
                           DataPath_RF_bus_reg_dataout_416_port, regs(415) => 
                           DataPath_RF_bus_reg_dataout_415_port, regs(414) => 
                           DataPath_RF_bus_reg_dataout_414_port, regs(413) => 
                           DataPath_RF_bus_reg_dataout_413_port, regs(412) => 
                           DataPath_RF_bus_reg_dataout_412_port, regs(411) => 
                           DataPath_RF_bus_reg_dataout_411_port, regs(410) => 
                           DataPath_RF_bus_reg_dataout_410_port, regs(409) => 
                           DataPath_RF_bus_reg_dataout_409_port, regs(408) => 
                           DataPath_RF_bus_reg_dataout_408_port, regs(407) => 
                           DataPath_RF_bus_reg_dataout_407_port, regs(406) => 
                           DataPath_RF_bus_reg_dataout_406_port, regs(405) => 
                           DataPath_RF_bus_reg_dataout_405_port, regs(404) => 
                           DataPath_RF_bus_reg_dataout_404_port, regs(403) => 
                           DataPath_RF_bus_reg_dataout_403_port, regs(402) => 
                           DataPath_RF_bus_reg_dataout_402_port, regs(401) => 
                           DataPath_RF_bus_reg_dataout_401_port, regs(400) => 
                           DataPath_RF_bus_reg_dataout_400_port, regs(399) => 
                           DataPath_RF_bus_reg_dataout_399_port, regs(398) => 
                           DataPath_RF_bus_reg_dataout_398_port, regs(397) => 
                           DataPath_RF_bus_reg_dataout_397_port, regs(396) => 
                           DataPath_RF_bus_reg_dataout_396_port, regs(395) => 
                           DataPath_RF_bus_reg_dataout_395_port, regs(394) => 
                           DataPath_RF_bus_reg_dataout_394_port, regs(393) => 
                           DataPath_RF_bus_reg_dataout_393_port, regs(392) => 
                           DataPath_RF_bus_reg_dataout_392_port, regs(391) => 
                           DataPath_RF_bus_reg_dataout_391_port, regs(390) => 
                           DataPath_RF_bus_reg_dataout_390_port, regs(389) => 
                           DataPath_RF_bus_reg_dataout_389_port, regs(388) => 
                           DataPath_RF_bus_reg_dataout_388_port, regs(387) => 
                           DataPath_RF_bus_reg_dataout_387_port, regs(386) => 
                           DataPath_RF_bus_reg_dataout_386_port, regs(385) => 
                           DataPath_RF_bus_reg_dataout_385_port, regs(384) => 
                           DataPath_RF_bus_reg_dataout_384_port, regs(383) => 
                           DataPath_RF_bus_reg_dataout_383_port, regs(382) => 
                           DataPath_RF_bus_reg_dataout_382_port, regs(381) => 
                           DataPath_RF_bus_reg_dataout_381_port, regs(380) => 
                           DataPath_RF_bus_reg_dataout_380_port, regs(379) => 
                           DataPath_RF_bus_reg_dataout_379_port, regs(378) => 
                           DataPath_RF_bus_reg_dataout_378_port, regs(377) => 
                           DataPath_RF_bus_reg_dataout_377_port, regs(376) => 
                           DataPath_RF_bus_reg_dataout_376_port, regs(375) => 
                           DataPath_RF_bus_reg_dataout_375_port, regs(374) => 
                           DataPath_RF_bus_reg_dataout_374_port, regs(373) => 
                           DataPath_RF_bus_reg_dataout_373_port, regs(372) => 
                           DataPath_RF_bus_reg_dataout_372_port, regs(371) => 
                           DataPath_RF_bus_reg_dataout_371_port, regs(370) => 
                           DataPath_RF_bus_reg_dataout_370_port, regs(369) => 
                           DataPath_RF_bus_reg_dataout_369_port, regs(368) => 
                           DataPath_RF_bus_reg_dataout_368_port, regs(367) => 
                           DataPath_RF_bus_reg_dataout_367_port, regs(366) => 
                           DataPath_RF_bus_reg_dataout_366_port, regs(365) => 
                           DataPath_RF_bus_reg_dataout_365_port, regs(364) => 
                           DataPath_RF_bus_reg_dataout_364_port, regs(363) => 
                           DataPath_RF_bus_reg_dataout_363_port, regs(362) => 
                           DataPath_RF_bus_reg_dataout_362_port, regs(361) => 
                           DataPath_RF_bus_reg_dataout_361_port, regs(360) => 
                           DataPath_RF_bus_reg_dataout_360_port, regs(359) => 
                           DataPath_RF_bus_reg_dataout_359_port, regs(358) => 
                           DataPath_RF_bus_reg_dataout_358_port, regs(357) => 
                           DataPath_RF_bus_reg_dataout_357_port, regs(356) => 
                           DataPath_RF_bus_reg_dataout_356_port, regs(355) => 
                           DataPath_RF_bus_reg_dataout_355_port, regs(354) => 
                           DataPath_RF_bus_reg_dataout_354_port, regs(353) => 
                           DataPath_RF_bus_reg_dataout_353_port, regs(352) => 
                           DataPath_RF_bus_reg_dataout_352_port, regs(351) => 
                           DataPath_RF_bus_reg_dataout_351_port, regs(350) => 
                           DataPath_RF_bus_reg_dataout_350_port, regs(349) => 
                           DataPath_RF_bus_reg_dataout_349_port, regs(348) => 
                           DataPath_RF_bus_reg_dataout_348_port, regs(347) => 
                           DataPath_RF_bus_reg_dataout_347_port, regs(346) => 
                           DataPath_RF_bus_reg_dataout_346_port, regs(345) => 
                           DataPath_RF_bus_reg_dataout_345_port, regs(344) => 
                           DataPath_RF_bus_reg_dataout_344_port, regs(343) => 
                           DataPath_RF_bus_reg_dataout_343_port, regs(342) => 
                           DataPath_RF_bus_reg_dataout_342_port, regs(341) => 
                           DataPath_RF_bus_reg_dataout_341_port, regs(340) => 
                           DataPath_RF_bus_reg_dataout_340_port, regs(339) => 
                           DataPath_RF_bus_reg_dataout_339_port, regs(338) => 
                           DataPath_RF_bus_reg_dataout_338_port, regs(337) => 
                           DataPath_RF_bus_reg_dataout_337_port, regs(336) => 
                           DataPath_RF_bus_reg_dataout_336_port, regs(335) => 
                           DataPath_RF_bus_reg_dataout_335_port, regs(334) => 
                           DataPath_RF_bus_reg_dataout_334_port, regs(333) => 
                           DataPath_RF_bus_reg_dataout_333_port, regs(332) => 
                           DataPath_RF_bus_reg_dataout_332_port, regs(331) => 
                           DataPath_RF_bus_reg_dataout_331_port, regs(330) => 
                           DataPath_RF_bus_reg_dataout_330_port, regs(329) => 
                           DataPath_RF_bus_reg_dataout_329_port, regs(328) => 
                           DataPath_RF_bus_reg_dataout_328_port, regs(327) => 
                           DataPath_RF_bus_reg_dataout_327_port, regs(326) => 
                           DataPath_RF_bus_reg_dataout_326_port, regs(325) => 
                           DataPath_RF_bus_reg_dataout_325_port, regs(324) => 
                           DataPath_RF_bus_reg_dataout_324_port, regs(323) => 
                           DataPath_RF_bus_reg_dataout_323_port, regs(322) => 
                           DataPath_RF_bus_reg_dataout_322_port, regs(321) => 
                           DataPath_RF_bus_reg_dataout_321_port, regs(320) => 
                           DataPath_RF_bus_reg_dataout_320_port, regs(319) => 
                           DataPath_RF_bus_reg_dataout_319_port, regs(318) => 
                           DataPath_RF_bus_reg_dataout_318_port, regs(317) => 
                           DataPath_RF_bus_reg_dataout_317_port, regs(316) => 
                           DataPath_RF_bus_reg_dataout_316_port, regs(315) => 
                           DataPath_RF_bus_reg_dataout_315_port, regs(314) => 
                           DataPath_RF_bus_reg_dataout_314_port, regs(313) => 
                           DataPath_RF_bus_reg_dataout_313_port, regs(312) => 
                           DataPath_RF_bus_reg_dataout_312_port, regs(311) => 
                           DataPath_RF_bus_reg_dataout_311_port, regs(310) => 
                           DataPath_RF_bus_reg_dataout_310_port, regs(309) => 
                           DataPath_RF_bus_reg_dataout_309_port, regs(308) => 
                           DataPath_RF_bus_reg_dataout_308_port, regs(307) => 
                           DataPath_RF_bus_reg_dataout_307_port, regs(306) => 
                           DataPath_RF_bus_reg_dataout_306_port, regs(305) => 
                           DataPath_RF_bus_reg_dataout_305_port, regs(304) => 
                           DataPath_RF_bus_reg_dataout_304_port, regs(303) => 
                           DataPath_RF_bus_reg_dataout_303_port, regs(302) => 
                           DataPath_RF_bus_reg_dataout_302_port, regs(301) => 
                           DataPath_RF_bus_reg_dataout_301_port, regs(300) => 
                           DataPath_RF_bus_reg_dataout_300_port, regs(299) => 
                           DataPath_RF_bus_reg_dataout_299_port, regs(298) => 
                           DataPath_RF_bus_reg_dataout_298_port, regs(297) => 
                           DataPath_RF_bus_reg_dataout_297_port, regs(296) => 
                           DataPath_RF_bus_reg_dataout_296_port, regs(295) => 
                           DataPath_RF_bus_reg_dataout_295_port, regs(294) => 
                           DataPath_RF_bus_reg_dataout_294_port, regs(293) => 
                           DataPath_RF_bus_reg_dataout_293_port, regs(292) => 
                           DataPath_RF_bus_reg_dataout_292_port, regs(291) => 
                           DataPath_RF_bus_reg_dataout_291_port, regs(290) => 
                           DataPath_RF_bus_reg_dataout_290_port, regs(289) => 
                           DataPath_RF_bus_reg_dataout_289_port, regs(288) => 
                           DataPath_RF_bus_reg_dataout_288_port, regs(287) => 
                           DataPath_RF_bus_reg_dataout_287_port, regs(286) => 
                           DataPath_RF_bus_reg_dataout_286_port, regs(285) => 
                           DataPath_RF_bus_reg_dataout_285_port, regs(284) => 
                           DataPath_RF_bus_reg_dataout_284_port, regs(283) => 
                           DataPath_RF_bus_reg_dataout_283_port, regs(282) => 
                           DataPath_RF_bus_reg_dataout_282_port, regs(281) => 
                           DataPath_RF_bus_reg_dataout_281_port, regs(280) => 
                           DataPath_RF_bus_reg_dataout_280_port, regs(279) => 
                           DataPath_RF_bus_reg_dataout_279_port, regs(278) => 
                           DataPath_RF_bus_reg_dataout_278_port, regs(277) => 
                           DataPath_RF_bus_reg_dataout_277_port, regs(276) => 
                           DataPath_RF_bus_reg_dataout_276_port, regs(275) => 
                           DataPath_RF_bus_reg_dataout_275_port, regs(274) => 
                           DataPath_RF_bus_reg_dataout_274_port, regs(273) => 
                           DataPath_RF_bus_reg_dataout_273_port, regs(272) => 
                           DataPath_RF_bus_reg_dataout_272_port, regs(271) => 
                           DataPath_RF_bus_reg_dataout_271_port, regs(270) => 
                           DataPath_RF_bus_reg_dataout_270_port, regs(269) => 
                           DataPath_RF_bus_reg_dataout_269_port, regs(268) => 
                           DataPath_RF_bus_reg_dataout_268_port, regs(267) => 
                           DataPath_RF_bus_reg_dataout_267_port, regs(266) => 
                           DataPath_RF_bus_reg_dataout_266_port, regs(265) => 
                           DataPath_RF_bus_reg_dataout_265_port, regs(264) => 
                           DataPath_RF_bus_reg_dataout_264_port, regs(263) => 
                           DataPath_RF_bus_reg_dataout_263_port, regs(262) => 
                           DataPath_RF_bus_reg_dataout_262_port, regs(261) => 
                           DataPath_RF_bus_reg_dataout_261_port, regs(260) => 
                           DataPath_RF_bus_reg_dataout_260_port, regs(259) => 
                           DataPath_RF_bus_reg_dataout_259_port, regs(258) => 
                           DataPath_RF_bus_reg_dataout_258_port, regs(257) => 
                           DataPath_RF_bus_reg_dataout_257_port, regs(256) => 
                           DataPath_RF_bus_reg_dataout_256_port, regs(255) => 
                           DataPath_RF_bus_reg_dataout_255_port, regs(254) => 
                           DataPath_RF_bus_reg_dataout_254_port, regs(253) => 
                           DataPath_RF_bus_reg_dataout_253_port, regs(252) => 
                           DataPath_RF_bus_reg_dataout_252_port, regs(251) => 
                           DataPath_RF_bus_reg_dataout_251_port, regs(250) => 
                           DataPath_RF_bus_reg_dataout_250_port, regs(249) => 
                           DataPath_RF_bus_reg_dataout_249_port, regs(248) => 
                           DataPath_RF_bus_reg_dataout_248_port, regs(247) => 
                           DataPath_RF_bus_reg_dataout_247_port, regs(246) => 
                           DataPath_RF_bus_reg_dataout_246_port, regs(245) => 
                           DataPath_RF_bus_reg_dataout_245_port, regs(244) => 
                           DataPath_RF_bus_reg_dataout_244_port, regs(243) => 
                           DataPath_RF_bus_reg_dataout_243_port, regs(242) => 
                           DataPath_RF_bus_reg_dataout_242_port, regs(241) => 
                           DataPath_RF_bus_reg_dataout_241_port, regs(240) => 
                           DataPath_RF_bus_reg_dataout_240_port, regs(239) => 
                           DataPath_RF_bus_reg_dataout_239_port, regs(238) => 
                           DataPath_RF_bus_reg_dataout_238_port, regs(237) => 
                           DataPath_RF_bus_reg_dataout_237_port, regs(236) => 
                           DataPath_RF_bus_reg_dataout_236_port, regs(235) => 
                           DataPath_RF_bus_reg_dataout_235_port, regs(234) => 
                           DataPath_RF_bus_reg_dataout_234_port, regs(233) => 
                           DataPath_RF_bus_reg_dataout_233_port, regs(232) => 
                           DataPath_RF_bus_reg_dataout_232_port, regs(231) => 
                           DataPath_RF_bus_reg_dataout_231_port, regs(230) => 
                           DataPath_RF_bus_reg_dataout_230_port, regs(229) => 
                           DataPath_RF_bus_reg_dataout_229_port, regs(228) => 
                           DataPath_RF_bus_reg_dataout_228_port, regs(227) => 
                           DataPath_RF_bus_reg_dataout_227_port, regs(226) => 
                           DataPath_RF_bus_reg_dataout_226_port, regs(225) => 
                           DataPath_RF_bus_reg_dataout_225_port, regs(224) => 
                           DataPath_RF_bus_reg_dataout_224_port, regs(223) => 
                           DataPath_RF_bus_reg_dataout_223_port, regs(222) => 
                           DataPath_RF_bus_reg_dataout_222_port, regs(221) => 
                           DataPath_RF_bus_reg_dataout_221_port, regs(220) => 
                           DataPath_RF_bus_reg_dataout_220_port, regs(219) => 
                           DataPath_RF_bus_reg_dataout_219_port, regs(218) => 
                           DataPath_RF_bus_reg_dataout_218_port, regs(217) => 
                           DataPath_RF_bus_reg_dataout_217_port, regs(216) => 
                           DataPath_RF_bus_reg_dataout_216_port, regs(215) => 
                           DataPath_RF_bus_reg_dataout_215_port, regs(214) => 
                           DataPath_RF_bus_reg_dataout_214_port, regs(213) => 
                           DataPath_RF_bus_reg_dataout_213_port, regs(212) => 
                           DataPath_RF_bus_reg_dataout_212_port, regs(211) => 
                           DataPath_RF_bus_reg_dataout_211_port, regs(210) => 
                           DataPath_RF_bus_reg_dataout_210_port, regs(209) => 
                           DataPath_RF_bus_reg_dataout_209_port, regs(208) => 
                           DataPath_RF_bus_reg_dataout_208_port, regs(207) => 
                           DataPath_RF_bus_reg_dataout_207_port, regs(206) => 
                           DataPath_RF_bus_reg_dataout_206_port, regs(205) => 
                           DataPath_RF_bus_reg_dataout_205_port, regs(204) => 
                           DataPath_RF_bus_reg_dataout_204_port, regs(203) => 
                           DataPath_RF_bus_reg_dataout_203_port, regs(202) => 
                           DataPath_RF_bus_reg_dataout_202_port, regs(201) => 
                           DataPath_RF_bus_reg_dataout_201_port, regs(200) => 
                           DataPath_RF_bus_reg_dataout_200_port, regs(199) => 
                           DataPath_RF_bus_reg_dataout_199_port, regs(198) => 
                           DataPath_RF_bus_reg_dataout_198_port, regs(197) => 
                           DataPath_RF_bus_reg_dataout_197_port, regs(196) => 
                           DataPath_RF_bus_reg_dataout_196_port, regs(195) => 
                           DataPath_RF_bus_reg_dataout_195_port, regs(194) => 
                           DataPath_RF_bus_reg_dataout_194_port, regs(193) => 
                           DataPath_RF_bus_reg_dataout_193_port, regs(192) => 
                           DataPath_RF_bus_reg_dataout_192_port, regs(191) => 
                           DataPath_RF_bus_reg_dataout_191_port, regs(190) => 
                           DataPath_RF_bus_reg_dataout_190_port, regs(189) => 
                           DataPath_RF_bus_reg_dataout_189_port, regs(188) => 
                           DataPath_RF_bus_reg_dataout_188_port, regs(187) => 
                           DataPath_RF_bus_reg_dataout_187_port, regs(186) => 
                           DataPath_RF_bus_reg_dataout_186_port, regs(185) => 
                           DataPath_RF_bus_reg_dataout_185_port, regs(184) => 
                           DataPath_RF_bus_reg_dataout_184_port, regs(183) => 
                           DataPath_RF_bus_reg_dataout_183_port, regs(182) => 
                           DataPath_RF_bus_reg_dataout_182_port, regs(181) => 
                           DataPath_RF_bus_reg_dataout_181_port, regs(180) => 
                           DataPath_RF_bus_reg_dataout_180_port, regs(179) => 
                           DataPath_RF_bus_reg_dataout_179_port, regs(178) => 
                           DataPath_RF_bus_reg_dataout_178_port, regs(177) => 
                           DataPath_RF_bus_reg_dataout_177_port, regs(176) => 
                           DataPath_RF_bus_reg_dataout_176_port, regs(175) => 
                           DataPath_RF_bus_reg_dataout_175_port, regs(174) => 
                           DataPath_RF_bus_reg_dataout_174_port, regs(173) => 
                           DataPath_RF_bus_reg_dataout_173_port, regs(172) => 
                           DataPath_RF_bus_reg_dataout_172_port, regs(171) => 
                           DataPath_RF_bus_reg_dataout_171_port, regs(170) => 
                           DataPath_RF_bus_reg_dataout_170_port, regs(169) => 
                           DataPath_RF_bus_reg_dataout_169_port, regs(168) => 
                           DataPath_RF_bus_reg_dataout_168_port, regs(167) => 
                           DataPath_RF_bus_reg_dataout_167_port, regs(166) => 
                           DataPath_RF_bus_reg_dataout_166_port, regs(165) => 
                           DataPath_RF_bus_reg_dataout_165_port, regs(164) => 
                           DataPath_RF_bus_reg_dataout_164_port, regs(163) => 
                           DataPath_RF_bus_reg_dataout_163_port, regs(162) => 
                           DataPath_RF_bus_reg_dataout_162_port, regs(161) => 
                           DataPath_RF_bus_reg_dataout_161_port, regs(160) => 
                           DataPath_RF_bus_reg_dataout_160_port, regs(159) => 
                           DataPath_RF_bus_reg_dataout_159_port, regs(158) => 
                           DataPath_RF_bus_reg_dataout_158_port, regs(157) => 
                           DataPath_RF_bus_reg_dataout_157_port, regs(156) => 
                           DataPath_RF_bus_reg_dataout_156_port, regs(155) => 
                           DataPath_RF_bus_reg_dataout_155_port, regs(154) => 
                           DataPath_RF_bus_reg_dataout_154_port, regs(153) => 
                           DataPath_RF_bus_reg_dataout_153_port, regs(152) => 
                           DataPath_RF_bus_reg_dataout_152_port, regs(151) => 
                           DataPath_RF_bus_reg_dataout_151_port, regs(150) => 
                           DataPath_RF_bus_reg_dataout_150_port, regs(149) => 
                           DataPath_RF_bus_reg_dataout_149_port, regs(148) => 
                           DataPath_RF_bus_reg_dataout_148_port, regs(147) => 
                           DataPath_RF_bus_reg_dataout_147_port, regs(146) => 
                           DataPath_RF_bus_reg_dataout_146_port, regs(145) => 
                           DataPath_RF_bus_reg_dataout_145_port, regs(144) => 
                           DataPath_RF_bus_reg_dataout_144_port, regs(143) => 
                           DataPath_RF_bus_reg_dataout_143_port, regs(142) => 
                           DataPath_RF_bus_reg_dataout_142_port, regs(141) => 
                           DataPath_RF_bus_reg_dataout_141_port, regs(140) => 
                           DataPath_RF_bus_reg_dataout_140_port, regs(139) => 
                           DataPath_RF_bus_reg_dataout_139_port, regs(138) => 
                           DataPath_RF_bus_reg_dataout_138_port, regs(137) => 
                           DataPath_RF_bus_reg_dataout_137_port, regs(136) => 
                           DataPath_RF_bus_reg_dataout_136_port, regs(135) => 
                           DataPath_RF_bus_reg_dataout_135_port, regs(134) => 
                           DataPath_RF_bus_reg_dataout_134_port, regs(133) => 
                           DataPath_RF_bus_reg_dataout_133_port, regs(132) => 
                           DataPath_RF_bus_reg_dataout_132_port, regs(131) => 
                           DataPath_RF_bus_reg_dataout_131_port, regs(130) => 
                           DataPath_RF_bus_reg_dataout_130_port, regs(129) => 
                           DataPath_RF_bus_reg_dataout_129_port, regs(128) => 
                           DataPath_RF_bus_reg_dataout_128_port, regs(127) => 
                           DataPath_RF_bus_reg_dataout_127_port, regs(126) => 
                           DataPath_RF_bus_reg_dataout_126_port, regs(125) => 
                           DataPath_RF_bus_reg_dataout_125_port, regs(124) => 
                           DataPath_RF_bus_reg_dataout_124_port, regs(123) => 
                           DataPath_RF_bus_reg_dataout_123_port, regs(122) => 
                           DataPath_RF_bus_reg_dataout_122_port, regs(121) => 
                           DataPath_RF_bus_reg_dataout_121_port, regs(120) => 
                           DataPath_RF_bus_reg_dataout_120_port, regs(119) => 
                           DataPath_RF_bus_reg_dataout_119_port, regs(118) => 
                           DataPath_RF_bus_reg_dataout_118_port, regs(117) => 
                           DataPath_RF_bus_reg_dataout_117_port, regs(116) => 
                           DataPath_RF_bus_reg_dataout_116_port, regs(115) => 
                           DataPath_RF_bus_reg_dataout_115_port, regs(114) => 
                           DataPath_RF_bus_reg_dataout_114_port, regs(113) => 
                           DataPath_RF_bus_reg_dataout_113_port, regs(112) => 
                           DataPath_RF_bus_reg_dataout_112_port, regs(111) => 
                           DataPath_RF_bus_reg_dataout_111_port, regs(110) => 
                           DataPath_RF_bus_reg_dataout_110_port, regs(109) => 
                           DataPath_RF_bus_reg_dataout_109_port, regs(108) => 
                           DataPath_RF_bus_reg_dataout_108_port, regs(107) => 
                           DataPath_RF_bus_reg_dataout_107_port, regs(106) => 
                           DataPath_RF_bus_reg_dataout_106_port, regs(105) => 
                           DataPath_RF_bus_reg_dataout_105_port, regs(104) => 
                           DataPath_RF_bus_reg_dataout_104_port, regs(103) => 
                           DataPath_RF_bus_reg_dataout_103_port, regs(102) => 
                           DataPath_RF_bus_reg_dataout_102_port, regs(101) => 
                           DataPath_RF_bus_reg_dataout_101_port, regs(100) => 
                           DataPath_RF_bus_reg_dataout_100_port, regs(99) => 
                           DataPath_RF_bus_reg_dataout_99_port, regs(98) => 
                           DataPath_RF_bus_reg_dataout_98_port, regs(97) => 
                           DataPath_RF_bus_reg_dataout_97_port, regs(96) => 
                           DataPath_RF_bus_reg_dataout_96_port, regs(95) => 
                           DataPath_RF_bus_reg_dataout_95_port, regs(94) => 
                           DataPath_RF_bus_reg_dataout_94_port, regs(93) => 
                           DataPath_RF_bus_reg_dataout_93_port, regs(92) => 
                           DataPath_RF_bus_reg_dataout_92_port, regs(91) => 
                           DataPath_RF_bus_reg_dataout_91_port, regs(90) => 
                           DataPath_RF_bus_reg_dataout_90_port, regs(89) => 
                           DataPath_RF_bus_reg_dataout_89_port, regs(88) => 
                           DataPath_RF_bus_reg_dataout_88_port, regs(87) => 
                           DataPath_RF_bus_reg_dataout_87_port, regs(86) => 
                           DataPath_RF_bus_reg_dataout_86_port, regs(85) => 
                           DataPath_RF_bus_reg_dataout_85_port, regs(84) => 
                           DataPath_RF_bus_reg_dataout_84_port, regs(83) => 
                           DataPath_RF_bus_reg_dataout_83_port, regs(82) => 
                           DataPath_RF_bus_reg_dataout_82_port, regs(81) => 
                           DataPath_RF_bus_reg_dataout_81_port, regs(80) => 
                           DataPath_RF_bus_reg_dataout_80_port, regs(79) => 
                           DataPath_RF_bus_reg_dataout_79_port, regs(78) => 
                           DataPath_RF_bus_reg_dataout_78_port, regs(77) => 
                           DataPath_RF_bus_reg_dataout_77_port, regs(76) => 
                           DataPath_RF_bus_reg_dataout_76_port, regs(75) => 
                           DataPath_RF_bus_reg_dataout_75_port, regs(74) => 
                           DataPath_RF_bus_reg_dataout_74_port, regs(73) => 
                           DataPath_RF_bus_reg_dataout_73_port, regs(72) => 
                           DataPath_RF_bus_reg_dataout_72_port, regs(71) => 
                           DataPath_RF_bus_reg_dataout_71_port, regs(70) => 
                           DataPath_RF_bus_reg_dataout_70_port, regs(69) => 
                           DataPath_RF_bus_reg_dataout_69_port, regs(68) => 
                           DataPath_RF_bus_reg_dataout_68_port, regs(67) => 
                           DataPath_RF_bus_reg_dataout_67_port, regs(66) => 
                           DataPath_RF_bus_reg_dataout_66_port, regs(65) => 
                           DataPath_RF_bus_reg_dataout_65_port, regs(64) => 
                           DataPath_RF_bus_reg_dataout_64_port, regs(63) => 
                           DataPath_RF_bus_reg_dataout_63_port, regs(62) => 
                           DataPath_RF_bus_reg_dataout_62_port, regs(61) => 
                           DataPath_RF_bus_reg_dataout_61_port, regs(60) => 
                           DataPath_RF_bus_reg_dataout_60_port, regs(59) => 
                           DataPath_RF_bus_reg_dataout_59_port, regs(58) => 
                           DataPath_RF_bus_reg_dataout_58_port, regs(57) => 
                           DataPath_RF_bus_reg_dataout_57_port, regs(56) => 
                           DataPath_RF_bus_reg_dataout_56_port, regs(55) => 
                           DataPath_RF_bus_reg_dataout_55_port, regs(54) => 
                           DataPath_RF_bus_reg_dataout_54_port, regs(53) => 
                           DataPath_RF_bus_reg_dataout_53_port, regs(52) => 
                           DataPath_RF_bus_reg_dataout_52_port, regs(51) => 
                           DataPath_RF_bus_reg_dataout_51_port, regs(50) => 
                           DataPath_RF_bus_reg_dataout_50_port, regs(49) => 
                           DataPath_RF_bus_reg_dataout_49_port, regs(48) => 
                           DataPath_RF_bus_reg_dataout_48_port, regs(47) => 
                           DataPath_RF_bus_reg_dataout_47_port, regs(46) => 
                           DataPath_RF_bus_reg_dataout_46_port, regs(45) => 
                           DataPath_RF_bus_reg_dataout_45_port, regs(44) => 
                           DataPath_RF_bus_reg_dataout_44_port, regs(43) => 
                           DataPath_RF_bus_reg_dataout_43_port, regs(42) => 
                           DataPath_RF_bus_reg_dataout_42_port, regs(41) => 
                           DataPath_RF_bus_reg_dataout_41_port, regs(40) => 
                           DataPath_RF_bus_reg_dataout_40_port, regs(39) => 
                           DataPath_RF_bus_reg_dataout_39_port, regs(38) => 
                           DataPath_RF_bus_reg_dataout_38_port, regs(37) => 
                           DataPath_RF_bus_reg_dataout_37_port, regs(36) => 
                           DataPath_RF_bus_reg_dataout_36_port, regs(35) => 
                           DataPath_RF_bus_reg_dataout_35_port, regs(34) => 
                           DataPath_RF_bus_reg_dataout_34_port, regs(33) => 
                           DataPath_RF_bus_reg_dataout_33_port, regs(32) => 
                           DataPath_RF_bus_reg_dataout_32_port, regs(31) => 
                           DataPath_RF_bus_reg_dataout_31_port, regs(30) => 
                           DataPath_RF_bus_reg_dataout_30_port, regs(29) => 
                           DataPath_RF_bus_reg_dataout_29_port, regs(28) => 
                           DataPath_RF_bus_reg_dataout_28_port, regs(27) => 
                           DataPath_RF_bus_reg_dataout_27_port, regs(26) => 
                           DataPath_RF_bus_reg_dataout_26_port, regs(25) => 
                           DataPath_RF_bus_reg_dataout_25_port, regs(24) => 
                           DataPath_RF_bus_reg_dataout_24_port, regs(23) => 
                           DataPath_RF_bus_reg_dataout_23_port, regs(22) => 
                           DataPath_RF_bus_reg_dataout_22_port, regs(21) => 
                           DataPath_RF_bus_reg_dataout_21_port, regs(20) => 
                           DataPath_RF_bus_reg_dataout_20_port, regs(19) => 
                           DataPath_RF_bus_reg_dataout_19_port, regs(18) => 
                           DataPath_RF_bus_reg_dataout_18_port, regs(17) => 
                           DataPath_RF_bus_reg_dataout_17_port, regs(16) => 
                           DataPath_RF_bus_reg_dataout_16_port, regs(15) => 
                           DataPath_RF_bus_reg_dataout_15_port, regs(14) => 
                           DataPath_RF_bus_reg_dataout_14_port, regs(13) => 
                           DataPath_RF_bus_reg_dataout_13_port, regs(12) => 
                           DataPath_RF_bus_reg_dataout_12_port, regs(11) => 
                           DataPath_RF_bus_reg_dataout_11_port, regs(10) => 
                           DataPath_RF_bus_reg_dataout_10_port, regs(9) => 
                           DataPath_RF_bus_reg_dataout_9_port, regs(8) => 
                           DataPath_RF_bus_reg_dataout_8_port, regs(7) => 
                           DataPath_RF_bus_reg_dataout_7_port, regs(6) => 
                           DataPath_RF_bus_reg_dataout_6_port, regs(5) => 
                           DataPath_RF_bus_reg_dataout_5_port, regs(4) => 
                           DataPath_RF_bus_reg_dataout_4_port, regs(3) => 
                           DataPath_RF_bus_reg_dataout_3_port, regs(2) => 
                           DataPath_RF_bus_reg_dataout_2_port, regs(1) => 
                           DataPath_RF_bus_reg_dataout_1_port, regs(0) => 
                           DataPath_RF_bus_reg_dataout_0_port, win(4) => n8678,
                           win(3) => DataPath_RF_c_win_3_port, win(2) => 
                           DataPath_RF_c_win_2_port, win(1) => 
                           DataPath_RF_c_win_1_port, win(0) => 
                           DataPath_RF_c_win_0_port, curr_proc_regs(767) => 
                           DataPath_RF_bus_selected_win_data_767_port, 
                           curr_proc_regs(766) => 
                           DataPath_RF_bus_selected_win_data_766_port, 
                           curr_proc_regs(765) => 
                           DataPath_RF_bus_selected_win_data_765_port, 
                           curr_proc_regs(764) => 
                           DataPath_RF_bus_selected_win_data_764_port, 
                           curr_proc_regs(763) => 
                           DataPath_RF_bus_selected_win_data_763_port, 
                           curr_proc_regs(762) => 
                           DataPath_RF_bus_selected_win_data_762_port, 
                           curr_proc_regs(761) => 
                           DataPath_RF_bus_selected_win_data_761_port, 
                           curr_proc_regs(760) => 
                           DataPath_RF_bus_selected_win_data_760_port, 
                           curr_proc_regs(759) => 
                           DataPath_RF_bus_selected_win_data_759_port, 
                           curr_proc_regs(758) => 
                           DataPath_RF_bus_selected_win_data_758_port, 
                           curr_proc_regs(757) => 
                           DataPath_RF_bus_selected_win_data_757_port, 
                           curr_proc_regs(756) => 
                           DataPath_RF_bus_selected_win_data_756_port, 
                           curr_proc_regs(755) => 
                           DataPath_RF_bus_selected_win_data_755_port, 
                           curr_proc_regs(754) => 
                           DataPath_RF_bus_selected_win_data_754_port, 
                           curr_proc_regs(753) => 
                           DataPath_RF_bus_selected_win_data_753_port, 
                           curr_proc_regs(752) => 
                           DataPath_RF_bus_selected_win_data_752_port, 
                           curr_proc_regs(751) => 
                           DataPath_RF_bus_selected_win_data_751_port, 
                           curr_proc_regs(750) => 
                           DataPath_RF_bus_selected_win_data_750_port, 
                           curr_proc_regs(749) => 
                           DataPath_RF_bus_selected_win_data_749_port, 
                           curr_proc_regs(748) => 
                           DataPath_RF_bus_selected_win_data_748_port, 
                           curr_proc_regs(747) => 
                           DataPath_RF_bus_selected_win_data_747_port, 
                           curr_proc_regs(746) => 
                           DataPath_RF_bus_selected_win_data_746_port, 
                           curr_proc_regs(745) => 
                           DataPath_RF_bus_selected_win_data_745_port, 
                           curr_proc_regs(744) => 
                           DataPath_RF_bus_selected_win_data_744_port, 
                           curr_proc_regs(743) => 
                           DataPath_RF_bus_selected_win_data_743_port, 
                           curr_proc_regs(742) => 
                           DataPath_RF_bus_selected_win_data_742_port, 
                           curr_proc_regs(741) => 
                           DataPath_RF_bus_selected_win_data_741_port, 
                           curr_proc_regs(740) => 
                           DataPath_RF_bus_selected_win_data_740_port, 
                           curr_proc_regs(739) => 
                           DataPath_RF_bus_selected_win_data_739_port, 
                           curr_proc_regs(738) => 
                           DataPath_RF_bus_selected_win_data_738_port, 
                           curr_proc_regs(737) => 
                           DataPath_RF_bus_selected_win_data_737_port, 
                           curr_proc_regs(736) => 
                           DataPath_RF_bus_selected_win_data_736_port, 
                           curr_proc_regs(735) => 
                           DataPath_RF_bus_selected_win_data_735_port, 
                           curr_proc_regs(734) => 
                           DataPath_RF_bus_selected_win_data_734_port, 
                           curr_proc_regs(733) => 
                           DataPath_RF_bus_selected_win_data_733_port, 
                           curr_proc_regs(732) => 
                           DataPath_RF_bus_selected_win_data_732_port, 
                           curr_proc_regs(731) => 
                           DataPath_RF_bus_selected_win_data_731_port, 
                           curr_proc_regs(730) => 
                           DataPath_RF_bus_selected_win_data_730_port, 
                           curr_proc_regs(729) => 
                           DataPath_RF_bus_selected_win_data_729_port, 
                           curr_proc_regs(728) => 
                           DataPath_RF_bus_selected_win_data_728_port, 
                           curr_proc_regs(727) => 
                           DataPath_RF_bus_selected_win_data_727_port, 
                           curr_proc_regs(726) => 
                           DataPath_RF_bus_selected_win_data_726_port, 
                           curr_proc_regs(725) => 
                           DataPath_RF_bus_selected_win_data_725_port, 
                           curr_proc_regs(724) => 
                           DataPath_RF_bus_selected_win_data_724_port, 
                           curr_proc_regs(723) => 
                           DataPath_RF_bus_selected_win_data_723_port, 
                           curr_proc_regs(722) => 
                           DataPath_RF_bus_selected_win_data_722_port, 
                           curr_proc_regs(721) => 
                           DataPath_RF_bus_selected_win_data_721_port, 
                           curr_proc_regs(720) => 
                           DataPath_RF_bus_selected_win_data_720_port, 
                           curr_proc_regs(719) => 
                           DataPath_RF_bus_selected_win_data_719_port, 
                           curr_proc_regs(718) => 
                           DataPath_RF_bus_selected_win_data_718_port, 
                           curr_proc_regs(717) => 
                           DataPath_RF_bus_selected_win_data_717_port, 
                           curr_proc_regs(716) => 
                           DataPath_RF_bus_selected_win_data_716_port, 
                           curr_proc_regs(715) => 
                           DataPath_RF_bus_selected_win_data_715_port, 
                           curr_proc_regs(714) => 
                           DataPath_RF_bus_selected_win_data_714_port, 
                           curr_proc_regs(713) => 
                           DataPath_RF_bus_selected_win_data_713_port, 
                           curr_proc_regs(712) => 
                           DataPath_RF_bus_selected_win_data_712_port, 
                           curr_proc_regs(711) => 
                           DataPath_RF_bus_selected_win_data_711_port, 
                           curr_proc_regs(710) => 
                           DataPath_RF_bus_selected_win_data_710_port, 
                           curr_proc_regs(709) => 
                           DataPath_RF_bus_selected_win_data_709_port, 
                           curr_proc_regs(708) => 
                           DataPath_RF_bus_selected_win_data_708_port, 
                           curr_proc_regs(707) => 
                           DataPath_RF_bus_selected_win_data_707_port, 
                           curr_proc_regs(706) => 
                           DataPath_RF_bus_selected_win_data_706_port, 
                           curr_proc_regs(705) => 
                           DataPath_RF_bus_selected_win_data_705_port, 
                           curr_proc_regs(704) => 
                           DataPath_RF_bus_selected_win_data_704_port, 
                           curr_proc_regs(703) => 
                           DataPath_RF_bus_selected_win_data_703_port, 
                           curr_proc_regs(702) => 
                           DataPath_RF_bus_selected_win_data_702_port, 
                           curr_proc_regs(701) => 
                           DataPath_RF_bus_selected_win_data_701_port, 
                           curr_proc_regs(700) => 
                           DataPath_RF_bus_selected_win_data_700_port, 
                           curr_proc_regs(699) => 
                           DataPath_RF_bus_selected_win_data_699_port, 
                           curr_proc_regs(698) => 
                           DataPath_RF_bus_selected_win_data_698_port, 
                           curr_proc_regs(697) => 
                           DataPath_RF_bus_selected_win_data_697_port, 
                           curr_proc_regs(696) => 
                           DataPath_RF_bus_selected_win_data_696_port, 
                           curr_proc_regs(695) => 
                           DataPath_RF_bus_selected_win_data_695_port, 
                           curr_proc_regs(694) => 
                           DataPath_RF_bus_selected_win_data_694_port, 
                           curr_proc_regs(693) => 
                           DataPath_RF_bus_selected_win_data_693_port, 
                           curr_proc_regs(692) => 
                           DataPath_RF_bus_selected_win_data_692_port, 
                           curr_proc_regs(691) => 
                           DataPath_RF_bus_selected_win_data_691_port, 
                           curr_proc_regs(690) => 
                           DataPath_RF_bus_selected_win_data_690_port, 
                           curr_proc_regs(689) => 
                           DataPath_RF_bus_selected_win_data_689_port, 
                           curr_proc_regs(688) => 
                           DataPath_RF_bus_selected_win_data_688_port, 
                           curr_proc_regs(687) => 
                           DataPath_RF_bus_selected_win_data_687_port, 
                           curr_proc_regs(686) => 
                           DataPath_RF_bus_selected_win_data_686_port, 
                           curr_proc_regs(685) => 
                           DataPath_RF_bus_selected_win_data_685_port, 
                           curr_proc_regs(684) => 
                           DataPath_RF_bus_selected_win_data_684_port, 
                           curr_proc_regs(683) => 
                           DataPath_RF_bus_selected_win_data_683_port, 
                           curr_proc_regs(682) => 
                           DataPath_RF_bus_selected_win_data_682_port, 
                           curr_proc_regs(681) => 
                           DataPath_RF_bus_selected_win_data_681_port, 
                           curr_proc_regs(680) => 
                           DataPath_RF_bus_selected_win_data_680_port, 
                           curr_proc_regs(679) => 
                           DataPath_RF_bus_selected_win_data_679_port, 
                           curr_proc_regs(678) => 
                           DataPath_RF_bus_selected_win_data_678_port, 
                           curr_proc_regs(677) => 
                           DataPath_RF_bus_selected_win_data_677_port, 
                           curr_proc_regs(676) => 
                           DataPath_RF_bus_selected_win_data_676_port, 
                           curr_proc_regs(675) => 
                           DataPath_RF_bus_selected_win_data_675_port, 
                           curr_proc_regs(674) => 
                           DataPath_RF_bus_selected_win_data_674_port, 
                           curr_proc_regs(673) => 
                           DataPath_RF_bus_selected_win_data_673_port, 
                           curr_proc_regs(672) => 
                           DataPath_RF_bus_selected_win_data_672_port, 
                           curr_proc_regs(671) => 
                           DataPath_RF_bus_selected_win_data_671_port, 
                           curr_proc_regs(670) => 
                           DataPath_RF_bus_selected_win_data_670_port, 
                           curr_proc_regs(669) => 
                           DataPath_RF_bus_selected_win_data_669_port, 
                           curr_proc_regs(668) => 
                           DataPath_RF_bus_selected_win_data_668_port, 
                           curr_proc_regs(667) => 
                           DataPath_RF_bus_selected_win_data_667_port, 
                           curr_proc_regs(666) => 
                           DataPath_RF_bus_selected_win_data_666_port, 
                           curr_proc_regs(665) => 
                           DataPath_RF_bus_selected_win_data_665_port, 
                           curr_proc_regs(664) => 
                           DataPath_RF_bus_selected_win_data_664_port, 
                           curr_proc_regs(663) => 
                           DataPath_RF_bus_selected_win_data_663_port, 
                           curr_proc_regs(662) => 
                           DataPath_RF_bus_selected_win_data_662_port, 
                           curr_proc_regs(661) => 
                           DataPath_RF_bus_selected_win_data_661_port, 
                           curr_proc_regs(660) => 
                           DataPath_RF_bus_selected_win_data_660_port, 
                           curr_proc_regs(659) => 
                           DataPath_RF_bus_selected_win_data_659_port, 
                           curr_proc_regs(658) => 
                           DataPath_RF_bus_selected_win_data_658_port, 
                           curr_proc_regs(657) => 
                           DataPath_RF_bus_selected_win_data_657_port, 
                           curr_proc_regs(656) => 
                           DataPath_RF_bus_selected_win_data_656_port, 
                           curr_proc_regs(655) => 
                           DataPath_RF_bus_selected_win_data_655_port, 
                           curr_proc_regs(654) => 
                           DataPath_RF_bus_selected_win_data_654_port, 
                           curr_proc_regs(653) => 
                           DataPath_RF_bus_selected_win_data_653_port, 
                           curr_proc_regs(652) => 
                           DataPath_RF_bus_selected_win_data_652_port, 
                           curr_proc_regs(651) => 
                           DataPath_RF_bus_selected_win_data_651_port, 
                           curr_proc_regs(650) => 
                           DataPath_RF_bus_selected_win_data_650_port, 
                           curr_proc_regs(649) => 
                           DataPath_RF_bus_selected_win_data_649_port, 
                           curr_proc_regs(648) => 
                           DataPath_RF_bus_selected_win_data_648_port, 
                           curr_proc_regs(647) => 
                           DataPath_RF_bus_selected_win_data_647_port, 
                           curr_proc_regs(646) => 
                           DataPath_RF_bus_selected_win_data_646_port, 
                           curr_proc_regs(645) => 
                           DataPath_RF_bus_selected_win_data_645_port, 
                           curr_proc_regs(644) => 
                           DataPath_RF_bus_selected_win_data_644_port, 
                           curr_proc_regs(643) => 
                           DataPath_RF_bus_selected_win_data_643_port, 
                           curr_proc_regs(642) => 
                           DataPath_RF_bus_selected_win_data_642_port, 
                           curr_proc_regs(641) => 
                           DataPath_RF_bus_selected_win_data_641_port, 
                           curr_proc_regs(640) => 
                           DataPath_RF_bus_selected_win_data_640_port, 
                           curr_proc_regs(639) => 
                           DataPath_RF_bus_selected_win_data_639_port, 
                           curr_proc_regs(638) => 
                           DataPath_RF_bus_selected_win_data_638_port, 
                           curr_proc_regs(637) => 
                           DataPath_RF_bus_selected_win_data_637_port, 
                           curr_proc_regs(636) => 
                           DataPath_RF_bus_selected_win_data_636_port, 
                           curr_proc_regs(635) => 
                           DataPath_RF_bus_selected_win_data_635_port, 
                           curr_proc_regs(634) => 
                           DataPath_RF_bus_selected_win_data_634_port, 
                           curr_proc_regs(633) => 
                           DataPath_RF_bus_selected_win_data_633_port, 
                           curr_proc_regs(632) => 
                           DataPath_RF_bus_selected_win_data_632_port, 
                           curr_proc_regs(631) => 
                           DataPath_RF_bus_selected_win_data_631_port, 
                           curr_proc_regs(630) => 
                           DataPath_RF_bus_selected_win_data_630_port, 
                           curr_proc_regs(629) => 
                           DataPath_RF_bus_selected_win_data_629_port, 
                           curr_proc_regs(628) => 
                           DataPath_RF_bus_selected_win_data_628_port, 
                           curr_proc_regs(627) => 
                           DataPath_RF_bus_selected_win_data_627_port, 
                           curr_proc_regs(626) => 
                           DataPath_RF_bus_selected_win_data_626_port, 
                           curr_proc_regs(625) => 
                           DataPath_RF_bus_selected_win_data_625_port, 
                           curr_proc_regs(624) => 
                           DataPath_RF_bus_selected_win_data_624_port, 
                           curr_proc_regs(623) => 
                           DataPath_RF_bus_selected_win_data_623_port, 
                           curr_proc_regs(622) => 
                           DataPath_RF_bus_selected_win_data_622_port, 
                           curr_proc_regs(621) => 
                           DataPath_RF_bus_selected_win_data_621_port, 
                           curr_proc_regs(620) => 
                           DataPath_RF_bus_selected_win_data_620_port, 
                           curr_proc_regs(619) => 
                           DataPath_RF_bus_selected_win_data_619_port, 
                           curr_proc_regs(618) => 
                           DataPath_RF_bus_selected_win_data_618_port, 
                           curr_proc_regs(617) => 
                           DataPath_RF_bus_selected_win_data_617_port, 
                           curr_proc_regs(616) => 
                           DataPath_RF_bus_selected_win_data_616_port, 
                           curr_proc_regs(615) => 
                           DataPath_RF_bus_selected_win_data_615_port, 
                           curr_proc_regs(614) => 
                           DataPath_RF_bus_selected_win_data_614_port, 
                           curr_proc_regs(613) => 
                           DataPath_RF_bus_selected_win_data_613_port, 
                           curr_proc_regs(612) => 
                           DataPath_RF_bus_selected_win_data_612_port, 
                           curr_proc_regs(611) => 
                           DataPath_RF_bus_selected_win_data_611_port, 
                           curr_proc_regs(610) => 
                           DataPath_RF_bus_selected_win_data_610_port, 
                           curr_proc_regs(609) => 
                           DataPath_RF_bus_selected_win_data_609_port, 
                           curr_proc_regs(608) => 
                           DataPath_RF_bus_selected_win_data_608_port, 
                           curr_proc_regs(607) => 
                           DataPath_RF_bus_selected_win_data_607_port, 
                           curr_proc_regs(606) => 
                           DataPath_RF_bus_selected_win_data_606_port, 
                           curr_proc_regs(605) => 
                           DataPath_RF_bus_selected_win_data_605_port, 
                           curr_proc_regs(604) => 
                           DataPath_RF_bus_selected_win_data_604_port, 
                           curr_proc_regs(603) => 
                           DataPath_RF_bus_selected_win_data_603_port, 
                           curr_proc_regs(602) => 
                           DataPath_RF_bus_selected_win_data_602_port, 
                           curr_proc_regs(601) => 
                           DataPath_RF_bus_selected_win_data_601_port, 
                           curr_proc_regs(600) => 
                           DataPath_RF_bus_selected_win_data_600_port, 
                           curr_proc_regs(599) => 
                           DataPath_RF_bus_selected_win_data_599_port, 
                           curr_proc_regs(598) => 
                           DataPath_RF_bus_selected_win_data_598_port, 
                           curr_proc_regs(597) => 
                           DataPath_RF_bus_selected_win_data_597_port, 
                           curr_proc_regs(596) => 
                           DataPath_RF_bus_selected_win_data_596_port, 
                           curr_proc_regs(595) => 
                           DataPath_RF_bus_selected_win_data_595_port, 
                           curr_proc_regs(594) => 
                           DataPath_RF_bus_selected_win_data_594_port, 
                           curr_proc_regs(593) => 
                           DataPath_RF_bus_selected_win_data_593_port, 
                           curr_proc_regs(592) => 
                           DataPath_RF_bus_selected_win_data_592_port, 
                           curr_proc_regs(591) => 
                           DataPath_RF_bus_selected_win_data_591_port, 
                           curr_proc_regs(590) => 
                           DataPath_RF_bus_selected_win_data_590_port, 
                           curr_proc_regs(589) => 
                           DataPath_RF_bus_selected_win_data_589_port, 
                           curr_proc_regs(588) => 
                           DataPath_RF_bus_selected_win_data_588_port, 
                           curr_proc_regs(587) => 
                           DataPath_RF_bus_selected_win_data_587_port, 
                           curr_proc_regs(586) => 
                           DataPath_RF_bus_selected_win_data_586_port, 
                           curr_proc_regs(585) => 
                           DataPath_RF_bus_selected_win_data_585_port, 
                           curr_proc_regs(584) => 
                           DataPath_RF_bus_selected_win_data_584_port, 
                           curr_proc_regs(583) => 
                           DataPath_RF_bus_selected_win_data_583_port, 
                           curr_proc_regs(582) => 
                           DataPath_RF_bus_selected_win_data_582_port, 
                           curr_proc_regs(581) => 
                           DataPath_RF_bus_selected_win_data_581_port, 
                           curr_proc_regs(580) => 
                           DataPath_RF_bus_selected_win_data_580_port, 
                           curr_proc_regs(579) => 
                           DataPath_RF_bus_selected_win_data_579_port, 
                           curr_proc_regs(578) => 
                           DataPath_RF_bus_selected_win_data_578_port, 
                           curr_proc_regs(577) => 
                           DataPath_RF_bus_selected_win_data_577_port, 
                           curr_proc_regs(576) => 
                           DataPath_RF_bus_selected_win_data_576_port, 
                           curr_proc_regs(575) => 
                           DataPath_RF_bus_selected_win_data_575_port, 
                           curr_proc_regs(574) => 
                           DataPath_RF_bus_selected_win_data_574_port, 
                           curr_proc_regs(573) => 
                           DataPath_RF_bus_selected_win_data_573_port, 
                           curr_proc_regs(572) => 
                           DataPath_RF_bus_selected_win_data_572_port, 
                           curr_proc_regs(571) => 
                           DataPath_RF_bus_selected_win_data_571_port, 
                           curr_proc_regs(570) => 
                           DataPath_RF_bus_selected_win_data_570_port, 
                           curr_proc_regs(569) => 
                           DataPath_RF_bus_selected_win_data_569_port, 
                           curr_proc_regs(568) => 
                           DataPath_RF_bus_selected_win_data_568_port, 
                           curr_proc_regs(567) => 
                           DataPath_RF_bus_selected_win_data_567_port, 
                           curr_proc_regs(566) => 
                           DataPath_RF_bus_selected_win_data_566_port, 
                           curr_proc_regs(565) => 
                           DataPath_RF_bus_selected_win_data_565_port, 
                           curr_proc_regs(564) => 
                           DataPath_RF_bus_selected_win_data_564_port, 
                           curr_proc_regs(563) => 
                           DataPath_RF_bus_selected_win_data_563_port, 
                           curr_proc_regs(562) => 
                           DataPath_RF_bus_selected_win_data_562_port, 
                           curr_proc_regs(561) => 
                           DataPath_RF_bus_selected_win_data_561_port, 
                           curr_proc_regs(560) => 
                           DataPath_RF_bus_selected_win_data_560_port, 
                           curr_proc_regs(559) => 
                           DataPath_RF_bus_selected_win_data_559_port, 
                           curr_proc_regs(558) => 
                           DataPath_RF_bus_selected_win_data_558_port, 
                           curr_proc_regs(557) => 
                           DataPath_RF_bus_selected_win_data_557_port, 
                           curr_proc_regs(556) => 
                           DataPath_RF_bus_selected_win_data_556_port, 
                           curr_proc_regs(555) => 
                           DataPath_RF_bus_selected_win_data_555_port, 
                           curr_proc_regs(554) => 
                           DataPath_RF_bus_selected_win_data_554_port, 
                           curr_proc_regs(553) => 
                           DataPath_RF_bus_selected_win_data_553_port, 
                           curr_proc_regs(552) => 
                           DataPath_RF_bus_selected_win_data_552_port, 
                           curr_proc_regs(551) => 
                           DataPath_RF_bus_selected_win_data_551_port, 
                           curr_proc_regs(550) => 
                           DataPath_RF_bus_selected_win_data_550_port, 
                           curr_proc_regs(549) => 
                           DataPath_RF_bus_selected_win_data_549_port, 
                           curr_proc_regs(548) => 
                           DataPath_RF_bus_selected_win_data_548_port, 
                           curr_proc_regs(547) => 
                           DataPath_RF_bus_selected_win_data_547_port, 
                           curr_proc_regs(546) => 
                           DataPath_RF_bus_selected_win_data_546_port, 
                           curr_proc_regs(545) => 
                           DataPath_RF_bus_selected_win_data_545_port, 
                           curr_proc_regs(544) => 
                           DataPath_RF_bus_selected_win_data_544_port, 
                           curr_proc_regs(543) => 
                           DataPath_RF_bus_selected_win_data_543_port, 
                           curr_proc_regs(542) => 
                           DataPath_RF_bus_selected_win_data_542_port, 
                           curr_proc_regs(541) => 
                           DataPath_RF_bus_selected_win_data_541_port, 
                           curr_proc_regs(540) => 
                           DataPath_RF_bus_selected_win_data_540_port, 
                           curr_proc_regs(539) => 
                           DataPath_RF_bus_selected_win_data_539_port, 
                           curr_proc_regs(538) => 
                           DataPath_RF_bus_selected_win_data_538_port, 
                           curr_proc_regs(537) => 
                           DataPath_RF_bus_selected_win_data_537_port, 
                           curr_proc_regs(536) => 
                           DataPath_RF_bus_selected_win_data_536_port, 
                           curr_proc_regs(535) => 
                           DataPath_RF_bus_selected_win_data_535_port, 
                           curr_proc_regs(534) => 
                           DataPath_RF_bus_selected_win_data_534_port, 
                           curr_proc_regs(533) => 
                           DataPath_RF_bus_selected_win_data_533_port, 
                           curr_proc_regs(532) => 
                           DataPath_RF_bus_selected_win_data_532_port, 
                           curr_proc_regs(531) => 
                           DataPath_RF_bus_selected_win_data_531_port, 
                           curr_proc_regs(530) => 
                           DataPath_RF_bus_selected_win_data_530_port, 
                           curr_proc_regs(529) => 
                           DataPath_RF_bus_selected_win_data_529_port, 
                           curr_proc_regs(528) => 
                           DataPath_RF_bus_selected_win_data_528_port, 
                           curr_proc_regs(527) => 
                           DataPath_RF_bus_selected_win_data_527_port, 
                           curr_proc_regs(526) => 
                           DataPath_RF_bus_selected_win_data_526_port, 
                           curr_proc_regs(525) => 
                           DataPath_RF_bus_selected_win_data_525_port, 
                           curr_proc_regs(524) => 
                           DataPath_RF_bus_selected_win_data_524_port, 
                           curr_proc_regs(523) => 
                           DataPath_RF_bus_selected_win_data_523_port, 
                           curr_proc_regs(522) => 
                           DataPath_RF_bus_selected_win_data_522_port, 
                           curr_proc_regs(521) => 
                           DataPath_RF_bus_selected_win_data_521_port, 
                           curr_proc_regs(520) => 
                           DataPath_RF_bus_selected_win_data_520_port, 
                           curr_proc_regs(519) => 
                           DataPath_RF_bus_selected_win_data_519_port, 
                           curr_proc_regs(518) => 
                           DataPath_RF_bus_selected_win_data_518_port, 
                           curr_proc_regs(517) => 
                           DataPath_RF_bus_selected_win_data_517_port, 
                           curr_proc_regs(516) => 
                           DataPath_RF_bus_selected_win_data_516_port, 
                           curr_proc_regs(515) => 
                           DataPath_RF_bus_selected_win_data_515_port, 
                           curr_proc_regs(514) => 
                           DataPath_RF_bus_selected_win_data_514_port, 
                           curr_proc_regs(513) => 
                           DataPath_RF_bus_selected_win_data_513_port, 
                           curr_proc_regs(512) => 
                           DataPath_RF_bus_selected_win_data_512_port, 
                           curr_proc_regs(511) => 
                           DataPath_RF_bus_selected_win_data_511_port, 
                           curr_proc_regs(510) => 
                           DataPath_RF_bus_selected_win_data_510_port, 
                           curr_proc_regs(509) => 
                           DataPath_RF_bus_selected_win_data_509_port, 
                           curr_proc_regs(508) => 
                           DataPath_RF_bus_selected_win_data_508_port, 
                           curr_proc_regs(507) => 
                           DataPath_RF_bus_selected_win_data_507_port, 
                           curr_proc_regs(506) => 
                           DataPath_RF_bus_selected_win_data_506_port, 
                           curr_proc_regs(505) => 
                           DataPath_RF_bus_selected_win_data_505_port, 
                           curr_proc_regs(504) => 
                           DataPath_RF_bus_selected_win_data_504_port, 
                           curr_proc_regs(503) => 
                           DataPath_RF_bus_selected_win_data_503_port, 
                           curr_proc_regs(502) => 
                           DataPath_RF_bus_selected_win_data_502_port, 
                           curr_proc_regs(501) => 
                           DataPath_RF_bus_selected_win_data_501_port, 
                           curr_proc_regs(500) => 
                           DataPath_RF_bus_selected_win_data_500_port, 
                           curr_proc_regs(499) => 
                           DataPath_RF_bus_selected_win_data_499_port, 
                           curr_proc_regs(498) => 
                           DataPath_RF_bus_selected_win_data_498_port, 
                           curr_proc_regs(497) => 
                           DataPath_RF_bus_selected_win_data_497_port, 
                           curr_proc_regs(496) => 
                           DataPath_RF_bus_selected_win_data_496_port, 
                           curr_proc_regs(495) => 
                           DataPath_RF_bus_selected_win_data_495_port, 
                           curr_proc_regs(494) => 
                           DataPath_RF_bus_selected_win_data_494_port, 
                           curr_proc_regs(493) => 
                           DataPath_RF_bus_selected_win_data_493_port, 
                           curr_proc_regs(492) => 
                           DataPath_RF_bus_selected_win_data_492_port, 
                           curr_proc_regs(491) => 
                           DataPath_RF_bus_selected_win_data_491_port, 
                           curr_proc_regs(490) => 
                           DataPath_RF_bus_selected_win_data_490_port, 
                           curr_proc_regs(489) => 
                           DataPath_RF_bus_selected_win_data_489_port, 
                           curr_proc_regs(488) => 
                           DataPath_RF_bus_selected_win_data_488_port, 
                           curr_proc_regs(487) => 
                           DataPath_RF_bus_selected_win_data_487_port, 
                           curr_proc_regs(486) => 
                           DataPath_RF_bus_selected_win_data_486_port, 
                           curr_proc_regs(485) => 
                           DataPath_RF_bus_selected_win_data_485_port, 
                           curr_proc_regs(484) => 
                           DataPath_RF_bus_selected_win_data_484_port, 
                           curr_proc_regs(483) => 
                           DataPath_RF_bus_selected_win_data_483_port, 
                           curr_proc_regs(482) => 
                           DataPath_RF_bus_selected_win_data_482_port, 
                           curr_proc_regs(481) => 
                           DataPath_RF_bus_selected_win_data_481_port, 
                           curr_proc_regs(480) => 
                           DataPath_RF_bus_selected_win_data_480_port, 
                           curr_proc_regs(479) => 
                           DataPath_RF_bus_selected_win_data_479_port, 
                           curr_proc_regs(478) => 
                           DataPath_RF_bus_selected_win_data_478_port, 
                           curr_proc_regs(477) => 
                           DataPath_RF_bus_selected_win_data_477_port, 
                           curr_proc_regs(476) => 
                           DataPath_RF_bus_selected_win_data_476_port, 
                           curr_proc_regs(475) => 
                           DataPath_RF_bus_selected_win_data_475_port, 
                           curr_proc_regs(474) => 
                           DataPath_RF_bus_selected_win_data_474_port, 
                           curr_proc_regs(473) => 
                           DataPath_RF_bus_selected_win_data_473_port, 
                           curr_proc_regs(472) => 
                           DataPath_RF_bus_selected_win_data_472_port, 
                           curr_proc_regs(471) => 
                           DataPath_RF_bus_selected_win_data_471_port, 
                           curr_proc_regs(470) => 
                           DataPath_RF_bus_selected_win_data_470_port, 
                           curr_proc_regs(469) => 
                           DataPath_RF_bus_selected_win_data_469_port, 
                           curr_proc_regs(468) => 
                           DataPath_RF_bus_selected_win_data_468_port, 
                           curr_proc_regs(467) => 
                           DataPath_RF_bus_selected_win_data_467_port, 
                           curr_proc_regs(466) => 
                           DataPath_RF_bus_selected_win_data_466_port, 
                           curr_proc_regs(465) => 
                           DataPath_RF_bus_selected_win_data_465_port, 
                           curr_proc_regs(464) => 
                           DataPath_RF_bus_selected_win_data_464_port, 
                           curr_proc_regs(463) => 
                           DataPath_RF_bus_selected_win_data_463_port, 
                           curr_proc_regs(462) => 
                           DataPath_RF_bus_selected_win_data_462_port, 
                           curr_proc_regs(461) => 
                           DataPath_RF_bus_selected_win_data_461_port, 
                           curr_proc_regs(460) => 
                           DataPath_RF_bus_selected_win_data_460_port, 
                           curr_proc_regs(459) => 
                           DataPath_RF_bus_selected_win_data_459_port, 
                           curr_proc_regs(458) => 
                           DataPath_RF_bus_selected_win_data_458_port, 
                           curr_proc_regs(457) => 
                           DataPath_RF_bus_selected_win_data_457_port, 
                           curr_proc_regs(456) => 
                           DataPath_RF_bus_selected_win_data_456_port, 
                           curr_proc_regs(455) => 
                           DataPath_RF_bus_selected_win_data_455_port, 
                           curr_proc_regs(454) => 
                           DataPath_RF_bus_selected_win_data_454_port, 
                           curr_proc_regs(453) => 
                           DataPath_RF_bus_selected_win_data_453_port, 
                           curr_proc_regs(452) => 
                           DataPath_RF_bus_selected_win_data_452_port, 
                           curr_proc_regs(451) => 
                           DataPath_RF_bus_selected_win_data_451_port, 
                           curr_proc_regs(450) => 
                           DataPath_RF_bus_selected_win_data_450_port, 
                           curr_proc_regs(449) => 
                           DataPath_RF_bus_selected_win_data_449_port, 
                           curr_proc_regs(448) => 
                           DataPath_RF_bus_selected_win_data_448_port, 
                           curr_proc_regs(447) => 
                           DataPath_RF_bus_selected_win_data_447_port, 
                           curr_proc_regs(446) => 
                           DataPath_RF_bus_selected_win_data_446_port, 
                           curr_proc_regs(445) => 
                           DataPath_RF_bus_selected_win_data_445_port, 
                           curr_proc_regs(444) => 
                           DataPath_RF_bus_selected_win_data_444_port, 
                           curr_proc_regs(443) => 
                           DataPath_RF_bus_selected_win_data_443_port, 
                           curr_proc_regs(442) => 
                           DataPath_RF_bus_selected_win_data_442_port, 
                           curr_proc_regs(441) => 
                           DataPath_RF_bus_selected_win_data_441_port, 
                           curr_proc_regs(440) => 
                           DataPath_RF_bus_selected_win_data_440_port, 
                           curr_proc_regs(439) => 
                           DataPath_RF_bus_selected_win_data_439_port, 
                           curr_proc_regs(438) => 
                           DataPath_RF_bus_selected_win_data_438_port, 
                           curr_proc_regs(437) => 
                           DataPath_RF_bus_selected_win_data_437_port, 
                           curr_proc_regs(436) => 
                           DataPath_RF_bus_selected_win_data_436_port, 
                           curr_proc_regs(435) => 
                           DataPath_RF_bus_selected_win_data_435_port, 
                           curr_proc_regs(434) => 
                           DataPath_RF_bus_selected_win_data_434_port, 
                           curr_proc_regs(433) => 
                           DataPath_RF_bus_selected_win_data_433_port, 
                           curr_proc_regs(432) => 
                           DataPath_RF_bus_selected_win_data_432_port, 
                           curr_proc_regs(431) => 
                           DataPath_RF_bus_selected_win_data_431_port, 
                           curr_proc_regs(430) => 
                           DataPath_RF_bus_selected_win_data_430_port, 
                           curr_proc_regs(429) => 
                           DataPath_RF_bus_selected_win_data_429_port, 
                           curr_proc_regs(428) => 
                           DataPath_RF_bus_selected_win_data_428_port, 
                           curr_proc_regs(427) => 
                           DataPath_RF_bus_selected_win_data_427_port, 
                           curr_proc_regs(426) => 
                           DataPath_RF_bus_selected_win_data_426_port, 
                           curr_proc_regs(425) => 
                           DataPath_RF_bus_selected_win_data_425_port, 
                           curr_proc_regs(424) => 
                           DataPath_RF_bus_selected_win_data_424_port, 
                           curr_proc_regs(423) => 
                           DataPath_RF_bus_selected_win_data_423_port, 
                           curr_proc_regs(422) => 
                           DataPath_RF_bus_selected_win_data_422_port, 
                           curr_proc_regs(421) => 
                           DataPath_RF_bus_selected_win_data_421_port, 
                           curr_proc_regs(420) => 
                           DataPath_RF_bus_selected_win_data_420_port, 
                           curr_proc_regs(419) => 
                           DataPath_RF_bus_selected_win_data_419_port, 
                           curr_proc_regs(418) => 
                           DataPath_RF_bus_selected_win_data_418_port, 
                           curr_proc_regs(417) => 
                           DataPath_RF_bus_selected_win_data_417_port, 
                           curr_proc_regs(416) => 
                           DataPath_RF_bus_selected_win_data_416_port, 
                           curr_proc_regs(415) => 
                           DataPath_RF_bus_selected_win_data_415_port, 
                           curr_proc_regs(414) => 
                           DataPath_RF_bus_selected_win_data_414_port, 
                           curr_proc_regs(413) => 
                           DataPath_RF_bus_selected_win_data_413_port, 
                           curr_proc_regs(412) => 
                           DataPath_RF_bus_selected_win_data_412_port, 
                           curr_proc_regs(411) => 
                           DataPath_RF_bus_selected_win_data_411_port, 
                           curr_proc_regs(410) => 
                           DataPath_RF_bus_selected_win_data_410_port, 
                           curr_proc_regs(409) => 
                           DataPath_RF_bus_selected_win_data_409_port, 
                           curr_proc_regs(408) => 
                           DataPath_RF_bus_selected_win_data_408_port, 
                           curr_proc_regs(407) => 
                           DataPath_RF_bus_selected_win_data_407_port, 
                           curr_proc_regs(406) => 
                           DataPath_RF_bus_selected_win_data_406_port, 
                           curr_proc_regs(405) => 
                           DataPath_RF_bus_selected_win_data_405_port, 
                           curr_proc_regs(404) => 
                           DataPath_RF_bus_selected_win_data_404_port, 
                           curr_proc_regs(403) => 
                           DataPath_RF_bus_selected_win_data_403_port, 
                           curr_proc_regs(402) => 
                           DataPath_RF_bus_selected_win_data_402_port, 
                           curr_proc_regs(401) => 
                           DataPath_RF_bus_selected_win_data_401_port, 
                           curr_proc_regs(400) => 
                           DataPath_RF_bus_selected_win_data_400_port, 
                           curr_proc_regs(399) => 
                           DataPath_RF_bus_selected_win_data_399_port, 
                           curr_proc_regs(398) => 
                           DataPath_RF_bus_selected_win_data_398_port, 
                           curr_proc_regs(397) => 
                           DataPath_RF_bus_selected_win_data_397_port, 
                           curr_proc_regs(396) => 
                           DataPath_RF_bus_selected_win_data_396_port, 
                           curr_proc_regs(395) => 
                           DataPath_RF_bus_selected_win_data_395_port, 
                           curr_proc_regs(394) => 
                           DataPath_RF_bus_selected_win_data_394_port, 
                           curr_proc_regs(393) => 
                           DataPath_RF_bus_selected_win_data_393_port, 
                           curr_proc_regs(392) => 
                           DataPath_RF_bus_selected_win_data_392_port, 
                           curr_proc_regs(391) => 
                           DataPath_RF_bus_selected_win_data_391_port, 
                           curr_proc_regs(390) => 
                           DataPath_RF_bus_selected_win_data_390_port, 
                           curr_proc_regs(389) => 
                           DataPath_RF_bus_selected_win_data_389_port, 
                           curr_proc_regs(388) => 
                           DataPath_RF_bus_selected_win_data_388_port, 
                           curr_proc_regs(387) => 
                           DataPath_RF_bus_selected_win_data_387_port, 
                           curr_proc_regs(386) => 
                           DataPath_RF_bus_selected_win_data_386_port, 
                           curr_proc_regs(385) => 
                           DataPath_RF_bus_selected_win_data_385_port, 
                           curr_proc_regs(384) => 
                           DataPath_RF_bus_selected_win_data_384_port, 
                           curr_proc_regs(383) => 
                           DataPath_RF_bus_selected_win_data_383_port, 
                           curr_proc_regs(382) => 
                           DataPath_RF_bus_selected_win_data_382_port, 
                           curr_proc_regs(381) => 
                           DataPath_RF_bus_selected_win_data_381_port, 
                           curr_proc_regs(380) => 
                           DataPath_RF_bus_selected_win_data_380_port, 
                           curr_proc_regs(379) => 
                           DataPath_RF_bus_selected_win_data_379_port, 
                           curr_proc_regs(378) => 
                           DataPath_RF_bus_selected_win_data_378_port, 
                           curr_proc_regs(377) => 
                           DataPath_RF_bus_selected_win_data_377_port, 
                           curr_proc_regs(376) => 
                           DataPath_RF_bus_selected_win_data_376_port, 
                           curr_proc_regs(375) => 
                           DataPath_RF_bus_selected_win_data_375_port, 
                           curr_proc_regs(374) => 
                           DataPath_RF_bus_selected_win_data_374_port, 
                           curr_proc_regs(373) => 
                           DataPath_RF_bus_selected_win_data_373_port, 
                           curr_proc_regs(372) => 
                           DataPath_RF_bus_selected_win_data_372_port, 
                           curr_proc_regs(371) => 
                           DataPath_RF_bus_selected_win_data_371_port, 
                           curr_proc_regs(370) => 
                           DataPath_RF_bus_selected_win_data_370_port, 
                           curr_proc_regs(369) => 
                           DataPath_RF_bus_selected_win_data_369_port, 
                           curr_proc_regs(368) => 
                           DataPath_RF_bus_selected_win_data_368_port, 
                           curr_proc_regs(367) => 
                           DataPath_RF_bus_selected_win_data_367_port, 
                           curr_proc_regs(366) => 
                           DataPath_RF_bus_selected_win_data_366_port, 
                           curr_proc_regs(365) => 
                           DataPath_RF_bus_selected_win_data_365_port, 
                           curr_proc_regs(364) => 
                           DataPath_RF_bus_selected_win_data_364_port, 
                           curr_proc_regs(363) => 
                           DataPath_RF_bus_selected_win_data_363_port, 
                           curr_proc_regs(362) => 
                           DataPath_RF_bus_selected_win_data_362_port, 
                           curr_proc_regs(361) => 
                           DataPath_RF_bus_selected_win_data_361_port, 
                           curr_proc_regs(360) => 
                           DataPath_RF_bus_selected_win_data_360_port, 
                           curr_proc_regs(359) => 
                           DataPath_RF_bus_selected_win_data_359_port, 
                           curr_proc_regs(358) => 
                           DataPath_RF_bus_selected_win_data_358_port, 
                           curr_proc_regs(357) => 
                           DataPath_RF_bus_selected_win_data_357_port, 
                           curr_proc_regs(356) => 
                           DataPath_RF_bus_selected_win_data_356_port, 
                           curr_proc_regs(355) => 
                           DataPath_RF_bus_selected_win_data_355_port, 
                           curr_proc_regs(354) => 
                           DataPath_RF_bus_selected_win_data_354_port, 
                           curr_proc_regs(353) => 
                           DataPath_RF_bus_selected_win_data_353_port, 
                           curr_proc_regs(352) => 
                           DataPath_RF_bus_selected_win_data_352_port, 
                           curr_proc_regs(351) => 
                           DataPath_RF_bus_selected_win_data_351_port, 
                           curr_proc_regs(350) => 
                           DataPath_RF_bus_selected_win_data_350_port, 
                           curr_proc_regs(349) => 
                           DataPath_RF_bus_selected_win_data_349_port, 
                           curr_proc_regs(348) => 
                           DataPath_RF_bus_selected_win_data_348_port, 
                           curr_proc_regs(347) => 
                           DataPath_RF_bus_selected_win_data_347_port, 
                           curr_proc_regs(346) => 
                           DataPath_RF_bus_selected_win_data_346_port, 
                           curr_proc_regs(345) => 
                           DataPath_RF_bus_selected_win_data_345_port, 
                           curr_proc_regs(344) => 
                           DataPath_RF_bus_selected_win_data_344_port, 
                           curr_proc_regs(343) => 
                           DataPath_RF_bus_selected_win_data_343_port, 
                           curr_proc_regs(342) => 
                           DataPath_RF_bus_selected_win_data_342_port, 
                           curr_proc_regs(341) => 
                           DataPath_RF_bus_selected_win_data_341_port, 
                           curr_proc_regs(340) => 
                           DataPath_RF_bus_selected_win_data_340_port, 
                           curr_proc_regs(339) => 
                           DataPath_RF_bus_selected_win_data_339_port, 
                           curr_proc_regs(338) => 
                           DataPath_RF_bus_selected_win_data_338_port, 
                           curr_proc_regs(337) => 
                           DataPath_RF_bus_selected_win_data_337_port, 
                           curr_proc_regs(336) => 
                           DataPath_RF_bus_selected_win_data_336_port, 
                           curr_proc_regs(335) => 
                           DataPath_RF_bus_selected_win_data_335_port, 
                           curr_proc_regs(334) => 
                           DataPath_RF_bus_selected_win_data_334_port, 
                           curr_proc_regs(333) => 
                           DataPath_RF_bus_selected_win_data_333_port, 
                           curr_proc_regs(332) => 
                           DataPath_RF_bus_selected_win_data_332_port, 
                           curr_proc_regs(331) => 
                           DataPath_RF_bus_selected_win_data_331_port, 
                           curr_proc_regs(330) => 
                           DataPath_RF_bus_selected_win_data_330_port, 
                           curr_proc_regs(329) => 
                           DataPath_RF_bus_selected_win_data_329_port, 
                           curr_proc_regs(328) => 
                           DataPath_RF_bus_selected_win_data_328_port, 
                           curr_proc_regs(327) => 
                           DataPath_RF_bus_selected_win_data_327_port, 
                           curr_proc_regs(326) => 
                           DataPath_RF_bus_selected_win_data_326_port, 
                           curr_proc_regs(325) => 
                           DataPath_RF_bus_selected_win_data_325_port, 
                           curr_proc_regs(324) => 
                           DataPath_RF_bus_selected_win_data_324_port, 
                           curr_proc_regs(323) => 
                           DataPath_RF_bus_selected_win_data_323_port, 
                           curr_proc_regs(322) => 
                           DataPath_RF_bus_selected_win_data_322_port, 
                           curr_proc_regs(321) => 
                           DataPath_RF_bus_selected_win_data_321_port, 
                           curr_proc_regs(320) => 
                           DataPath_RF_bus_selected_win_data_320_port, 
                           curr_proc_regs(319) => 
                           DataPath_RF_bus_selected_win_data_319_port, 
                           curr_proc_regs(318) => 
                           DataPath_RF_bus_selected_win_data_318_port, 
                           curr_proc_regs(317) => 
                           DataPath_RF_bus_selected_win_data_317_port, 
                           curr_proc_regs(316) => 
                           DataPath_RF_bus_selected_win_data_316_port, 
                           curr_proc_regs(315) => 
                           DataPath_RF_bus_selected_win_data_315_port, 
                           curr_proc_regs(314) => 
                           DataPath_RF_bus_selected_win_data_314_port, 
                           curr_proc_regs(313) => 
                           DataPath_RF_bus_selected_win_data_313_port, 
                           curr_proc_regs(312) => 
                           DataPath_RF_bus_selected_win_data_312_port, 
                           curr_proc_regs(311) => 
                           DataPath_RF_bus_selected_win_data_311_port, 
                           curr_proc_regs(310) => 
                           DataPath_RF_bus_selected_win_data_310_port, 
                           curr_proc_regs(309) => 
                           DataPath_RF_bus_selected_win_data_309_port, 
                           curr_proc_regs(308) => 
                           DataPath_RF_bus_selected_win_data_308_port, 
                           curr_proc_regs(307) => 
                           DataPath_RF_bus_selected_win_data_307_port, 
                           curr_proc_regs(306) => 
                           DataPath_RF_bus_selected_win_data_306_port, 
                           curr_proc_regs(305) => 
                           DataPath_RF_bus_selected_win_data_305_port, 
                           curr_proc_regs(304) => 
                           DataPath_RF_bus_selected_win_data_304_port, 
                           curr_proc_regs(303) => 
                           DataPath_RF_bus_selected_win_data_303_port, 
                           curr_proc_regs(302) => 
                           DataPath_RF_bus_selected_win_data_302_port, 
                           curr_proc_regs(301) => 
                           DataPath_RF_bus_selected_win_data_301_port, 
                           curr_proc_regs(300) => 
                           DataPath_RF_bus_selected_win_data_300_port, 
                           curr_proc_regs(299) => 
                           DataPath_RF_bus_selected_win_data_299_port, 
                           curr_proc_regs(298) => 
                           DataPath_RF_bus_selected_win_data_298_port, 
                           curr_proc_regs(297) => 
                           DataPath_RF_bus_selected_win_data_297_port, 
                           curr_proc_regs(296) => 
                           DataPath_RF_bus_selected_win_data_296_port, 
                           curr_proc_regs(295) => 
                           DataPath_RF_bus_selected_win_data_295_port, 
                           curr_proc_regs(294) => 
                           DataPath_RF_bus_selected_win_data_294_port, 
                           curr_proc_regs(293) => 
                           DataPath_RF_bus_selected_win_data_293_port, 
                           curr_proc_regs(292) => 
                           DataPath_RF_bus_selected_win_data_292_port, 
                           curr_proc_regs(291) => 
                           DataPath_RF_bus_selected_win_data_291_port, 
                           curr_proc_regs(290) => 
                           DataPath_RF_bus_selected_win_data_290_port, 
                           curr_proc_regs(289) => 
                           DataPath_RF_bus_selected_win_data_289_port, 
                           curr_proc_regs(288) => 
                           DataPath_RF_bus_selected_win_data_288_port, 
                           curr_proc_regs(287) => 
                           DataPath_RF_bus_selected_win_data_287_port, 
                           curr_proc_regs(286) => 
                           DataPath_RF_bus_selected_win_data_286_port, 
                           curr_proc_regs(285) => 
                           DataPath_RF_bus_selected_win_data_285_port, 
                           curr_proc_regs(284) => 
                           DataPath_RF_bus_selected_win_data_284_port, 
                           curr_proc_regs(283) => 
                           DataPath_RF_bus_selected_win_data_283_port, 
                           curr_proc_regs(282) => 
                           DataPath_RF_bus_selected_win_data_282_port, 
                           curr_proc_regs(281) => 
                           DataPath_RF_bus_selected_win_data_281_port, 
                           curr_proc_regs(280) => 
                           DataPath_RF_bus_selected_win_data_280_port, 
                           curr_proc_regs(279) => 
                           DataPath_RF_bus_selected_win_data_279_port, 
                           curr_proc_regs(278) => 
                           DataPath_RF_bus_selected_win_data_278_port, 
                           curr_proc_regs(277) => 
                           DataPath_RF_bus_selected_win_data_277_port, 
                           curr_proc_regs(276) => 
                           DataPath_RF_bus_selected_win_data_276_port, 
                           curr_proc_regs(275) => 
                           DataPath_RF_bus_selected_win_data_275_port, 
                           curr_proc_regs(274) => 
                           DataPath_RF_bus_selected_win_data_274_port, 
                           curr_proc_regs(273) => 
                           DataPath_RF_bus_selected_win_data_273_port, 
                           curr_proc_regs(272) => 
                           DataPath_RF_bus_selected_win_data_272_port, 
                           curr_proc_regs(271) => 
                           DataPath_RF_bus_selected_win_data_271_port, 
                           curr_proc_regs(270) => 
                           DataPath_RF_bus_selected_win_data_270_port, 
                           curr_proc_regs(269) => 
                           DataPath_RF_bus_selected_win_data_269_port, 
                           curr_proc_regs(268) => 
                           DataPath_RF_bus_selected_win_data_268_port, 
                           curr_proc_regs(267) => 
                           DataPath_RF_bus_selected_win_data_267_port, 
                           curr_proc_regs(266) => 
                           DataPath_RF_bus_selected_win_data_266_port, 
                           curr_proc_regs(265) => 
                           DataPath_RF_bus_selected_win_data_265_port, 
                           curr_proc_regs(264) => 
                           DataPath_RF_bus_selected_win_data_264_port, 
                           curr_proc_regs(263) => 
                           DataPath_RF_bus_selected_win_data_263_port, 
                           curr_proc_regs(262) => 
                           DataPath_RF_bus_selected_win_data_262_port, 
                           curr_proc_regs(261) => 
                           DataPath_RF_bus_selected_win_data_261_port, 
                           curr_proc_regs(260) => 
                           DataPath_RF_bus_selected_win_data_260_port, 
                           curr_proc_regs(259) => 
                           DataPath_RF_bus_selected_win_data_259_port, 
                           curr_proc_regs(258) => 
                           DataPath_RF_bus_selected_win_data_258_port, 
                           curr_proc_regs(257) => 
                           DataPath_RF_bus_selected_win_data_257_port, 
                           curr_proc_regs(256) => 
                           DataPath_RF_bus_selected_win_data_256_port, 
                           curr_proc_regs(255) => 
                           DataPath_RF_bus_selected_win_data_255_port, 
                           curr_proc_regs(254) => 
                           DataPath_RF_bus_selected_win_data_254_port, 
                           curr_proc_regs(253) => 
                           DataPath_RF_bus_selected_win_data_253_port, 
                           curr_proc_regs(252) => 
                           DataPath_RF_bus_selected_win_data_252_port, 
                           curr_proc_regs(251) => 
                           DataPath_RF_bus_selected_win_data_251_port, 
                           curr_proc_regs(250) => 
                           DataPath_RF_bus_selected_win_data_250_port, 
                           curr_proc_regs(249) => 
                           DataPath_RF_bus_selected_win_data_249_port, 
                           curr_proc_regs(248) => 
                           DataPath_RF_bus_selected_win_data_248_port, 
                           curr_proc_regs(247) => 
                           DataPath_RF_bus_selected_win_data_247_port, 
                           curr_proc_regs(246) => 
                           DataPath_RF_bus_selected_win_data_246_port, 
                           curr_proc_regs(245) => 
                           DataPath_RF_bus_selected_win_data_245_port, 
                           curr_proc_regs(244) => 
                           DataPath_RF_bus_selected_win_data_244_port, 
                           curr_proc_regs(243) => 
                           DataPath_RF_bus_selected_win_data_243_port, 
                           curr_proc_regs(242) => 
                           DataPath_RF_bus_selected_win_data_242_port, 
                           curr_proc_regs(241) => 
                           DataPath_RF_bus_selected_win_data_241_port, 
                           curr_proc_regs(240) => 
                           DataPath_RF_bus_selected_win_data_240_port, 
                           curr_proc_regs(239) => 
                           DataPath_RF_bus_selected_win_data_239_port, 
                           curr_proc_regs(238) => 
                           DataPath_RF_bus_selected_win_data_238_port, 
                           curr_proc_regs(237) => 
                           DataPath_RF_bus_selected_win_data_237_port, 
                           curr_proc_regs(236) => 
                           DataPath_RF_bus_selected_win_data_236_port, 
                           curr_proc_regs(235) => 
                           DataPath_RF_bus_selected_win_data_235_port, 
                           curr_proc_regs(234) => 
                           DataPath_RF_bus_selected_win_data_234_port, 
                           curr_proc_regs(233) => 
                           DataPath_RF_bus_selected_win_data_233_port, 
                           curr_proc_regs(232) => 
                           DataPath_RF_bus_selected_win_data_232_port, 
                           curr_proc_regs(231) => 
                           DataPath_RF_bus_selected_win_data_231_port, 
                           curr_proc_regs(230) => 
                           DataPath_RF_bus_selected_win_data_230_port, 
                           curr_proc_regs(229) => 
                           DataPath_RF_bus_selected_win_data_229_port, 
                           curr_proc_regs(228) => 
                           DataPath_RF_bus_selected_win_data_228_port, 
                           curr_proc_regs(227) => 
                           DataPath_RF_bus_selected_win_data_227_port, 
                           curr_proc_regs(226) => 
                           DataPath_RF_bus_selected_win_data_226_port, 
                           curr_proc_regs(225) => 
                           DataPath_RF_bus_selected_win_data_225_port, 
                           curr_proc_regs(224) => 
                           DataPath_RF_bus_selected_win_data_224_port, 
                           curr_proc_regs(223) => 
                           DataPath_RF_bus_selected_win_data_223_port, 
                           curr_proc_regs(222) => 
                           DataPath_RF_bus_selected_win_data_222_port, 
                           curr_proc_regs(221) => 
                           DataPath_RF_bus_selected_win_data_221_port, 
                           curr_proc_regs(220) => 
                           DataPath_RF_bus_selected_win_data_220_port, 
                           curr_proc_regs(219) => 
                           DataPath_RF_bus_selected_win_data_219_port, 
                           curr_proc_regs(218) => 
                           DataPath_RF_bus_selected_win_data_218_port, 
                           curr_proc_regs(217) => 
                           DataPath_RF_bus_selected_win_data_217_port, 
                           curr_proc_regs(216) => 
                           DataPath_RF_bus_selected_win_data_216_port, 
                           curr_proc_regs(215) => 
                           DataPath_RF_bus_selected_win_data_215_port, 
                           curr_proc_regs(214) => 
                           DataPath_RF_bus_selected_win_data_214_port, 
                           curr_proc_regs(213) => 
                           DataPath_RF_bus_selected_win_data_213_port, 
                           curr_proc_regs(212) => 
                           DataPath_RF_bus_selected_win_data_212_port, 
                           curr_proc_regs(211) => 
                           DataPath_RF_bus_selected_win_data_211_port, 
                           curr_proc_regs(210) => 
                           DataPath_RF_bus_selected_win_data_210_port, 
                           curr_proc_regs(209) => 
                           DataPath_RF_bus_selected_win_data_209_port, 
                           curr_proc_regs(208) => 
                           DataPath_RF_bus_selected_win_data_208_port, 
                           curr_proc_regs(207) => 
                           DataPath_RF_bus_selected_win_data_207_port, 
                           curr_proc_regs(206) => 
                           DataPath_RF_bus_selected_win_data_206_port, 
                           curr_proc_regs(205) => 
                           DataPath_RF_bus_selected_win_data_205_port, 
                           curr_proc_regs(204) => 
                           DataPath_RF_bus_selected_win_data_204_port, 
                           curr_proc_regs(203) => 
                           DataPath_RF_bus_selected_win_data_203_port, 
                           curr_proc_regs(202) => 
                           DataPath_RF_bus_selected_win_data_202_port, 
                           curr_proc_regs(201) => 
                           DataPath_RF_bus_selected_win_data_201_port, 
                           curr_proc_regs(200) => 
                           DataPath_RF_bus_selected_win_data_200_port, 
                           curr_proc_regs(199) => 
                           DataPath_RF_bus_selected_win_data_199_port, 
                           curr_proc_regs(198) => 
                           DataPath_RF_bus_selected_win_data_198_port, 
                           curr_proc_regs(197) => 
                           DataPath_RF_bus_selected_win_data_197_port, 
                           curr_proc_regs(196) => 
                           DataPath_RF_bus_selected_win_data_196_port, 
                           curr_proc_regs(195) => 
                           DataPath_RF_bus_selected_win_data_195_port, 
                           curr_proc_regs(194) => 
                           DataPath_RF_bus_selected_win_data_194_port, 
                           curr_proc_regs(193) => 
                           DataPath_RF_bus_selected_win_data_193_port, 
                           curr_proc_regs(192) => 
                           DataPath_RF_bus_selected_win_data_192_port, 
                           curr_proc_regs(191) => 
                           DataPath_RF_bus_selected_win_data_191_port, 
                           curr_proc_regs(190) => 
                           DataPath_RF_bus_selected_win_data_190_port, 
                           curr_proc_regs(189) => 
                           DataPath_RF_bus_selected_win_data_189_port, 
                           curr_proc_regs(188) => 
                           DataPath_RF_bus_selected_win_data_188_port, 
                           curr_proc_regs(187) => 
                           DataPath_RF_bus_selected_win_data_187_port, 
                           curr_proc_regs(186) => 
                           DataPath_RF_bus_selected_win_data_186_port, 
                           curr_proc_regs(185) => 
                           DataPath_RF_bus_selected_win_data_185_port, 
                           curr_proc_regs(184) => 
                           DataPath_RF_bus_selected_win_data_184_port, 
                           curr_proc_regs(183) => 
                           DataPath_RF_bus_selected_win_data_183_port, 
                           curr_proc_regs(182) => 
                           DataPath_RF_bus_selected_win_data_182_port, 
                           curr_proc_regs(181) => 
                           DataPath_RF_bus_selected_win_data_181_port, 
                           curr_proc_regs(180) => 
                           DataPath_RF_bus_selected_win_data_180_port, 
                           curr_proc_regs(179) => 
                           DataPath_RF_bus_selected_win_data_179_port, 
                           curr_proc_regs(178) => 
                           DataPath_RF_bus_selected_win_data_178_port, 
                           curr_proc_regs(177) => 
                           DataPath_RF_bus_selected_win_data_177_port, 
                           curr_proc_regs(176) => 
                           DataPath_RF_bus_selected_win_data_176_port, 
                           curr_proc_regs(175) => 
                           DataPath_RF_bus_selected_win_data_175_port, 
                           curr_proc_regs(174) => 
                           DataPath_RF_bus_selected_win_data_174_port, 
                           curr_proc_regs(173) => 
                           DataPath_RF_bus_selected_win_data_173_port, 
                           curr_proc_regs(172) => 
                           DataPath_RF_bus_selected_win_data_172_port, 
                           curr_proc_regs(171) => 
                           DataPath_RF_bus_selected_win_data_171_port, 
                           curr_proc_regs(170) => 
                           DataPath_RF_bus_selected_win_data_170_port, 
                           curr_proc_regs(169) => 
                           DataPath_RF_bus_selected_win_data_169_port, 
                           curr_proc_regs(168) => 
                           DataPath_RF_bus_selected_win_data_168_port, 
                           curr_proc_regs(167) => 
                           DataPath_RF_bus_selected_win_data_167_port, 
                           curr_proc_regs(166) => 
                           DataPath_RF_bus_selected_win_data_166_port, 
                           curr_proc_regs(165) => 
                           DataPath_RF_bus_selected_win_data_165_port, 
                           curr_proc_regs(164) => 
                           DataPath_RF_bus_selected_win_data_164_port, 
                           curr_proc_regs(163) => 
                           DataPath_RF_bus_selected_win_data_163_port, 
                           curr_proc_regs(162) => 
                           DataPath_RF_bus_selected_win_data_162_port, 
                           curr_proc_regs(161) => 
                           DataPath_RF_bus_selected_win_data_161_port, 
                           curr_proc_regs(160) => 
                           DataPath_RF_bus_selected_win_data_160_port, 
                           curr_proc_regs(159) => 
                           DataPath_RF_bus_selected_win_data_159_port, 
                           curr_proc_regs(158) => 
                           DataPath_RF_bus_selected_win_data_158_port, 
                           curr_proc_regs(157) => 
                           DataPath_RF_bus_selected_win_data_157_port, 
                           curr_proc_regs(156) => 
                           DataPath_RF_bus_selected_win_data_156_port, 
                           curr_proc_regs(155) => 
                           DataPath_RF_bus_selected_win_data_155_port, 
                           curr_proc_regs(154) => 
                           DataPath_RF_bus_selected_win_data_154_port, 
                           curr_proc_regs(153) => 
                           DataPath_RF_bus_selected_win_data_153_port, 
                           curr_proc_regs(152) => 
                           DataPath_RF_bus_selected_win_data_152_port, 
                           curr_proc_regs(151) => 
                           DataPath_RF_bus_selected_win_data_151_port, 
                           curr_proc_regs(150) => 
                           DataPath_RF_bus_selected_win_data_150_port, 
                           curr_proc_regs(149) => 
                           DataPath_RF_bus_selected_win_data_149_port, 
                           curr_proc_regs(148) => 
                           DataPath_RF_bus_selected_win_data_148_port, 
                           curr_proc_regs(147) => 
                           DataPath_RF_bus_selected_win_data_147_port, 
                           curr_proc_regs(146) => 
                           DataPath_RF_bus_selected_win_data_146_port, 
                           curr_proc_regs(145) => 
                           DataPath_RF_bus_selected_win_data_145_port, 
                           curr_proc_regs(144) => 
                           DataPath_RF_bus_selected_win_data_144_port, 
                           curr_proc_regs(143) => 
                           DataPath_RF_bus_selected_win_data_143_port, 
                           curr_proc_regs(142) => 
                           DataPath_RF_bus_selected_win_data_142_port, 
                           curr_proc_regs(141) => 
                           DataPath_RF_bus_selected_win_data_141_port, 
                           curr_proc_regs(140) => 
                           DataPath_RF_bus_selected_win_data_140_port, 
                           curr_proc_regs(139) => 
                           DataPath_RF_bus_selected_win_data_139_port, 
                           curr_proc_regs(138) => 
                           DataPath_RF_bus_selected_win_data_138_port, 
                           curr_proc_regs(137) => 
                           DataPath_RF_bus_selected_win_data_137_port, 
                           curr_proc_regs(136) => 
                           DataPath_RF_bus_selected_win_data_136_port, 
                           curr_proc_regs(135) => 
                           DataPath_RF_bus_selected_win_data_135_port, 
                           curr_proc_regs(134) => 
                           DataPath_RF_bus_selected_win_data_134_port, 
                           curr_proc_regs(133) => 
                           DataPath_RF_bus_selected_win_data_133_port, 
                           curr_proc_regs(132) => 
                           DataPath_RF_bus_selected_win_data_132_port, 
                           curr_proc_regs(131) => 
                           DataPath_RF_bus_selected_win_data_131_port, 
                           curr_proc_regs(130) => 
                           DataPath_RF_bus_selected_win_data_130_port, 
                           curr_proc_regs(129) => 
                           DataPath_RF_bus_selected_win_data_129_port, 
                           curr_proc_regs(128) => 
                           DataPath_RF_bus_selected_win_data_128_port, 
                           curr_proc_regs(127) => 
                           DataPath_RF_bus_selected_win_data_127_port, 
                           curr_proc_regs(126) => 
                           DataPath_RF_bus_selected_win_data_126_port, 
                           curr_proc_regs(125) => 
                           DataPath_RF_bus_selected_win_data_125_port, 
                           curr_proc_regs(124) => 
                           DataPath_RF_bus_selected_win_data_124_port, 
                           curr_proc_regs(123) => 
                           DataPath_RF_bus_selected_win_data_123_port, 
                           curr_proc_regs(122) => 
                           DataPath_RF_bus_selected_win_data_122_port, 
                           curr_proc_regs(121) => 
                           DataPath_RF_bus_selected_win_data_121_port, 
                           curr_proc_regs(120) => 
                           DataPath_RF_bus_selected_win_data_120_port, 
                           curr_proc_regs(119) => 
                           DataPath_RF_bus_selected_win_data_119_port, 
                           curr_proc_regs(118) => 
                           DataPath_RF_bus_selected_win_data_118_port, 
                           curr_proc_regs(117) => 
                           DataPath_RF_bus_selected_win_data_117_port, 
                           curr_proc_regs(116) => 
                           DataPath_RF_bus_selected_win_data_116_port, 
                           curr_proc_regs(115) => 
                           DataPath_RF_bus_selected_win_data_115_port, 
                           curr_proc_regs(114) => 
                           DataPath_RF_bus_selected_win_data_114_port, 
                           curr_proc_regs(113) => 
                           DataPath_RF_bus_selected_win_data_113_port, 
                           curr_proc_regs(112) => 
                           DataPath_RF_bus_selected_win_data_112_port, 
                           curr_proc_regs(111) => 
                           DataPath_RF_bus_selected_win_data_111_port, 
                           curr_proc_regs(110) => 
                           DataPath_RF_bus_selected_win_data_110_port, 
                           curr_proc_regs(109) => 
                           DataPath_RF_bus_selected_win_data_109_port, 
                           curr_proc_regs(108) => 
                           DataPath_RF_bus_selected_win_data_108_port, 
                           curr_proc_regs(107) => 
                           DataPath_RF_bus_selected_win_data_107_port, 
                           curr_proc_regs(106) => 
                           DataPath_RF_bus_selected_win_data_106_port, 
                           curr_proc_regs(105) => 
                           DataPath_RF_bus_selected_win_data_105_port, 
                           curr_proc_regs(104) => 
                           DataPath_RF_bus_selected_win_data_104_port, 
                           curr_proc_regs(103) => 
                           DataPath_RF_bus_selected_win_data_103_port, 
                           curr_proc_regs(102) => 
                           DataPath_RF_bus_selected_win_data_102_port, 
                           curr_proc_regs(101) => 
                           DataPath_RF_bus_selected_win_data_101_port, 
                           curr_proc_regs(100) => 
                           DataPath_RF_bus_selected_win_data_100_port, 
                           curr_proc_regs(99) => 
                           DataPath_RF_bus_selected_win_data_99_port, 
                           curr_proc_regs(98) => 
                           DataPath_RF_bus_selected_win_data_98_port, 
                           curr_proc_regs(97) => 
                           DataPath_RF_bus_selected_win_data_97_port, 
                           curr_proc_regs(96) => 
                           DataPath_RF_bus_selected_win_data_96_port, 
                           curr_proc_regs(95) => 
                           DataPath_RF_bus_selected_win_data_95_port, 
                           curr_proc_regs(94) => 
                           DataPath_RF_bus_selected_win_data_94_port, 
                           curr_proc_regs(93) => 
                           DataPath_RF_bus_selected_win_data_93_port, 
                           curr_proc_regs(92) => 
                           DataPath_RF_bus_selected_win_data_92_port, 
                           curr_proc_regs(91) => 
                           DataPath_RF_bus_selected_win_data_91_port, 
                           curr_proc_regs(90) => 
                           DataPath_RF_bus_selected_win_data_90_port, 
                           curr_proc_regs(89) => 
                           DataPath_RF_bus_selected_win_data_89_port, 
                           curr_proc_regs(88) => 
                           DataPath_RF_bus_selected_win_data_88_port, 
                           curr_proc_regs(87) => 
                           DataPath_RF_bus_selected_win_data_87_port, 
                           curr_proc_regs(86) => 
                           DataPath_RF_bus_selected_win_data_86_port, 
                           curr_proc_regs(85) => 
                           DataPath_RF_bus_selected_win_data_85_port, 
                           curr_proc_regs(84) => 
                           DataPath_RF_bus_selected_win_data_84_port, 
                           curr_proc_regs(83) => 
                           DataPath_RF_bus_selected_win_data_83_port, 
                           curr_proc_regs(82) => 
                           DataPath_RF_bus_selected_win_data_82_port, 
                           curr_proc_regs(81) => 
                           DataPath_RF_bus_selected_win_data_81_port, 
                           curr_proc_regs(80) => 
                           DataPath_RF_bus_selected_win_data_80_port, 
                           curr_proc_regs(79) => 
                           DataPath_RF_bus_selected_win_data_79_port, 
                           curr_proc_regs(78) => 
                           DataPath_RF_bus_selected_win_data_78_port, 
                           curr_proc_regs(77) => 
                           DataPath_RF_bus_selected_win_data_77_port, 
                           curr_proc_regs(76) => 
                           DataPath_RF_bus_selected_win_data_76_port, 
                           curr_proc_regs(75) => 
                           DataPath_RF_bus_selected_win_data_75_port, 
                           curr_proc_regs(74) => 
                           DataPath_RF_bus_selected_win_data_74_port, 
                           curr_proc_regs(73) => 
                           DataPath_RF_bus_selected_win_data_73_port, 
                           curr_proc_regs(72) => 
                           DataPath_RF_bus_selected_win_data_72_port, 
                           curr_proc_regs(71) => 
                           DataPath_RF_bus_selected_win_data_71_port, 
                           curr_proc_regs(70) => 
                           DataPath_RF_bus_selected_win_data_70_port, 
                           curr_proc_regs(69) => 
                           DataPath_RF_bus_selected_win_data_69_port, 
                           curr_proc_regs(68) => 
                           DataPath_RF_bus_selected_win_data_68_port, 
                           curr_proc_regs(67) => 
                           DataPath_RF_bus_selected_win_data_67_port, 
                           curr_proc_regs(66) => 
                           DataPath_RF_bus_selected_win_data_66_port, 
                           curr_proc_regs(65) => 
                           DataPath_RF_bus_selected_win_data_65_port, 
                           curr_proc_regs(64) => 
                           DataPath_RF_bus_selected_win_data_64_port, 
                           curr_proc_regs(63) => 
                           DataPath_RF_bus_selected_win_data_63_port, 
                           curr_proc_regs(62) => 
                           DataPath_RF_bus_selected_win_data_62_port, 
                           curr_proc_regs(61) => 
                           DataPath_RF_bus_selected_win_data_61_port, 
                           curr_proc_regs(60) => 
                           DataPath_RF_bus_selected_win_data_60_port, 
                           curr_proc_regs(59) => 
                           DataPath_RF_bus_selected_win_data_59_port, 
                           curr_proc_regs(58) => 
                           DataPath_RF_bus_selected_win_data_58_port, 
                           curr_proc_regs(57) => 
                           DataPath_RF_bus_selected_win_data_57_port, 
                           curr_proc_regs(56) => 
                           DataPath_RF_bus_selected_win_data_56_port, 
                           curr_proc_regs(55) => 
                           DataPath_RF_bus_selected_win_data_55_port, 
                           curr_proc_regs(54) => 
                           DataPath_RF_bus_selected_win_data_54_port, 
                           curr_proc_regs(53) => 
                           DataPath_RF_bus_selected_win_data_53_port, 
                           curr_proc_regs(52) => 
                           DataPath_RF_bus_selected_win_data_52_port, 
                           curr_proc_regs(51) => 
                           DataPath_RF_bus_selected_win_data_51_port, 
                           curr_proc_regs(50) => 
                           DataPath_RF_bus_selected_win_data_50_port, 
                           curr_proc_regs(49) => 
                           DataPath_RF_bus_selected_win_data_49_port, 
                           curr_proc_regs(48) => 
                           DataPath_RF_bus_selected_win_data_48_port, 
                           curr_proc_regs(47) => 
                           DataPath_RF_bus_selected_win_data_47_port, 
                           curr_proc_regs(46) => 
                           DataPath_RF_bus_selected_win_data_46_port, 
                           curr_proc_regs(45) => 
                           DataPath_RF_bus_selected_win_data_45_port, 
                           curr_proc_regs(44) => 
                           DataPath_RF_bus_selected_win_data_44_port, 
                           curr_proc_regs(43) => 
                           DataPath_RF_bus_selected_win_data_43_port, 
                           curr_proc_regs(42) => 
                           DataPath_RF_bus_selected_win_data_42_port, 
                           curr_proc_regs(41) => 
                           DataPath_RF_bus_selected_win_data_41_port, 
                           curr_proc_regs(40) => 
                           DataPath_RF_bus_selected_win_data_40_port, 
                           curr_proc_regs(39) => 
                           DataPath_RF_bus_selected_win_data_39_port, 
                           curr_proc_regs(38) => 
                           DataPath_RF_bus_selected_win_data_38_port, 
                           curr_proc_regs(37) => 
                           DataPath_RF_bus_selected_win_data_37_port, 
                           curr_proc_regs(36) => 
                           DataPath_RF_bus_selected_win_data_36_port, 
                           curr_proc_regs(35) => 
                           DataPath_RF_bus_selected_win_data_35_port, 
                           curr_proc_regs(34) => 
                           DataPath_RF_bus_selected_win_data_34_port, 
                           curr_proc_regs(33) => 
                           DataPath_RF_bus_selected_win_data_33_port, 
                           curr_proc_regs(32) => 
                           DataPath_RF_bus_selected_win_data_32_port, 
                           curr_proc_regs(31) => 
                           DataPath_RF_bus_selected_win_data_31_port, 
                           curr_proc_regs(30) => 
                           DataPath_RF_bus_selected_win_data_30_port, 
                           curr_proc_regs(29) => 
                           DataPath_RF_bus_selected_win_data_29_port, 
                           curr_proc_regs(28) => 
                           DataPath_RF_bus_selected_win_data_28_port, 
                           curr_proc_regs(27) => 
                           DataPath_RF_bus_selected_win_data_27_port, 
                           curr_proc_regs(26) => 
                           DataPath_RF_bus_selected_win_data_26_port, 
                           curr_proc_regs(25) => 
                           DataPath_RF_bus_selected_win_data_25_port, 
                           curr_proc_regs(24) => 
                           DataPath_RF_bus_selected_win_data_24_port, 
                           curr_proc_regs(23) => 
                           DataPath_RF_bus_selected_win_data_23_port, 
                           curr_proc_regs(22) => 
                           DataPath_RF_bus_selected_win_data_22_port, 
                           curr_proc_regs(21) => 
                           DataPath_RF_bus_selected_win_data_21_port, 
                           curr_proc_regs(20) => 
                           DataPath_RF_bus_selected_win_data_20_port, 
                           curr_proc_regs(19) => 
                           DataPath_RF_bus_selected_win_data_19_port, 
                           curr_proc_regs(18) => 
                           DataPath_RF_bus_selected_win_data_18_port, 
                           curr_proc_regs(17) => 
                           DataPath_RF_bus_selected_win_data_17_port, 
                           curr_proc_regs(16) => 
                           DataPath_RF_bus_selected_win_data_16_port, 
                           curr_proc_regs(15) => 
                           DataPath_RF_bus_selected_win_data_15_port, 
                           curr_proc_regs(14) => 
                           DataPath_RF_bus_selected_win_data_14_port, 
                           curr_proc_regs(13) => 
                           DataPath_RF_bus_selected_win_data_13_port, 
                           curr_proc_regs(12) => 
                           DataPath_RF_bus_selected_win_data_12_port, 
                           curr_proc_regs(11) => 
                           DataPath_RF_bus_selected_win_data_11_port, 
                           curr_proc_regs(10) => 
                           DataPath_RF_bus_selected_win_data_10_port, 
                           curr_proc_regs(9) => 
                           DataPath_RF_bus_selected_win_data_9_port, 
                           curr_proc_regs(8) => 
                           DataPath_RF_bus_selected_win_data_8_port, 
                           curr_proc_regs(7) => 
                           DataPath_RF_bus_selected_win_data_7_port, 
                           curr_proc_regs(6) => 
                           DataPath_RF_bus_selected_win_data_6_port, 
                           curr_proc_regs(5) => 
                           DataPath_RF_bus_selected_win_data_5_port, 
                           curr_proc_regs(4) => 
                           DataPath_RF_bus_selected_win_data_4_port, 
                           curr_proc_regs(3) => 
                           DataPath_RF_bus_selected_win_data_3_port, 
                           curr_proc_regs(2) => 
                           DataPath_RF_bus_selected_win_data_2_port, 
                           curr_proc_regs(1) => 
                           DataPath_RF_bus_selected_win_data_1_port, 
                           curr_proc_regs(0) => 
                           DataPath_RF_bus_selected_win_data_0_port);
   DataPath_WRF_CUhw_curr_data_reg_0_inst : DFF_X1 port map( D => n3357, CK => 
                           CLK, Q => n_1064, QN => 
                           DataPath_WRF_CUhw_curr_data_0_port);
   DataPath_WRF_CUhw_curr_data_reg_1_inst : DFF_X1 port map( D => n3356, CK => 
                           CLK, Q => n_1065, QN => 
                           DataPath_WRF_CUhw_curr_data_1_port);
   DataPath_WRF_CUhw_curr_data_reg_2_inst : DFF_X1 port map( D => n3355, CK => 
                           CLK, Q => n_1066, QN => 
                           DataPath_WRF_CUhw_curr_data_2_port);
   DataPath_WRF_CUhw_curr_data_reg_3_inst : DFF_X1 port map( D => n3354, CK => 
                           CLK, Q => n_1067, QN => 
                           DataPath_WRF_CUhw_curr_data_3_port);
   DataPath_WRF_CUhw_curr_data_reg_4_inst : DFF_X1 port map( D => n3353, CK => 
                           CLK, Q => n_1068, QN => 
                           DataPath_WRF_CUhw_curr_data_4_port);
   DataPath_WRF_CUhw_curr_data_reg_5_inst : DFF_X1 port map( D => n3352, CK => 
                           CLK, Q => n_1069, QN => 
                           DataPath_WRF_CUhw_curr_data_5_port);
   DataPath_WRF_CUhw_curr_data_reg_6_inst : DFF_X1 port map( D => n3351, CK => 
                           CLK, Q => n_1070, QN => 
                           DataPath_WRF_CUhw_curr_data_6_port);
   DataPath_WRF_CUhw_curr_data_reg_7_inst : DFF_X1 port map( D => n3350, CK => 
                           CLK, Q => n_1071, QN => 
                           DataPath_WRF_CUhw_curr_data_7_port);
   DataPath_WRF_CUhw_curr_data_reg_8_inst : DFF_X1 port map( D => n3349, CK => 
                           CLK, Q => n_1072, QN => 
                           DataPath_WRF_CUhw_curr_data_8_port);
   DataPath_WRF_CUhw_curr_data_reg_9_inst : DFF_X1 port map( D => n3348, CK => 
                           CLK, Q => n_1073, QN => 
                           DataPath_WRF_CUhw_curr_data_9_port);
   DataPath_WRF_CUhw_curr_data_reg_10_inst : DFF_X1 port map( D => n3347, CK =>
                           CLK, Q => n_1074, QN => 
                           DataPath_WRF_CUhw_curr_data_10_port);
   DataPath_WRF_CUhw_curr_data_reg_11_inst : DFF_X1 port map( D => n3346, CK =>
                           CLK, Q => n_1075, QN => 
                           DataPath_WRF_CUhw_curr_data_11_port);
   DataPath_WRF_CUhw_curr_data_reg_12_inst : DFF_X1 port map( D => n3345, CK =>
                           CLK, Q => n_1076, QN => 
                           DataPath_WRF_CUhw_curr_data_12_port);
   DataPath_WRF_CUhw_curr_data_reg_13_inst : DFF_X1 port map( D => n3344, CK =>
                           CLK, Q => n_1077, QN => 
                           DataPath_WRF_CUhw_curr_data_13_port);
   DataPath_WRF_CUhw_curr_data_reg_14_inst : DFF_X1 port map( D => n3343, CK =>
                           CLK, Q => n_1078, QN => 
                           DataPath_WRF_CUhw_curr_data_14_port);
   DataPath_WRF_CUhw_curr_data_reg_15_inst : DFF_X1 port map( D => n3342, CK =>
                           CLK, Q => n_1079, QN => 
                           DataPath_WRF_CUhw_curr_data_15_port);
   DataPath_WRF_CUhw_curr_data_reg_16_inst : DFF_X1 port map( D => n3341, CK =>
                           CLK, Q => n_1080, QN => 
                           DataPath_WRF_CUhw_curr_data_16_port);
   DataPath_WRF_CUhw_curr_data_reg_17_inst : DFF_X1 port map( D => n3340, CK =>
                           CLK, Q => n_1081, QN => 
                           DataPath_WRF_CUhw_curr_data_17_port);
   DataPath_WRF_CUhw_curr_data_reg_18_inst : DFF_X1 port map( D => n3339, CK =>
                           CLK, Q => n_1082, QN => 
                           DataPath_WRF_CUhw_curr_data_18_port);
   DataPath_WRF_CUhw_curr_data_reg_19_inst : DFF_X1 port map( D => n3338, CK =>
                           CLK, Q => n_1083, QN => 
                           DataPath_WRF_CUhw_curr_data_19_port);
   DataPath_WRF_CUhw_curr_data_reg_20_inst : DFF_X1 port map( D => n3337, CK =>
                           CLK, Q => n_1084, QN => 
                           DataPath_WRF_CUhw_curr_data_20_port);
   DataPath_WRF_CUhw_curr_data_reg_21_inst : DFF_X1 port map( D => n3336, CK =>
                           CLK, Q => n_1085, QN => 
                           DataPath_WRF_CUhw_curr_data_21_port);
   DataPath_WRF_CUhw_curr_data_reg_22_inst : DFF_X1 port map( D => n3335, CK =>
                           CLK, Q => n_1086, QN => 
                           DataPath_WRF_CUhw_curr_data_22_port);
   DataPath_WRF_CUhw_curr_data_reg_23_inst : DFF_X1 port map( D => n3334, CK =>
                           CLK, Q => n_1087, QN => 
                           DataPath_WRF_CUhw_curr_data_23_port);
   DataPath_WRF_CUhw_curr_data_reg_24_inst : DFF_X1 port map( D => n3333, CK =>
                           CLK, Q => n_1088, QN => 
                           DataPath_WRF_CUhw_curr_data_24_port);
   DataPath_WRF_CUhw_curr_data_reg_25_inst : DFF_X1 port map( D => n3332, CK =>
                           CLK, Q => n_1089, QN => 
                           DataPath_WRF_CUhw_curr_data_25_port);
   DataPath_WRF_CUhw_curr_data_reg_26_inst : DFF_X1 port map( D => n3331, CK =>
                           CLK, Q => n_1090, QN => 
                           DataPath_WRF_CUhw_curr_data_26_port);
   DataPath_WRF_CUhw_curr_data_reg_27_inst : DFF_X1 port map( D => n3330, CK =>
                           CLK, Q => n_1091, QN => 
                           DataPath_WRF_CUhw_curr_data_27_port);
   DataPath_WRF_CUhw_curr_data_reg_28_inst : DFF_X1 port map( D => n3329, CK =>
                           CLK, Q => n_1092, QN => 
                           DataPath_WRF_CUhw_curr_data_28_port);
   DataPath_WRF_CUhw_curr_data_reg_29_inst : DFF_X1 port map( D => n3328, CK =>
                           CLK, Q => n_1093, QN => 
                           DataPath_WRF_CUhw_curr_data_29_port);
   DataPath_WRF_CUhw_curr_data_reg_30_inst : DFF_X1 port map( D => n3327, CK =>
                           CLK, Q => n_1094, QN => 
                           DataPath_WRF_CUhw_curr_data_30_port);
   DataPath_WRF_CUhw_curr_data_reg_31_inst : DFF_X1 port map( D => n3324, CK =>
                           CLK, Q => n_1095, QN => 
                           DataPath_WRF_CUhw_curr_data_31_port);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_0_inst : DFF_X1 port map( D => 
                           n7152, CK => CLK, Q => n8328, QN => n543);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_1_inst : DFF_X1 port map( D => 
                           n7151, CK => CLK, Q => n_1096, QN => n544);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_3_inst : DFF_X1 port map( D => 
                           n7149, CK => CLK, Q => n_1097, QN => n546);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_4_inst : DFF_X1 port map( D => 
                           n7148, CK => CLK, Q => DECODEhw_i_tickcounter_4_port
                           , QN => n_1098);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_5_inst : DFF_X1 port map( D => 
                           n7147, CK => CLK, Q => n_1099, QN => n548);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_6_inst : DFF_X1 port map( D => 
                           n7146, CK => CLK, Q => DECODEhw_i_tickcounter_6_port
                           , QN => n_1100);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_7_inst : DFF_X1 port map( D => 
                           n7145, CK => CLK, Q => n_1101, QN => n550);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_8_inst : DFF_X1 port map( D => 
                           n7144, CK => CLK, Q => DECODEhw_i_tickcounter_8_port
                           , QN => n_1102);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_9_inst : DFF_X1 port map( D => 
                           n7143, CK => CLK, Q => n_1103, QN => n552);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_10_inst : DFF_X1 port map( D => 
                           n7142, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_10_port, QN => n_1104);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_11_inst : DFF_X1 port map( D => 
                           n7141, CK => CLK, Q => n8330, QN => n554);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_12_inst : DFF_X1 port map( D => 
                           n7140, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_12_port, QN => n_1105);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_13_inst : DFF_X1 port map( D => 
                           n7139, CK => CLK, Q => n_1106, QN => n556);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_14_inst : DFF_X1 port map( D => 
                           n7138, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_14_port, QN => n_1107);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_15_inst : DFF_X1 port map( D => 
                           n7137, CK => CLK, Q => n8331, QN => n558);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_16_inst : DFF_X1 port map( D => 
                           n7136, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_16_port, QN => n8368);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_17_inst : DFF_X1 port map( D => 
                           n7135, CK => CLK, Q => n_1108, QN => n560);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_18_inst : DFF_X1 port map( D => 
                           n7134, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_18_port, QN => n8375);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_19_inst : DFF_X1 port map( D => 
                           n7133, CK => CLK, Q => n_1109, QN => n562);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_20_inst : DFF_X1 port map( D => 
                           n7132, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_20_port, QN => n8369);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_21_inst : DFF_X1 port map( D => 
                           n7131, CK => CLK, Q => n_1110, QN => n564);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_22_inst : DFF_X1 port map( D => 
                           n7130, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_22_port, QN => n8374);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_23_inst : DFF_X1 port map( D => 
                           n7129, CK => CLK, Q => n_1111, QN => n566);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_24_inst : DFF_X1 port map( D => 
                           n7128, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_24_port, QN => n8373);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_25_inst : DFF_X1 port map( D => 
                           n7127, CK => CLK, Q => n_1112, QN => n568);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_26_inst : DFF_X1 port map( D => 
                           n7126, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_26_port, QN => n8370);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_27_inst : DFF_X1 port map( D => 
                           n7125, CK => CLK, Q => n_1113, QN => n570);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_28_inst : DFF_X1 port map( D => 
                           n7124, CK => CLK, Q => n_1114, QN => n571);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_29_inst : DFF_X1 port map( D => 
                           n3280, CK => CLK, Q => n8334, QN => 
                           DECODEhw_i_tickcounter_29_port);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_30_inst : DFF_X1 port map( D => 
                           n7123, CK => CLK, Q => n_1115, QN => n572);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_31_inst : DFF_X1 port map( D => 
                           n7153, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_31_port, QN => n8372);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_15_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N61, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_15_port, QN => 
                           n_1116);
   DataPath_RF_BLOCKi_72_Q_reg_0_inst : DFF_X1 port map( D => n5900, CK => CLK,
                           Q => n_1117, QN => 
                           DataPath_RF_bus_reg_dataout_2048_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_31_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N35, Q => i_RD2_31_port
                           );
   DataPath_REG_B_Q_reg_31_inst : DFF_X1 port map( D => n2844, CK => CLK, Q => 
                           n8404, QN => DataPath_i_PIPLIN_B_31_port);
   DataPath_REG_ME_Q_reg_31_inst : DFF_X1 port map( D => n2813, CK => CLK, Q =>
                           n_1118, QN => DataPath_i_REG_ME_DATA_DATAMEM_31_port
                           );
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_10_inst : DFF_X1 port map( D => n2308, CK 
                           => CLK, Q => n_1119, QN => 
                           DataPath_i_REG_LDSTR_OUT_10_port);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_10_inst : DFF_X1 port map( D => n6981, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_234_port
                           , QN => n798);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_31_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N35, Q => i_RD1_31_port
                           );
   CU_I_CW_ID_reg_24_inst : DLL_X1 port map( D => CU_I_CW_24_port, GN => n7768,
                           Q => i_RF2);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_0_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N4, Q => i_RD2_0_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_1_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N5, Q => i_RD2_1_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_2_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N6, Q => i_RD2_2_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_3_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N7, Q => i_RD2_3_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_4_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N8, Q => i_RD2_4_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_5_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N9, Q => i_RD2_5_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_6_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N10, Q => i_RD2_6_port)
                           ;
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_7_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N11, Q => i_RD2_7_port)
                           ;
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_8_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N12, Q => i_RD2_8_port)
                           ;
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_9_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N13, Q => i_RD2_9_port)
                           ;
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_10_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N14, Q => i_RD2_10_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_11_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N15, Q => i_RD2_11_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_12_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N16, Q => i_RD2_12_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_13_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N17, Q => i_RD2_13_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_14_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N18, Q => i_RD2_14_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_15_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N19, Q => i_RD2_15_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_16_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N20, Q => i_RD2_16_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_17_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N21, Q => i_RD2_17_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_18_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N22, Q => i_RD2_18_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_19_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N23, Q => i_RD2_19_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_20_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N24, Q => i_RD2_20_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_21_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N25, Q => i_RD2_21_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_22_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N26, Q => i_RD2_22_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_23_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N27, Q => i_RD2_23_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_24_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N28, Q => i_RD2_24_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_25_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N29, Q => i_RD2_25_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_26_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N30, Q => i_RD2_26_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_27_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N31, Q => i_RD2_27_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_28_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N32, Q => i_RD2_28_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_29_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N33, Q => i_RD2_29_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_30_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N34, Q => i_RD2_30_port
                           );
   IR_reg_20_inst : DFFR_X1 port map( D => n7115, CK => CLK, RN => n8694, Q => 
                           n_1120, QN => n189);
   IR_reg_19_inst : DFFR_X1 port map( D => n7116, CK => CLK, RN => n8691, Q => 
                           n_1121, QN => n190);
   IR_reg_18_inst : DFFR_X1 port map( D => n7117, CK => CLK, RN => n8691, Q => 
                           n_1122, QN => n191);
   IR_reg_17_inst : DFFR_X1 port map( D => n7118, CK => CLK, RN => n8691, Q => 
                           n_1123, QN => n192);
   IR_reg_16_inst : DFFR_X1 port map( D => n7119, CK => CLK, RN => n8691, Q => 
                           n_1124, QN => n193);
   IR_reg_8_inst : DFFS_X1 port map( D => n3010, CK => CLK, SN => n8693, Q => 
                           n8324, QN => IR_8_port);
   IR_reg_10_inst : DFFS_X1 port map( D => n3009, CK => CLK, SN => n8693, Q => 
                           n8323, QN => IR_10_port);
   IR_reg_13_inst : DFFS_X1 port map( D => n3006, CK => CLK, SN => n8693, Q => 
                           n8406, QN => IR_13_port);
   CU_I_CW_ID_reg_2_inst : DLL_X1 port map( D => n10836, GN => n7768, Q => 
                           CU_I_CW_ID_2_port);
   CU_I_CW_EX_reg_2_inst : DFF_X1 port map( D => n2960, CK => CLK, Q => n_1125,
                           QN => CU_I_CW_EX_2_port);
   CU_I_CW_MEM_reg_2_inst : DFF_X1 port map( D => n2953, CK => CLK, Q => n_1126
                           , QN => CU_I_CW_MEM_2_port);
   CU_I_setcmp_1_reg_2_inst : DFF_X1 port map( D => n7080, CK => CLK, Q => 
                           n_1127, QN => n235);
   CU_I_aluOpcode1_reg_0_inst : DFF_X1 port map( D => n7087, CK => CLK, Q => 
                           i_ALU_OP_0_port, QN => n8400);
   CU_I_aluOpcode1_reg_1_inst : DFF_X1 port map( D => n7086, CK => CLK, Q => 
                           i_ALU_OP_1_port, QN => n_1128);
   CU_I_aluOpcode1_reg_3_inst : DFF_X1 port map( D => n7084, CK => CLK, Q => 
                           i_ALU_OP_3_port, QN => n8319);
   CU_I_setcmp_1_reg_0_inst : DFF_X1 port map( D => n7082, CK => CLK, Q => 
                           i_SEL_LGET_0_port, QN => n8438);
   CU_I_setcmp_1_reg_1_inst : DFF_X1 port map( D => n7081, CK => CLK, Q => 
                           i_SEL_LGET_1_port, QN => n8378);
   CU_I_sel_alu_setcmp_1_reg : DFF_X1 port map( D => n7079, CK => CLK, Q => 
                           n_1129, QN => n8380);
   CU_I_i_FILL_delay_reg : DFF_X1 port map( D => n10845, CK => CLK, Q => 
                           CU_I_i_FILL_delay, QN => n_1130);
   DataPath_RF_POP_ADDRGEN_curr_state_reg_0_inst : DFF_X1 port map( D => n7061,
                           CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_state_0_port, QN => 
                           n_1131);
   DataPath_RF_POP_ADDRGEN_curr_state_reg_1_inst : DFF_X1 port map( D => n10844
                           , CK => CLK, Q => n_1132, QN => n851);
   DataPath_RF_CWP_Q_reg_4_inst : DFF_X1 port map( D => n7069, CK => CLK, Q => 
                           DataPath_RF_c_win_4_port, QN => n8441);
   CU_I_i_SPILL_delay_reg : DFF_X1 port map( D => CU_I_N184, CK => CLK, Q => 
                           CU_I_i_SPILL_delay, QN => n_1133);
   DataPath_RF_PUSH_ADDRGEN_curr_state_reg_1_inst : DFF_X1 port map( D => n7067
                           , CK => CLK, Q => n_1134, QN => n838);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_0_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N46, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, QN => 
                           n8437);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_1_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N47, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, QN => 
                           n_1135);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_2_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N48, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, QN => 
                           n_1136);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_3_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N49, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, QN => 
                           n_1137);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_4_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N50, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, QN => 
                           n_1138);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_5_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N51, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, QN => 
                           n_1139);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_6_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N52, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, QN => 
                           n_1140);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_7_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N53, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, QN => 
                           n_1141);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_8_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N54, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, QN => 
                           n_1142);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_9_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N55, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, QN => 
                           n_1143);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_10_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N56, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, QN => 
                           n_1144);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_11_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N57, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, QN => 
                           n_1145);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_12_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N58, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, QN => 
                           n_1146);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_13_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N59, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, QN => 
                           n_1147);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_14_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N60, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_14_port, QN => 
                           n_1148);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_15_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N61, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_15_port, QN => 
                           n8413);
   DataPath_RF_PUSH_ADDRGEN_curr_state_reg_0_inst : DFF_X1 port map( D => n7068
                           , CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_state_0_port, QN => 
                           n_1149);
   DataPath_RF_SWP_Q_reg_3_inst : DFF_X1 port map( D => n7063, CK => CLK, Q => 
                           DataPath_RF_c_swin_3_port, QN => n823);
   DataPath_RF_SWP_Q_reg_2_inst : DFF_X1 port map( D => n7064, CK => CLK, Q => 
                           DataPath_RF_c_swin_2_port, QN => n822);
   DataPath_RF_SWP_Q_reg_1_inst : DFF_X1 port map( D => n7065, CK => CLK, Q => 
                           DataPath_RF_c_swin_1_port, QN => n821);
   DataPath_RF_SWP_Q_reg_0_inst : DFF_X1 port map( D => n7066, CK => CLK, Q => 
                           DataPath_RF_c_swin_0_port, QN => n8327);
   DataPath_WRF_CUhw_curr_state_reg_1_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N145, CK => CLK, Q => n_1150, QN 
                           => n477);
   DataPath_WRF_CUhw_curr_state_reg_0_inst : DFF_X1 port map( D => n104, CK => 
                           CLK, Q => n8313, QN => n476);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_0_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N46, CK => CLK, Q => n8410, 
                           QN => n852);
   CU_I_CW_ID_reg_25_inst : DLL_X1 port map( D => CU_I_CW_25_port, GN => n7768,
                           Q => i_RF1);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_0_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N4, Q => i_RD1_0_port);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_1_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N5, Q => i_RD1_1_port);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_2_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N6, Q => i_RD1_2_port);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_3_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N7, Q => i_RD1_3_port);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_4_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N8, Q => i_RD1_4_port);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_5_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N9, Q => i_RD1_5_port);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_6_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N10, Q => i_RD1_6_port)
                           ;
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_7_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N11, Q => i_RD1_7_port)
                           ;
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_8_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N12, Q => i_RD1_8_port)
                           ;
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_9_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N13, Q => i_RD1_9_port)
                           ;
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_10_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N14, Q => i_RD1_10_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_11_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N15, Q => i_RD1_11_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_12_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N16, Q => i_RD1_12_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_13_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N17, Q => i_RD1_13_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_14_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N18, Q => i_RD1_14_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_15_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N19, Q => i_RD1_15_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_16_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N20, Q => i_RD1_16_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_17_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N21, Q => i_RD1_17_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_18_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N22, Q => i_RD1_18_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_19_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N23, Q => i_RD1_19_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_20_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N24, Q => i_RD1_20_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_21_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N25, Q => i_RD1_21_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_22_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N26, Q => i_RD1_22_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_23_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N27, Q => i_RD1_23_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_24_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N28, Q => i_RD1_24_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_25_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N29, Q => i_RD1_25_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_26_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N30, Q => i_RD1_26_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_27_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N31, Q => i_RD1_27_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_28_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N32, Q => i_RD1_28_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_29_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N33, Q => i_RD1_29_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_30_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N34, Q => i_RD1_30_port
                           );
   CU_I_CW_ID_reg_23_inst : DLL_X1 port map( D => CU_I_CW_23_port, GN => n7768,
                           Q => i_SEL_CMPB);
   CU_I_CW_ID_reg_22_inst : DLL_X1 port map( D => CU_I_CW_22_port, GN => n7768,
                           Q => CU_I_CW_ID_22);
   CU_I_unsigned_1_reg : DFF_X1 port map( D => n2876, CK => CLK, Q => n_1151, 
                           QN => CU_I_unsigned_1);
   CU_I_unsigned_2_reg : DFF_X1 port map( D => n2874, CK => CLK, Q => n8382, QN
                           => i_UNSIG_SIGN_N);
   CU_I_CW_ID_reg_21_inst : DLL_X1 port map( D => CU_I_CW_21_port, GN => n7768,
                           Q => i_NPC_SEL);
   PC_reg_7_inst : DFFR_X1 port map( D => n7052, CK => CLK, RN => n8690, Q => 
                           IRAM_ADDRESS_7_port, QN => n_1152);
   PC_reg_8_inst : DFFR_X1 port map( D => n7051, CK => CLK, RN => n8690, Q => 
                           IRAM_ADDRESS_8_port, QN => n_1153);
   PC_reg_17_inst : DFFR_X1 port map( D => n7042, CK => CLK, RN => n8690, Q => 
                           IRAM_ADDRESS_17_port, QN => n_1154);
   PC_reg_18_inst : DFFR_X1 port map( D => n7041, CK => CLK, RN => n8689, Q => 
                           IRAM_ADDRESS_18_port, QN => n_1155);
   PC_reg_25_inst : DFFR_X1 port map( D => n7034, CK => CLK, RN => n8689, Q => 
                           IRAM_ADDRESS_25_port, QN => n_1156);
   PC_reg_26_inst : DFFR_X1 port map( D => n7033, CK => CLK, RN => n8689, Q => 
                           IRAM_ADDRESS_26_port, QN => n_1157);
   PC_reg_27_inst : DFFR_X1 port map( D => n7032, CK => CLK, RN => n8689, Q => 
                           IRAM_ADDRESS_27_port, QN => n_1158);
   CU_I_CW_ID_reg_20_inst : DLL_X1 port map( D => n8440, GN => n7768, Q => n473
                           );
   CU_I_CW_ID_reg_17_inst : DLL_X1 port map( D => n10843, GN => n7768, Q => 
                           CU_I_CW_ID_17);
   CU_I_CW_EX_reg_17_inst : DFF_X1 port map( D => n7077, CK => CLK, Q => n8314,
                           QN => n472);
   CU_I_CW_ID_reg_16_inst : DLL_X1 port map( D => CU_I_CW_16_port, GN => n7768,
                           Q => CU_I_CW_ID_16);
   CU_I_CW_ID_reg_6_inst : DLL_X1 port map( D => CU_I_CW_6_port, GN => n7768, Q
                           => CU_I_CW_ID_6_port);
   CU_I_CW_EX_reg_6_inst : DFF_X1 port map( D => n2992, CK => CLK, Q => n_1159,
                           QN => CU_I_CW_EX_6_port);
   CU_I_CW_MEM_reg_6_inst : DFF_X1 port map( D => n382, CK => CLK, Q => 
                           i_DATAMEM_WM, QN => DRAM_READNOTWRITE);
   CU_I_CW_ID_reg_5_inst : DLL_X1 port map( D => CU_I_CW_5_port, GN => n7768, Q
                           => CU_I_CW_ID_5_port);
   CU_I_CW_EX_reg_5_inst : DFF_X1 port map( D => n2957, CK => CLK, Q => n_1160,
                           QN => CU_I_CW_EX_5_port);
   CU_I_CW_ID_reg_4_inst : DLL_X1 port map( D => CU_I_CW_4_port, GN => n7768, Q
                           => CU_I_CW_ID_4_port);
   CU_I_CW_EX_reg_4_inst : DFF_X1 port map( D => n2958, CK => CLK, Q => n_1161,
                           QN => CU_I_CW_EX_4_port);
   CU_I_CW_MEM_reg_4_inst : DFF_X1 port map( D => n384, CK => CLK, Q => 
                           DATA_SIZE_1_port, QN => n393);
   CU_I_CW_ID_reg_3_inst : DLL_X1 port map( D => CU_I_CW_3_port, GN => n7768, Q
                           => CU_I_CW_ID_3_port);
   CU_I_CW_EX_reg_3_inst : DFF_X1 port map( D => n2959, CK => CLK, Q => n_1162,
                           QN => CU_I_CW_EX_3_port);
   CU_I_CW_MEM_reg_3_inst : DFF_X1 port map( D => n383, CK => CLK, Q => 
                           DATA_SIZE_0_port, QN => n392);
   CU_I_CW_ID_reg_1_inst : DLL_X1 port map( D => CU_I_CW_5_port, GN => n7768, Q
                           => CU_I_CW_ID_1_port);
   CU_I_CW_EX_reg_1_inst : DFF_X1 port map( D => n2961, CK => CLK, Q => n_1163,
                           QN => CU_I_CW_EX_1_port);
   CU_I_CW_MEM_reg_1_inst : DFF_X1 port map( D => n2955, CK => CLK, Q => n_1164
                           , QN => CU_I_CW_MEM_1_port);
   CU_I_CW_WB_reg_1_inst : DFF_X1 port map( D => CU_I_N171, CK => CLK, Q => 
                           n8301, QN => n8411);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_7_inst : DFF_X1 port map( D => n2311, CK =>
                           CLK, Q => n_1165, QN => 
                           DataPath_i_REG_LDSTR_OUT_7_port);
   CU_I_CW_ID_reg_18_inst : DLL_X1 port map( D => n10836, GN => n7768, Q => 
                           CU_I_CW_ID_18);
   CU_I_CW_EX_reg_18_inst : DFF_X1 port map( D => n2887, CK => CLK, Q => n_1166
                           , QN => CU_I_CW_EX_18);
   CU_I_CW_ID_reg_19_inst : DLL_X1 port map( D => n10836, GN => n7768, Q => 
                           CU_I_CW_ID_19);
   DataPath_REG_IN2_Q_reg_16_inst : DFF_X1 port map( D => n7021, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_16_port, QN => n_1167);
   DataPath_REG_IN2_Q_reg_14_inst : DFF_X1 port map( D => n7022, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_14_port, QN => n8432);
   DataPath_REG_IN2_Q_reg_13_inst : DFF_X1 port map( D => n7023, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_13_port, QN => n_1168);
   DataPath_REG_IN2_Q_reg_10_inst : DFF_X1 port map( D => n7024, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_10_port, QN => n_1169);
   DataPath_REG_IN2_Q_reg_8_inst : DFF_X1 port map( D => n7025, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_8_port, QN => n8431);
   DataPath_REG_IN2_Q_reg_6_inst : DFF_X1 port map( D => n7026, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_6_port, QN => n_1170);
   DataPath_REG_IN2_Q_reg_3_inst : DFF_X1 port map( D => n7027, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_3_port, QN => n_1171);
   DataPath_REG_B_Q_reg_16_inst : DFF_X1 port map( D => n7075, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_16_port, QN => n_1172);
   DataPath_REG_ME_Q_reg_16_inst : DFF_X1 port map( D => n2828, CK => CLK, Q =>
                           n_1173, QN => DataPath_i_REG_ME_DATA_DATAMEM_16_port
                           );
   DataPath_REG_B_Q_reg_6_inst : DFF_X1 port map( D => n7076, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_6_port, QN => n_1174);
   DataPath_REG_ME_Q_reg_6_inst : DFF_X1 port map( D => n7074, CK => CLK, Q => 
                           DataPath_i_REG_ME_DATA_DATAMEM_6_port, QN => n_1175)
                           ;
   DataPath_REG_CMP_Q_reg_1_inst : DFF_X1 port map( D => n7104, CK => CLK, Q =>
                           n_1176, QN => n494);
   DataPath_REG_A_Q_reg_20_inst : DFF_X1 port map( D => n6730, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_20_port, QN => n8439);
   DataPath_REG_A_Q_reg_14_inst : DFF_X1 port map( D => n6731, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_14_port, QN => n_1177);
   DataPath_REG_A_Q_reg_13_inst : DFF_X1 port map( D => n6732, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_13_port, QN => n_1178);
   DataPath_REG_A_Q_reg_8_inst : DFF_X1 port map( D => n6733, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_8_port, QN => n_1179);
   DataPath_REG_A_Q_reg_3_inst : DFF_X1 port map( D => n6734, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_3_port, QN => n_1180);
   DataPath_REG_A_Q_reg_1_inst : DFF_X1 port map( D => n6735, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_1_port, QN => n_1181);
   DataPath_REG_A_Q_reg_0_inst : DFF_X1 port map( D => n3383, CK => CLK, Q => 
                           n_1182, QN => DataPath_i_PIPLIN_A_0_port);
   DataPath_REG_A_Q_reg_2_inst : DFF_X1 port map( D => n3382, CK => CLK, Q => 
                           n_1183, QN => DataPath_i_PIPLIN_A_2_port);
   DataPath_REG_A_Q_reg_4_inst : DFF_X1 port map( D => n3381, CK => CLK, Q => 
                           n_1184, QN => DataPath_i_PIPLIN_A_4_port);
   DataPath_REG_A_Q_reg_5_inst : DFF_X1 port map( D => n3380, CK => CLK, Q => 
                           n_1185, QN => DataPath_i_PIPLIN_A_5_port);
   DataPath_REG_A_Q_reg_6_inst : DFF_X1 port map( D => n3379, CK => CLK, Q => 
                           n_1186, QN => DataPath_i_PIPLIN_A_6_port);
   DataPath_REG_A_Q_reg_7_inst : DFF_X1 port map( D => n3378, CK => CLK, Q => 
                           n_1187, QN => DataPath_i_PIPLIN_A_7_port);
   DataPath_REG_A_Q_reg_9_inst : DFF_X1 port map( D => n3377, CK => CLK, Q => 
                           n_1188, QN => DataPath_i_PIPLIN_A_9_port);
   DataPath_REG_A_Q_reg_10_inst : DFF_X1 port map( D => n3376, CK => CLK, Q => 
                           n_1189, QN => DataPath_i_PIPLIN_A_10_port);
   DataPath_REG_A_Q_reg_11_inst : DFF_X1 port map( D => n3375, CK => CLK, Q => 
                           n_1190, QN => DataPath_i_PIPLIN_A_11_port);
   DataPath_REG_A_Q_reg_12_inst : DFF_X1 port map( D => n3374, CK => CLK, Q => 
                           n_1191, QN => DataPath_i_PIPLIN_A_12_port);
   DataPath_REG_A_Q_reg_15_inst : DFF_X1 port map( D => n3373, CK => CLK, Q => 
                           n_1192, QN => DataPath_i_PIPLIN_A_15_port);
   DataPath_REG_A_Q_reg_16_inst : DFF_X1 port map( D => n3372, CK => CLK, Q => 
                           n_1193, QN => DataPath_i_PIPLIN_A_16_port);
   DataPath_REG_A_Q_reg_17_inst : DFF_X1 port map( D => n3371, CK => CLK, Q => 
                           n_1194, QN => DataPath_i_PIPLIN_A_17_port);
   DataPath_REG_A_Q_reg_18_inst : DFF_X1 port map( D => n3370, CK => CLK, Q => 
                           n_1195, QN => DataPath_i_PIPLIN_A_18_port);
   DataPath_REG_A_Q_reg_19_inst : DFF_X1 port map( D => n3369, CK => CLK, Q => 
                           n_1196, QN => DataPath_i_PIPLIN_A_19_port);
   DataPath_REG_A_Q_reg_21_inst : DFF_X1 port map( D => n3368, CK => CLK, Q => 
                           n_1197, QN => DataPath_i_PIPLIN_A_21_port);
   DataPath_REG_A_Q_reg_22_inst : DFF_X1 port map( D => n3367, CK => CLK, Q => 
                           n_1198, QN => DataPath_i_PIPLIN_A_22_port);
   DataPath_REG_A_Q_reg_23_inst : DFF_X1 port map( D => n3366, CK => CLK, Q => 
                           n_1199, QN => DataPath_i_PIPLIN_A_23_port);
   DataPath_REG_A_Q_reg_24_inst : DFF_X1 port map( D => n3365, CK => CLK, Q => 
                           n_1200, QN => DataPath_i_PIPLIN_A_24_port);
   DataPath_REG_A_Q_reg_25_inst : DFF_X1 port map( D => n3364, CK => CLK, Q => 
                           n_1201, QN => DataPath_i_PIPLIN_A_25_port);
   DataPath_REG_A_Q_reg_26_inst : DFF_X1 port map( D => n3363, CK => CLK, Q => 
                           n_1202, QN => DataPath_i_PIPLIN_A_26_port);
   DataPath_REG_A_Q_reg_27_inst : DFF_X1 port map( D => n3362, CK => CLK, Q => 
                           n_1203, QN => DataPath_i_PIPLIN_A_27_port);
   DataPath_REG_A_Q_reg_28_inst : DFF_X1 port map( D => n3361, CK => CLK, Q => 
                           n_1204, QN => DataPath_i_PIPLIN_A_28_port);
   DataPath_REG_A_Q_reg_29_inst : DFF_X1 port map( D => n3360, CK => CLK, Q => 
                           n_1205, QN => DataPath_i_PIPLIN_A_29_port);
   DataPath_REG_A_Q_reg_30_inst : DFF_X1 port map( D => n3359, CK => CLK, Q => 
                           n_1206, QN => DataPath_i_PIPLIN_A_30_port);
   DataPath_REG_A_Q_reg_31_inst : DFF_X1 port map( D => n3358, CK => CLK, Q => 
                           n_1207, QN => DataPath_i_PIPLIN_A_31_port);
   DataPath_WRB1_Q_reg_0_inst : DFF_X1 port map( D => n2990, CK => CLK, Q => 
                           n_1208, QN => DataPath_i_PIPLIN_WRB1_0_port);
   DataPath_WRB2_Q_reg_0_inst : DFF_X1 port map( D => n2886, CK => CLK, Q => 
                           n_1209, QN => DataPath_i_PIPLIN_WRB2_0_port);
   DataPath_WRB3_Q_reg_0_inst : DFF_X1 port map( D => n372, CK => CLK, Q => 
                           i_ADD_WB_0_port, QN => n525);
   DataPath_WRB1_Q_reg_1_inst : DFF_X1 port map( D => n2989, CK => CLK, Q => 
                           n_1210, QN => DataPath_i_PIPLIN_WRB1_1_port);
   DataPath_WRB2_Q_reg_1_inst : DFF_X1 port map( D => n2885, CK => CLK, Q => 
                           n_1211, QN => DataPath_i_PIPLIN_WRB2_1_port);
   DataPath_WRB3_Q_reg_1_inst : DFF_X1 port map( D => n373, CK => CLK, Q => 
                           i_ADD_WB_1_port, QN => n526);
   DataPath_WRB1_Q_reg_2_inst : DFF_X1 port map( D => n2988, CK => CLK, Q => 
                           n_1212, QN => DataPath_i_PIPLIN_WRB1_2_port);
   DataPath_WRB2_Q_reg_2_inst : DFF_X1 port map( D => n2884, CK => CLK, Q => 
                           n_1213, QN => DataPath_i_PIPLIN_WRB2_2_port);
   DataPath_WRB3_Q_reg_2_inst : DFF_X1 port map( D => n374, CK => CLK, Q => 
                           i_ADD_WB_2_port, QN => n527);
   DataPath_WRB1_Q_reg_3_inst : DFF_X1 port map( D => n2987, CK => CLK, Q => 
                           n_1214, QN => DataPath_i_PIPLIN_WRB1_3_port);
   DataPath_WRB2_Q_reg_3_inst : DFF_X1 port map( D => n2883, CK => CLK, Q => 
                           n_1215, QN => DataPath_i_PIPLIN_WRB2_3_port);
   DataPath_WRB3_Q_reg_3_inst : DFF_X1 port map( D => n375, CK => CLK, Q => 
                           i_ADD_WB_3_port, QN => n_1216);
   DataPath_WRB1_Q_reg_4_inst : DFF_X1 port map( D => n2986, CK => CLK, Q => 
                           n_1217, QN => DataPath_i_PIPLIN_WRB1_4_port);
   DataPath_WRB2_Q_reg_4_inst : DFF_X1 port map( D => n2882, CK => CLK, Q => 
                           n_1218, QN => DataPath_i_PIPLIN_WRB2_4_port);
   DataPath_WRB3_Q_reg_4_inst : DFF_X1 port map( D => n376, CK => CLK, Q => 
                           i_ADD_WB_4_port, QN => n8310);
   DataPath_REG_CMP_Q_reg_0_inst : DFF_X1 port map( D => n116, CK => CLK, Q => 
                           DataPath_i_LGET_0_port, QN => n8386);
   DataPath_REG_IN1_Q_reg_0_inst : DFF_X1 port map( D => n2982, CK => CLK, Q =>
                           n8365, QN => DataPath_i_PIPLIN_IN1_0_port);
   DataPath_REG_IN1_Q_reg_1_inst : DFF_X1 port map( D => n2981, CK => CLK, Q =>
                           n_1219, QN => DataPath_i_PIPLIN_IN1_1_port);
   DataPath_REG_IN1_Q_reg_2_inst : DFF_X1 port map( D => n2977, CK => CLK, Q =>
                           n8436, QN => DataPath_i_PIPLIN_IN1_2_port);
   DataPath_REG_IN1_Q_reg_3_inst : DFF_X1 port map( D => n2976, CK => CLK, Q =>
                           n_1220, QN => DataPath_i_PIPLIN_IN1_3_port);
   DataPath_REG_IN1_Q_reg_4_inst : DFF_X1 port map( D => n2975, CK => CLK, Q =>
                           n8364, QN => DataPath_i_PIPLIN_IN1_4_port);
   DataPath_REG_IN1_Q_reg_5_inst : DFF_X1 port map( D => n2974, CK => CLK, Q =>
                           n8362, QN => DataPath_i_PIPLIN_IN1_5_port);
   DataPath_REG_IN1_Q_reg_6_inst : DFF_X1 port map( D => n2973, CK => CLK, Q =>
                           n8360, QN => DataPath_i_PIPLIN_IN1_6_port);
   DataPath_REG_IN1_Q_reg_7_inst : DFF_X1 port map( D => n2972, CK => CLK, Q =>
                           n8361, QN => DataPath_i_PIPLIN_IN1_7_port);
   DataPath_REG_IN1_Q_reg_8_inst : DFF_X1 port map( D => n2971, CK => CLK, Q =>
                           n_1221, QN => DataPath_i_PIPLIN_IN1_8_port);
   DataPath_REG_IN1_Q_reg_9_inst : DFF_X1 port map( D => n2970, CK => CLK, Q =>
                           n8357, QN => DataPath_i_PIPLIN_IN1_9_port);
   DataPath_REG_IN1_Q_reg_10_inst : DFF_X1 port map( D => n2969, CK => CLK, Q 
                           => n8358, QN => DataPath_i_PIPLIN_IN1_10_port);
   DataPath_REG_IN1_Q_reg_11_inst : DFF_X1 port map( D => n2968, CK => CLK, Q 
                           => n8359, QN => DataPath_i_PIPLIN_IN1_11_port);
   DataPath_REG_IN1_Q_reg_12_inst : DFF_X1 port map( D => n2967, CK => CLK, Q 
                           => n8363, QN => DataPath_i_PIPLIN_IN1_12_port);
   DataPath_REG_IN1_Q_reg_13_inst : DFF_X1 port map( D => n2966, CK => CLK, Q 
                           => n_1222, QN => DataPath_i_PIPLIN_IN1_13_port);
   DataPath_REG_IN1_Q_reg_14_inst : DFF_X1 port map( D => n2965, CK => CLK, Q 
                           => n_1223, QN => DataPath_i_PIPLIN_IN1_14_port);
   DataPath_REG_IN1_Q_reg_15_inst : DFF_X1 port map( D => n2963, CK => CLK, Q 
                           => n_1224, QN => DataPath_i_PIPLIN_IN1_15_port);
   DataPath_REG_B_Q_reg_0_inst : DFF_X1 port map( D => n2873, CK => CLK, Q => 
                           n8337, QN => DataPath_i_PIPLIN_B_0_port);
   DataPath_REG_ME_Q_reg_0_inst : DFF_X1 port map( D => n2843, CK => CLK, Q => 
                           n_1225, QN => DataPath_i_REG_ME_DATA_DATAMEM_0_port)
                           ;
   DataPath_REG_B_Q_reg_1_inst : DFF_X1 port map( D => n2872, CK => CLK, Q => 
                           n_1226, QN => DataPath_i_PIPLIN_B_1_port);
   DataPath_REG_ME_Q_reg_1_inst : DFF_X1 port map( D => n2842, CK => CLK, Q => 
                           n_1227, QN => DataPath_i_REG_ME_DATA_DATAMEM_1_port)
                           ;
   DataPath_REG_B_Q_reg_2_inst : DFF_X1 port map( D => n2871, CK => CLK, Q => 
                           n8336, QN => DataPath_i_PIPLIN_B_2_port);
   DataPath_REG_ME_Q_reg_2_inst : DFF_X1 port map( D => n2841, CK => CLK, Q => 
                           n_1228, QN => DataPath_i_REG_ME_DATA_DATAMEM_2_port)
                           ;
   DataPath_REG_B_Q_reg_3_inst : DFF_X1 port map( D => n2870, CK => CLK, Q => 
                           n_1229, QN => DataPath_i_PIPLIN_B_3_port);
   DataPath_REG_ME_Q_reg_3_inst : DFF_X1 port map( D => n2840, CK => CLK, Q => 
                           n_1230, QN => DataPath_i_REG_ME_DATA_DATAMEM_3_port)
                           ;
   DataPath_REG_B_Q_reg_4_inst : DFF_X1 port map( D => n2869, CK => CLK, Q => 
                           n8335, QN => DataPath_i_PIPLIN_B_4_port);
   DataPath_REG_ME_Q_reg_4_inst : DFF_X1 port map( D => n2839, CK => CLK, Q => 
                           n_1231, QN => DataPath_i_REG_ME_DATA_DATAMEM_4_port)
                           ;
   DataPath_REG_B_Q_reg_5_inst : DFF_X1 port map( D => n2868, CK => CLK, Q => 
                           n8338, QN => DataPath_i_PIPLIN_B_5_port);
   DataPath_REG_ME_Q_reg_5_inst : DFF_X1 port map( D => n2838, CK => CLK, Q => 
                           n_1232, QN => DataPath_i_REG_ME_DATA_DATAMEM_5_port)
                           ;
   DataPath_REG_B_Q_reg_7_inst : DFF_X1 port map( D => n2867, CK => CLK, Q => 
                           n8339, QN => DataPath_i_PIPLIN_B_7_port);
   DataPath_REG_ME_Q_reg_7_inst : DFF_X1 port map( D => n2837, CK => CLK, Q => 
                           n_1233, QN => DataPath_i_REG_ME_DATA_DATAMEM_7_port)
                           ;
   DataPath_REG_B_Q_reg_8_inst : DFF_X1 port map( D => n2866, CK => CLK, Q => 
                           n8341, QN => DataPath_i_PIPLIN_B_8_port);
   DataPath_REG_ME_Q_reg_8_inst : DFF_X1 port map( D => n2836, CK => CLK, Q => 
                           n_1234, QN => DataPath_i_REG_ME_DATA_DATAMEM_8_port)
                           ;
   DataPath_REG_B_Q_reg_9_inst : DFF_X1 port map( D => n2865, CK => CLK, Q => 
                           n8340, QN => DataPath_i_PIPLIN_B_9_port);
   DataPath_REG_ME_Q_reg_9_inst : DFF_X1 port map( D => n2835, CK => CLK, Q => 
                           n_1235, QN => DataPath_i_REG_ME_DATA_DATAMEM_9_port)
                           ;
   DataPath_REG_B_Q_reg_10_inst : DFF_X1 port map( D => n2864, CK => CLK, Q => 
                           n8343, QN => DataPath_i_PIPLIN_B_10_port);
   DataPath_REG_ME_Q_reg_10_inst : DFF_X1 port map( D => n2834, CK => CLK, Q =>
                           n_1236, QN => DataPath_i_REG_ME_DATA_DATAMEM_10_port
                           );
   DataPath_REG_B_Q_reg_11_inst : DFF_X1 port map( D => n2863, CK => CLK, Q => 
                           n8342, QN => DataPath_i_PIPLIN_B_11_port);
   DataPath_REG_ME_Q_reg_11_inst : DFF_X1 port map( D => n2833, CK => CLK, Q =>
                           n_1237, QN => DataPath_i_REG_ME_DATA_DATAMEM_11_port
                           );
   DataPath_REG_B_Q_reg_12_inst : DFF_X1 port map( D => n2862, CK => CLK, Q => 
                           n8345, QN => DataPath_i_PIPLIN_B_12_port);
   DataPath_REG_ME_Q_reg_12_inst : DFF_X1 port map( D => n2832, CK => CLK, Q =>
                           n_1238, QN => DataPath_i_REG_ME_DATA_DATAMEM_12_port
                           );
   DataPath_REG_B_Q_reg_13_inst : DFF_X1 port map( D => n2861, CK => CLK, Q => 
                           n8344, QN => DataPath_i_PIPLIN_B_13_port);
   DataPath_REG_ME_Q_reg_13_inst : DFF_X1 port map( D => n2831, CK => CLK, Q =>
                           n_1239, QN => DataPath_i_REG_ME_DATA_DATAMEM_13_port
                           );
   DataPath_REG_B_Q_reg_14_inst : DFF_X1 port map( D => n2860, CK => CLK, Q => 
                           n8347, QN => DataPath_i_PIPLIN_B_14_port);
   DataPath_REG_ME_Q_reg_14_inst : DFF_X1 port map( D => n2830, CK => CLK, Q =>
                           n_1240, QN => DataPath_i_REG_ME_DATA_DATAMEM_14_port
                           );
   DataPath_REG_B_Q_reg_15_inst : DFF_X1 port map( D => n2859, CK => CLK, Q => 
                           n8346, QN => DataPath_i_PIPLIN_B_15_port);
   DataPath_REG_ME_Q_reg_15_inst : DFF_X1 port map( D => n2829, CK => CLK, Q =>
                           n_1241, QN => DataPath_i_REG_ME_DATA_DATAMEM_15_port
                           );
   DataPath_REG_B_Q_reg_17_inst : DFF_X1 port map( D => n2858, CK => CLK, Q => 
                           n8348, QN => DataPath_i_PIPLIN_B_17_port);
   DataPath_REG_ME_Q_reg_17_inst : DFF_X1 port map( D => n2827, CK => CLK, Q =>
                           n_1242, QN => DataPath_i_REG_ME_DATA_DATAMEM_17_port
                           );
   DataPath_REG_B_Q_reg_18_inst : DFF_X1 port map( D => n2857, CK => CLK, Q => 
                           n8350, QN => DataPath_i_PIPLIN_B_18_port);
   DataPath_REG_ME_Q_reg_18_inst : DFF_X1 port map( D => n2826, CK => CLK, Q =>
                           n_1243, QN => DataPath_i_REG_ME_DATA_DATAMEM_18_port
                           );
   DataPath_REG_B_Q_reg_19_inst : DFF_X1 port map( D => n2856, CK => CLK, Q => 
                           n8349, QN => DataPath_i_PIPLIN_B_19_port);
   DataPath_REG_ME_Q_reg_19_inst : DFF_X1 port map( D => n2825, CK => CLK, Q =>
                           n_1244, QN => DataPath_i_REG_ME_DATA_DATAMEM_19_port
                           );
   DataPath_REG_B_Q_reg_20_inst : DFF_X1 port map( D => n2855, CK => CLK, Q => 
                           n8351, QN => DataPath_i_PIPLIN_B_20_port);
   DataPath_REG_ME_Q_reg_20_inst : DFF_X1 port map( D => n2824, CK => CLK, Q =>
                           n_1245, QN => DataPath_i_REG_ME_DATA_DATAMEM_20_port
                           );
   DataPath_REG_B_Q_reg_21_inst : DFF_X1 port map( D => n2854, CK => CLK, Q => 
                           n8321, QN => DataPath_i_PIPLIN_B_21_port);
   DataPath_REG_ME_Q_reg_21_inst : DFF_X1 port map( D => n2823, CK => CLK, Q =>
                           n_1246, QN => DataPath_i_REG_ME_DATA_DATAMEM_21_port
                           );
   DataPath_REG_B_Q_reg_22_inst : DFF_X1 port map( D => n2853, CK => CLK, Q => 
                           n8353, QN => DataPath_i_PIPLIN_B_22_port);
   DataPath_REG_ME_Q_reg_22_inst : DFF_X1 port map( D => n2822, CK => CLK, Q =>
                           n_1247, QN => DataPath_i_REG_ME_DATA_DATAMEM_22_port
                           );
   DataPath_REG_B_Q_reg_23_inst : DFF_X1 port map( D => n2852, CK => CLK, Q => 
                           n8352, QN => DataPath_i_PIPLIN_B_23_port);
   DataPath_REG_ME_Q_reg_23_inst : DFF_X1 port map( D => n2821, CK => CLK, Q =>
                           n_1248, QN => DataPath_i_REG_ME_DATA_DATAMEM_23_port
                           );
   DataPath_REG_B_Q_reg_24_inst : DFF_X1 port map( D => n2851, CK => CLK, Q => 
                           n8354, QN => DataPath_i_PIPLIN_B_24_port);
   DataPath_REG_ME_Q_reg_24_inst : DFF_X1 port map( D => n2820, CK => CLK, Q =>
                           n_1249, QN => DataPath_i_REG_ME_DATA_DATAMEM_24_port
                           );
   DataPath_REG_B_Q_reg_25_inst : DFF_X1 port map( D => n2850, CK => CLK, Q => 
                           n8322, QN => DataPath_i_PIPLIN_B_25_port);
   DataPath_REG_ME_Q_reg_25_inst : DFF_X1 port map( D => n2819, CK => CLK, Q =>
                           n_1250, QN => DataPath_i_REG_ME_DATA_DATAMEM_25_port
                           );
   DataPath_REG_B_Q_reg_26_inst : DFF_X1 port map( D => n2849, CK => CLK, Q => 
                           n8356, QN => DataPath_i_PIPLIN_B_26_port);
   DataPath_REG_ME_Q_reg_26_inst : DFF_X1 port map( D => n2818, CK => CLK, Q =>
                           n_1251, QN => DataPath_i_REG_ME_DATA_DATAMEM_26_port
                           );
   DataPath_REG_B_Q_reg_27_inst : DFF_X1 port map( D => n2848, CK => CLK, Q => 
                           n8355, QN => DataPath_i_PIPLIN_B_27_port);
   DataPath_REG_ME_Q_reg_27_inst : DFF_X1 port map( D => n2817, CK => CLK, Q =>
                           n_1252, QN => DataPath_i_REG_ME_DATA_DATAMEM_27_port
                           );
   DataPath_REG_B_Q_reg_28_inst : DFF_X1 port map( D => n2847, CK => CLK, Q => 
                           n8403, QN => DataPath_i_PIPLIN_B_28_port);
   DataPath_REG_ME_Q_reg_28_inst : DFF_X1 port map( D => n2816, CK => CLK, Q =>
                           n_1253, QN => DataPath_i_REG_ME_DATA_DATAMEM_28_port
                           );
   DataPath_REG_B_Q_reg_29_inst : DFF_X1 port map( D => n2846, CK => CLK, Q => 
                           n8402, QN => DataPath_i_PIPLIN_B_29_port);
   DataPath_REG_ME_Q_reg_29_inst : DFF_X1 port map( D => n2815, CK => CLK, Q =>
                           n_1254, QN => DataPath_i_REG_ME_DATA_DATAMEM_29_port
                           );
   DataPath_REG_B_Q_reg_30_inst : DFF_X1 port map( D => n2845, CK => CLK, Q => 
                           n8405, QN => DataPath_i_PIPLIN_B_30_port);
   DataPath_REG_ME_Q_reg_30_inst : DFF_X1 port map( D => n2814, CK => CLK, Q =>
                           n_1255, QN => DataPath_i_REG_ME_DATA_DATAMEM_30_port
                           );
   DataPath_REG_IN2_Q_reg_0_inst : DFF_X1 port map( D => n2498, CK => CLK, Q =>
                           n_1256, QN => DataPath_i_PIPLIN_IN2_0_port);
   DataPath_REG_IN2_Q_reg_1_inst : DFF_X1 port map( D => n2496, CK => CLK, Q =>
                           n8333, QN => DataPath_i_PIPLIN_IN2_1_port);
   DataPath_REG_IN2_Q_reg_2_inst : DFF_X1 port map( D => n2494, CK => CLK, Q =>
                           n_1257, QN => DataPath_i_PIPLIN_IN2_2_port);
   DataPath_REG_IN2_Q_reg_4_inst : DFF_X1 port map( D => n2491, CK => CLK, Q =>
                           n8435, QN => DataPath_i_PIPLIN_IN2_4_port);
   DataPath_REG_ALU_OUT_Q_reg_0_inst : DFF_X1 port map( D => n7020, CK => CLK, 
                           Q => n8388, QN => n495);
   DataPath_REG_MEM_ALUOUT_Q_reg_0_inst : DFF_X1 port map( D => n1258, CK => 
                           CLK, Q => n_1258, QN => 
                           DataPath_i_REG_MEM_ALUOUT_0_port);
   DataPath_REG_ALU_OUT_Q_reg_1_inst : DFF_X1 port map( D => n7019, CK => CLK, 
                           Q => n8376, QN => n496);
   DataPath_REG_MEM_ALUOUT_Q_reg_1_inst : DFF_X1 port map( D => n1257, CK => 
                           CLK, Q => n_1259, QN => 
                           DataPath_i_REG_MEM_ALUOUT_1_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_23_inst : DFF_X1 port map( D => n2295, CK 
                           => CLK, Q => n_1260, QN => 
                           DataPath_i_REG_LDSTR_OUT_23_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_31_inst : DFF_X1 port map( D => n2287, CK 
                           => CLK, Q => n_1261, QN => 
                           DataPath_i_REG_LDSTR_OUT_31_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_15_inst : DFF_X1 port map( D => n2303, CK 
                           => CLK, Q => n_1262, QN => 
                           DataPath_i_REG_LDSTR_OUT_15_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_17_inst : DFF_X1 port map( D => n2301, CK 
                           => CLK, Q => n_1263, QN => 
                           DataPath_i_REG_LDSTR_OUT_17_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_25_inst : DFF_X1 port map( D => n2293, CK 
                           => CLK, Q => n_1264, QN => 
                           DataPath_i_REG_LDSTR_OUT_25_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_9_inst : DFF_X1 port map( D => n2309, CK =>
                           CLK, Q => n_1265, QN => 
                           DataPath_i_REG_LDSTR_OUT_9_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_1_inst : DFF_X1 port map( D => n2317, CK =>
                           CLK, Q => n_1266, QN => 
                           DataPath_i_REG_LDSTR_OUT_1_port);
   DataPath_RF_BLOCKi_72_Q_reg_1_inst : DFF_X1 port map( D => n5899, CK => CLK,
                           Q => n_1267, QN => 
                           DataPath_RF_bus_reg_dataout_2049_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_14_inst : DFF_X1 port map( D => n2304, CK 
                           => CLK, Q => n_1268, QN => 
                           DataPath_i_REG_LDSTR_OUT_14_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_22_inst : DFF_X1 port map( D => n2296, CK 
                           => CLK, Q => n_1269, QN => 
                           DataPath_i_REG_LDSTR_OUT_22_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_30_inst : DFF_X1 port map( D => n2288, CK 
                           => CLK, Q => n_1270, QN => 
                           DataPath_i_REG_LDSTR_OUT_30_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_6_inst : DFF_X1 port map( D => n2312, CK =>
                           CLK, Q => n_1271, QN => 
                           DataPath_i_REG_LDSTR_OUT_6_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_13_inst : DFF_X1 port map( D => n2305, CK 
                           => CLK, Q => n_1272, QN => 
                           DataPath_i_REG_LDSTR_OUT_13_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_21_inst : DFF_X1 port map( D => n2297, CK 
                           => CLK, Q => n_1273, QN => 
                           DataPath_i_REG_LDSTR_OUT_21_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_29_inst : DFF_X1 port map( D => n2289, CK 
                           => CLK, Q => n_1274, QN => 
                           DataPath_i_REG_LDSTR_OUT_29_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_5_inst : DFF_X1 port map( D => n2313, CK =>
                           CLK, Q => n_1275, QN => 
                           DataPath_i_REG_LDSTR_OUT_5_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_12_inst : DFF_X1 port map( D => n2306, CK 
                           => CLK, Q => n_1276, QN => 
                           DataPath_i_REG_LDSTR_OUT_12_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_20_inst : DFF_X1 port map( D => n2298, CK 
                           => CLK, Q => n_1277, QN => 
                           DataPath_i_REG_LDSTR_OUT_20_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_28_inst : DFF_X1 port map( D => n2290, CK 
                           => CLK, Q => n_1278, QN => 
                           DataPath_i_REG_LDSTR_OUT_28_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_4_inst : DFF_X1 port map( D => n2314, CK =>
                           CLK, Q => n_1279, QN => 
                           DataPath_i_REG_LDSTR_OUT_4_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_11_inst : DFF_X1 port map( D => n2307, CK 
                           => CLK, Q => n_1280, QN => 
                           DataPath_i_REG_LDSTR_OUT_11_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_19_inst : DFF_X1 port map( D => n2299, CK 
                           => CLK, Q => n_1281, QN => 
                           DataPath_i_REG_LDSTR_OUT_19_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_27_inst : DFF_X1 port map( D => n2291, CK 
                           => CLK, Q => n_1282, QN => 
                           DataPath_i_REG_LDSTR_OUT_27_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_3_inst : DFF_X1 port map( D => n2315, CK =>
                           CLK, Q => n_1283, QN => 
                           DataPath_i_REG_LDSTR_OUT_3_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_18_inst : DFF_X1 port map( D => n2300, CK 
                           => CLK, Q => n_1284, QN => 
                           DataPath_i_REG_LDSTR_OUT_18_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_26_inst : DFF_X1 port map( D => n2292, CK 
                           => CLK, Q => n_1285, QN => 
                           DataPath_i_REG_LDSTR_OUT_26_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_2_inst : DFF_X1 port map( D => n2316, CK =>
                           CLK, Q => n_1286, QN => 
                           DataPath_i_REG_LDSTR_OUT_2_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_16_inst : DFF_X1 port map( D => n2302, CK 
                           => CLK, Q => n_1287, QN => 
                           DataPath_i_REG_LDSTR_OUT_16_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_24_inst : DFF_X1 port map( D => n2294, CK 
                           => CLK, Q => n_1288, QN => 
                           DataPath_i_REG_LDSTR_OUT_24_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_8_inst : DFF_X1 port map( D => n2310, CK =>
                           CLK, Q => n_1289, QN => 
                           DataPath_i_REG_LDSTR_OUT_8_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_0_inst : DFF_X1 port map( D => n2318, CK =>
                           CLK, Q => n_1290, QN => 
                           DataPath_i_REG_LDSTR_OUT_0_port);
   DataPath_REG_ALU_OUT_Q_reg_3_inst : DFF_X1 port map( D => n2228, CK => CLK, 
                           Q => n_1291, QN => DRAM_ADDRESS_3_port);
   DataPath_REG_MEM_ALUOUT_Q_reg_3_inst : DFF_X1 port map( D => n1255, CK => 
                           CLK, Q => n_1292, QN => 
                           DataPath_i_REG_MEM_ALUOUT_3_port);
   DataPath_RF_BLOCKi_72_Q_reg_3_inst : DFF_X1 port map( D => n5897, CK => CLK,
                           Q => n_1293, QN => 
                           DataPath_RF_bus_reg_dataout_2051_port);
   DataPath_REG_ALU_OUT_Q_reg_2_inst : DFF_X1 port map( D => n2260, CK => CLK, 
                           Q => n_1294, QN => DRAM_ADDRESS_2_port);
   DataPath_REG_MEM_ALUOUT_Q_reg_2_inst : DFF_X1 port map( D => n1256, CK => 
                           CLK, Q => n_1295, QN => 
                           DataPath_i_REG_MEM_ALUOUT_2_port);
   DataPath_RF_BLOCKi_72_Q_reg_2_inst : DFF_X1 port map( D => n5898, CK => CLK,
                           Q => n_1296, QN => 
                           DataPath_RF_bus_reg_dataout_2050_port);
   DataPath_REG_ALU_OUT_Q_reg_4_inst : DFF_X1 port map( D => n7018, CK => CLK, 
                           Q => DRAM_ADDRESS_4_port, QN => n497);
   DataPath_REG_MEM_ALUOUT_Q_reg_4_inst : DFF_X1 port map( D => n1254, CK => 
                           CLK, Q => n_1297, QN => 
                           DataPath_i_REG_MEM_ALUOUT_4_port);
   DataPath_RF_BLOCKi_72_Q_reg_4_inst : DFF_X1 port map( D => n5896, CK => CLK,
                           Q => n_1298, QN => 
                           DataPath_RF_bus_reg_dataout_2052_port);
   DataPath_REG_IN2_Q_reg_5_inst : DFF_X1 port map( D => n2489, CK => CLK, Q =>
                           n_1299, QN => DataPath_i_PIPLIN_IN2_5_port);
   DataPath_REG_ALU_OUT_Q_reg_6_inst : DFF_X1 port map( D => n7016, CK => CLK, 
                           Q => DRAM_ADDRESS_6_port, QN => n498);
   DataPath_REG_MEM_ALUOUT_Q_reg_6_inst : DFF_X1 port map( D => n1252, CK => 
                           CLK, Q => n_1300, QN => 
                           DataPath_i_REG_MEM_ALUOUT_6_port);
   DataPath_RF_BLOCKi_72_Q_reg_6_inst : DFF_X1 port map( D => n5894, CK => CLK,
                           Q => n_1301, QN => 
                           DataPath_RF_bus_reg_dataout_2054_port);
   DataPath_REG_ALU_OUT_Q_reg_5_inst : DFF_X1 port map( D => n7017, CK => CLK, 
                           Q => DRAM_ADDRESS_5_port, QN => n8434);
   DataPath_REG_MEM_ALUOUT_Q_reg_5_inst : DFF_X1 port map( D => n1253, CK => 
                           CLK, Q => n_1302, QN => 
                           DataPath_i_REG_MEM_ALUOUT_5_port);
   DataPath_RF_BLOCKi_72_Q_reg_5_inst : DFF_X1 port map( D => n5895, CK => CLK,
                           Q => n_1303, QN => 
                           DataPath_RF_bus_reg_dataout_2053_port);
   DataPath_REG_IN2_Q_reg_7_inst : DFF_X1 port map( D => n2486, CK => CLK, Q =>
                           n_1304, QN => DataPath_i_PIPLIN_IN2_7_port);
   DataPath_REG_ALU_OUT_Q_reg_8_inst : DFF_X1 port map( D => n7015, CK => CLK, 
                           Q => DRAM_ADDRESS_8_port, QN => n499);
   DataPath_REG_MEM_ALUOUT_Q_reg_8_inst : DFF_X1 port map( D => n1250, CK => 
                           CLK, Q => n_1305, QN => 
                           DataPath_i_REG_MEM_ALUOUT_8_port);
   DataPath_RF_BLOCKi_72_Q_reg_8_inst : DFF_X1 port map( D => n5892, CK => CLK,
                           Q => n_1306, QN => 
                           DataPath_RF_bus_reg_dataout_2056_port);
   DataPath_REG_ALU_OUT_Q_reg_7_inst : DFF_X1 port map( D => n2106, CK => CLK, 
                           Q => n_1307, QN => DRAM_ADDRESS_7_port);
   DataPath_REG_MEM_ALUOUT_Q_reg_7_inst : DFF_X1 port map( D => n1251, CK => 
                           CLK, Q => n_1308, QN => 
                           DataPath_i_REG_MEM_ALUOUT_7_port);
   DataPath_RF_BLOCKi_72_Q_reg_7_inst : DFF_X1 port map( D => n5893, CK => CLK,
                           Q => n_1309, QN => 
                           DataPath_RF_bus_reg_dataout_2055_port);
   DataPath_REG_IN2_Q_reg_9_inst : DFF_X1 port map( D => n2483, CK => CLK, Q =>
                           n_1310, QN => DataPath_i_PIPLIN_IN2_9_port);
   DataPath_REG_ALU_OUT_Q_reg_10_inst : DFF_X1 port map( D => n7013, CK => CLK,
                           Q => DRAM_ADDRESS_10_port, QN => n500);
   DataPath_REG_MEM_ALUOUT_Q_reg_10_inst : DFF_X1 port map( D => n1248, CK => 
                           CLK, Q => n_1311, QN => 
                           DataPath_i_REG_MEM_ALUOUT_10_port);
   DataPath_REG_ALU_OUT_Q_reg_9_inst : DFF_X1 port map( D => n7014, CK => CLK, 
                           Q => DRAM_ADDRESS_9_port, QN => n8433);
   DataPath_REG_MEM_ALUOUT_Q_reg_9_inst : DFF_X1 port map( D => n1249, CK => 
                           CLK, Q => n_1312, QN => 
                           DataPath_i_REG_MEM_ALUOUT_9_port);
   DataPath_RF_BLOCKi_72_Q_reg_9_inst : DFF_X1 port map( D => n5891, CK => CLK,
                           Q => n_1313, QN => 
                           DataPath_RF_bus_reg_dataout_2057_port);
   DataPath_REG_IN2_Q_reg_11_inst : DFF_X1 port map( D => n2480, CK => CLK, Q 
                           => n_1314, QN => DataPath_i_PIPLIN_IN2_11_port);
   DataPath_REG_ALU_OUT_Q_reg_11_inst : DFF_X1 port map( D => n7012, CK => CLK,
                           Q => DRAM_ADDRESS_11_port, QN => n501);
   DataPath_REG_MEM_ALUOUT_Q_reg_11_inst : DFF_X1 port map( D => n1247, CK => 
                           CLK, Q => n_1315, QN => 
                           DataPath_i_REG_MEM_ALUOUT_11_port);
   DataPath_RF_BLOCKi_72_Q_reg_11_inst : DFF_X1 port map( D => n5889, CK => CLK
                           , Q => n_1316, QN => 
                           DataPath_RF_bus_reg_dataout_2059_port);
   DataPath_REG_IN2_Q_reg_12_inst : DFF_X1 port map( D => n2478, CK => CLK, Q 
                           => n_1317, QN => DataPath_i_PIPLIN_IN2_12_port);
   DataPath_REG_ALU_OUT_Q_reg_14_inst : DFF_X1 port map( D => n7009, CK => CLK,
                           Q => DRAM_ADDRESS_14_port, QN => n503);
   DataPath_REG_MEM_ALUOUT_Q_reg_14_inst : DFF_X1 port map( D => n1244, CK => 
                           CLK, Q => n_1318, QN => 
                           DataPath_i_REG_MEM_ALUOUT_14_port);
   DataPath_RF_BLOCKi_72_Q_reg_14_inst : DFF_X1 port map( D => n5886, CK => CLK
                           , Q => n_1319, QN => 
                           DataPath_RF_bus_reg_dataout_2062_port);
   DataPath_REG_ALU_OUT_Q_reg_13_inst : DFF_X1 port map( D => n7010, CK => CLK,
                           Q => DRAM_ADDRESS_13_port, QN => n_1320);
   DataPath_REG_MEM_ALUOUT_Q_reg_13_inst : DFF_X1 port map( D => n1245, CK => 
                           CLK, Q => n_1321, QN => 
                           DataPath_i_REG_MEM_ALUOUT_13_port);
   DataPath_RF_BLOCKi_72_Q_reg_13_inst : DFF_X1 port map( D => n5887, CK => CLK
                           , Q => n_1322, QN => 
                           DataPath_RF_bus_reg_dataout_2061_port);
   DataPath_REG_ALU_OUT_Q_reg_12_inst : DFF_X1 port map( D => n7011, CK => CLK,
                           Q => DRAM_ADDRESS_12_port, QN => n502);
   DataPath_REG_MEM_ALUOUT_Q_reg_12_inst : DFF_X1 port map( D => n1246, CK => 
                           CLK, Q => n_1323, QN => 
                           DataPath_i_REG_MEM_ALUOUT_12_port);
   DataPath_RF_BLOCKi_72_Q_reg_12_inst : DFF_X1 port map( D => n5888, CK => CLK
                           , Q => n_1324, QN => 
                           DataPath_RF_bus_reg_dataout_2060_port);
   DataPath_REG_IN2_Q_reg_15_inst : DFF_X1 port map( D => n2474, CK => CLK, Q 
                           => n_1325, QN => DataPath_i_PIPLIN_IN2_15_port);
   DataPath_REG_ALU_OUT_Q_reg_16_inst : DFF_X1 port map( D => n7007, CK => CLK,
                           Q => DRAM_ADDRESS_16_port, QN => n505);
   DataPath_REG_MEM_ALUOUT_Q_reg_16_inst : DFF_X1 port map( D => n1242, CK => 
                           CLK, Q => n_1326, QN => 
                           DataPath_i_REG_MEM_ALUOUT_16_port);
   DataPath_RF_BLOCKi_72_Q_reg_16_inst : DFF_X1 port map( D => n5884, CK => CLK
                           , Q => n_1327, QN => 
                           DataPath_RF_bus_reg_dataout_2064_port);
   DataPath_REG_ALU_OUT_Q_reg_15_inst : DFF_X1 port map( D => n7008, CK => CLK,
                           Q => DRAM_ADDRESS_15_port, QN => n504);
   DataPath_REG_MEM_ALUOUT_Q_reg_15_inst : DFF_X1 port map( D => n1243, CK => 
                           CLK, Q => n_1328, QN => 
                           DataPath_i_REG_MEM_ALUOUT_15_port);
   DataPath_RF_BLOCKi_72_Q_reg_15_inst : DFF_X1 port map( D => n5885, CK => CLK
                           , Q => n_1329, QN => 
                           DataPath_RF_bus_reg_dataout_2063_port);
   DataPath_REG_IN2_Q_reg_17_inst : DFF_X1 port map( D => n2469, CK => CLK, Q 
                           => n_1330, QN => DataPath_i_PIPLIN_IN2_17_port);
   DataPath_REG_ALU_OUT_Q_reg_17_inst : DFF_X1 port map( D => n7006, CK => CLK,
                           Q => DRAM_ADDRESS_17_port, QN => n_1331);
   DataPath_REG_MEM_ALUOUT_Q_reg_17_inst : DFF_X1 port map( D => n1241, CK => 
                           CLK, Q => n_1332, QN => 
                           DataPath_i_REG_MEM_ALUOUT_17_port);
   DataPath_RF_BLOCKi_72_Q_reg_17_inst : DFF_X1 port map( D => n5883, CK => CLK
                           , Q => n_1333, QN => 
                           DataPath_RF_bus_reg_dataout_2065_port);
   DataPath_REG_IN2_Q_reg_18_inst : DFF_X1 port map( D => n2467, CK => CLK, Q 
                           => n_1334, QN => DataPath_i_PIPLIN_IN2_18_port);
   DataPath_REG_ALU_OUT_Q_reg_18_inst : DFF_X1 port map( D => n7005, CK => CLK,
                           Q => DRAM_ADDRESS_18_port, QN => n506);
   DataPath_REG_MEM_ALUOUT_Q_reg_18_inst : DFF_X1 port map( D => n1240, CK => 
                           CLK, Q => n_1335, QN => 
                           DataPath_i_REG_MEM_ALUOUT_18_port);
   DataPath_RF_BLOCKi_72_Q_reg_18_inst : DFF_X1 port map( D => n5882, CK => CLK
                           , Q => n_1336, QN => 
                           DataPath_RF_bus_reg_dataout_2066_port);
   DataPath_REG_IN2_Q_reg_19_inst : DFF_X1 port map( D => n2465, CK => CLK, Q 
                           => n_1337, QN => DataPath_i_PIPLIN_IN2_19_port);
   DataPath_REG_ALU_OUT_Q_reg_19_inst : DFF_X1 port map( D => n7004, CK => CLK,
                           Q => DRAM_ADDRESS_19_port, QN => n507);
   DataPath_REG_MEM_ALUOUT_Q_reg_19_inst : DFF_X1 port map( D => n1239, CK => 
                           CLK, Q => n_1338, QN => 
                           DataPath_i_REG_MEM_ALUOUT_19_port);
   DataPath_RF_BLOCKi_72_Q_reg_19_inst : DFF_X1 port map( D => n5881, CK => CLK
                           , Q => n_1339, QN => 
                           DataPath_RF_bus_reg_dataout_2067_port);
   DataPath_REG_IN2_Q_reg_20_inst : DFF_X1 port map( D => n2463, CK => CLK, Q 
                           => n_1340, QN => DataPath_i_PIPLIN_IN2_20_port);
   DataPath_REG_ALU_OUT_Q_reg_20_inst : DFF_X1 port map( D => n7003, CK => CLK,
                           Q => DRAM_ADDRESS_20_port, QN => n508);
   DataPath_REG_MEM_ALUOUT_Q_reg_20_inst : DFF_X1 port map( D => n1238, CK => 
                           CLK, Q => n_1341, QN => 
                           DataPath_i_REG_MEM_ALUOUT_20_port);
   DataPath_RF_BLOCKi_72_Q_reg_20_inst : DFF_X1 port map( D => n5880, CK => CLK
                           , Q => n_1342, QN => 
                           DataPath_RF_bus_reg_dataout_2068_port);
   DataPath_REG_IN2_Q_reg_21_inst : DFF_X1 port map( D => n2461, CK => CLK, Q 
                           => n_1343, QN => DataPath_i_PIPLIN_IN2_21_port);
   DataPath_REG_ALU_OUT_Q_reg_21_inst : DFF_X1 port map( D => n7002, CK => CLK,
                           Q => DRAM_ADDRESS_21_port, QN => n_1344);
   DataPath_REG_MEM_ALUOUT_Q_reg_21_inst : DFF_X1 port map( D => n1237, CK => 
                           CLK, Q => n_1345, QN => 
                           DataPath_i_REG_MEM_ALUOUT_21_port);
   DataPath_RF_BLOCKi_72_Q_reg_21_inst : DFF_X1 port map( D => n5879, CK => CLK
                           , Q => n_1346, QN => 
                           DataPath_RF_bus_reg_dataout_2069_port);
   DataPath_REG_IN2_Q_reg_22_inst : DFF_X1 port map( D => n2459, CK => CLK, Q 
                           => n_1347, QN => DataPath_i_PIPLIN_IN2_22_port);
   DataPath_REG_ALU_OUT_Q_reg_22_inst : DFF_X1 port map( D => n7001, CK => CLK,
                           Q => DRAM_ADDRESS_22_port, QN => n509);
   DataPath_REG_MEM_ALUOUT_Q_reg_22_inst : DFF_X1 port map( D => n1236, CK => 
                           CLK, Q => n_1348, QN => 
                           DataPath_i_REG_MEM_ALUOUT_22_port);
   DataPath_RF_BLOCKi_72_Q_reg_22_inst : DFF_X1 port map( D => n5878, CK => CLK
                           , Q => n_1349, QN => 
                           DataPath_RF_bus_reg_dataout_2070_port);
   DataPath_REG_IN2_Q_reg_23_inst : DFF_X1 port map( D => n2457, CK => CLK, Q 
                           => n_1350, QN => DataPath_i_PIPLIN_IN2_23_port);
   DataPath_REG_ALU_OUT_Q_reg_23_inst : DFF_X1 port map( D => n7000, CK => CLK,
                           Q => DRAM_ADDRESS_23_port, QN => n510);
   DataPath_REG_MEM_ALUOUT_Q_reg_23_inst : DFF_X1 port map( D => n1235, CK => 
                           CLK, Q => n_1351, QN => 
                           DataPath_i_REG_MEM_ALUOUT_23_port);
   DataPath_RF_BLOCKi_72_Q_reg_23_inst : DFF_X1 port map( D => n5877, CK => CLK
                           , Q => n_1352, QN => 
                           DataPath_RF_bus_reg_dataout_2071_port);
   DataPath_REG_IN2_Q_reg_24_inst : DFF_X1 port map( D => n2455, CK => CLK, Q 
                           => n_1353, QN => DataPath_i_PIPLIN_IN2_24_port);
   DataPath_REG_ALU_OUT_Q_reg_24_inst : DFF_X1 port map( D => n6999, CK => CLK,
                           Q => DRAM_ADDRESS_24_port, QN => n511);
   DataPath_REG_MEM_ALUOUT_Q_reg_24_inst : DFF_X1 port map( D => n1234, CK => 
                           CLK, Q => n_1354, QN => 
                           DataPath_i_REG_MEM_ALUOUT_24_port);
   DataPath_RF_BLOCKi_72_Q_reg_24_inst : DFF_X1 port map( D => n5876, CK => CLK
                           , Q => n_1355, QN => 
                           DataPath_RF_bus_reg_dataout_2072_port);
   DataPath_REG_IN2_Q_reg_25_inst : DFF_X1 port map( D => n2453, CK => CLK, Q 
                           => n_1356, QN => DataPath_i_PIPLIN_IN2_25_port);
   DataPath_REG_ALU_OUT_Q_reg_25_inst : DFF_X1 port map( D => n6998, CK => CLK,
                           Q => DRAM_ADDRESS_25_port, QN => n_1357);
   DataPath_REG_MEM_ALUOUT_Q_reg_25_inst : DFF_X1 port map( D => n1233, CK => 
                           CLK, Q => n_1358, QN => 
                           DataPath_i_REG_MEM_ALUOUT_25_port);
   DataPath_RF_BLOCKi_72_Q_reg_25_inst : DFF_X1 port map( D => n5875, CK => CLK
                           , Q => n_1359, QN => 
                           DataPath_RF_bus_reg_dataout_2073_port);
   DataPath_REG_IN2_Q_reg_26_inst : DFF_X1 port map( D => n2451, CK => CLK, Q 
                           => n_1360, QN => DataPath_i_PIPLIN_IN2_26_port);
   DataPath_REG_ALU_OUT_Q_reg_26_inst : DFF_X1 port map( D => n6997, CK => CLK,
                           Q => DRAM_ADDRESS_26_port, QN => n512);
   DataPath_REG_MEM_ALUOUT_Q_reg_26_inst : DFF_X1 port map( D => n1232, CK => 
                           CLK, Q => n_1361, QN => 
                           DataPath_i_REG_MEM_ALUOUT_26_port);
   DataPath_RF_BLOCKi_72_Q_reg_26_inst : DFF_X1 port map( D => n5874, CK => CLK
                           , Q => n_1362, QN => 
                           DataPath_RF_bus_reg_dataout_2074_port);
   DataPath_REG_IN2_Q_reg_27_inst : DFF_X1 port map( D => n2449, CK => CLK, Q 
                           => n_1363, QN => DataPath_i_PIPLIN_IN2_27_port);
   DataPath_REG_ALU_OUT_Q_reg_27_inst : DFF_X1 port map( D => n6996, CK => CLK,
                           Q => DRAM_ADDRESS_27_port, QN => n513);
   DataPath_REG_MEM_ALUOUT_Q_reg_27_inst : DFF_X1 port map( D => n1231, CK => 
                           CLK, Q => n_1364, QN => 
                           DataPath_i_REG_MEM_ALUOUT_27_port);
   DataPath_RF_BLOCKi_72_Q_reg_27_inst : DFF_X1 port map( D => n5873, CK => CLK
                           , Q => n_1365, QN => 
                           DataPath_RF_bus_reg_dataout_2075_port);
   DataPath_REG_IN2_Q_reg_28_inst : DFF_X1 port map( D => n2447, CK => CLK, Q 
                           => n_1366, QN => DataPath_i_PIPLIN_IN2_28_port);
   DataPath_REG_ALU_OUT_Q_reg_28_inst : DFF_X1 port map( D => n6995, CK => CLK,
                           Q => DRAM_ADDRESS_28_port, QN => n514);
   DataPath_REG_MEM_ALUOUT_Q_reg_28_inst : DFF_X1 port map( D => n1230, CK => 
                           CLK, Q => n_1367, QN => 
                           DataPath_i_REG_MEM_ALUOUT_28_port);
   DataPath_RF_BLOCKi_72_Q_reg_28_inst : DFF_X1 port map( D => n5872, CK => CLK
                           , Q => n_1368, QN => 
                           DataPath_RF_bus_reg_dataout_2076_port);
   DataPath_REG_IN2_Q_reg_29_inst : DFF_X1 port map( D => n2445, CK => CLK, Q 
                           => n_1369, QN => DataPath_i_PIPLIN_IN2_29_port);
   DataPath_REG_ALU_OUT_Q_reg_29_inst : DFF_X1 port map( D => n6994, CK => CLK,
                           Q => DRAM_ADDRESS_29_port, QN => n_1370);
   DataPath_REG_MEM_ALUOUT_Q_reg_29_inst : DFF_X1 port map( D => n1229, CK => 
                           CLK, Q => n_1371, QN => 
                           DataPath_i_REG_MEM_ALUOUT_29_port);
   DataPath_RF_BLOCKi_72_Q_reg_29_inst : DFF_X1 port map( D => n5871, CK => CLK
                           , Q => n_1372, QN => 
                           DataPath_RF_bus_reg_dataout_2077_port);
   DataPath_REG_IN2_Q_reg_30_inst : DFF_X1 port map( D => n2443, CK => CLK, Q 
                           => n_1373, QN => DataPath_i_PIPLIN_IN2_30_port);
   DataPath_REG_ALU_OUT_Q_reg_30_inst : DFF_X1 port map( D => n6993, CK => CLK,
                           Q => DRAM_ADDRESS_30_port, QN => n515);
   DataPath_REG_MEM_ALUOUT_Q_reg_30_inst : DFF_X1 port map( D => n1228, CK => 
                           CLK, Q => n_1374, QN => 
                           DataPath_i_REG_MEM_ALUOUT_30_port);
   DataPath_RF_BLOCKi_72_Q_reg_30_inst : DFF_X1 port map( D => n5870, CK => CLK
                           , Q => n_1375, QN => 
                           DataPath_RF_bus_reg_dataout_2078_port);
   DataPath_REG_IN2_Q_reg_31_inst : DFF_X1 port map( D => n2441, CK => CLK, Q 
                           => n_1376, QN => DataPath_i_PIPLIN_IN2_31_port);
   DataPath_REG_MEM_ALUOUT_Q_reg_31_inst : DFF_X1 port map( D => n1225, CK => 
                           CLK, Q => n_1377, QN => 
                           DataPath_i_REG_MEM_ALUOUT_31_port);
   DataPath_RF_BLOCKi_72_Q_reg_31_inst : DFF_X1 port map( D => n5867, CK => CLK
                           , Q => n_1378, QN => 
                           DataPath_RF_bus_reg_dataout_2079_port);
   CU_I_CW_ID_reg_0_inst : DLL_X1 port map( D => CU_I_CW_IF_0, GN => n7768, Q 
                           => CU_I_CW_ID_0_port);
   CU_I_CW_EX_reg_0_inst : DFF_X1 port map( D => n2962, CK => CLK, Q => n_1379,
                           QN => CU_I_CW_EX_0_port);
   CU_I_CW_MEM_reg_0_inst : DFF_X1 port map( D => n2956, CK => CLK, Q => n_1380
                           , QN => CU_I_CW_MEM_0_port);
   CU_I_CW_WB_reg_0_inst : DFF_X1 port map( D => CU_I_N170, CK => CLK, Q => 
                           i_WF, QN => n8409);
   DataPath_RF_BLOCKi_8_Q_reg_31_inst : DFF_X1 port map( D => n3274, CK => CLK,
                           Q => n_1381, QN => 
                           DataPath_RF_bus_reg_dataout_31_port);
   DataPath_RF_BLOCKi_8_Q_reg_30_inst : DFF_X1 port map( D => n3432, CK => CLK,
                           Q => n_1382, QN => 
                           DataPath_RF_bus_reg_dataout_30_port);
   DataPath_RF_BLOCKi_8_Q_reg_29_inst : DFF_X1 port map( D => n3434, CK => CLK,
                           Q => n_1383, QN => 
                           DataPath_RF_bus_reg_dataout_29_port);
   DataPath_RF_BLOCKi_8_Q_reg_28_inst : DFF_X1 port map( D => n3436, CK => CLK,
                           Q => n_1384, QN => 
                           DataPath_RF_bus_reg_dataout_28_port);
   DataPath_RF_BLOCKi_8_Q_reg_27_inst : DFF_X1 port map( D => n3438, CK => CLK,
                           Q => n_1385, QN => 
                           DataPath_RF_bus_reg_dataout_27_port);
   DataPath_RF_BLOCKi_8_Q_reg_26_inst : DFF_X1 port map( D => n3440, CK => CLK,
                           Q => n_1386, QN => 
                           DataPath_RF_bus_reg_dataout_26_port);
   DataPath_RF_BLOCKi_8_Q_reg_25_inst : DFF_X1 port map( D => n3442, CK => CLK,
                           Q => n_1387, QN => 
                           DataPath_RF_bus_reg_dataout_25_port);
   DataPath_RF_BLOCKi_8_Q_reg_24_inst : DFF_X1 port map( D => n3444, CK => CLK,
                           Q => n_1388, QN => 
                           DataPath_RF_bus_reg_dataout_24_port);
   DataPath_RF_BLOCKi_8_Q_reg_23_inst : DFF_X1 port map( D => n3446, CK => CLK,
                           Q => n_1389, QN => 
                           DataPath_RF_bus_reg_dataout_23_port);
   DataPath_RF_BLOCKi_8_Q_reg_22_inst : DFF_X1 port map( D => n3448, CK => CLK,
                           Q => n_1390, QN => 
                           DataPath_RF_bus_reg_dataout_22_port);
   DataPath_RF_BLOCKi_8_Q_reg_21_inst : DFF_X1 port map( D => n3450, CK => CLK,
                           Q => n_1391, QN => 
                           DataPath_RF_bus_reg_dataout_21_port);
   DataPath_RF_BLOCKi_8_Q_reg_20_inst : DFF_X1 port map( D => n3452, CK => CLK,
                           Q => n_1392, QN => 
                           DataPath_RF_bus_reg_dataout_20_port);
   DataPath_RF_BLOCKi_8_Q_reg_19_inst : DFF_X1 port map( D => n3454, CK => CLK,
                           Q => n_1393, QN => 
                           DataPath_RF_bus_reg_dataout_19_port);
   DataPath_RF_BLOCKi_8_Q_reg_18_inst : DFF_X1 port map( D => n3456, CK => CLK,
                           Q => n_1394, QN => 
                           DataPath_RF_bus_reg_dataout_18_port);
   DataPath_RF_BLOCKi_8_Q_reg_17_inst : DFF_X1 port map( D => n3458, CK => CLK,
                           Q => n_1395, QN => 
                           DataPath_RF_bus_reg_dataout_17_port);
   DataPath_RF_BLOCKi_8_Q_reg_16_inst : DFF_X1 port map( D => n3460, CK => CLK,
                           Q => n_1396, QN => 
                           DataPath_RF_bus_reg_dataout_16_port);
   DataPath_RF_BLOCKi_8_Q_reg_15_inst : DFF_X1 port map( D => n3462, CK => CLK,
                           Q => n_1397, QN => 
                           DataPath_RF_bus_reg_dataout_15_port);
   DataPath_RF_BLOCKi_8_Q_reg_14_inst : DFF_X1 port map( D => n3464, CK => CLK,
                           Q => n_1398, QN => 
                           DataPath_RF_bus_reg_dataout_14_port);
   DataPath_RF_BLOCKi_8_Q_reg_13_inst : DFF_X1 port map( D => n3466, CK => CLK,
                           Q => n_1399, QN => 
                           DataPath_RF_bus_reg_dataout_13_port);
   DataPath_RF_BLOCKi_8_Q_reg_12_inst : DFF_X1 port map( D => n3468, CK => CLK,
                           Q => n_1400, QN => 
                           DataPath_RF_bus_reg_dataout_12_port);
   DataPath_RF_BLOCKi_8_Q_reg_11_inst : DFF_X1 port map( D => n3470, CK => CLK,
                           Q => n_1401, QN => 
                           DataPath_RF_bus_reg_dataout_11_port);
   DataPath_RF_BLOCKi_8_Q_reg_9_inst : DFF_X1 port map( D => n3474, CK => CLK, 
                           Q => n_1402, QN => 
                           DataPath_RF_bus_reg_dataout_9_port);
   DataPath_RF_BLOCKi_8_Q_reg_8_inst : DFF_X1 port map( D => n3476, CK => CLK, 
                           Q => n_1403, QN => 
                           DataPath_RF_bus_reg_dataout_8_port);
   DataPath_RF_BLOCKi_8_Q_reg_7_inst : DFF_X1 port map( D => n3478, CK => CLK, 
                           Q => n_1404, QN => 
                           DataPath_RF_bus_reg_dataout_7_port);
   DataPath_RF_BLOCKi_8_Q_reg_6_inst : DFF_X1 port map( D => n3480, CK => CLK, 
                           Q => n_1405, QN => 
                           DataPath_RF_bus_reg_dataout_6_port);
   DataPath_RF_BLOCKi_8_Q_reg_5_inst : DFF_X1 port map( D => n3482, CK => CLK, 
                           Q => n_1406, QN => 
                           DataPath_RF_bus_reg_dataout_5_port);
   DataPath_RF_BLOCKi_8_Q_reg_4_inst : DFF_X1 port map( D => n3484, CK => CLK, 
                           Q => n_1407, QN => 
                           DataPath_RF_bus_reg_dataout_4_port);
   DataPath_RF_BLOCKi_8_Q_reg_3_inst : DFF_X1 port map( D => n3486, CK => CLK, 
                           Q => n_1408, QN => 
                           DataPath_RF_bus_reg_dataout_3_port);
   DataPath_RF_BLOCKi_8_Q_reg_2_inst : DFF_X1 port map( D => n3488, CK => CLK, 
                           Q => n_1409, QN => 
                           DataPath_RF_bus_reg_dataout_2_port);
   DataPath_RF_BLOCKi_8_Q_reg_1_inst : DFF_X1 port map( D => n3490, CK => CLK, 
                           Q => n_1410, QN => 
                           DataPath_RF_bus_reg_dataout_1_port);
   DataPath_RF_BLOCKi_8_Q_reg_0_inst : DFF_X1 port map( D => n3492, CK => CLK, 
                           Q => n_1411, QN => 
                           DataPath_RF_bus_reg_dataout_0_port);
   DataPath_RF_BLOCKi_24_Q_reg_31_inst : DFF_X1 port map( D => n4077, CK => CLK
                           , Q => n_1412, QN => 
                           DataPath_RF_bus_reg_dataout_543_port);
   DataPath_RF_BLOCKi_24_Q_reg_30_inst : DFF_X1 port map( D => n4081, CK => CLK
                           , Q => n_1413, QN => 
                           DataPath_RF_bus_reg_dataout_542_port);
   DataPath_RF_BLOCKi_24_Q_reg_29_inst : DFF_X1 port map( D => n4083, CK => CLK
                           , Q => n_1414, QN => 
                           DataPath_RF_bus_reg_dataout_541_port);
   DataPath_RF_BLOCKi_24_Q_reg_28_inst : DFF_X1 port map( D => n4085, CK => CLK
                           , Q => n_1415, QN => 
                           DataPath_RF_bus_reg_dataout_540_port);
   DataPath_RF_BLOCKi_24_Q_reg_27_inst : DFF_X1 port map( D => n4087, CK => CLK
                           , Q => n_1416, QN => 
                           DataPath_RF_bus_reg_dataout_539_port);
   DataPath_RF_BLOCKi_24_Q_reg_26_inst : DFF_X1 port map( D => n4089, CK => CLK
                           , Q => n_1417, QN => 
                           DataPath_RF_bus_reg_dataout_538_port);
   DataPath_RF_BLOCKi_24_Q_reg_25_inst : DFF_X1 port map( D => n4091, CK => CLK
                           , Q => n_1418, QN => 
                           DataPath_RF_bus_reg_dataout_537_port);
   DataPath_RF_BLOCKi_24_Q_reg_24_inst : DFF_X1 port map( D => n4093, CK => CLK
                           , Q => n_1419, QN => 
                           DataPath_RF_bus_reg_dataout_536_port);
   DataPath_RF_BLOCKi_24_Q_reg_23_inst : DFF_X1 port map( D => n4095, CK => CLK
                           , Q => n_1420, QN => 
                           DataPath_RF_bus_reg_dataout_535_port);
   DataPath_RF_BLOCKi_24_Q_reg_22_inst : DFF_X1 port map( D => n4097, CK => CLK
                           , Q => n_1421, QN => 
                           DataPath_RF_bus_reg_dataout_534_port);
   DataPath_RF_BLOCKi_24_Q_reg_21_inst : DFF_X1 port map( D => n4099, CK => CLK
                           , Q => n_1422, QN => 
                           DataPath_RF_bus_reg_dataout_533_port);
   DataPath_RF_BLOCKi_24_Q_reg_20_inst : DFF_X1 port map( D => n4101, CK => CLK
                           , Q => n_1423, QN => 
                           DataPath_RF_bus_reg_dataout_532_port);
   DataPath_RF_BLOCKi_24_Q_reg_19_inst : DFF_X1 port map( D => n4103, CK => CLK
                           , Q => n_1424, QN => 
                           DataPath_RF_bus_reg_dataout_531_port);
   DataPath_RF_BLOCKi_24_Q_reg_18_inst : DFF_X1 port map( D => n4105, CK => CLK
                           , Q => n_1425, QN => 
                           DataPath_RF_bus_reg_dataout_530_port);
   DataPath_RF_BLOCKi_24_Q_reg_17_inst : DFF_X1 port map( D => n4107, CK => CLK
                           , Q => n_1426, QN => 
                           DataPath_RF_bus_reg_dataout_529_port);
   DataPath_RF_BLOCKi_24_Q_reg_16_inst : DFF_X1 port map( D => n4109, CK => CLK
                           , Q => n_1427, QN => 
                           DataPath_RF_bus_reg_dataout_528_port);
   DataPath_RF_BLOCKi_24_Q_reg_15_inst : DFF_X1 port map( D => n4111, CK => CLK
                           , Q => n_1428, QN => 
                           DataPath_RF_bus_reg_dataout_527_port);
   DataPath_RF_BLOCKi_24_Q_reg_14_inst : DFF_X1 port map( D => n4113, CK => CLK
                           , Q => n_1429, QN => 
                           DataPath_RF_bus_reg_dataout_526_port);
   DataPath_RF_BLOCKi_24_Q_reg_13_inst : DFF_X1 port map( D => n4115, CK => CLK
                           , Q => n_1430, QN => 
                           DataPath_RF_bus_reg_dataout_525_port);
   DataPath_RF_BLOCKi_24_Q_reg_12_inst : DFF_X1 port map( D => n4117, CK => CLK
                           , Q => n_1431, QN => 
                           DataPath_RF_bus_reg_dataout_524_port);
   DataPath_RF_BLOCKi_24_Q_reg_11_inst : DFF_X1 port map( D => n4119, CK => CLK
                           , Q => n_1432, QN => 
                           DataPath_RF_bus_reg_dataout_523_port);
   DataPath_RF_BLOCKi_24_Q_reg_9_inst : DFF_X1 port map( D => n4123, CK => CLK,
                           Q => n_1433, QN => 
                           DataPath_RF_bus_reg_dataout_521_port);
   DataPath_RF_BLOCKi_24_Q_reg_8_inst : DFF_X1 port map( D => n4125, CK => CLK,
                           Q => n_1434, QN => 
                           DataPath_RF_bus_reg_dataout_520_port);
   DataPath_RF_BLOCKi_24_Q_reg_7_inst : DFF_X1 port map( D => n4127, CK => CLK,
                           Q => n_1435, QN => 
                           DataPath_RF_bus_reg_dataout_519_port);
   DataPath_RF_BLOCKi_24_Q_reg_6_inst : DFF_X1 port map( D => n4129, CK => CLK,
                           Q => n_1436, QN => 
                           DataPath_RF_bus_reg_dataout_518_port);
   DataPath_RF_BLOCKi_24_Q_reg_5_inst : DFF_X1 port map( D => n4131, CK => CLK,
                           Q => n_1437, QN => 
                           DataPath_RF_bus_reg_dataout_517_port);
   DataPath_RF_BLOCKi_24_Q_reg_4_inst : DFF_X1 port map( D => n4133, CK => CLK,
                           Q => n_1438, QN => 
                           DataPath_RF_bus_reg_dataout_516_port);
   DataPath_RF_BLOCKi_24_Q_reg_3_inst : DFF_X1 port map( D => n4135, CK => CLK,
                           Q => n_1439, QN => 
                           DataPath_RF_bus_reg_dataout_515_port);
   DataPath_RF_BLOCKi_24_Q_reg_2_inst : DFF_X1 port map( D => n4137, CK => CLK,
                           Q => n_1440, QN => 
                           DataPath_RF_bus_reg_dataout_514_port);
   DataPath_RF_BLOCKi_24_Q_reg_1_inst : DFF_X1 port map( D => n4139, CK => CLK,
                           Q => n_1441, QN => 
                           DataPath_RF_bus_reg_dataout_513_port);
   DataPath_RF_BLOCKi_24_Q_reg_0_inst : DFF_X1 port map( D => n4141, CK => CLK,
                           Q => n_1442, QN => 
                           DataPath_RF_bus_reg_dataout_512_port);
   DataPath_RF_BLOCKi_40_Q_reg_31_inst : DFF_X1 port map( D => n4670, CK => CLK
                           , Q => n_1443, QN => 
                           DataPath_RF_bus_reg_dataout_1055_port);
   DataPath_RF_BLOCKi_40_Q_reg_30_inst : DFF_X1 port map( D => n4674, CK => CLK
                           , Q => n_1444, QN => 
                           DataPath_RF_bus_reg_dataout_1054_port);
   DataPath_RF_BLOCKi_40_Q_reg_29_inst : DFF_X1 port map( D => n4676, CK => CLK
                           , Q => n_1445, QN => 
                           DataPath_RF_bus_reg_dataout_1053_port);
   DataPath_RF_BLOCKi_40_Q_reg_28_inst : DFF_X1 port map( D => n4678, CK => CLK
                           , Q => n_1446, QN => 
                           DataPath_RF_bus_reg_dataout_1052_port);
   DataPath_RF_BLOCKi_40_Q_reg_27_inst : DFF_X1 port map( D => n4680, CK => CLK
                           , Q => n_1447, QN => 
                           DataPath_RF_bus_reg_dataout_1051_port);
   DataPath_RF_BLOCKi_40_Q_reg_26_inst : DFF_X1 port map( D => n4682, CK => CLK
                           , Q => n_1448, QN => 
                           DataPath_RF_bus_reg_dataout_1050_port);
   DataPath_RF_BLOCKi_40_Q_reg_25_inst : DFF_X1 port map( D => n4684, CK => CLK
                           , Q => n_1449, QN => 
                           DataPath_RF_bus_reg_dataout_1049_port);
   DataPath_RF_BLOCKi_40_Q_reg_24_inst : DFF_X1 port map( D => n4686, CK => CLK
                           , Q => n_1450, QN => 
                           DataPath_RF_bus_reg_dataout_1048_port);
   DataPath_RF_BLOCKi_40_Q_reg_23_inst : DFF_X1 port map( D => n4688, CK => CLK
                           , Q => n_1451, QN => 
                           DataPath_RF_bus_reg_dataout_1047_port);
   DataPath_RF_BLOCKi_40_Q_reg_22_inst : DFF_X1 port map( D => n4690, CK => CLK
                           , Q => n_1452, QN => 
                           DataPath_RF_bus_reg_dataout_1046_port);
   DataPath_RF_BLOCKi_40_Q_reg_21_inst : DFF_X1 port map( D => n4692, CK => CLK
                           , Q => n_1453, QN => 
                           DataPath_RF_bus_reg_dataout_1045_port);
   DataPath_RF_BLOCKi_40_Q_reg_20_inst : DFF_X1 port map( D => n4694, CK => CLK
                           , Q => n_1454, QN => 
                           DataPath_RF_bus_reg_dataout_1044_port);
   DataPath_RF_BLOCKi_40_Q_reg_19_inst : DFF_X1 port map( D => n4696, CK => CLK
                           , Q => n_1455, QN => 
                           DataPath_RF_bus_reg_dataout_1043_port);
   DataPath_RF_BLOCKi_40_Q_reg_18_inst : DFF_X1 port map( D => n4698, CK => CLK
                           , Q => n_1456, QN => 
                           DataPath_RF_bus_reg_dataout_1042_port);
   DataPath_RF_BLOCKi_40_Q_reg_17_inst : DFF_X1 port map( D => n4700, CK => CLK
                           , Q => n_1457, QN => 
                           DataPath_RF_bus_reg_dataout_1041_port);
   DataPath_RF_BLOCKi_40_Q_reg_16_inst : DFF_X1 port map( D => n4702, CK => CLK
                           , Q => n_1458, QN => 
                           DataPath_RF_bus_reg_dataout_1040_port);
   DataPath_RF_BLOCKi_40_Q_reg_15_inst : DFF_X1 port map( D => n4704, CK => CLK
                           , Q => n_1459, QN => 
                           DataPath_RF_bus_reg_dataout_1039_port);
   DataPath_RF_BLOCKi_40_Q_reg_14_inst : DFF_X1 port map( D => n4706, CK => CLK
                           , Q => n_1460, QN => 
                           DataPath_RF_bus_reg_dataout_1038_port);
   DataPath_RF_BLOCKi_40_Q_reg_13_inst : DFF_X1 port map( D => n4708, CK => CLK
                           , Q => n_1461, QN => 
                           DataPath_RF_bus_reg_dataout_1037_port);
   DataPath_RF_BLOCKi_40_Q_reg_12_inst : DFF_X1 port map( D => n4710, CK => CLK
                           , Q => n_1462, QN => 
                           DataPath_RF_bus_reg_dataout_1036_port);
   DataPath_RF_BLOCKi_40_Q_reg_11_inst : DFF_X1 port map( D => n4712, CK => CLK
                           , Q => n_1463, QN => 
                           DataPath_RF_bus_reg_dataout_1035_port);
   DataPath_RF_BLOCKi_40_Q_reg_9_inst : DFF_X1 port map( D => n4716, CK => CLK,
                           Q => n_1464, QN => 
                           DataPath_RF_bus_reg_dataout_1033_port);
   DataPath_RF_BLOCKi_40_Q_reg_8_inst : DFF_X1 port map( D => n4718, CK => CLK,
                           Q => n_1465, QN => 
                           DataPath_RF_bus_reg_dataout_1032_port);
   DataPath_RF_BLOCKi_40_Q_reg_7_inst : DFF_X1 port map( D => n4720, CK => CLK,
                           Q => n_1466, QN => 
                           DataPath_RF_bus_reg_dataout_1031_port);
   DataPath_RF_BLOCKi_40_Q_reg_6_inst : DFF_X1 port map( D => n4722, CK => CLK,
                           Q => n_1467, QN => 
                           DataPath_RF_bus_reg_dataout_1030_port);
   DataPath_RF_BLOCKi_40_Q_reg_5_inst : DFF_X1 port map( D => n4724, CK => CLK,
                           Q => n_1468, QN => 
                           DataPath_RF_bus_reg_dataout_1029_port);
   DataPath_RF_BLOCKi_40_Q_reg_4_inst : DFF_X1 port map( D => n4726, CK => CLK,
                           Q => n_1469, QN => 
                           DataPath_RF_bus_reg_dataout_1028_port);
   DataPath_RF_BLOCKi_40_Q_reg_3_inst : DFF_X1 port map( D => n4728, CK => CLK,
                           Q => n_1470, QN => 
                           DataPath_RF_bus_reg_dataout_1027_port);
   DataPath_RF_BLOCKi_40_Q_reg_2_inst : DFF_X1 port map( D => n4730, CK => CLK,
                           Q => n_1471, QN => 
                           DataPath_RF_bus_reg_dataout_1026_port);
   DataPath_RF_BLOCKi_40_Q_reg_1_inst : DFF_X1 port map( D => n4732, CK => CLK,
                           Q => n_1472, QN => 
                           DataPath_RF_bus_reg_dataout_1025_port);
   DataPath_RF_BLOCKi_40_Q_reg_0_inst : DFF_X1 port map( D => n4734, CK => CLK,
                           Q => n_1473, QN => 
                           DataPath_RF_bus_reg_dataout_1024_port);
   DataPath_RF_BLOCKi_56_Q_reg_31_inst : DFF_X1 port map( D => n5263, CK => CLK
                           , Q => n_1474, QN => 
                           DataPath_RF_bus_reg_dataout_1567_port);
   DataPath_RF_BLOCKi_56_Q_reg_30_inst : DFF_X1 port map( D => n5267, CK => CLK
                           , Q => n_1475, QN => 
                           DataPath_RF_bus_reg_dataout_1566_port);
   DataPath_RF_BLOCKi_56_Q_reg_29_inst : DFF_X1 port map( D => n5269, CK => CLK
                           , Q => n_1476, QN => 
                           DataPath_RF_bus_reg_dataout_1565_port);
   DataPath_RF_BLOCKi_56_Q_reg_28_inst : DFF_X1 port map( D => n5271, CK => CLK
                           , Q => n_1477, QN => 
                           DataPath_RF_bus_reg_dataout_1564_port);
   DataPath_RF_BLOCKi_56_Q_reg_27_inst : DFF_X1 port map( D => n5273, CK => CLK
                           , Q => n_1478, QN => 
                           DataPath_RF_bus_reg_dataout_1563_port);
   DataPath_RF_BLOCKi_56_Q_reg_26_inst : DFF_X1 port map( D => n5275, CK => CLK
                           , Q => n_1479, QN => 
                           DataPath_RF_bus_reg_dataout_1562_port);
   DataPath_RF_BLOCKi_56_Q_reg_25_inst : DFF_X1 port map( D => n5277, CK => CLK
                           , Q => n_1480, QN => 
                           DataPath_RF_bus_reg_dataout_1561_port);
   DataPath_RF_BLOCKi_56_Q_reg_24_inst : DFF_X1 port map( D => n5279, CK => CLK
                           , Q => n_1481, QN => 
                           DataPath_RF_bus_reg_dataout_1560_port);
   DataPath_RF_BLOCKi_56_Q_reg_23_inst : DFF_X1 port map( D => n5281, CK => CLK
                           , Q => n_1482, QN => 
                           DataPath_RF_bus_reg_dataout_1559_port);
   DataPath_RF_BLOCKi_56_Q_reg_22_inst : DFF_X1 port map( D => n5283, CK => CLK
                           , Q => n_1483, QN => 
                           DataPath_RF_bus_reg_dataout_1558_port);
   DataPath_RF_BLOCKi_56_Q_reg_21_inst : DFF_X1 port map( D => n5285, CK => CLK
                           , Q => n_1484, QN => 
                           DataPath_RF_bus_reg_dataout_1557_port);
   DataPath_RF_BLOCKi_56_Q_reg_20_inst : DFF_X1 port map( D => n5287, CK => CLK
                           , Q => n_1485, QN => 
                           DataPath_RF_bus_reg_dataout_1556_port);
   DataPath_RF_BLOCKi_56_Q_reg_19_inst : DFF_X1 port map( D => n5289, CK => CLK
                           , Q => n_1486, QN => 
                           DataPath_RF_bus_reg_dataout_1555_port);
   DataPath_RF_BLOCKi_56_Q_reg_18_inst : DFF_X1 port map( D => n5291, CK => CLK
                           , Q => n_1487, QN => 
                           DataPath_RF_bus_reg_dataout_1554_port);
   DataPath_RF_BLOCKi_56_Q_reg_17_inst : DFF_X1 port map( D => n5293, CK => CLK
                           , Q => n_1488, QN => 
                           DataPath_RF_bus_reg_dataout_1553_port);
   DataPath_RF_BLOCKi_56_Q_reg_16_inst : DFF_X1 port map( D => n5295, CK => CLK
                           , Q => n_1489, QN => 
                           DataPath_RF_bus_reg_dataout_1552_port);
   DataPath_RF_BLOCKi_56_Q_reg_15_inst : DFF_X1 port map( D => n5297, CK => CLK
                           , Q => n_1490, QN => 
                           DataPath_RF_bus_reg_dataout_1551_port);
   DataPath_RF_BLOCKi_56_Q_reg_14_inst : DFF_X1 port map( D => n5299, CK => CLK
                           , Q => n_1491, QN => 
                           DataPath_RF_bus_reg_dataout_1550_port);
   DataPath_RF_BLOCKi_56_Q_reg_13_inst : DFF_X1 port map( D => n5301, CK => CLK
                           , Q => n_1492, QN => 
                           DataPath_RF_bus_reg_dataout_1549_port);
   DataPath_RF_BLOCKi_56_Q_reg_12_inst : DFF_X1 port map( D => n5303, CK => CLK
                           , Q => n_1493, QN => 
                           DataPath_RF_bus_reg_dataout_1548_port);
   DataPath_RF_BLOCKi_56_Q_reg_11_inst : DFF_X1 port map( D => n5305, CK => CLK
                           , Q => n_1494, QN => 
                           DataPath_RF_bus_reg_dataout_1547_port);
   DataPath_RF_BLOCKi_56_Q_reg_9_inst : DFF_X1 port map( D => n5309, CK => CLK,
                           Q => n_1495, QN => 
                           DataPath_RF_bus_reg_dataout_1545_port);
   DataPath_RF_BLOCKi_56_Q_reg_8_inst : DFF_X1 port map( D => n5311, CK => CLK,
                           Q => n_1496, QN => 
                           DataPath_RF_bus_reg_dataout_1544_port);
   DataPath_RF_BLOCKi_56_Q_reg_7_inst : DFF_X1 port map( D => n5313, CK => CLK,
                           Q => n_1497, QN => 
                           DataPath_RF_bus_reg_dataout_1543_port);
   DataPath_RF_BLOCKi_56_Q_reg_6_inst : DFF_X1 port map( D => n5315, CK => CLK,
                           Q => n_1498, QN => 
                           DataPath_RF_bus_reg_dataout_1542_port);
   DataPath_RF_BLOCKi_56_Q_reg_5_inst : DFF_X1 port map( D => n5317, CK => CLK,
                           Q => n_1499, QN => 
                           DataPath_RF_bus_reg_dataout_1541_port);
   DataPath_RF_BLOCKi_56_Q_reg_4_inst : DFF_X1 port map( D => n5319, CK => CLK,
                           Q => n_1500, QN => 
                           DataPath_RF_bus_reg_dataout_1540_port);
   DataPath_RF_BLOCKi_56_Q_reg_3_inst : DFF_X1 port map( D => n5321, CK => CLK,
                           Q => n_1501, QN => 
                           DataPath_RF_bus_reg_dataout_1539_port);
   DataPath_RF_BLOCKi_56_Q_reg_2_inst : DFF_X1 port map( D => n5323, CK => CLK,
                           Q => n_1502, QN => 
                           DataPath_RF_bus_reg_dataout_1538_port);
   DataPath_RF_BLOCKi_56_Q_reg_1_inst : DFF_X1 port map( D => n5325, CK => CLK,
                           Q => n_1503, QN => 
                           DataPath_RF_bus_reg_dataout_1537_port);
   DataPath_RF_BLOCKi_56_Q_reg_0_inst : DFF_X1 port map( D => n5327, CK => CLK,
                           Q => n_1504, QN => 
                           DataPath_RF_bus_reg_dataout_1536_port);
   DataPath_RF_BLOCKi_9_Q_reg_31_inst : DFF_X1 port map( D => n3499, CK => CLK,
                           Q => n_1505, QN => 
                           DataPath_RF_bus_reg_dataout_63_port);
   DataPath_RF_BLOCKi_9_Q_reg_30_inst : DFF_X1 port map( D => n3502, CK => CLK,
                           Q => n_1506, QN => 
                           DataPath_RF_bus_reg_dataout_62_port);
   DataPath_RF_BLOCKi_9_Q_reg_29_inst : DFF_X1 port map( D => n3503, CK => CLK,
                           Q => n_1507, QN => 
                           DataPath_RF_bus_reg_dataout_61_port);
   DataPath_RF_BLOCKi_9_Q_reg_28_inst : DFF_X1 port map( D => n3504, CK => CLK,
                           Q => n_1508, QN => 
                           DataPath_RF_bus_reg_dataout_60_port);
   DataPath_RF_BLOCKi_9_Q_reg_27_inst : DFF_X1 port map( D => n3505, CK => CLK,
                           Q => n_1509, QN => 
                           DataPath_RF_bus_reg_dataout_59_port);
   DataPath_RF_BLOCKi_9_Q_reg_26_inst : DFF_X1 port map( D => n3506, CK => CLK,
                           Q => n_1510, QN => 
                           DataPath_RF_bus_reg_dataout_58_port);
   DataPath_RF_BLOCKi_9_Q_reg_25_inst : DFF_X1 port map( D => n3507, CK => CLK,
                           Q => n_1511, QN => 
                           DataPath_RF_bus_reg_dataout_57_port);
   DataPath_RF_BLOCKi_9_Q_reg_24_inst : DFF_X1 port map( D => n3508, CK => CLK,
                           Q => n_1512, QN => 
                           DataPath_RF_bus_reg_dataout_56_port);
   DataPath_RF_BLOCKi_9_Q_reg_23_inst : DFF_X1 port map( D => n3509, CK => CLK,
                           Q => n_1513, QN => 
                           DataPath_RF_bus_reg_dataout_55_port);
   DataPath_RF_BLOCKi_9_Q_reg_22_inst : DFF_X1 port map( D => n3510, CK => CLK,
                           Q => n_1514, QN => 
                           DataPath_RF_bus_reg_dataout_54_port);
   DataPath_RF_BLOCKi_9_Q_reg_21_inst : DFF_X1 port map( D => n3511, CK => CLK,
                           Q => n_1515, QN => 
                           DataPath_RF_bus_reg_dataout_53_port);
   DataPath_RF_BLOCKi_9_Q_reg_20_inst : DFF_X1 port map( D => n3512, CK => CLK,
                           Q => n_1516, QN => 
                           DataPath_RF_bus_reg_dataout_52_port);
   DataPath_RF_BLOCKi_9_Q_reg_19_inst : DFF_X1 port map( D => n3513, CK => CLK,
                           Q => n_1517, QN => 
                           DataPath_RF_bus_reg_dataout_51_port);
   DataPath_RF_BLOCKi_9_Q_reg_18_inst : DFF_X1 port map( D => n3514, CK => CLK,
                           Q => n_1518, QN => 
                           DataPath_RF_bus_reg_dataout_50_port);
   DataPath_RF_BLOCKi_9_Q_reg_17_inst : DFF_X1 port map( D => n3515, CK => CLK,
                           Q => n_1519, QN => 
                           DataPath_RF_bus_reg_dataout_49_port);
   DataPath_RF_BLOCKi_9_Q_reg_16_inst : DFF_X1 port map( D => n3516, CK => CLK,
                           Q => n_1520, QN => 
                           DataPath_RF_bus_reg_dataout_48_port);
   DataPath_RF_BLOCKi_9_Q_reg_15_inst : DFF_X1 port map( D => n3517, CK => CLK,
                           Q => n_1521, QN => 
                           DataPath_RF_bus_reg_dataout_47_port);
   DataPath_RF_BLOCKi_9_Q_reg_14_inst : DFF_X1 port map( D => n3518, CK => CLK,
                           Q => n_1522, QN => 
                           DataPath_RF_bus_reg_dataout_46_port);
   DataPath_RF_BLOCKi_9_Q_reg_13_inst : DFF_X1 port map( D => n3519, CK => CLK,
                           Q => n_1523, QN => 
                           DataPath_RF_bus_reg_dataout_45_port);
   DataPath_RF_BLOCKi_9_Q_reg_12_inst : DFF_X1 port map( D => n3520, CK => CLK,
                           Q => n_1524, QN => 
                           DataPath_RF_bus_reg_dataout_44_port);
   DataPath_RF_BLOCKi_9_Q_reg_11_inst : DFF_X1 port map( D => n3521, CK => CLK,
                           Q => n_1525, QN => 
                           DataPath_RF_bus_reg_dataout_43_port);
   DataPath_RF_BLOCKi_9_Q_reg_9_inst : DFF_X1 port map( D => n3523, CK => CLK, 
                           Q => n_1526, QN => 
                           DataPath_RF_bus_reg_dataout_41_port);
   DataPath_RF_BLOCKi_9_Q_reg_8_inst : DFF_X1 port map( D => n3524, CK => CLK, 
                           Q => n_1527, QN => 
                           DataPath_RF_bus_reg_dataout_40_port);
   DataPath_RF_BLOCKi_9_Q_reg_7_inst : DFF_X1 port map( D => n3525, CK => CLK, 
                           Q => n_1528, QN => 
                           DataPath_RF_bus_reg_dataout_39_port);
   DataPath_RF_BLOCKi_9_Q_reg_6_inst : DFF_X1 port map( D => n3526, CK => CLK, 
                           Q => n_1529, QN => 
                           DataPath_RF_bus_reg_dataout_38_port);
   DataPath_RF_BLOCKi_9_Q_reg_5_inst : DFF_X1 port map( D => n3527, CK => CLK, 
                           Q => n_1530, QN => 
                           DataPath_RF_bus_reg_dataout_37_port);
   DataPath_RF_BLOCKi_9_Q_reg_4_inst : DFF_X1 port map( D => n3528, CK => CLK, 
                           Q => n_1531, QN => 
                           DataPath_RF_bus_reg_dataout_36_port);
   DataPath_RF_BLOCKi_9_Q_reg_3_inst : DFF_X1 port map( D => n3529, CK => CLK, 
                           Q => n_1532, QN => 
                           DataPath_RF_bus_reg_dataout_35_port);
   DataPath_RF_BLOCKi_9_Q_reg_2_inst : DFF_X1 port map( D => n3530, CK => CLK, 
                           Q => n_1533, QN => 
                           DataPath_RF_bus_reg_dataout_34_port);
   DataPath_RF_BLOCKi_9_Q_reg_1_inst : DFF_X1 port map( D => n3531, CK => CLK, 
                           Q => n_1534, QN => 
                           DataPath_RF_bus_reg_dataout_33_port);
   DataPath_RF_BLOCKi_9_Q_reg_0_inst : DFF_X1 port map( D => n3532, CK => CLK, 
                           Q => n_1535, QN => 
                           DataPath_RF_bus_reg_dataout_32_port);
   DataPath_RF_BLOCKi_25_Q_reg_31_inst : DFF_X1 port map( D => n4145, CK => CLK
                           , Q => n_1536, QN => 
                           DataPath_RF_bus_reg_dataout_575_port);
   DataPath_RF_BLOCKi_25_Q_reg_30_inst : DFF_X1 port map( D => n4148, CK => CLK
                           , Q => n_1537, QN => 
                           DataPath_RF_bus_reg_dataout_574_port);
   DataPath_RF_BLOCKi_25_Q_reg_29_inst : DFF_X1 port map( D => n4149, CK => CLK
                           , Q => n_1538, QN => 
                           DataPath_RF_bus_reg_dataout_573_port);
   DataPath_RF_BLOCKi_25_Q_reg_28_inst : DFF_X1 port map( D => n4150, CK => CLK
                           , Q => n_1539, QN => 
                           DataPath_RF_bus_reg_dataout_572_port);
   DataPath_RF_BLOCKi_25_Q_reg_27_inst : DFF_X1 port map( D => n4151, CK => CLK
                           , Q => n_1540, QN => 
                           DataPath_RF_bus_reg_dataout_571_port);
   DataPath_RF_BLOCKi_25_Q_reg_26_inst : DFF_X1 port map( D => n4152, CK => CLK
                           , Q => n_1541, QN => 
                           DataPath_RF_bus_reg_dataout_570_port);
   DataPath_RF_BLOCKi_25_Q_reg_25_inst : DFF_X1 port map( D => n4153, CK => CLK
                           , Q => n_1542, QN => 
                           DataPath_RF_bus_reg_dataout_569_port);
   DataPath_RF_BLOCKi_25_Q_reg_24_inst : DFF_X1 port map( D => n4154, CK => CLK
                           , Q => n_1543, QN => 
                           DataPath_RF_bus_reg_dataout_568_port);
   DataPath_RF_BLOCKi_25_Q_reg_23_inst : DFF_X1 port map( D => n4155, CK => CLK
                           , Q => n_1544, QN => 
                           DataPath_RF_bus_reg_dataout_567_port);
   DataPath_RF_BLOCKi_25_Q_reg_22_inst : DFF_X1 port map( D => n4156, CK => CLK
                           , Q => n_1545, QN => 
                           DataPath_RF_bus_reg_dataout_566_port);
   DataPath_RF_BLOCKi_25_Q_reg_21_inst : DFF_X1 port map( D => n4157, CK => CLK
                           , Q => n_1546, QN => 
                           DataPath_RF_bus_reg_dataout_565_port);
   DataPath_RF_BLOCKi_25_Q_reg_20_inst : DFF_X1 port map( D => n4158, CK => CLK
                           , Q => n_1547, QN => 
                           DataPath_RF_bus_reg_dataout_564_port);
   DataPath_RF_BLOCKi_25_Q_reg_19_inst : DFF_X1 port map( D => n4159, CK => CLK
                           , Q => n_1548, QN => 
                           DataPath_RF_bus_reg_dataout_563_port);
   DataPath_RF_BLOCKi_25_Q_reg_18_inst : DFF_X1 port map( D => n4160, CK => CLK
                           , Q => n_1549, QN => 
                           DataPath_RF_bus_reg_dataout_562_port);
   DataPath_RF_BLOCKi_25_Q_reg_17_inst : DFF_X1 port map( D => n4161, CK => CLK
                           , Q => n_1550, QN => 
                           DataPath_RF_bus_reg_dataout_561_port);
   DataPath_RF_BLOCKi_25_Q_reg_16_inst : DFF_X1 port map( D => n4162, CK => CLK
                           , Q => n_1551, QN => 
                           DataPath_RF_bus_reg_dataout_560_port);
   DataPath_RF_BLOCKi_25_Q_reg_15_inst : DFF_X1 port map( D => n4163, CK => CLK
                           , Q => n_1552, QN => 
                           DataPath_RF_bus_reg_dataout_559_port);
   DataPath_RF_BLOCKi_25_Q_reg_14_inst : DFF_X1 port map( D => n4164, CK => CLK
                           , Q => n_1553, QN => 
                           DataPath_RF_bus_reg_dataout_558_port);
   DataPath_RF_BLOCKi_25_Q_reg_13_inst : DFF_X1 port map( D => n4165, CK => CLK
                           , Q => n_1554, QN => 
                           DataPath_RF_bus_reg_dataout_557_port);
   DataPath_RF_BLOCKi_25_Q_reg_12_inst : DFF_X1 port map( D => n4166, CK => CLK
                           , Q => n_1555, QN => 
                           DataPath_RF_bus_reg_dataout_556_port);
   DataPath_RF_BLOCKi_25_Q_reg_11_inst : DFF_X1 port map( D => n4167, CK => CLK
                           , Q => n_1556, QN => 
                           DataPath_RF_bus_reg_dataout_555_port);
   DataPath_RF_BLOCKi_25_Q_reg_9_inst : DFF_X1 port map( D => n4169, CK => CLK,
                           Q => n_1557, QN => 
                           DataPath_RF_bus_reg_dataout_553_port);
   DataPath_RF_BLOCKi_25_Q_reg_8_inst : DFF_X1 port map( D => n4170, CK => CLK,
                           Q => n_1558, QN => 
                           DataPath_RF_bus_reg_dataout_552_port);
   DataPath_RF_BLOCKi_25_Q_reg_7_inst : DFF_X1 port map( D => n4171, CK => CLK,
                           Q => n_1559, QN => 
                           DataPath_RF_bus_reg_dataout_551_port);
   DataPath_RF_BLOCKi_25_Q_reg_6_inst : DFF_X1 port map( D => n4172, CK => CLK,
                           Q => n_1560, QN => 
                           DataPath_RF_bus_reg_dataout_550_port);
   DataPath_RF_BLOCKi_25_Q_reg_5_inst : DFF_X1 port map( D => n4173, CK => CLK,
                           Q => n_1561, QN => 
                           DataPath_RF_bus_reg_dataout_549_port);
   DataPath_RF_BLOCKi_25_Q_reg_4_inst : DFF_X1 port map( D => n4174, CK => CLK,
                           Q => n_1562, QN => 
                           DataPath_RF_bus_reg_dataout_548_port);
   DataPath_RF_BLOCKi_25_Q_reg_3_inst : DFF_X1 port map( D => n4175, CK => CLK,
                           Q => n_1563, QN => 
                           DataPath_RF_bus_reg_dataout_547_port);
   DataPath_RF_BLOCKi_25_Q_reg_2_inst : DFF_X1 port map( D => n4176, CK => CLK,
                           Q => n_1564, QN => 
                           DataPath_RF_bus_reg_dataout_546_port);
   DataPath_RF_BLOCKi_25_Q_reg_1_inst : DFF_X1 port map( D => n4177, CK => CLK,
                           Q => n_1565, QN => 
                           DataPath_RF_bus_reg_dataout_545_port);
   DataPath_RF_BLOCKi_25_Q_reg_0_inst : DFF_X1 port map( D => n4178, CK => CLK,
                           Q => n_1566, QN => 
                           DataPath_RF_bus_reg_dataout_544_port);
   DataPath_RF_BLOCKi_41_Q_reg_31_inst : DFF_X1 port map( D => n4738, CK => CLK
                           , Q => n_1567, QN => 
                           DataPath_RF_bus_reg_dataout_1087_port);
   DataPath_RF_BLOCKi_41_Q_reg_30_inst : DFF_X1 port map( D => n4741, CK => CLK
                           , Q => n_1568, QN => 
                           DataPath_RF_bus_reg_dataout_1086_port);
   DataPath_RF_BLOCKi_41_Q_reg_29_inst : DFF_X1 port map( D => n4742, CK => CLK
                           , Q => n_1569, QN => 
                           DataPath_RF_bus_reg_dataout_1085_port);
   DataPath_RF_BLOCKi_41_Q_reg_28_inst : DFF_X1 port map( D => n4743, CK => CLK
                           , Q => n_1570, QN => 
                           DataPath_RF_bus_reg_dataout_1084_port);
   DataPath_RF_BLOCKi_41_Q_reg_27_inst : DFF_X1 port map( D => n4744, CK => CLK
                           , Q => n_1571, QN => 
                           DataPath_RF_bus_reg_dataout_1083_port);
   DataPath_RF_BLOCKi_41_Q_reg_26_inst : DFF_X1 port map( D => n4745, CK => CLK
                           , Q => n_1572, QN => 
                           DataPath_RF_bus_reg_dataout_1082_port);
   DataPath_RF_BLOCKi_41_Q_reg_25_inst : DFF_X1 port map( D => n4746, CK => CLK
                           , Q => n_1573, QN => 
                           DataPath_RF_bus_reg_dataout_1081_port);
   DataPath_RF_BLOCKi_41_Q_reg_24_inst : DFF_X1 port map( D => n4747, CK => CLK
                           , Q => n_1574, QN => 
                           DataPath_RF_bus_reg_dataout_1080_port);
   DataPath_RF_BLOCKi_41_Q_reg_23_inst : DFF_X1 port map( D => n4748, CK => CLK
                           , Q => n_1575, QN => 
                           DataPath_RF_bus_reg_dataout_1079_port);
   DataPath_RF_BLOCKi_41_Q_reg_22_inst : DFF_X1 port map( D => n4749, CK => CLK
                           , Q => n_1576, QN => 
                           DataPath_RF_bus_reg_dataout_1078_port);
   DataPath_RF_BLOCKi_41_Q_reg_21_inst : DFF_X1 port map( D => n4750, CK => CLK
                           , Q => n_1577, QN => 
                           DataPath_RF_bus_reg_dataout_1077_port);
   DataPath_RF_BLOCKi_41_Q_reg_20_inst : DFF_X1 port map( D => n4751, CK => CLK
                           , Q => n_1578, QN => 
                           DataPath_RF_bus_reg_dataout_1076_port);
   DataPath_RF_BLOCKi_41_Q_reg_19_inst : DFF_X1 port map( D => n4752, CK => CLK
                           , Q => n_1579, QN => 
                           DataPath_RF_bus_reg_dataout_1075_port);
   DataPath_RF_BLOCKi_41_Q_reg_18_inst : DFF_X1 port map( D => n4753, CK => CLK
                           , Q => n_1580, QN => 
                           DataPath_RF_bus_reg_dataout_1074_port);
   DataPath_RF_BLOCKi_41_Q_reg_17_inst : DFF_X1 port map( D => n4754, CK => CLK
                           , Q => n_1581, QN => 
                           DataPath_RF_bus_reg_dataout_1073_port);
   DataPath_RF_BLOCKi_41_Q_reg_16_inst : DFF_X1 port map( D => n4755, CK => CLK
                           , Q => n_1582, QN => 
                           DataPath_RF_bus_reg_dataout_1072_port);
   DataPath_RF_BLOCKi_41_Q_reg_15_inst : DFF_X1 port map( D => n4756, CK => CLK
                           , Q => n_1583, QN => 
                           DataPath_RF_bus_reg_dataout_1071_port);
   DataPath_RF_BLOCKi_41_Q_reg_14_inst : DFF_X1 port map( D => n4757, CK => CLK
                           , Q => n_1584, QN => 
                           DataPath_RF_bus_reg_dataout_1070_port);
   DataPath_RF_BLOCKi_41_Q_reg_13_inst : DFF_X1 port map( D => n4758, CK => CLK
                           , Q => n_1585, QN => 
                           DataPath_RF_bus_reg_dataout_1069_port);
   DataPath_RF_BLOCKi_41_Q_reg_12_inst : DFF_X1 port map( D => n4759, CK => CLK
                           , Q => n_1586, QN => 
                           DataPath_RF_bus_reg_dataout_1068_port);
   DataPath_RF_BLOCKi_41_Q_reg_11_inst : DFF_X1 port map( D => n4760, CK => CLK
                           , Q => n_1587, QN => 
                           DataPath_RF_bus_reg_dataout_1067_port);
   DataPath_RF_BLOCKi_41_Q_reg_9_inst : DFF_X1 port map( D => n4762, CK => CLK,
                           Q => n_1588, QN => 
                           DataPath_RF_bus_reg_dataout_1065_port);
   DataPath_RF_BLOCKi_41_Q_reg_8_inst : DFF_X1 port map( D => n4763, CK => CLK,
                           Q => n_1589, QN => 
                           DataPath_RF_bus_reg_dataout_1064_port);
   DataPath_RF_BLOCKi_41_Q_reg_7_inst : DFF_X1 port map( D => n4764, CK => CLK,
                           Q => n_1590, QN => 
                           DataPath_RF_bus_reg_dataout_1063_port);
   DataPath_RF_BLOCKi_41_Q_reg_6_inst : DFF_X1 port map( D => n4765, CK => CLK,
                           Q => n_1591, QN => 
                           DataPath_RF_bus_reg_dataout_1062_port);
   DataPath_RF_BLOCKi_41_Q_reg_5_inst : DFF_X1 port map( D => n4766, CK => CLK,
                           Q => n_1592, QN => 
                           DataPath_RF_bus_reg_dataout_1061_port);
   DataPath_RF_BLOCKi_41_Q_reg_4_inst : DFF_X1 port map( D => n4767, CK => CLK,
                           Q => n_1593, QN => 
                           DataPath_RF_bus_reg_dataout_1060_port);
   DataPath_RF_BLOCKi_41_Q_reg_3_inst : DFF_X1 port map( D => n4768, CK => CLK,
                           Q => n_1594, QN => 
                           DataPath_RF_bus_reg_dataout_1059_port);
   DataPath_RF_BLOCKi_41_Q_reg_2_inst : DFF_X1 port map( D => n4769, CK => CLK,
                           Q => n_1595, QN => 
                           DataPath_RF_bus_reg_dataout_1058_port);
   DataPath_RF_BLOCKi_41_Q_reg_1_inst : DFF_X1 port map( D => n4770, CK => CLK,
                           Q => n_1596, QN => 
                           DataPath_RF_bus_reg_dataout_1057_port);
   DataPath_RF_BLOCKi_41_Q_reg_0_inst : DFF_X1 port map( D => n4771, CK => CLK,
                           Q => n_1597, QN => 
                           DataPath_RF_bus_reg_dataout_1056_port);
   DataPath_RF_BLOCKi_57_Q_reg_31_inst : DFF_X1 port map( D => n5331, CK => CLK
                           , Q => n_1598, QN => 
                           DataPath_RF_bus_reg_dataout_1599_port);
   DataPath_RF_BLOCKi_57_Q_reg_30_inst : DFF_X1 port map( D => n5334, CK => CLK
                           , Q => n_1599, QN => 
                           DataPath_RF_bus_reg_dataout_1598_port);
   DataPath_RF_BLOCKi_57_Q_reg_29_inst : DFF_X1 port map( D => n5335, CK => CLK
                           , Q => n_1600, QN => 
                           DataPath_RF_bus_reg_dataout_1597_port);
   DataPath_RF_BLOCKi_57_Q_reg_28_inst : DFF_X1 port map( D => n5336, CK => CLK
                           , Q => n_1601, QN => 
                           DataPath_RF_bus_reg_dataout_1596_port);
   DataPath_RF_BLOCKi_57_Q_reg_27_inst : DFF_X1 port map( D => n5337, CK => CLK
                           , Q => n_1602, QN => 
                           DataPath_RF_bus_reg_dataout_1595_port);
   DataPath_RF_BLOCKi_57_Q_reg_26_inst : DFF_X1 port map( D => n5338, CK => CLK
                           , Q => n_1603, QN => 
                           DataPath_RF_bus_reg_dataout_1594_port);
   DataPath_RF_BLOCKi_57_Q_reg_25_inst : DFF_X1 port map( D => n5339, CK => CLK
                           , Q => n_1604, QN => 
                           DataPath_RF_bus_reg_dataout_1593_port);
   DataPath_RF_BLOCKi_57_Q_reg_24_inst : DFF_X1 port map( D => n5340, CK => CLK
                           , Q => n_1605, QN => 
                           DataPath_RF_bus_reg_dataout_1592_port);
   DataPath_RF_BLOCKi_57_Q_reg_23_inst : DFF_X1 port map( D => n5341, CK => CLK
                           , Q => n_1606, QN => 
                           DataPath_RF_bus_reg_dataout_1591_port);
   DataPath_RF_BLOCKi_57_Q_reg_22_inst : DFF_X1 port map( D => n5342, CK => CLK
                           , Q => n_1607, QN => 
                           DataPath_RF_bus_reg_dataout_1590_port);
   DataPath_RF_BLOCKi_57_Q_reg_21_inst : DFF_X1 port map( D => n5343, CK => CLK
                           , Q => n_1608, QN => 
                           DataPath_RF_bus_reg_dataout_1589_port);
   DataPath_RF_BLOCKi_57_Q_reg_20_inst : DFF_X1 port map( D => n5344, CK => CLK
                           , Q => n_1609, QN => 
                           DataPath_RF_bus_reg_dataout_1588_port);
   DataPath_RF_BLOCKi_57_Q_reg_19_inst : DFF_X1 port map( D => n5345, CK => CLK
                           , Q => n_1610, QN => 
                           DataPath_RF_bus_reg_dataout_1587_port);
   DataPath_RF_BLOCKi_57_Q_reg_18_inst : DFF_X1 port map( D => n5346, CK => CLK
                           , Q => n_1611, QN => 
                           DataPath_RF_bus_reg_dataout_1586_port);
   DataPath_RF_BLOCKi_57_Q_reg_17_inst : DFF_X1 port map( D => n5347, CK => CLK
                           , Q => n_1612, QN => 
                           DataPath_RF_bus_reg_dataout_1585_port);
   DataPath_RF_BLOCKi_57_Q_reg_16_inst : DFF_X1 port map( D => n5348, CK => CLK
                           , Q => n_1613, QN => 
                           DataPath_RF_bus_reg_dataout_1584_port);
   DataPath_RF_BLOCKi_57_Q_reg_15_inst : DFF_X1 port map( D => n5349, CK => CLK
                           , Q => n_1614, QN => 
                           DataPath_RF_bus_reg_dataout_1583_port);
   DataPath_RF_BLOCKi_57_Q_reg_14_inst : DFF_X1 port map( D => n5350, CK => CLK
                           , Q => n_1615, QN => 
                           DataPath_RF_bus_reg_dataout_1582_port);
   DataPath_RF_BLOCKi_57_Q_reg_13_inst : DFF_X1 port map( D => n5351, CK => CLK
                           , Q => n_1616, QN => 
                           DataPath_RF_bus_reg_dataout_1581_port);
   DataPath_RF_BLOCKi_57_Q_reg_12_inst : DFF_X1 port map( D => n5352, CK => CLK
                           , Q => n_1617, QN => 
                           DataPath_RF_bus_reg_dataout_1580_port);
   DataPath_RF_BLOCKi_57_Q_reg_11_inst : DFF_X1 port map( D => n5353, CK => CLK
                           , Q => n_1618, QN => 
                           DataPath_RF_bus_reg_dataout_1579_port);
   DataPath_RF_BLOCKi_57_Q_reg_9_inst : DFF_X1 port map( D => n5355, CK => CLK,
                           Q => n_1619, QN => 
                           DataPath_RF_bus_reg_dataout_1577_port);
   DataPath_RF_BLOCKi_57_Q_reg_8_inst : DFF_X1 port map( D => n5356, CK => CLK,
                           Q => n_1620, QN => 
                           DataPath_RF_bus_reg_dataout_1576_port);
   DataPath_RF_BLOCKi_57_Q_reg_7_inst : DFF_X1 port map( D => n5357, CK => CLK,
                           Q => n_1621, QN => 
                           DataPath_RF_bus_reg_dataout_1575_port);
   DataPath_RF_BLOCKi_57_Q_reg_6_inst : DFF_X1 port map( D => n5358, CK => CLK,
                           Q => n_1622, QN => 
                           DataPath_RF_bus_reg_dataout_1574_port);
   DataPath_RF_BLOCKi_57_Q_reg_5_inst : DFF_X1 port map( D => n5359, CK => CLK,
                           Q => n_1623, QN => 
                           DataPath_RF_bus_reg_dataout_1573_port);
   DataPath_RF_BLOCKi_57_Q_reg_4_inst : DFF_X1 port map( D => n5360, CK => CLK,
                           Q => n_1624, QN => 
                           DataPath_RF_bus_reg_dataout_1572_port);
   DataPath_RF_BLOCKi_57_Q_reg_3_inst : DFF_X1 port map( D => n5361, CK => CLK,
                           Q => n_1625, QN => 
                           DataPath_RF_bus_reg_dataout_1571_port);
   DataPath_RF_BLOCKi_57_Q_reg_2_inst : DFF_X1 port map( D => n5362, CK => CLK,
                           Q => n_1626, QN => 
                           DataPath_RF_bus_reg_dataout_1570_port);
   DataPath_RF_BLOCKi_57_Q_reg_1_inst : DFF_X1 port map( D => n5363, CK => CLK,
                           Q => n_1627, QN => 
                           DataPath_RF_bus_reg_dataout_1569_port);
   DataPath_RF_BLOCKi_57_Q_reg_0_inst : DFF_X1 port map( D => n5364, CK => CLK,
                           Q => n_1628, QN => 
                           DataPath_RF_bus_reg_dataout_1568_port);
   DataPath_RF_BLOCKi_73_Q_reg_31_inst : DFF_X1 port map( D => n5905, CK => CLK
                           , Q => n_1629, QN => 
                           DataPath_RF_bus_reg_dataout_2111_port);
   DataPath_RF_BLOCKi_73_Q_reg_30_inst : DFF_X1 port map( D => n5908, CK => CLK
                           , Q => n_1630, QN => 
                           DataPath_RF_bus_reg_dataout_2110_port);
   DataPath_RF_BLOCKi_73_Q_reg_29_inst : DFF_X1 port map( D => n5909, CK => CLK
                           , Q => n_1631, QN => 
                           DataPath_RF_bus_reg_dataout_2109_port);
   DataPath_RF_BLOCKi_73_Q_reg_28_inst : DFF_X1 port map( D => n5910, CK => CLK
                           , Q => n_1632, QN => 
                           DataPath_RF_bus_reg_dataout_2108_port);
   DataPath_RF_BLOCKi_73_Q_reg_27_inst : DFF_X1 port map( D => n5911, CK => CLK
                           , Q => n_1633, QN => 
                           DataPath_RF_bus_reg_dataout_2107_port);
   DataPath_RF_BLOCKi_73_Q_reg_26_inst : DFF_X1 port map( D => n5912, CK => CLK
                           , Q => n_1634, QN => 
                           DataPath_RF_bus_reg_dataout_2106_port);
   DataPath_RF_BLOCKi_73_Q_reg_25_inst : DFF_X1 port map( D => n5913, CK => CLK
                           , Q => n_1635, QN => 
                           DataPath_RF_bus_reg_dataout_2105_port);
   DataPath_RF_BLOCKi_73_Q_reg_24_inst : DFF_X1 port map( D => n5914, CK => CLK
                           , Q => n_1636, QN => 
                           DataPath_RF_bus_reg_dataout_2104_port);
   DataPath_RF_BLOCKi_73_Q_reg_23_inst : DFF_X1 port map( D => n5915, CK => CLK
                           , Q => n_1637, QN => 
                           DataPath_RF_bus_reg_dataout_2103_port);
   DataPath_RF_BLOCKi_73_Q_reg_22_inst : DFF_X1 port map( D => n5916, CK => CLK
                           , Q => n_1638, QN => 
                           DataPath_RF_bus_reg_dataout_2102_port);
   DataPath_RF_BLOCKi_73_Q_reg_21_inst : DFF_X1 port map( D => n5917, CK => CLK
                           , Q => n_1639, QN => 
                           DataPath_RF_bus_reg_dataout_2101_port);
   DataPath_RF_BLOCKi_73_Q_reg_20_inst : DFF_X1 port map( D => n5918, CK => CLK
                           , Q => n_1640, QN => 
                           DataPath_RF_bus_reg_dataout_2100_port);
   DataPath_RF_BLOCKi_73_Q_reg_19_inst : DFF_X1 port map( D => n5919, CK => CLK
                           , Q => n_1641, QN => 
                           DataPath_RF_bus_reg_dataout_2099_port);
   DataPath_RF_BLOCKi_73_Q_reg_18_inst : DFF_X1 port map( D => n5920, CK => CLK
                           , Q => n_1642, QN => 
                           DataPath_RF_bus_reg_dataout_2098_port);
   DataPath_RF_BLOCKi_73_Q_reg_17_inst : DFF_X1 port map( D => n5921, CK => CLK
                           , Q => n_1643, QN => 
                           DataPath_RF_bus_reg_dataout_2097_port);
   DataPath_RF_BLOCKi_73_Q_reg_16_inst : DFF_X1 port map( D => n5922, CK => CLK
                           , Q => n_1644, QN => 
                           DataPath_RF_bus_reg_dataout_2096_port);
   DataPath_RF_BLOCKi_73_Q_reg_15_inst : DFF_X1 port map( D => n5923, CK => CLK
                           , Q => n_1645, QN => 
                           DataPath_RF_bus_reg_dataout_2095_port);
   DataPath_RF_BLOCKi_73_Q_reg_14_inst : DFF_X1 port map( D => n5924, CK => CLK
                           , Q => n_1646, QN => 
                           DataPath_RF_bus_reg_dataout_2094_port);
   DataPath_RF_BLOCKi_73_Q_reg_13_inst : DFF_X1 port map( D => n5925, CK => CLK
                           , Q => n_1647, QN => 
                           DataPath_RF_bus_reg_dataout_2093_port);
   DataPath_RF_BLOCKi_73_Q_reg_12_inst : DFF_X1 port map( D => n5926, CK => CLK
                           , Q => n_1648, QN => 
                           DataPath_RF_bus_reg_dataout_2092_port);
   DataPath_RF_BLOCKi_73_Q_reg_11_inst : DFF_X1 port map( D => n5927, CK => CLK
                           , Q => n_1649, QN => 
                           DataPath_RF_bus_reg_dataout_2091_port);
   DataPath_RF_BLOCKi_73_Q_reg_9_inst : DFF_X1 port map( D => n5929, CK => CLK,
                           Q => n_1650, QN => 
                           DataPath_RF_bus_reg_dataout_2089_port);
   DataPath_RF_BLOCKi_73_Q_reg_8_inst : DFF_X1 port map( D => n5930, CK => CLK,
                           Q => n_1651, QN => 
                           DataPath_RF_bus_reg_dataout_2088_port);
   DataPath_RF_BLOCKi_73_Q_reg_7_inst : DFF_X1 port map( D => n5931, CK => CLK,
                           Q => n_1652, QN => 
                           DataPath_RF_bus_reg_dataout_2087_port);
   DataPath_RF_BLOCKi_73_Q_reg_6_inst : DFF_X1 port map( D => n5932, CK => CLK,
                           Q => n_1653, QN => 
                           DataPath_RF_bus_reg_dataout_2086_port);
   DataPath_RF_BLOCKi_73_Q_reg_5_inst : DFF_X1 port map( D => n5933, CK => CLK,
                           Q => n_1654, QN => 
                           DataPath_RF_bus_reg_dataout_2085_port);
   DataPath_RF_BLOCKi_73_Q_reg_4_inst : DFF_X1 port map( D => n5934, CK => CLK,
                           Q => n_1655, QN => 
                           DataPath_RF_bus_reg_dataout_2084_port);
   DataPath_RF_BLOCKi_73_Q_reg_3_inst : DFF_X1 port map( D => n5935, CK => CLK,
                           Q => n_1656, QN => 
                           DataPath_RF_bus_reg_dataout_2083_port);
   DataPath_RF_BLOCKi_73_Q_reg_2_inst : DFF_X1 port map( D => n5936, CK => CLK,
                           Q => n_1657, QN => 
                           DataPath_RF_bus_reg_dataout_2082_port);
   DataPath_RF_BLOCKi_73_Q_reg_1_inst : DFF_X1 port map( D => n5937, CK => CLK,
                           Q => n_1658, QN => 
                           DataPath_RF_bus_reg_dataout_2081_port);
   DataPath_RF_BLOCKi_73_Q_reg_0_inst : DFF_X1 port map( D => n5938, CK => CLK,
                           Q => n_1659, QN => 
                           DataPath_RF_bus_reg_dataout_2080_port);
   DataPath_RF_BLOCKi_10_Q_reg_31_inst : DFF_X1 port map( D => n3537, CK => CLK
                           , Q => n_1660, QN => 
                           DataPath_RF_bus_reg_dataout_95_port);
   DataPath_RF_BLOCKi_10_Q_reg_30_inst : DFF_X1 port map( D => n3540, CK => CLK
                           , Q => n_1661, QN => 
                           DataPath_RF_bus_reg_dataout_94_port);
   DataPath_RF_BLOCKi_10_Q_reg_29_inst : DFF_X1 port map( D => n3541, CK => CLK
                           , Q => n_1662, QN => 
                           DataPath_RF_bus_reg_dataout_93_port);
   DataPath_RF_BLOCKi_10_Q_reg_28_inst : DFF_X1 port map( D => n3542, CK => CLK
                           , Q => n_1663, QN => 
                           DataPath_RF_bus_reg_dataout_92_port);
   DataPath_RF_BLOCKi_10_Q_reg_27_inst : DFF_X1 port map( D => n3543, CK => CLK
                           , Q => n_1664, QN => 
                           DataPath_RF_bus_reg_dataout_91_port);
   DataPath_RF_BLOCKi_10_Q_reg_26_inst : DFF_X1 port map( D => n3544, CK => CLK
                           , Q => n_1665, QN => 
                           DataPath_RF_bus_reg_dataout_90_port);
   DataPath_RF_BLOCKi_10_Q_reg_25_inst : DFF_X1 port map( D => n3545, CK => CLK
                           , Q => n_1666, QN => 
                           DataPath_RF_bus_reg_dataout_89_port);
   DataPath_RF_BLOCKi_10_Q_reg_24_inst : DFF_X1 port map( D => n3546, CK => CLK
                           , Q => n_1667, QN => 
                           DataPath_RF_bus_reg_dataout_88_port);
   DataPath_RF_BLOCKi_10_Q_reg_23_inst : DFF_X1 port map( D => n3547, CK => CLK
                           , Q => n_1668, QN => 
                           DataPath_RF_bus_reg_dataout_87_port);
   DataPath_RF_BLOCKi_10_Q_reg_22_inst : DFF_X1 port map( D => n3548, CK => CLK
                           , Q => n_1669, QN => 
                           DataPath_RF_bus_reg_dataout_86_port);
   DataPath_RF_BLOCKi_10_Q_reg_21_inst : DFF_X1 port map( D => n3549, CK => CLK
                           , Q => n_1670, QN => 
                           DataPath_RF_bus_reg_dataout_85_port);
   DataPath_RF_BLOCKi_10_Q_reg_20_inst : DFF_X1 port map( D => n3550, CK => CLK
                           , Q => n_1671, QN => 
                           DataPath_RF_bus_reg_dataout_84_port);
   DataPath_RF_BLOCKi_10_Q_reg_19_inst : DFF_X1 port map( D => n3551, CK => CLK
                           , Q => n_1672, QN => 
                           DataPath_RF_bus_reg_dataout_83_port);
   DataPath_RF_BLOCKi_10_Q_reg_18_inst : DFF_X1 port map( D => n3552, CK => CLK
                           , Q => n_1673, QN => 
                           DataPath_RF_bus_reg_dataout_82_port);
   DataPath_RF_BLOCKi_10_Q_reg_17_inst : DFF_X1 port map( D => n3553, CK => CLK
                           , Q => n_1674, QN => 
                           DataPath_RF_bus_reg_dataout_81_port);
   DataPath_RF_BLOCKi_10_Q_reg_16_inst : DFF_X1 port map( D => n3554, CK => CLK
                           , Q => n_1675, QN => 
                           DataPath_RF_bus_reg_dataout_80_port);
   DataPath_RF_BLOCKi_10_Q_reg_15_inst : DFF_X1 port map( D => n3555, CK => CLK
                           , Q => n_1676, QN => 
                           DataPath_RF_bus_reg_dataout_79_port);
   DataPath_RF_BLOCKi_10_Q_reg_14_inst : DFF_X1 port map( D => n3556, CK => CLK
                           , Q => n_1677, QN => 
                           DataPath_RF_bus_reg_dataout_78_port);
   DataPath_RF_BLOCKi_10_Q_reg_13_inst : DFF_X1 port map( D => n3557, CK => CLK
                           , Q => n_1678, QN => 
                           DataPath_RF_bus_reg_dataout_77_port);
   DataPath_RF_BLOCKi_10_Q_reg_12_inst : DFF_X1 port map( D => n3558, CK => CLK
                           , Q => n_1679, QN => 
                           DataPath_RF_bus_reg_dataout_76_port);
   DataPath_RF_BLOCKi_10_Q_reg_11_inst : DFF_X1 port map( D => n3559, CK => CLK
                           , Q => n_1680, QN => 
                           DataPath_RF_bus_reg_dataout_75_port);
   DataPath_RF_BLOCKi_10_Q_reg_9_inst : DFF_X1 port map( D => n3561, CK => CLK,
                           Q => n_1681, QN => 
                           DataPath_RF_bus_reg_dataout_73_port);
   DataPath_RF_BLOCKi_10_Q_reg_8_inst : DFF_X1 port map( D => n3562, CK => CLK,
                           Q => n_1682, QN => 
                           DataPath_RF_bus_reg_dataout_72_port);
   DataPath_RF_BLOCKi_10_Q_reg_7_inst : DFF_X1 port map( D => n3563, CK => CLK,
                           Q => n_1683, QN => 
                           DataPath_RF_bus_reg_dataout_71_port);
   DataPath_RF_BLOCKi_10_Q_reg_6_inst : DFF_X1 port map( D => n3564, CK => CLK,
                           Q => n_1684, QN => 
                           DataPath_RF_bus_reg_dataout_70_port);
   DataPath_RF_BLOCKi_10_Q_reg_5_inst : DFF_X1 port map( D => n3565, CK => CLK,
                           Q => n_1685, QN => 
                           DataPath_RF_bus_reg_dataout_69_port);
   DataPath_RF_BLOCKi_10_Q_reg_4_inst : DFF_X1 port map( D => n3566, CK => CLK,
                           Q => n_1686, QN => 
                           DataPath_RF_bus_reg_dataout_68_port);
   DataPath_RF_BLOCKi_10_Q_reg_3_inst : DFF_X1 port map( D => n3567, CK => CLK,
                           Q => n_1687, QN => 
                           DataPath_RF_bus_reg_dataout_67_port);
   DataPath_RF_BLOCKi_10_Q_reg_2_inst : DFF_X1 port map( D => n3568, CK => CLK,
                           Q => n_1688, QN => 
                           DataPath_RF_bus_reg_dataout_66_port);
   DataPath_RF_BLOCKi_10_Q_reg_1_inst : DFF_X1 port map( D => n3569, CK => CLK,
                           Q => n_1689, QN => 
                           DataPath_RF_bus_reg_dataout_65_port);
   DataPath_RF_BLOCKi_10_Q_reg_0_inst : DFF_X1 port map( D => n3570, CK => CLK,
                           Q => n_1690, QN => 
                           DataPath_RF_bus_reg_dataout_64_port);
   DataPath_RF_BLOCKi_26_Q_reg_31_inst : DFF_X1 port map( D => n4180, CK => CLK
                           , Q => n_1691, QN => 
                           DataPath_RF_bus_reg_dataout_607_port);
   DataPath_RF_BLOCKi_26_Q_reg_30_inst : DFF_X1 port map( D => n4183, CK => CLK
                           , Q => n_1692, QN => 
                           DataPath_RF_bus_reg_dataout_606_port);
   DataPath_RF_BLOCKi_26_Q_reg_29_inst : DFF_X1 port map( D => n4184, CK => CLK
                           , Q => n_1693, QN => 
                           DataPath_RF_bus_reg_dataout_605_port);
   DataPath_RF_BLOCKi_26_Q_reg_28_inst : DFF_X1 port map( D => n4185, CK => CLK
                           , Q => n_1694, QN => 
                           DataPath_RF_bus_reg_dataout_604_port);
   DataPath_RF_BLOCKi_26_Q_reg_27_inst : DFF_X1 port map( D => n4186, CK => CLK
                           , Q => n_1695, QN => 
                           DataPath_RF_bus_reg_dataout_603_port);
   DataPath_RF_BLOCKi_26_Q_reg_26_inst : DFF_X1 port map( D => n4187, CK => CLK
                           , Q => n_1696, QN => 
                           DataPath_RF_bus_reg_dataout_602_port);
   DataPath_RF_BLOCKi_26_Q_reg_25_inst : DFF_X1 port map( D => n4188, CK => CLK
                           , Q => n_1697, QN => 
                           DataPath_RF_bus_reg_dataout_601_port);
   DataPath_RF_BLOCKi_26_Q_reg_24_inst : DFF_X1 port map( D => n4189, CK => CLK
                           , Q => n_1698, QN => 
                           DataPath_RF_bus_reg_dataout_600_port);
   DataPath_RF_BLOCKi_26_Q_reg_23_inst : DFF_X1 port map( D => n4190, CK => CLK
                           , Q => n_1699, QN => 
                           DataPath_RF_bus_reg_dataout_599_port);
   DataPath_RF_BLOCKi_26_Q_reg_22_inst : DFF_X1 port map( D => n4191, CK => CLK
                           , Q => n_1700, QN => 
                           DataPath_RF_bus_reg_dataout_598_port);
   DataPath_RF_BLOCKi_26_Q_reg_21_inst : DFF_X1 port map( D => n4192, CK => CLK
                           , Q => n_1701, QN => 
                           DataPath_RF_bus_reg_dataout_597_port);
   DataPath_RF_BLOCKi_26_Q_reg_20_inst : DFF_X1 port map( D => n4193, CK => CLK
                           , Q => n_1702, QN => 
                           DataPath_RF_bus_reg_dataout_596_port);
   DataPath_RF_BLOCKi_26_Q_reg_19_inst : DFF_X1 port map( D => n4194, CK => CLK
                           , Q => n_1703, QN => 
                           DataPath_RF_bus_reg_dataout_595_port);
   DataPath_RF_BLOCKi_26_Q_reg_18_inst : DFF_X1 port map( D => n4195, CK => CLK
                           , Q => n_1704, QN => 
                           DataPath_RF_bus_reg_dataout_594_port);
   DataPath_RF_BLOCKi_26_Q_reg_17_inst : DFF_X1 port map( D => n4196, CK => CLK
                           , Q => n_1705, QN => 
                           DataPath_RF_bus_reg_dataout_593_port);
   DataPath_RF_BLOCKi_26_Q_reg_16_inst : DFF_X1 port map( D => n4197, CK => CLK
                           , Q => n_1706, QN => 
                           DataPath_RF_bus_reg_dataout_592_port);
   DataPath_RF_BLOCKi_26_Q_reg_15_inst : DFF_X1 port map( D => n4198, CK => CLK
                           , Q => n_1707, QN => 
                           DataPath_RF_bus_reg_dataout_591_port);
   DataPath_RF_BLOCKi_26_Q_reg_14_inst : DFF_X1 port map( D => n4199, CK => CLK
                           , Q => n_1708, QN => 
                           DataPath_RF_bus_reg_dataout_590_port);
   DataPath_RF_BLOCKi_26_Q_reg_13_inst : DFF_X1 port map( D => n4200, CK => CLK
                           , Q => n_1709, QN => 
                           DataPath_RF_bus_reg_dataout_589_port);
   DataPath_RF_BLOCKi_26_Q_reg_12_inst : DFF_X1 port map( D => n4201, CK => CLK
                           , Q => n_1710, QN => 
                           DataPath_RF_bus_reg_dataout_588_port);
   DataPath_RF_BLOCKi_26_Q_reg_11_inst : DFF_X1 port map( D => n4202, CK => CLK
                           , Q => n_1711, QN => 
                           DataPath_RF_bus_reg_dataout_587_port);
   DataPath_RF_BLOCKi_26_Q_reg_9_inst : DFF_X1 port map( D => n4204, CK => CLK,
                           Q => n_1712, QN => 
                           DataPath_RF_bus_reg_dataout_585_port);
   DataPath_RF_BLOCKi_26_Q_reg_8_inst : DFF_X1 port map( D => n4205, CK => CLK,
                           Q => n_1713, QN => 
                           DataPath_RF_bus_reg_dataout_584_port);
   DataPath_RF_BLOCKi_26_Q_reg_7_inst : DFF_X1 port map( D => n4206, CK => CLK,
                           Q => n_1714, QN => 
                           DataPath_RF_bus_reg_dataout_583_port);
   DataPath_RF_BLOCKi_26_Q_reg_6_inst : DFF_X1 port map( D => n4207, CK => CLK,
                           Q => n_1715, QN => 
                           DataPath_RF_bus_reg_dataout_582_port);
   DataPath_RF_BLOCKi_26_Q_reg_5_inst : DFF_X1 port map( D => n4208, CK => CLK,
                           Q => n_1716, QN => 
                           DataPath_RF_bus_reg_dataout_581_port);
   DataPath_RF_BLOCKi_26_Q_reg_4_inst : DFF_X1 port map( D => n4209, CK => CLK,
                           Q => n_1717, QN => 
                           DataPath_RF_bus_reg_dataout_580_port);
   DataPath_RF_BLOCKi_26_Q_reg_3_inst : DFF_X1 port map( D => n4210, CK => CLK,
                           Q => n_1718, QN => 
                           DataPath_RF_bus_reg_dataout_579_port);
   DataPath_RF_BLOCKi_26_Q_reg_2_inst : DFF_X1 port map( D => n4211, CK => CLK,
                           Q => n_1719, QN => 
                           DataPath_RF_bus_reg_dataout_578_port);
   DataPath_RF_BLOCKi_26_Q_reg_1_inst : DFF_X1 port map( D => n4212, CK => CLK,
                           Q => n_1720, QN => 
                           DataPath_RF_bus_reg_dataout_577_port);
   DataPath_RF_BLOCKi_26_Q_reg_0_inst : DFF_X1 port map( D => n4213, CK => CLK,
                           Q => n_1721, QN => 
                           DataPath_RF_bus_reg_dataout_576_port);
   DataPath_RF_BLOCKi_42_Q_reg_31_inst : DFF_X1 port map( D => n4773, CK => CLK
                           , Q => n_1722, QN => 
                           DataPath_RF_bus_reg_dataout_1119_port);
   DataPath_RF_BLOCKi_42_Q_reg_30_inst : DFF_X1 port map( D => n4776, CK => CLK
                           , Q => n_1723, QN => 
                           DataPath_RF_bus_reg_dataout_1118_port);
   DataPath_RF_BLOCKi_42_Q_reg_29_inst : DFF_X1 port map( D => n4777, CK => CLK
                           , Q => n_1724, QN => 
                           DataPath_RF_bus_reg_dataout_1117_port);
   DataPath_RF_BLOCKi_42_Q_reg_28_inst : DFF_X1 port map( D => n4778, CK => CLK
                           , Q => n_1725, QN => 
                           DataPath_RF_bus_reg_dataout_1116_port);
   DataPath_RF_BLOCKi_42_Q_reg_27_inst : DFF_X1 port map( D => n4779, CK => CLK
                           , Q => n_1726, QN => 
                           DataPath_RF_bus_reg_dataout_1115_port);
   DataPath_RF_BLOCKi_42_Q_reg_26_inst : DFF_X1 port map( D => n4780, CK => CLK
                           , Q => n_1727, QN => 
                           DataPath_RF_bus_reg_dataout_1114_port);
   DataPath_RF_BLOCKi_42_Q_reg_25_inst : DFF_X1 port map( D => n4781, CK => CLK
                           , Q => n_1728, QN => 
                           DataPath_RF_bus_reg_dataout_1113_port);
   DataPath_RF_BLOCKi_42_Q_reg_24_inst : DFF_X1 port map( D => n4782, CK => CLK
                           , Q => n_1729, QN => 
                           DataPath_RF_bus_reg_dataout_1112_port);
   DataPath_RF_BLOCKi_42_Q_reg_23_inst : DFF_X1 port map( D => n4783, CK => CLK
                           , Q => n_1730, QN => 
                           DataPath_RF_bus_reg_dataout_1111_port);
   DataPath_RF_BLOCKi_42_Q_reg_22_inst : DFF_X1 port map( D => n4784, CK => CLK
                           , Q => n_1731, QN => 
                           DataPath_RF_bus_reg_dataout_1110_port);
   DataPath_RF_BLOCKi_42_Q_reg_21_inst : DFF_X1 port map( D => n4785, CK => CLK
                           , Q => n_1732, QN => 
                           DataPath_RF_bus_reg_dataout_1109_port);
   DataPath_RF_BLOCKi_42_Q_reg_20_inst : DFF_X1 port map( D => n4786, CK => CLK
                           , Q => n_1733, QN => 
                           DataPath_RF_bus_reg_dataout_1108_port);
   DataPath_RF_BLOCKi_42_Q_reg_19_inst : DFF_X1 port map( D => n4787, CK => CLK
                           , Q => n_1734, QN => 
                           DataPath_RF_bus_reg_dataout_1107_port);
   DataPath_RF_BLOCKi_42_Q_reg_18_inst : DFF_X1 port map( D => n4788, CK => CLK
                           , Q => n_1735, QN => 
                           DataPath_RF_bus_reg_dataout_1106_port);
   DataPath_RF_BLOCKi_42_Q_reg_17_inst : DFF_X1 port map( D => n4789, CK => CLK
                           , Q => n_1736, QN => 
                           DataPath_RF_bus_reg_dataout_1105_port);
   DataPath_RF_BLOCKi_42_Q_reg_16_inst : DFF_X1 port map( D => n4790, CK => CLK
                           , Q => n_1737, QN => 
                           DataPath_RF_bus_reg_dataout_1104_port);
   DataPath_RF_BLOCKi_42_Q_reg_15_inst : DFF_X1 port map( D => n4791, CK => CLK
                           , Q => n_1738, QN => 
                           DataPath_RF_bus_reg_dataout_1103_port);
   DataPath_RF_BLOCKi_42_Q_reg_14_inst : DFF_X1 port map( D => n4792, CK => CLK
                           , Q => n_1739, QN => 
                           DataPath_RF_bus_reg_dataout_1102_port);
   DataPath_RF_BLOCKi_42_Q_reg_13_inst : DFF_X1 port map( D => n4793, CK => CLK
                           , Q => n_1740, QN => 
                           DataPath_RF_bus_reg_dataout_1101_port);
   DataPath_RF_BLOCKi_42_Q_reg_12_inst : DFF_X1 port map( D => n4794, CK => CLK
                           , Q => n_1741, QN => 
                           DataPath_RF_bus_reg_dataout_1100_port);
   DataPath_RF_BLOCKi_42_Q_reg_11_inst : DFF_X1 port map( D => n4795, CK => CLK
                           , Q => n_1742, QN => 
                           DataPath_RF_bus_reg_dataout_1099_port);
   DataPath_RF_BLOCKi_42_Q_reg_9_inst : DFF_X1 port map( D => n4797, CK => CLK,
                           Q => n_1743, QN => 
                           DataPath_RF_bus_reg_dataout_1097_port);
   DataPath_RF_BLOCKi_42_Q_reg_8_inst : DFF_X1 port map( D => n4798, CK => CLK,
                           Q => n_1744, QN => 
                           DataPath_RF_bus_reg_dataout_1096_port);
   DataPath_RF_BLOCKi_42_Q_reg_7_inst : DFF_X1 port map( D => n4799, CK => CLK,
                           Q => n_1745, QN => 
                           DataPath_RF_bus_reg_dataout_1095_port);
   DataPath_RF_BLOCKi_42_Q_reg_6_inst : DFF_X1 port map( D => n4800, CK => CLK,
                           Q => n_1746, QN => 
                           DataPath_RF_bus_reg_dataout_1094_port);
   DataPath_RF_BLOCKi_42_Q_reg_5_inst : DFF_X1 port map( D => n4801, CK => CLK,
                           Q => n_1747, QN => 
                           DataPath_RF_bus_reg_dataout_1093_port);
   DataPath_RF_BLOCKi_42_Q_reg_4_inst : DFF_X1 port map( D => n4802, CK => CLK,
                           Q => n_1748, QN => 
                           DataPath_RF_bus_reg_dataout_1092_port);
   DataPath_RF_BLOCKi_42_Q_reg_3_inst : DFF_X1 port map( D => n4803, CK => CLK,
                           Q => n_1749, QN => 
                           DataPath_RF_bus_reg_dataout_1091_port);
   DataPath_RF_BLOCKi_42_Q_reg_2_inst : DFF_X1 port map( D => n4804, CK => CLK,
                           Q => n_1750, QN => 
                           DataPath_RF_bus_reg_dataout_1090_port);
   DataPath_RF_BLOCKi_42_Q_reg_1_inst : DFF_X1 port map( D => n4805, CK => CLK,
                           Q => n_1751, QN => 
                           DataPath_RF_bus_reg_dataout_1089_port);
   DataPath_RF_BLOCKi_42_Q_reg_0_inst : DFF_X1 port map( D => n4806, CK => CLK,
                           Q => n_1752, QN => 
                           DataPath_RF_bus_reg_dataout_1088_port);
   DataPath_RF_BLOCKi_58_Q_reg_31_inst : DFF_X1 port map( D => n5366, CK => CLK
                           , Q => n_1753, QN => 
                           DataPath_RF_bus_reg_dataout_1631_port);
   DataPath_RF_BLOCKi_58_Q_reg_30_inst : DFF_X1 port map( D => n5369, CK => CLK
                           , Q => n_1754, QN => 
                           DataPath_RF_bus_reg_dataout_1630_port);
   DataPath_RF_BLOCKi_58_Q_reg_29_inst : DFF_X1 port map( D => n5370, CK => CLK
                           , Q => n_1755, QN => 
                           DataPath_RF_bus_reg_dataout_1629_port);
   DataPath_RF_BLOCKi_58_Q_reg_28_inst : DFF_X1 port map( D => n5371, CK => CLK
                           , Q => n_1756, QN => 
                           DataPath_RF_bus_reg_dataout_1628_port);
   DataPath_RF_BLOCKi_58_Q_reg_27_inst : DFF_X1 port map( D => n5372, CK => CLK
                           , Q => n_1757, QN => 
                           DataPath_RF_bus_reg_dataout_1627_port);
   DataPath_RF_BLOCKi_58_Q_reg_26_inst : DFF_X1 port map( D => n5373, CK => CLK
                           , Q => n_1758, QN => 
                           DataPath_RF_bus_reg_dataout_1626_port);
   DataPath_RF_BLOCKi_58_Q_reg_25_inst : DFF_X1 port map( D => n5374, CK => CLK
                           , Q => n_1759, QN => 
                           DataPath_RF_bus_reg_dataout_1625_port);
   DataPath_RF_BLOCKi_58_Q_reg_24_inst : DFF_X1 port map( D => n5375, CK => CLK
                           , Q => n_1760, QN => 
                           DataPath_RF_bus_reg_dataout_1624_port);
   DataPath_RF_BLOCKi_58_Q_reg_23_inst : DFF_X1 port map( D => n5376, CK => CLK
                           , Q => n_1761, QN => 
                           DataPath_RF_bus_reg_dataout_1623_port);
   DataPath_RF_BLOCKi_58_Q_reg_22_inst : DFF_X1 port map( D => n5377, CK => CLK
                           , Q => n_1762, QN => 
                           DataPath_RF_bus_reg_dataout_1622_port);
   DataPath_RF_BLOCKi_58_Q_reg_21_inst : DFF_X1 port map( D => n5378, CK => CLK
                           , Q => n_1763, QN => 
                           DataPath_RF_bus_reg_dataout_1621_port);
   DataPath_RF_BLOCKi_58_Q_reg_20_inst : DFF_X1 port map( D => n5379, CK => CLK
                           , Q => n_1764, QN => 
                           DataPath_RF_bus_reg_dataout_1620_port);
   DataPath_RF_BLOCKi_58_Q_reg_19_inst : DFF_X1 port map( D => n5380, CK => CLK
                           , Q => n_1765, QN => 
                           DataPath_RF_bus_reg_dataout_1619_port);
   DataPath_RF_BLOCKi_58_Q_reg_18_inst : DFF_X1 port map( D => n5381, CK => CLK
                           , Q => n_1766, QN => 
                           DataPath_RF_bus_reg_dataout_1618_port);
   DataPath_RF_BLOCKi_58_Q_reg_17_inst : DFF_X1 port map( D => n5382, CK => CLK
                           , Q => n_1767, QN => 
                           DataPath_RF_bus_reg_dataout_1617_port);
   DataPath_RF_BLOCKi_58_Q_reg_16_inst : DFF_X1 port map( D => n5383, CK => CLK
                           , Q => n_1768, QN => 
                           DataPath_RF_bus_reg_dataout_1616_port);
   DataPath_RF_BLOCKi_58_Q_reg_15_inst : DFF_X1 port map( D => n5384, CK => CLK
                           , Q => n_1769, QN => 
                           DataPath_RF_bus_reg_dataout_1615_port);
   DataPath_RF_BLOCKi_58_Q_reg_14_inst : DFF_X1 port map( D => n5385, CK => CLK
                           , Q => n_1770, QN => 
                           DataPath_RF_bus_reg_dataout_1614_port);
   DataPath_RF_BLOCKi_58_Q_reg_13_inst : DFF_X1 port map( D => n5386, CK => CLK
                           , Q => n_1771, QN => 
                           DataPath_RF_bus_reg_dataout_1613_port);
   DataPath_RF_BLOCKi_58_Q_reg_12_inst : DFF_X1 port map( D => n5387, CK => CLK
                           , Q => n_1772, QN => 
                           DataPath_RF_bus_reg_dataout_1612_port);
   DataPath_RF_BLOCKi_58_Q_reg_11_inst : DFF_X1 port map( D => n5388, CK => CLK
                           , Q => n_1773, QN => 
                           DataPath_RF_bus_reg_dataout_1611_port);
   DataPath_RF_BLOCKi_58_Q_reg_9_inst : DFF_X1 port map( D => n5390, CK => CLK,
                           Q => n_1774, QN => 
                           DataPath_RF_bus_reg_dataout_1609_port);
   DataPath_RF_BLOCKi_58_Q_reg_8_inst : DFF_X1 port map( D => n5391, CK => CLK,
                           Q => n_1775, QN => 
                           DataPath_RF_bus_reg_dataout_1608_port);
   DataPath_RF_BLOCKi_58_Q_reg_7_inst : DFF_X1 port map( D => n5392, CK => CLK,
                           Q => n_1776, QN => 
                           DataPath_RF_bus_reg_dataout_1607_port);
   DataPath_RF_BLOCKi_58_Q_reg_6_inst : DFF_X1 port map( D => n5393, CK => CLK,
                           Q => n_1777, QN => 
                           DataPath_RF_bus_reg_dataout_1606_port);
   DataPath_RF_BLOCKi_58_Q_reg_5_inst : DFF_X1 port map( D => n5394, CK => CLK,
                           Q => n_1778, QN => 
                           DataPath_RF_bus_reg_dataout_1605_port);
   DataPath_RF_BLOCKi_58_Q_reg_4_inst : DFF_X1 port map( D => n5395, CK => CLK,
                           Q => n_1779, QN => 
                           DataPath_RF_bus_reg_dataout_1604_port);
   DataPath_RF_BLOCKi_58_Q_reg_3_inst : DFF_X1 port map( D => n5396, CK => CLK,
                           Q => n_1780, QN => 
                           DataPath_RF_bus_reg_dataout_1603_port);
   DataPath_RF_BLOCKi_58_Q_reg_2_inst : DFF_X1 port map( D => n5397, CK => CLK,
                           Q => n_1781, QN => 
                           DataPath_RF_bus_reg_dataout_1602_port);
   DataPath_RF_BLOCKi_58_Q_reg_1_inst : DFF_X1 port map( D => n5398, CK => CLK,
                           Q => n_1782, QN => 
                           DataPath_RF_bus_reg_dataout_1601_port);
   DataPath_RF_BLOCKi_58_Q_reg_0_inst : DFF_X1 port map( D => n5399, CK => CLK,
                           Q => n_1783, QN => 
                           DataPath_RF_bus_reg_dataout_1600_port);
   DataPath_RF_BLOCKi_74_Q_reg_31_inst : DFF_X1 port map( D => n5942, CK => CLK
                           , Q => n_1784, QN => 
                           DataPath_RF_bus_reg_dataout_2143_port);
   DataPath_RF_BLOCKi_74_Q_reg_30_inst : DFF_X1 port map( D => n5945, CK => CLK
                           , Q => n_1785, QN => 
                           DataPath_RF_bus_reg_dataout_2142_port);
   DataPath_RF_BLOCKi_74_Q_reg_29_inst : DFF_X1 port map( D => n5946, CK => CLK
                           , Q => n_1786, QN => 
                           DataPath_RF_bus_reg_dataout_2141_port);
   DataPath_RF_BLOCKi_74_Q_reg_28_inst : DFF_X1 port map( D => n5947, CK => CLK
                           , Q => n_1787, QN => 
                           DataPath_RF_bus_reg_dataout_2140_port);
   DataPath_RF_BLOCKi_74_Q_reg_27_inst : DFF_X1 port map( D => n5948, CK => CLK
                           , Q => n_1788, QN => 
                           DataPath_RF_bus_reg_dataout_2139_port);
   DataPath_RF_BLOCKi_74_Q_reg_26_inst : DFF_X1 port map( D => n5949, CK => CLK
                           , Q => n_1789, QN => 
                           DataPath_RF_bus_reg_dataout_2138_port);
   DataPath_RF_BLOCKi_74_Q_reg_25_inst : DFF_X1 port map( D => n5950, CK => CLK
                           , Q => n_1790, QN => 
                           DataPath_RF_bus_reg_dataout_2137_port);
   DataPath_RF_BLOCKi_74_Q_reg_24_inst : DFF_X1 port map( D => n5951, CK => CLK
                           , Q => n_1791, QN => 
                           DataPath_RF_bus_reg_dataout_2136_port);
   DataPath_RF_BLOCKi_74_Q_reg_23_inst : DFF_X1 port map( D => n5952, CK => CLK
                           , Q => n_1792, QN => 
                           DataPath_RF_bus_reg_dataout_2135_port);
   DataPath_RF_BLOCKi_74_Q_reg_22_inst : DFF_X1 port map( D => n5953, CK => CLK
                           , Q => n_1793, QN => 
                           DataPath_RF_bus_reg_dataout_2134_port);
   DataPath_RF_BLOCKi_74_Q_reg_21_inst : DFF_X1 port map( D => n5954, CK => CLK
                           , Q => n_1794, QN => 
                           DataPath_RF_bus_reg_dataout_2133_port);
   DataPath_RF_BLOCKi_74_Q_reg_20_inst : DFF_X1 port map( D => n5955, CK => CLK
                           , Q => n_1795, QN => 
                           DataPath_RF_bus_reg_dataout_2132_port);
   DataPath_RF_BLOCKi_74_Q_reg_19_inst : DFF_X1 port map( D => n5956, CK => CLK
                           , Q => n_1796, QN => 
                           DataPath_RF_bus_reg_dataout_2131_port);
   DataPath_RF_BLOCKi_74_Q_reg_18_inst : DFF_X1 port map( D => n5957, CK => CLK
                           , Q => n_1797, QN => 
                           DataPath_RF_bus_reg_dataout_2130_port);
   DataPath_RF_BLOCKi_74_Q_reg_17_inst : DFF_X1 port map( D => n5958, CK => CLK
                           , Q => n_1798, QN => 
                           DataPath_RF_bus_reg_dataout_2129_port);
   DataPath_RF_BLOCKi_74_Q_reg_16_inst : DFF_X1 port map( D => n5959, CK => CLK
                           , Q => n_1799, QN => 
                           DataPath_RF_bus_reg_dataout_2128_port);
   DataPath_RF_BLOCKi_74_Q_reg_15_inst : DFF_X1 port map( D => n5960, CK => CLK
                           , Q => n_1800, QN => 
                           DataPath_RF_bus_reg_dataout_2127_port);
   DataPath_RF_BLOCKi_74_Q_reg_14_inst : DFF_X1 port map( D => n5961, CK => CLK
                           , Q => n_1801, QN => 
                           DataPath_RF_bus_reg_dataout_2126_port);
   DataPath_RF_BLOCKi_74_Q_reg_13_inst : DFF_X1 port map( D => n5962, CK => CLK
                           , Q => n_1802, QN => 
                           DataPath_RF_bus_reg_dataout_2125_port);
   DataPath_RF_BLOCKi_74_Q_reg_12_inst : DFF_X1 port map( D => n5963, CK => CLK
                           , Q => n_1803, QN => 
                           DataPath_RF_bus_reg_dataout_2124_port);
   DataPath_RF_BLOCKi_74_Q_reg_11_inst : DFF_X1 port map( D => n5964, CK => CLK
                           , Q => n_1804, QN => 
                           DataPath_RF_bus_reg_dataout_2123_port);
   DataPath_RF_BLOCKi_74_Q_reg_9_inst : DFF_X1 port map( D => n5966, CK => CLK,
                           Q => n_1805, QN => 
                           DataPath_RF_bus_reg_dataout_2121_port);
   DataPath_RF_BLOCKi_74_Q_reg_8_inst : DFF_X1 port map( D => n5967, CK => CLK,
                           Q => n_1806, QN => 
                           DataPath_RF_bus_reg_dataout_2120_port);
   DataPath_RF_BLOCKi_74_Q_reg_7_inst : DFF_X1 port map( D => n5968, CK => CLK,
                           Q => n_1807, QN => 
                           DataPath_RF_bus_reg_dataout_2119_port);
   DataPath_RF_BLOCKi_74_Q_reg_6_inst : DFF_X1 port map( D => n5969, CK => CLK,
                           Q => n_1808, QN => 
                           DataPath_RF_bus_reg_dataout_2118_port);
   DataPath_RF_BLOCKi_74_Q_reg_5_inst : DFF_X1 port map( D => n5970, CK => CLK,
                           Q => n_1809, QN => 
                           DataPath_RF_bus_reg_dataout_2117_port);
   DataPath_RF_BLOCKi_74_Q_reg_4_inst : DFF_X1 port map( D => n5971, CK => CLK,
                           Q => n_1810, QN => 
                           DataPath_RF_bus_reg_dataout_2116_port);
   DataPath_RF_BLOCKi_74_Q_reg_3_inst : DFF_X1 port map( D => n5972, CK => CLK,
                           Q => n_1811, QN => 
                           DataPath_RF_bus_reg_dataout_2115_port);
   DataPath_RF_BLOCKi_74_Q_reg_2_inst : DFF_X1 port map( D => n5973, CK => CLK,
                           Q => n_1812, QN => 
                           DataPath_RF_bus_reg_dataout_2114_port);
   DataPath_RF_BLOCKi_74_Q_reg_1_inst : DFF_X1 port map( D => n5974, CK => CLK,
                           Q => n_1813, QN => 
                           DataPath_RF_bus_reg_dataout_2113_port);
   DataPath_RF_BLOCKi_74_Q_reg_0_inst : DFF_X1 port map( D => n5975, CK => CLK,
                           Q => n_1814, QN => 
                           DataPath_RF_bus_reg_dataout_2112_port);
   DataPath_RF_BLOCKi_11_Q_reg_31_inst : DFF_X1 port map( D => n3575, CK => CLK
                           , Q => n_1815, QN => 
                           DataPath_RF_bus_reg_dataout_127_port);
   DataPath_RF_BLOCKi_11_Q_reg_30_inst : DFF_X1 port map( D => n3578, CK => CLK
                           , Q => n_1816, QN => 
                           DataPath_RF_bus_reg_dataout_126_port);
   DataPath_RF_BLOCKi_11_Q_reg_29_inst : DFF_X1 port map( D => n3579, CK => CLK
                           , Q => n_1817, QN => 
                           DataPath_RF_bus_reg_dataout_125_port);
   DataPath_RF_BLOCKi_11_Q_reg_28_inst : DFF_X1 port map( D => n3580, CK => CLK
                           , Q => n_1818, QN => 
                           DataPath_RF_bus_reg_dataout_124_port);
   DataPath_RF_BLOCKi_11_Q_reg_27_inst : DFF_X1 port map( D => n3581, CK => CLK
                           , Q => n_1819, QN => 
                           DataPath_RF_bus_reg_dataout_123_port);
   DataPath_RF_BLOCKi_11_Q_reg_26_inst : DFF_X1 port map( D => n3582, CK => CLK
                           , Q => n_1820, QN => 
                           DataPath_RF_bus_reg_dataout_122_port);
   DataPath_RF_BLOCKi_11_Q_reg_25_inst : DFF_X1 port map( D => n3583, CK => CLK
                           , Q => n_1821, QN => 
                           DataPath_RF_bus_reg_dataout_121_port);
   DataPath_RF_BLOCKi_11_Q_reg_24_inst : DFF_X1 port map( D => n3584, CK => CLK
                           , Q => n_1822, QN => 
                           DataPath_RF_bus_reg_dataout_120_port);
   DataPath_RF_BLOCKi_11_Q_reg_23_inst : DFF_X1 port map( D => n3585, CK => CLK
                           , Q => n_1823, QN => 
                           DataPath_RF_bus_reg_dataout_119_port);
   DataPath_RF_BLOCKi_11_Q_reg_22_inst : DFF_X1 port map( D => n3586, CK => CLK
                           , Q => n_1824, QN => 
                           DataPath_RF_bus_reg_dataout_118_port);
   DataPath_RF_BLOCKi_11_Q_reg_21_inst : DFF_X1 port map( D => n3587, CK => CLK
                           , Q => n_1825, QN => 
                           DataPath_RF_bus_reg_dataout_117_port);
   DataPath_RF_BLOCKi_11_Q_reg_20_inst : DFF_X1 port map( D => n3588, CK => CLK
                           , Q => n_1826, QN => 
                           DataPath_RF_bus_reg_dataout_116_port);
   DataPath_RF_BLOCKi_11_Q_reg_19_inst : DFF_X1 port map( D => n3589, CK => CLK
                           , Q => n_1827, QN => 
                           DataPath_RF_bus_reg_dataout_115_port);
   DataPath_RF_BLOCKi_11_Q_reg_18_inst : DFF_X1 port map( D => n3590, CK => CLK
                           , Q => n_1828, QN => 
                           DataPath_RF_bus_reg_dataout_114_port);
   DataPath_RF_BLOCKi_11_Q_reg_17_inst : DFF_X1 port map( D => n3591, CK => CLK
                           , Q => n_1829, QN => 
                           DataPath_RF_bus_reg_dataout_113_port);
   DataPath_RF_BLOCKi_11_Q_reg_16_inst : DFF_X1 port map( D => n3592, CK => CLK
                           , Q => n_1830, QN => 
                           DataPath_RF_bus_reg_dataout_112_port);
   DataPath_RF_BLOCKi_11_Q_reg_15_inst : DFF_X1 port map( D => n3593, CK => CLK
                           , Q => n_1831, QN => 
                           DataPath_RF_bus_reg_dataout_111_port);
   DataPath_RF_BLOCKi_11_Q_reg_14_inst : DFF_X1 port map( D => n3594, CK => CLK
                           , Q => n_1832, QN => 
                           DataPath_RF_bus_reg_dataout_110_port);
   DataPath_RF_BLOCKi_11_Q_reg_13_inst : DFF_X1 port map( D => n3595, CK => CLK
                           , Q => n_1833, QN => 
                           DataPath_RF_bus_reg_dataout_109_port);
   DataPath_RF_BLOCKi_11_Q_reg_12_inst : DFF_X1 port map( D => n3596, CK => CLK
                           , Q => n_1834, QN => 
                           DataPath_RF_bus_reg_dataout_108_port);
   DataPath_RF_BLOCKi_11_Q_reg_11_inst : DFF_X1 port map( D => n3597, CK => CLK
                           , Q => n_1835, QN => 
                           DataPath_RF_bus_reg_dataout_107_port);
   DataPath_RF_BLOCKi_11_Q_reg_9_inst : DFF_X1 port map( D => n3599, CK => CLK,
                           Q => n_1836, QN => 
                           DataPath_RF_bus_reg_dataout_105_port);
   DataPath_RF_BLOCKi_11_Q_reg_8_inst : DFF_X1 port map( D => n3600, CK => CLK,
                           Q => n_1837, QN => 
                           DataPath_RF_bus_reg_dataout_104_port);
   DataPath_RF_BLOCKi_11_Q_reg_7_inst : DFF_X1 port map( D => n3601, CK => CLK,
                           Q => n_1838, QN => 
                           DataPath_RF_bus_reg_dataout_103_port);
   DataPath_RF_BLOCKi_11_Q_reg_6_inst : DFF_X1 port map( D => n3602, CK => CLK,
                           Q => n_1839, QN => 
                           DataPath_RF_bus_reg_dataout_102_port);
   DataPath_RF_BLOCKi_11_Q_reg_5_inst : DFF_X1 port map( D => n3603, CK => CLK,
                           Q => n_1840, QN => 
                           DataPath_RF_bus_reg_dataout_101_port);
   DataPath_RF_BLOCKi_11_Q_reg_4_inst : DFF_X1 port map( D => n3604, CK => CLK,
                           Q => n_1841, QN => 
                           DataPath_RF_bus_reg_dataout_100_port);
   DataPath_RF_BLOCKi_11_Q_reg_3_inst : DFF_X1 port map( D => n3605, CK => CLK,
                           Q => n_1842, QN => 
                           DataPath_RF_bus_reg_dataout_99_port);
   DataPath_RF_BLOCKi_11_Q_reg_2_inst : DFF_X1 port map( D => n3606, CK => CLK,
                           Q => n_1843, QN => 
                           DataPath_RF_bus_reg_dataout_98_port);
   DataPath_RF_BLOCKi_11_Q_reg_1_inst : DFF_X1 port map( D => n3607, CK => CLK,
                           Q => n_1844, QN => 
                           DataPath_RF_bus_reg_dataout_97_port);
   DataPath_RF_BLOCKi_11_Q_reg_0_inst : DFF_X1 port map( D => n3608, CK => CLK,
                           Q => n_1845, QN => 
                           DataPath_RF_bus_reg_dataout_96_port);
   DataPath_RF_BLOCKi_27_Q_reg_31_inst : DFF_X1 port map( D => n4215, CK => CLK
                           , Q => n_1846, QN => 
                           DataPath_RF_bus_reg_dataout_639_port);
   DataPath_RF_BLOCKi_27_Q_reg_30_inst : DFF_X1 port map( D => n4218, CK => CLK
                           , Q => n_1847, QN => 
                           DataPath_RF_bus_reg_dataout_638_port);
   DataPath_RF_BLOCKi_27_Q_reg_29_inst : DFF_X1 port map( D => n4219, CK => CLK
                           , Q => n_1848, QN => 
                           DataPath_RF_bus_reg_dataout_637_port);
   DataPath_RF_BLOCKi_27_Q_reg_28_inst : DFF_X1 port map( D => n4220, CK => CLK
                           , Q => n_1849, QN => 
                           DataPath_RF_bus_reg_dataout_636_port);
   DataPath_RF_BLOCKi_27_Q_reg_27_inst : DFF_X1 port map( D => n4221, CK => CLK
                           , Q => n_1850, QN => 
                           DataPath_RF_bus_reg_dataout_635_port);
   DataPath_RF_BLOCKi_27_Q_reg_26_inst : DFF_X1 port map( D => n4222, CK => CLK
                           , Q => n_1851, QN => 
                           DataPath_RF_bus_reg_dataout_634_port);
   DataPath_RF_BLOCKi_27_Q_reg_25_inst : DFF_X1 port map( D => n4223, CK => CLK
                           , Q => n_1852, QN => 
                           DataPath_RF_bus_reg_dataout_633_port);
   DataPath_RF_BLOCKi_27_Q_reg_24_inst : DFF_X1 port map( D => n4224, CK => CLK
                           , Q => n_1853, QN => 
                           DataPath_RF_bus_reg_dataout_632_port);
   DataPath_RF_BLOCKi_27_Q_reg_23_inst : DFF_X1 port map( D => n4225, CK => CLK
                           , Q => n_1854, QN => 
                           DataPath_RF_bus_reg_dataout_631_port);
   DataPath_RF_BLOCKi_27_Q_reg_22_inst : DFF_X1 port map( D => n4226, CK => CLK
                           , Q => n_1855, QN => 
                           DataPath_RF_bus_reg_dataout_630_port);
   DataPath_RF_BLOCKi_27_Q_reg_21_inst : DFF_X1 port map( D => n4227, CK => CLK
                           , Q => n_1856, QN => 
                           DataPath_RF_bus_reg_dataout_629_port);
   DataPath_RF_BLOCKi_27_Q_reg_20_inst : DFF_X1 port map( D => n4228, CK => CLK
                           , Q => n_1857, QN => 
                           DataPath_RF_bus_reg_dataout_628_port);
   DataPath_RF_BLOCKi_27_Q_reg_19_inst : DFF_X1 port map( D => n4229, CK => CLK
                           , Q => n_1858, QN => 
                           DataPath_RF_bus_reg_dataout_627_port);
   DataPath_RF_BLOCKi_27_Q_reg_18_inst : DFF_X1 port map( D => n4230, CK => CLK
                           , Q => n_1859, QN => 
                           DataPath_RF_bus_reg_dataout_626_port);
   DataPath_RF_BLOCKi_27_Q_reg_17_inst : DFF_X1 port map( D => n4231, CK => CLK
                           , Q => n_1860, QN => 
                           DataPath_RF_bus_reg_dataout_625_port);
   DataPath_RF_BLOCKi_27_Q_reg_16_inst : DFF_X1 port map( D => n4232, CK => CLK
                           , Q => n_1861, QN => 
                           DataPath_RF_bus_reg_dataout_624_port);
   DataPath_RF_BLOCKi_27_Q_reg_15_inst : DFF_X1 port map( D => n4233, CK => CLK
                           , Q => n_1862, QN => 
                           DataPath_RF_bus_reg_dataout_623_port);
   DataPath_RF_BLOCKi_27_Q_reg_14_inst : DFF_X1 port map( D => n4234, CK => CLK
                           , Q => n_1863, QN => 
                           DataPath_RF_bus_reg_dataout_622_port);
   DataPath_RF_BLOCKi_27_Q_reg_13_inst : DFF_X1 port map( D => n4235, CK => CLK
                           , Q => n_1864, QN => 
                           DataPath_RF_bus_reg_dataout_621_port);
   DataPath_RF_BLOCKi_27_Q_reg_12_inst : DFF_X1 port map( D => n4236, CK => CLK
                           , Q => n_1865, QN => 
                           DataPath_RF_bus_reg_dataout_620_port);
   DataPath_RF_BLOCKi_27_Q_reg_11_inst : DFF_X1 port map( D => n4237, CK => CLK
                           , Q => n_1866, QN => 
                           DataPath_RF_bus_reg_dataout_619_port);
   DataPath_RF_BLOCKi_27_Q_reg_9_inst : DFF_X1 port map( D => n4239, CK => CLK,
                           Q => n_1867, QN => 
                           DataPath_RF_bus_reg_dataout_617_port);
   DataPath_RF_BLOCKi_27_Q_reg_8_inst : DFF_X1 port map( D => n4240, CK => CLK,
                           Q => n_1868, QN => 
                           DataPath_RF_bus_reg_dataout_616_port);
   DataPath_RF_BLOCKi_27_Q_reg_7_inst : DFF_X1 port map( D => n4241, CK => CLK,
                           Q => n_1869, QN => 
                           DataPath_RF_bus_reg_dataout_615_port);
   DataPath_RF_BLOCKi_27_Q_reg_6_inst : DFF_X1 port map( D => n4242, CK => CLK,
                           Q => n_1870, QN => 
                           DataPath_RF_bus_reg_dataout_614_port);
   DataPath_RF_BLOCKi_27_Q_reg_5_inst : DFF_X1 port map( D => n4243, CK => CLK,
                           Q => n_1871, QN => 
                           DataPath_RF_bus_reg_dataout_613_port);
   DataPath_RF_BLOCKi_27_Q_reg_4_inst : DFF_X1 port map( D => n4244, CK => CLK,
                           Q => n_1872, QN => 
                           DataPath_RF_bus_reg_dataout_612_port);
   DataPath_RF_BLOCKi_27_Q_reg_3_inst : DFF_X1 port map( D => n4245, CK => CLK,
                           Q => n_1873, QN => 
                           DataPath_RF_bus_reg_dataout_611_port);
   DataPath_RF_BLOCKi_27_Q_reg_2_inst : DFF_X1 port map( D => n4246, CK => CLK,
                           Q => n_1874, QN => 
                           DataPath_RF_bus_reg_dataout_610_port);
   DataPath_RF_BLOCKi_27_Q_reg_1_inst : DFF_X1 port map( D => n4247, CK => CLK,
                           Q => n_1875, QN => 
                           DataPath_RF_bus_reg_dataout_609_port);
   DataPath_RF_BLOCKi_27_Q_reg_0_inst : DFF_X1 port map( D => n4248, CK => CLK,
                           Q => n_1876, QN => 
                           DataPath_RF_bus_reg_dataout_608_port);
   DataPath_RF_BLOCKi_43_Q_reg_31_inst : DFF_X1 port map( D => n4808, CK => CLK
                           , Q => n_1877, QN => 
                           DataPath_RF_bus_reg_dataout_1151_port);
   DataPath_RF_BLOCKi_43_Q_reg_30_inst : DFF_X1 port map( D => n4811, CK => CLK
                           , Q => n_1878, QN => 
                           DataPath_RF_bus_reg_dataout_1150_port);
   DataPath_RF_BLOCKi_43_Q_reg_29_inst : DFF_X1 port map( D => n4812, CK => CLK
                           , Q => n_1879, QN => 
                           DataPath_RF_bus_reg_dataout_1149_port);
   DataPath_RF_BLOCKi_43_Q_reg_28_inst : DFF_X1 port map( D => n4813, CK => CLK
                           , Q => n_1880, QN => 
                           DataPath_RF_bus_reg_dataout_1148_port);
   DataPath_RF_BLOCKi_43_Q_reg_27_inst : DFF_X1 port map( D => n4814, CK => CLK
                           , Q => n_1881, QN => 
                           DataPath_RF_bus_reg_dataout_1147_port);
   DataPath_RF_BLOCKi_43_Q_reg_26_inst : DFF_X1 port map( D => n4815, CK => CLK
                           , Q => n_1882, QN => 
                           DataPath_RF_bus_reg_dataout_1146_port);
   DataPath_RF_BLOCKi_43_Q_reg_25_inst : DFF_X1 port map( D => n4816, CK => CLK
                           , Q => n_1883, QN => 
                           DataPath_RF_bus_reg_dataout_1145_port);
   DataPath_RF_BLOCKi_43_Q_reg_24_inst : DFF_X1 port map( D => n4817, CK => CLK
                           , Q => n_1884, QN => 
                           DataPath_RF_bus_reg_dataout_1144_port);
   DataPath_RF_BLOCKi_43_Q_reg_23_inst : DFF_X1 port map( D => n4818, CK => CLK
                           , Q => n_1885, QN => 
                           DataPath_RF_bus_reg_dataout_1143_port);
   DataPath_RF_BLOCKi_43_Q_reg_22_inst : DFF_X1 port map( D => n4819, CK => CLK
                           , Q => n_1886, QN => 
                           DataPath_RF_bus_reg_dataout_1142_port);
   DataPath_RF_BLOCKi_43_Q_reg_21_inst : DFF_X1 port map( D => n4820, CK => CLK
                           , Q => n_1887, QN => 
                           DataPath_RF_bus_reg_dataout_1141_port);
   DataPath_RF_BLOCKi_43_Q_reg_20_inst : DFF_X1 port map( D => n4821, CK => CLK
                           , Q => n_1888, QN => 
                           DataPath_RF_bus_reg_dataout_1140_port);
   DataPath_RF_BLOCKi_43_Q_reg_19_inst : DFF_X1 port map( D => n4822, CK => CLK
                           , Q => n_1889, QN => 
                           DataPath_RF_bus_reg_dataout_1139_port);
   DataPath_RF_BLOCKi_43_Q_reg_18_inst : DFF_X1 port map( D => n4823, CK => CLK
                           , Q => n_1890, QN => 
                           DataPath_RF_bus_reg_dataout_1138_port);
   DataPath_RF_BLOCKi_43_Q_reg_17_inst : DFF_X1 port map( D => n4824, CK => CLK
                           , Q => n_1891, QN => 
                           DataPath_RF_bus_reg_dataout_1137_port);
   DataPath_RF_BLOCKi_43_Q_reg_16_inst : DFF_X1 port map( D => n4825, CK => CLK
                           , Q => n_1892, QN => 
                           DataPath_RF_bus_reg_dataout_1136_port);
   DataPath_RF_BLOCKi_43_Q_reg_15_inst : DFF_X1 port map( D => n4826, CK => CLK
                           , Q => n_1893, QN => 
                           DataPath_RF_bus_reg_dataout_1135_port);
   DataPath_RF_BLOCKi_43_Q_reg_14_inst : DFF_X1 port map( D => n4827, CK => CLK
                           , Q => n_1894, QN => 
                           DataPath_RF_bus_reg_dataout_1134_port);
   DataPath_RF_BLOCKi_43_Q_reg_13_inst : DFF_X1 port map( D => n4828, CK => CLK
                           , Q => n_1895, QN => 
                           DataPath_RF_bus_reg_dataout_1133_port);
   DataPath_RF_BLOCKi_43_Q_reg_12_inst : DFF_X1 port map( D => n4829, CK => CLK
                           , Q => n_1896, QN => 
                           DataPath_RF_bus_reg_dataout_1132_port);
   DataPath_RF_BLOCKi_43_Q_reg_11_inst : DFF_X1 port map( D => n4830, CK => CLK
                           , Q => n_1897, QN => 
                           DataPath_RF_bus_reg_dataout_1131_port);
   DataPath_RF_BLOCKi_43_Q_reg_9_inst : DFF_X1 port map( D => n4832, CK => CLK,
                           Q => n_1898, QN => 
                           DataPath_RF_bus_reg_dataout_1129_port);
   DataPath_RF_BLOCKi_43_Q_reg_8_inst : DFF_X1 port map( D => n4833, CK => CLK,
                           Q => n_1899, QN => 
                           DataPath_RF_bus_reg_dataout_1128_port);
   DataPath_RF_BLOCKi_43_Q_reg_7_inst : DFF_X1 port map( D => n4834, CK => CLK,
                           Q => n_1900, QN => 
                           DataPath_RF_bus_reg_dataout_1127_port);
   DataPath_RF_BLOCKi_43_Q_reg_6_inst : DFF_X1 port map( D => n4835, CK => CLK,
                           Q => n_1901, QN => 
                           DataPath_RF_bus_reg_dataout_1126_port);
   DataPath_RF_BLOCKi_43_Q_reg_5_inst : DFF_X1 port map( D => n4836, CK => CLK,
                           Q => n_1902, QN => 
                           DataPath_RF_bus_reg_dataout_1125_port);
   DataPath_RF_BLOCKi_43_Q_reg_4_inst : DFF_X1 port map( D => n4837, CK => CLK,
                           Q => n_1903, QN => 
                           DataPath_RF_bus_reg_dataout_1124_port);
   DataPath_RF_BLOCKi_43_Q_reg_3_inst : DFF_X1 port map( D => n4838, CK => CLK,
                           Q => n_1904, QN => 
                           DataPath_RF_bus_reg_dataout_1123_port);
   DataPath_RF_BLOCKi_43_Q_reg_2_inst : DFF_X1 port map( D => n4839, CK => CLK,
                           Q => n_1905, QN => 
                           DataPath_RF_bus_reg_dataout_1122_port);
   DataPath_RF_BLOCKi_43_Q_reg_1_inst : DFF_X1 port map( D => n4840, CK => CLK,
                           Q => n_1906, QN => 
                           DataPath_RF_bus_reg_dataout_1121_port);
   DataPath_RF_BLOCKi_43_Q_reg_0_inst : DFF_X1 port map( D => n4841, CK => CLK,
                           Q => n_1907, QN => 
                           DataPath_RF_bus_reg_dataout_1120_port);
   DataPath_RF_BLOCKi_59_Q_reg_31_inst : DFF_X1 port map( D => n5401, CK => CLK
                           , Q => n_1908, QN => 
                           DataPath_RF_bus_reg_dataout_1663_port);
   DataPath_RF_BLOCKi_59_Q_reg_30_inst : DFF_X1 port map( D => n5404, CK => CLK
                           , Q => n_1909, QN => 
                           DataPath_RF_bus_reg_dataout_1662_port);
   DataPath_RF_BLOCKi_59_Q_reg_29_inst : DFF_X1 port map( D => n5405, CK => CLK
                           , Q => n_1910, QN => 
                           DataPath_RF_bus_reg_dataout_1661_port);
   DataPath_RF_BLOCKi_59_Q_reg_28_inst : DFF_X1 port map( D => n5406, CK => CLK
                           , Q => n_1911, QN => 
                           DataPath_RF_bus_reg_dataout_1660_port);
   DataPath_RF_BLOCKi_59_Q_reg_27_inst : DFF_X1 port map( D => n5407, CK => CLK
                           , Q => n_1912, QN => 
                           DataPath_RF_bus_reg_dataout_1659_port);
   DataPath_RF_BLOCKi_59_Q_reg_26_inst : DFF_X1 port map( D => n5408, CK => CLK
                           , Q => n_1913, QN => 
                           DataPath_RF_bus_reg_dataout_1658_port);
   DataPath_RF_BLOCKi_59_Q_reg_25_inst : DFF_X1 port map( D => n5409, CK => CLK
                           , Q => n_1914, QN => 
                           DataPath_RF_bus_reg_dataout_1657_port);
   DataPath_RF_BLOCKi_59_Q_reg_24_inst : DFF_X1 port map( D => n5410, CK => CLK
                           , Q => n_1915, QN => 
                           DataPath_RF_bus_reg_dataout_1656_port);
   DataPath_RF_BLOCKi_59_Q_reg_23_inst : DFF_X1 port map( D => n5411, CK => CLK
                           , Q => n_1916, QN => 
                           DataPath_RF_bus_reg_dataout_1655_port);
   DataPath_RF_BLOCKi_59_Q_reg_22_inst : DFF_X1 port map( D => n5412, CK => CLK
                           , Q => n_1917, QN => 
                           DataPath_RF_bus_reg_dataout_1654_port);
   DataPath_RF_BLOCKi_59_Q_reg_21_inst : DFF_X1 port map( D => n5413, CK => CLK
                           , Q => n_1918, QN => 
                           DataPath_RF_bus_reg_dataout_1653_port);
   DataPath_RF_BLOCKi_59_Q_reg_20_inst : DFF_X1 port map( D => n5414, CK => CLK
                           , Q => n_1919, QN => 
                           DataPath_RF_bus_reg_dataout_1652_port);
   DataPath_RF_BLOCKi_59_Q_reg_19_inst : DFF_X1 port map( D => n5415, CK => CLK
                           , Q => n_1920, QN => 
                           DataPath_RF_bus_reg_dataout_1651_port);
   DataPath_RF_BLOCKi_59_Q_reg_18_inst : DFF_X1 port map( D => n5416, CK => CLK
                           , Q => n_1921, QN => 
                           DataPath_RF_bus_reg_dataout_1650_port);
   DataPath_RF_BLOCKi_59_Q_reg_17_inst : DFF_X1 port map( D => n5417, CK => CLK
                           , Q => n_1922, QN => 
                           DataPath_RF_bus_reg_dataout_1649_port);
   DataPath_RF_BLOCKi_59_Q_reg_16_inst : DFF_X1 port map( D => n5418, CK => CLK
                           , Q => n_1923, QN => 
                           DataPath_RF_bus_reg_dataout_1648_port);
   DataPath_RF_BLOCKi_59_Q_reg_15_inst : DFF_X1 port map( D => n5419, CK => CLK
                           , Q => n_1924, QN => 
                           DataPath_RF_bus_reg_dataout_1647_port);
   DataPath_RF_BLOCKi_59_Q_reg_14_inst : DFF_X1 port map( D => n5420, CK => CLK
                           , Q => n_1925, QN => 
                           DataPath_RF_bus_reg_dataout_1646_port);
   DataPath_RF_BLOCKi_59_Q_reg_13_inst : DFF_X1 port map( D => n5421, CK => CLK
                           , Q => n_1926, QN => 
                           DataPath_RF_bus_reg_dataout_1645_port);
   DataPath_RF_BLOCKi_59_Q_reg_12_inst : DFF_X1 port map( D => n5422, CK => CLK
                           , Q => n_1927, QN => 
                           DataPath_RF_bus_reg_dataout_1644_port);
   DataPath_RF_BLOCKi_59_Q_reg_11_inst : DFF_X1 port map( D => n5423, CK => CLK
                           , Q => n_1928, QN => 
                           DataPath_RF_bus_reg_dataout_1643_port);
   DataPath_RF_BLOCKi_59_Q_reg_9_inst : DFF_X1 port map( D => n5425, CK => CLK,
                           Q => n_1929, QN => 
                           DataPath_RF_bus_reg_dataout_1641_port);
   DataPath_RF_BLOCKi_59_Q_reg_8_inst : DFF_X1 port map( D => n5426, CK => CLK,
                           Q => n_1930, QN => 
                           DataPath_RF_bus_reg_dataout_1640_port);
   DataPath_RF_BLOCKi_59_Q_reg_7_inst : DFF_X1 port map( D => n5427, CK => CLK,
                           Q => n_1931, QN => 
                           DataPath_RF_bus_reg_dataout_1639_port);
   DataPath_RF_BLOCKi_59_Q_reg_6_inst : DFF_X1 port map( D => n5428, CK => CLK,
                           Q => n_1932, QN => 
                           DataPath_RF_bus_reg_dataout_1638_port);
   DataPath_RF_BLOCKi_59_Q_reg_5_inst : DFF_X1 port map( D => n5429, CK => CLK,
                           Q => n_1933, QN => 
                           DataPath_RF_bus_reg_dataout_1637_port);
   DataPath_RF_BLOCKi_59_Q_reg_4_inst : DFF_X1 port map( D => n5430, CK => CLK,
                           Q => n_1934, QN => 
                           DataPath_RF_bus_reg_dataout_1636_port);
   DataPath_RF_BLOCKi_59_Q_reg_3_inst : DFF_X1 port map( D => n5431, CK => CLK,
                           Q => n_1935, QN => 
                           DataPath_RF_bus_reg_dataout_1635_port);
   DataPath_RF_BLOCKi_59_Q_reg_2_inst : DFF_X1 port map( D => n5432, CK => CLK,
                           Q => n_1936, QN => 
                           DataPath_RF_bus_reg_dataout_1634_port);
   DataPath_RF_BLOCKi_59_Q_reg_1_inst : DFF_X1 port map( D => n5433, CK => CLK,
                           Q => n_1937, QN => 
                           DataPath_RF_bus_reg_dataout_1633_port);
   DataPath_RF_BLOCKi_59_Q_reg_0_inst : DFF_X1 port map( D => n5434, CK => CLK,
                           Q => n_1938, QN => 
                           DataPath_RF_bus_reg_dataout_1632_port);
   DataPath_RF_BLOCKi_75_Q_reg_31_inst : DFF_X1 port map( D => n5979, CK => CLK
                           , Q => n_1939, QN => 
                           DataPath_RF_bus_reg_dataout_2175_port);
   DataPath_RF_BLOCKi_75_Q_reg_30_inst : DFF_X1 port map( D => n5982, CK => CLK
                           , Q => n_1940, QN => 
                           DataPath_RF_bus_reg_dataout_2174_port);
   DataPath_RF_BLOCKi_75_Q_reg_29_inst : DFF_X1 port map( D => n5983, CK => CLK
                           , Q => n_1941, QN => 
                           DataPath_RF_bus_reg_dataout_2173_port);
   DataPath_RF_BLOCKi_75_Q_reg_28_inst : DFF_X1 port map( D => n5984, CK => CLK
                           , Q => n_1942, QN => 
                           DataPath_RF_bus_reg_dataout_2172_port);
   DataPath_RF_BLOCKi_75_Q_reg_27_inst : DFF_X1 port map( D => n5985, CK => CLK
                           , Q => n_1943, QN => 
                           DataPath_RF_bus_reg_dataout_2171_port);
   DataPath_RF_BLOCKi_75_Q_reg_26_inst : DFF_X1 port map( D => n5986, CK => CLK
                           , Q => n_1944, QN => 
                           DataPath_RF_bus_reg_dataout_2170_port);
   DataPath_RF_BLOCKi_75_Q_reg_25_inst : DFF_X1 port map( D => n5987, CK => CLK
                           , Q => n_1945, QN => 
                           DataPath_RF_bus_reg_dataout_2169_port);
   DataPath_RF_BLOCKi_75_Q_reg_24_inst : DFF_X1 port map( D => n5988, CK => CLK
                           , Q => n_1946, QN => 
                           DataPath_RF_bus_reg_dataout_2168_port);
   DataPath_RF_BLOCKi_75_Q_reg_23_inst : DFF_X1 port map( D => n5989, CK => CLK
                           , Q => n_1947, QN => 
                           DataPath_RF_bus_reg_dataout_2167_port);
   DataPath_RF_BLOCKi_75_Q_reg_22_inst : DFF_X1 port map( D => n5990, CK => CLK
                           , Q => n_1948, QN => 
                           DataPath_RF_bus_reg_dataout_2166_port);
   DataPath_RF_BLOCKi_75_Q_reg_21_inst : DFF_X1 port map( D => n5991, CK => CLK
                           , Q => n_1949, QN => 
                           DataPath_RF_bus_reg_dataout_2165_port);
   DataPath_RF_BLOCKi_75_Q_reg_20_inst : DFF_X1 port map( D => n5992, CK => CLK
                           , Q => n_1950, QN => 
                           DataPath_RF_bus_reg_dataout_2164_port);
   DataPath_RF_BLOCKi_75_Q_reg_19_inst : DFF_X1 port map( D => n5993, CK => CLK
                           , Q => n_1951, QN => 
                           DataPath_RF_bus_reg_dataout_2163_port);
   DataPath_RF_BLOCKi_75_Q_reg_18_inst : DFF_X1 port map( D => n5994, CK => CLK
                           , Q => n_1952, QN => 
                           DataPath_RF_bus_reg_dataout_2162_port);
   DataPath_RF_BLOCKi_75_Q_reg_17_inst : DFF_X1 port map( D => n5995, CK => CLK
                           , Q => n_1953, QN => 
                           DataPath_RF_bus_reg_dataout_2161_port);
   DataPath_RF_BLOCKi_75_Q_reg_16_inst : DFF_X1 port map( D => n5996, CK => CLK
                           , Q => n_1954, QN => 
                           DataPath_RF_bus_reg_dataout_2160_port);
   DataPath_RF_BLOCKi_75_Q_reg_15_inst : DFF_X1 port map( D => n5997, CK => CLK
                           , Q => n_1955, QN => 
                           DataPath_RF_bus_reg_dataout_2159_port);
   DataPath_RF_BLOCKi_75_Q_reg_14_inst : DFF_X1 port map( D => n5998, CK => CLK
                           , Q => n_1956, QN => 
                           DataPath_RF_bus_reg_dataout_2158_port);
   DataPath_RF_BLOCKi_75_Q_reg_13_inst : DFF_X1 port map( D => n5999, CK => CLK
                           , Q => n_1957, QN => 
                           DataPath_RF_bus_reg_dataout_2157_port);
   DataPath_RF_BLOCKi_75_Q_reg_12_inst : DFF_X1 port map( D => n6000, CK => CLK
                           , Q => n_1958, QN => 
                           DataPath_RF_bus_reg_dataout_2156_port);
   DataPath_RF_BLOCKi_75_Q_reg_11_inst : DFF_X1 port map( D => n6001, CK => CLK
                           , Q => n_1959, QN => 
                           DataPath_RF_bus_reg_dataout_2155_port);
   DataPath_RF_BLOCKi_75_Q_reg_9_inst : DFF_X1 port map( D => n6003, CK => CLK,
                           Q => n_1960, QN => 
                           DataPath_RF_bus_reg_dataout_2153_port);
   DataPath_RF_BLOCKi_75_Q_reg_8_inst : DFF_X1 port map( D => n6004, CK => CLK,
                           Q => n_1961, QN => 
                           DataPath_RF_bus_reg_dataout_2152_port);
   DataPath_RF_BLOCKi_75_Q_reg_7_inst : DFF_X1 port map( D => n6005, CK => CLK,
                           Q => n_1962, QN => 
                           DataPath_RF_bus_reg_dataout_2151_port);
   DataPath_RF_BLOCKi_75_Q_reg_6_inst : DFF_X1 port map( D => n6006, CK => CLK,
                           Q => n_1963, QN => 
                           DataPath_RF_bus_reg_dataout_2150_port);
   DataPath_RF_BLOCKi_75_Q_reg_5_inst : DFF_X1 port map( D => n6007, CK => CLK,
                           Q => n_1964, QN => 
                           DataPath_RF_bus_reg_dataout_2149_port);
   DataPath_RF_BLOCKi_75_Q_reg_4_inst : DFF_X1 port map( D => n6008, CK => CLK,
                           Q => n_1965, QN => 
                           DataPath_RF_bus_reg_dataout_2148_port);
   DataPath_RF_BLOCKi_75_Q_reg_3_inst : DFF_X1 port map( D => n6009, CK => CLK,
                           Q => n_1966, QN => 
                           DataPath_RF_bus_reg_dataout_2147_port);
   DataPath_RF_BLOCKi_75_Q_reg_2_inst : DFF_X1 port map( D => n6010, CK => CLK,
                           Q => n_1967, QN => 
                           DataPath_RF_bus_reg_dataout_2146_port);
   DataPath_RF_BLOCKi_75_Q_reg_1_inst : DFF_X1 port map( D => n6011, CK => CLK,
                           Q => n_1968, QN => 
                           DataPath_RF_bus_reg_dataout_2145_port);
   DataPath_RF_BLOCKi_75_Q_reg_0_inst : DFF_X1 port map( D => n6012, CK => CLK,
                           Q => n_1969, QN => 
                           DataPath_RF_bus_reg_dataout_2144_port);
   DataPath_RF_BLOCKi_12_Q_reg_31_inst : DFF_X1 port map( D => n3613, CK => CLK
                           , Q => n_1970, QN => 
                           DataPath_RF_bus_reg_dataout_159_port);
   DataPath_RF_BLOCKi_12_Q_reg_30_inst : DFF_X1 port map( D => n3616, CK => CLK
                           , Q => n_1971, QN => 
                           DataPath_RF_bus_reg_dataout_158_port);
   DataPath_RF_BLOCKi_12_Q_reg_29_inst : DFF_X1 port map( D => n3617, CK => CLK
                           , Q => n_1972, QN => 
                           DataPath_RF_bus_reg_dataout_157_port);
   DataPath_RF_BLOCKi_12_Q_reg_28_inst : DFF_X1 port map( D => n3618, CK => CLK
                           , Q => n_1973, QN => 
                           DataPath_RF_bus_reg_dataout_156_port);
   DataPath_RF_BLOCKi_12_Q_reg_27_inst : DFF_X1 port map( D => n3619, CK => CLK
                           , Q => n_1974, QN => 
                           DataPath_RF_bus_reg_dataout_155_port);
   DataPath_RF_BLOCKi_12_Q_reg_26_inst : DFF_X1 port map( D => n3620, CK => CLK
                           , Q => n_1975, QN => 
                           DataPath_RF_bus_reg_dataout_154_port);
   DataPath_RF_BLOCKi_12_Q_reg_25_inst : DFF_X1 port map( D => n3621, CK => CLK
                           , Q => n_1976, QN => 
                           DataPath_RF_bus_reg_dataout_153_port);
   DataPath_RF_BLOCKi_12_Q_reg_24_inst : DFF_X1 port map( D => n3622, CK => CLK
                           , Q => n_1977, QN => 
                           DataPath_RF_bus_reg_dataout_152_port);
   DataPath_RF_BLOCKi_12_Q_reg_23_inst : DFF_X1 port map( D => n3623, CK => CLK
                           , Q => n_1978, QN => 
                           DataPath_RF_bus_reg_dataout_151_port);
   DataPath_RF_BLOCKi_12_Q_reg_22_inst : DFF_X1 port map( D => n3624, CK => CLK
                           , Q => n_1979, QN => 
                           DataPath_RF_bus_reg_dataout_150_port);
   DataPath_RF_BLOCKi_12_Q_reg_21_inst : DFF_X1 port map( D => n3625, CK => CLK
                           , Q => n_1980, QN => 
                           DataPath_RF_bus_reg_dataout_149_port);
   DataPath_RF_BLOCKi_12_Q_reg_20_inst : DFF_X1 port map( D => n3626, CK => CLK
                           , Q => n_1981, QN => 
                           DataPath_RF_bus_reg_dataout_148_port);
   DataPath_RF_BLOCKi_12_Q_reg_19_inst : DFF_X1 port map( D => n3627, CK => CLK
                           , Q => n_1982, QN => 
                           DataPath_RF_bus_reg_dataout_147_port);
   DataPath_RF_BLOCKi_12_Q_reg_18_inst : DFF_X1 port map( D => n3628, CK => CLK
                           , Q => n_1983, QN => 
                           DataPath_RF_bus_reg_dataout_146_port);
   DataPath_RF_BLOCKi_12_Q_reg_17_inst : DFF_X1 port map( D => n3629, CK => CLK
                           , Q => n_1984, QN => 
                           DataPath_RF_bus_reg_dataout_145_port);
   DataPath_RF_BLOCKi_12_Q_reg_16_inst : DFF_X1 port map( D => n3630, CK => CLK
                           , Q => n_1985, QN => 
                           DataPath_RF_bus_reg_dataout_144_port);
   DataPath_RF_BLOCKi_12_Q_reg_15_inst : DFF_X1 port map( D => n3631, CK => CLK
                           , Q => n_1986, QN => 
                           DataPath_RF_bus_reg_dataout_143_port);
   DataPath_RF_BLOCKi_12_Q_reg_14_inst : DFF_X1 port map( D => n3632, CK => CLK
                           , Q => n_1987, QN => 
                           DataPath_RF_bus_reg_dataout_142_port);
   DataPath_RF_BLOCKi_12_Q_reg_13_inst : DFF_X1 port map( D => n3633, CK => CLK
                           , Q => n_1988, QN => 
                           DataPath_RF_bus_reg_dataout_141_port);
   DataPath_RF_BLOCKi_12_Q_reg_12_inst : DFF_X1 port map( D => n3634, CK => CLK
                           , Q => n_1989, QN => 
                           DataPath_RF_bus_reg_dataout_140_port);
   DataPath_RF_BLOCKi_12_Q_reg_11_inst : DFF_X1 port map( D => n3635, CK => CLK
                           , Q => n_1990, QN => 
                           DataPath_RF_bus_reg_dataout_139_port);
   DataPath_RF_BLOCKi_12_Q_reg_9_inst : DFF_X1 port map( D => n3637, CK => CLK,
                           Q => n_1991, QN => 
                           DataPath_RF_bus_reg_dataout_137_port);
   DataPath_RF_BLOCKi_12_Q_reg_8_inst : DFF_X1 port map( D => n3638, CK => CLK,
                           Q => n_1992, QN => 
                           DataPath_RF_bus_reg_dataout_136_port);
   DataPath_RF_BLOCKi_12_Q_reg_7_inst : DFF_X1 port map( D => n3639, CK => CLK,
                           Q => n_1993, QN => 
                           DataPath_RF_bus_reg_dataout_135_port);
   DataPath_RF_BLOCKi_12_Q_reg_6_inst : DFF_X1 port map( D => n3640, CK => CLK,
                           Q => n_1994, QN => 
                           DataPath_RF_bus_reg_dataout_134_port);
   DataPath_RF_BLOCKi_12_Q_reg_5_inst : DFF_X1 port map( D => n3641, CK => CLK,
                           Q => n_1995, QN => 
                           DataPath_RF_bus_reg_dataout_133_port);
   DataPath_RF_BLOCKi_12_Q_reg_4_inst : DFF_X1 port map( D => n3642, CK => CLK,
                           Q => n_1996, QN => 
                           DataPath_RF_bus_reg_dataout_132_port);
   DataPath_RF_BLOCKi_12_Q_reg_3_inst : DFF_X1 port map( D => n3643, CK => CLK,
                           Q => n_1997, QN => 
                           DataPath_RF_bus_reg_dataout_131_port);
   DataPath_RF_BLOCKi_12_Q_reg_2_inst : DFF_X1 port map( D => n3644, CK => CLK,
                           Q => n_1998, QN => 
                           DataPath_RF_bus_reg_dataout_130_port);
   DataPath_RF_BLOCKi_12_Q_reg_1_inst : DFF_X1 port map( D => n3645, CK => CLK,
                           Q => n_1999, QN => 
                           DataPath_RF_bus_reg_dataout_129_port);
   DataPath_RF_BLOCKi_12_Q_reg_0_inst : DFF_X1 port map( D => n3646, CK => CLK,
                           Q => n_2000, QN => 
                           DataPath_RF_bus_reg_dataout_128_port);
   DataPath_RF_BLOCKi_28_Q_reg_31_inst : DFF_X1 port map( D => n4250, CK => CLK
                           , Q => n_2001, QN => 
                           DataPath_RF_bus_reg_dataout_671_port);
   DataPath_RF_BLOCKi_28_Q_reg_30_inst : DFF_X1 port map( D => n4253, CK => CLK
                           , Q => n_2002, QN => 
                           DataPath_RF_bus_reg_dataout_670_port);
   DataPath_RF_BLOCKi_28_Q_reg_29_inst : DFF_X1 port map( D => n4254, CK => CLK
                           , Q => n_2003, QN => 
                           DataPath_RF_bus_reg_dataout_669_port);
   DataPath_RF_BLOCKi_28_Q_reg_28_inst : DFF_X1 port map( D => n4255, CK => CLK
                           , Q => n_2004, QN => 
                           DataPath_RF_bus_reg_dataout_668_port);
   DataPath_RF_BLOCKi_28_Q_reg_27_inst : DFF_X1 port map( D => n4256, CK => CLK
                           , Q => n_2005, QN => 
                           DataPath_RF_bus_reg_dataout_667_port);
   DataPath_RF_BLOCKi_28_Q_reg_26_inst : DFF_X1 port map( D => n4257, CK => CLK
                           , Q => n_2006, QN => 
                           DataPath_RF_bus_reg_dataout_666_port);
   DataPath_RF_BLOCKi_28_Q_reg_25_inst : DFF_X1 port map( D => n4258, CK => CLK
                           , Q => n_2007, QN => 
                           DataPath_RF_bus_reg_dataout_665_port);
   DataPath_RF_BLOCKi_28_Q_reg_24_inst : DFF_X1 port map( D => n4259, CK => CLK
                           , Q => n_2008, QN => 
                           DataPath_RF_bus_reg_dataout_664_port);
   DataPath_RF_BLOCKi_28_Q_reg_23_inst : DFF_X1 port map( D => n4260, CK => CLK
                           , Q => n_2009, QN => 
                           DataPath_RF_bus_reg_dataout_663_port);
   DataPath_RF_BLOCKi_28_Q_reg_22_inst : DFF_X1 port map( D => n4261, CK => CLK
                           , Q => n_2010, QN => 
                           DataPath_RF_bus_reg_dataout_662_port);
   DataPath_RF_BLOCKi_28_Q_reg_21_inst : DFF_X1 port map( D => n4262, CK => CLK
                           , Q => n_2011, QN => 
                           DataPath_RF_bus_reg_dataout_661_port);
   DataPath_RF_BLOCKi_28_Q_reg_20_inst : DFF_X1 port map( D => n4263, CK => CLK
                           , Q => n_2012, QN => 
                           DataPath_RF_bus_reg_dataout_660_port);
   DataPath_RF_BLOCKi_28_Q_reg_19_inst : DFF_X1 port map( D => n4264, CK => CLK
                           , Q => n_2013, QN => 
                           DataPath_RF_bus_reg_dataout_659_port);
   DataPath_RF_BLOCKi_28_Q_reg_18_inst : DFF_X1 port map( D => n4265, CK => CLK
                           , Q => n_2014, QN => 
                           DataPath_RF_bus_reg_dataout_658_port);
   DataPath_RF_BLOCKi_28_Q_reg_17_inst : DFF_X1 port map( D => n4266, CK => CLK
                           , Q => n_2015, QN => 
                           DataPath_RF_bus_reg_dataout_657_port);
   DataPath_RF_BLOCKi_28_Q_reg_16_inst : DFF_X1 port map( D => n4267, CK => CLK
                           , Q => n_2016, QN => 
                           DataPath_RF_bus_reg_dataout_656_port);
   DataPath_RF_BLOCKi_28_Q_reg_15_inst : DFF_X1 port map( D => n4268, CK => CLK
                           , Q => n_2017, QN => 
                           DataPath_RF_bus_reg_dataout_655_port);
   DataPath_RF_BLOCKi_28_Q_reg_14_inst : DFF_X1 port map( D => n4269, CK => CLK
                           , Q => n_2018, QN => 
                           DataPath_RF_bus_reg_dataout_654_port);
   DataPath_RF_BLOCKi_28_Q_reg_13_inst : DFF_X1 port map( D => n4270, CK => CLK
                           , Q => n_2019, QN => 
                           DataPath_RF_bus_reg_dataout_653_port);
   DataPath_RF_BLOCKi_28_Q_reg_12_inst : DFF_X1 port map( D => n4271, CK => CLK
                           , Q => n_2020, QN => 
                           DataPath_RF_bus_reg_dataout_652_port);
   DataPath_RF_BLOCKi_28_Q_reg_11_inst : DFF_X1 port map( D => n4272, CK => CLK
                           , Q => n_2021, QN => 
                           DataPath_RF_bus_reg_dataout_651_port);
   DataPath_RF_BLOCKi_28_Q_reg_9_inst : DFF_X1 port map( D => n4274, CK => CLK,
                           Q => n_2022, QN => 
                           DataPath_RF_bus_reg_dataout_649_port);
   DataPath_RF_BLOCKi_28_Q_reg_8_inst : DFF_X1 port map( D => n4275, CK => CLK,
                           Q => n_2023, QN => 
                           DataPath_RF_bus_reg_dataout_648_port);
   DataPath_RF_BLOCKi_28_Q_reg_7_inst : DFF_X1 port map( D => n4276, CK => CLK,
                           Q => n_2024, QN => 
                           DataPath_RF_bus_reg_dataout_647_port);
   DataPath_RF_BLOCKi_28_Q_reg_6_inst : DFF_X1 port map( D => n4277, CK => CLK,
                           Q => n_2025, QN => 
                           DataPath_RF_bus_reg_dataout_646_port);
   DataPath_RF_BLOCKi_28_Q_reg_5_inst : DFF_X1 port map( D => n4278, CK => CLK,
                           Q => n_2026, QN => 
                           DataPath_RF_bus_reg_dataout_645_port);
   DataPath_RF_BLOCKi_28_Q_reg_4_inst : DFF_X1 port map( D => n4279, CK => CLK,
                           Q => n_2027, QN => 
                           DataPath_RF_bus_reg_dataout_644_port);
   DataPath_RF_BLOCKi_28_Q_reg_3_inst : DFF_X1 port map( D => n4280, CK => CLK,
                           Q => n_2028, QN => 
                           DataPath_RF_bus_reg_dataout_643_port);
   DataPath_RF_BLOCKi_28_Q_reg_2_inst : DFF_X1 port map( D => n4281, CK => CLK,
                           Q => n_2029, QN => 
                           DataPath_RF_bus_reg_dataout_642_port);
   DataPath_RF_BLOCKi_28_Q_reg_1_inst : DFF_X1 port map( D => n4282, CK => CLK,
                           Q => n_2030, QN => 
                           DataPath_RF_bus_reg_dataout_641_port);
   DataPath_RF_BLOCKi_28_Q_reg_0_inst : DFF_X1 port map( D => n4283, CK => CLK,
                           Q => n_2031, QN => 
                           DataPath_RF_bus_reg_dataout_640_port);
   DataPath_RF_BLOCKi_44_Q_reg_31_inst : DFF_X1 port map( D => n4843, CK => CLK
                           , Q => n_2032, QN => 
                           DataPath_RF_bus_reg_dataout_1183_port);
   DataPath_RF_BLOCKi_44_Q_reg_30_inst : DFF_X1 port map( D => n4846, CK => CLK
                           , Q => n_2033, QN => 
                           DataPath_RF_bus_reg_dataout_1182_port);
   DataPath_RF_BLOCKi_44_Q_reg_29_inst : DFF_X1 port map( D => n4847, CK => CLK
                           , Q => n_2034, QN => 
                           DataPath_RF_bus_reg_dataout_1181_port);
   DataPath_RF_BLOCKi_44_Q_reg_28_inst : DFF_X1 port map( D => n4848, CK => CLK
                           , Q => n_2035, QN => 
                           DataPath_RF_bus_reg_dataout_1180_port);
   DataPath_RF_BLOCKi_44_Q_reg_27_inst : DFF_X1 port map( D => n4849, CK => CLK
                           , Q => n_2036, QN => 
                           DataPath_RF_bus_reg_dataout_1179_port);
   DataPath_RF_BLOCKi_44_Q_reg_26_inst : DFF_X1 port map( D => n4850, CK => CLK
                           , Q => n_2037, QN => 
                           DataPath_RF_bus_reg_dataout_1178_port);
   DataPath_RF_BLOCKi_44_Q_reg_25_inst : DFF_X1 port map( D => n4851, CK => CLK
                           , Q => n_2038, QN => 
                           DataPath_RF_bus_reg_dataout_1177_port);
   DataPath_RF_BLOCKi_44_Q_reg_24_inst : DFF_X1 port map( D => n4852, CK => CLK
                           , Q => n_2039, QN => 
                           DataPath_RF_bus_reg_dataout_1176_port);
   DataPath_RF_BLOCKi_44_Q_reg_23_inst : DFF_X1 port map( D => n4853, CK => CLK
                           , Q => n_2040, QN => 
                           DataPath_RF_bus_reg_dataout_1175_port);
   DataPath_RF_BLOCKi_44_Q_reg_22_inst : DFF_X1 port map( D => n4854, CK => CLK
                           , Q => n_2041, QN => 
                           DataPath_RF_bus_reg_dataout_1174_port);
   DataPath_RF_BLOCKi_44_Q_reg_21_inst : DFF_X1 port map( D => n4855, CK => CLK
                           , Q => n_2042, QN => 
                           DataPath_RF_bus_reg_dataout_1173_port);
   DataPath_RF_BLOCKi_44_Q_reg_20_inst : DFF_X1 port map( D => n4856, CK => CLK
                           , Q => n_2043, QN => 
                           DataPath_RF_bus_reg_dataout_1172_port);
   DataPath_RF_BLOCKi_44_Q_reg_19_inst : DFF_X1 port map( D => n4857, CK => CLK
                           , Q => n_2044, QN => 
                           DataPath_RF_bus_reg_dataout_1171_port);
   DataPath_RF_BLOCKi_44_Q_reg_18_inst : DFF_X1 port map( D => n4858, CK => CLK
                           , Q => n_2045, QN => 
                           DataPath_RF_bus_reg_dataout_1170_port);
   DataPath_RF_BLOCKi_44_Q_reg_17_inst : DFF_X1 port map( D => n4859, CK => CLK
                           , Q => n_2046, QN => 
                           DataPath_RF_bus_reg_dataout_1169_port);
   DataPath_RF_BLOCKi_44_Q_reg_16_inst : DFF_X1 port map( D => n4860, CK => CLK
                           , Q => n_2047, QN => 
                           DataPath_RF_bus_reg_dataout_1168_port);
   DataPath_RF_BLOCKi_44_Q_reg_15_inst : DFF_X1 port map( D => n4861, CK => CLK
                           , Q => n_2048, QN => 
                           DataPath_RF_bus_reg_dataout_1167_port);
   DataPath_RF_BLOCKi_44_Q_reg_14_inst : DFF_X1 port map( D => n4862, CK => CLK
                           , Q => n_2049, QN => 
                           DataPath_RF_bus_reg_dataout_1166_port);
   DataPath_RF_BLOCKi_44_Q_reg_13_inst : DFF_X1 port map( D => n4863, CK => CLK
                           , Q => n_2050, QN => 
                           DataPath_RF_bus_reg_dataout_1165_port);
   DataPath_RF_BLOCKi_44_Q_reg_12_inst : DFF_X1 port map( D => n4864, CK => CLK
                           , Q => n_2051, QN => 
                           DataPath_RF_bus_reg_dataout_1164_port);
   DataPath_RF_BLOCKi_44_Q_reg_11_inst : DFF_X1 port map( D => n4865, CK => CLK
                           , Q => n_2052, QN => 
                           DataPath_RF_bus_reg_dataout_1163_port);
   DataPath_RF_BLOCKi_44_Q_reg_9_inst : DFF_X1 port map( D => n4867, CK => CLK,
                           Q => n_2053, QN => 
                           DataPath_RF_bus_reg_dataout_1161_port);
   DataPath_RF_BLOCKi_44_Q_reg_8_inst : DFF_X1 port map( D => n4868, CK => CLK,
                           Q => n_2054, QN => 
                           DataPath_RF_bus_reg_dataout_1160_port);
   DataPath_RF_BLOCKi_44_Q_reg_7_inst : DFF_X1 port map( D => n4869, CK => CLK,
                           Q => n_2055, QN => 
                           DataPath_RF_bus_reg_dataout_1159_port);
   DataPath_RF_BLOCKi_44_Q_reg_6_inst : DFF_X1 port map( D => n4870, CK => CLK,
                           Q => n_2056, QN => 
                           DataPath_RF_bus_reg_dataout_1158_port);
   DataPath_RF_BLOCKi_44_Q_reg_5_inst : DFF_X1 port map( D => n4871, CK => CLK,
                           Q => n_2057, QN => 
                           DataPath_RF_bus_reg_dataout_1157_port);
   DataPath_RF_BLOCKi_44_Q_reg_4_inst : DFF_X1 port map( D => n4872, CK => CLK,
                           Q => n_2058, QN => 
                           DataPath_RF_bus_reg_dataout_1156_port);
   DataPath_RF_BLOCKi_44_Q_reg_3_inst : DFF_X1 port map( D => n4873, CK => CLK,
                           Q => n_2059, QN => 
                           DataPath_RF_bus_reg_dataout_1155_port);
   DataPath_RF_BLOCKi_44_Q_reg_2_inst : DFF_X1 port map( D => n4874, CK => CLK,
                           Q => n_2060, QN => 
                           DataPath_RF_bus_reg_dataout_1154_port);
   DataPath_RF_BLOCKi_44_Q_reg_1_inst : DFF_X1 port map( D => n4875, CK => CLK,
                           Q => n_2061, QN => 
                           DataPath_RF_bus_reg_dataout_1153_port);
   DataPath_RF_BLOCKi_44_Q_reg_0_inst : DFF_X1 port map( D => n4876, CK => CLK,
                           Q => n_2062, QN => 
                           DataPath_RF_bus_reg_dataout_1152_port);
   DataPath_RF_BLOCKi_60_Q_reg_31_inst : DFF_X1 port map( D => n5436, CK => CLK
                           , Q => n_2063, QN => 
                           DataPath_RF_bus_reg_dataout_1695_port);
   DataPath_RF_BLOCKi_60_Q_reg_30_inst : DFF_X1 port map( D => n5439, CK => CLK
                           , Q => n_2064, QN => 
                           DataPath_RF_bus_reg_dataout_1694_port);
   DataPath_RF_BLOCKi_60_Q_reg_29_inst : DFF_X1 port map( D => n5440, CK => CLK
                           , Q => n_2065, QN => 
                           DataPath_RF_bus_reg_dataout_1693_port);
   DataPath_RF_BLOCKi_60_Q_reg_28_inst : DFF_X1 port map( D => n5441, CK => CLK
                           , Q => n_2066, QN => 
                           DataPath_RF_bus_reg_dataout_1692_port);
   DataPath_RF_BLOCKi_60_Q_reg_27_inst : DFF_X1 port map( D => n5442, CK => CLK
                           , Q => n_2067, QN => 
                           DataPath_RF_bus_reg_dataout_1691_port);
   DataPath_RF_BLOCKi_60_Q_reg_26_inst : DFF_X1 port map( D => n5443, CK => CLK
                           , Q => n_2068, QN => 
                           DataPath_RF_bus_reg_dataout_1690_port);
   DataPath_RF_BLOCKi_60_Q_reg_25_inst : DFF_X1 port map( D => n5444, CK => CLK
                           , Q => n_2069, QN => 
                           DataPath_RF_bus_reg_dataout_1689_port);
   DataPath_RF_BLOCKi_60_Q_reg_24_inst : DFF_X1 port map( D => n5445, CK => CLK
                           , Q => n_2070, QN => 
                           DataPath_RF_bus_reg_dataout_1688_port);
   DataPath_RF_BLOCKi_60_Q_reg_23_inst : DFF_X1 port map( D => n5446, CK => CLK
                           , Q => n_2071, QN => 
                           DataPath_RF_bus_reg_dataout_1687_port);
   DataPath_RF_BLOCKi_60_Q_reg_22_inst : DFF_X1 port map( D => n5447, CK => CLK
                           , Q => n_2072, QN => 
                           DataPath_RF_bus_reg_dataout_1686_port);
   DataPath_RF_BLOCKi_60_Q_reg_21_inst : DFF_X1 port map( D => n5448, CK => CLK
                           , Q => n_2073, QN => 
                           DataPath_RF_bus_reg_dataout_1685_port);
   DataPath_RF_BLOCKi_60_Q_reg_20_inst : DFF_X1 port map( D => n5449, CK => CLK
                           , Q => n_2074, QN => 
                           DataPath_RF_bus_reg_dataout_1684_port);
   DataPath_RF_BLOCKi_60_Q_reg_19_inst : DFF_X1 port map( D => n5450, CK => CLK
                           , Q => n_2075, QN => 
                           DataPath_RF_bus_reg_dataout_1683_port);
   DataPath_RF_BLOCKi_60_Q_reg_18_inst : DFF_X1 port map( D => n5451, CK => CLK
                           , Q => n_2076, QN => 
                           DataPath_RF_bus_reg_dataout_1682_port);
   DataPath_RF_BLOCKi_60_Q_reg_17_inst : DFF_X1 port map( D => n5452, CK => CLK
                           , Q => n_2077, QN => 
                           DataPath_RF_bus_reg_dataout_1681_port);
   DataPath_RF_BLOCKi_60_Q_reg_16_inst : DFF_X1 port map( D => n5453, CK => CLK
                           , Q => n_2078, QN => 
                           DataPath_RF_bus_reg_dataout_1680_port);
   DataPath_RF_BLOCKi_60_Q_reg_15_inst : DFF_X1 port map( D => n5454, CK => CLK
                           , Q => n_2079, QN => 
                           DataPath_RF_bus_reg_dataout_1679_port);
   DataPath_RF_BLOCKi_60_Q_reg_14_inst : DFF_X1 port map( D => n5455, CK => CLK
                           , Q => n_2080, QN => 
                           DataPath_RF_bus_reg_dataout_1678_port);
   DataPath_RF_BLOCKi_60_Q_reg_13_inst : DFF_X1 port map( D => n5456, CK => CLK
                           , Q => n_2081, QN => 
                           DataPath_RF_bus_reg_dataout_1677_port);
   DataPath_RF_BLOCKi_60_Q_reg_12_inst : DFF_X1 port map( D => n5457, CK => CLK
                           , Q => n_2082, QN => 
                           DataPath_RF_bus_reg_dataout_1676_port);
   DataPath_RF_BLOCKi_60_Q_reg_11_inst : DFF_X1 port map( D => n5458, CK => CLK
                           , Q => n_2083, QN => 
                           DataPath_RF_bus_reg_dataout_1675_port);
   DataPath_RF_BLOCKi_60_Q_reg_9_inst : DFF_X1 port map( D => n5460, CK => CLK,
                           Q => n_2084, QN => 
                           DataPath_RF_bus_reg_dataout_1673_port);
   DataPath_RF_BLOCKi_60_Q_reg_8_inst : DFF_X1 port map( D => n5461, CK => CLK,
                           Q => n_2085, QN => 
                           DataPath_RF_bus_reg_dataout_1672_port);
   DataPath_RF_BLOCKi_60_Q_reg_7_inst : DFF_X1 port map( D => n5462, CK => CLK,
                           Q => n_2086, QN => 
                           DataPath_RF_bus_reg_dataout_1671_port);
   DataPath_RF_BLOCKi_60_Q_reg_6_inst : DFF_X1 port map( D => n5463, CK => CLK,
                           Q => n_2087, QN => 
                           DataPath_RF_bus_reg_dataout_1670_port);
   DataPath_RF_BLOCKi_60_Q_reg_5_inst : DFF_X1 port map( D => n5464, CK => CLK,
                           Q => n_2088, QN => 
                           DataPath_RF_bus_reg_dataout_1669_port);
   DataPath_RF_BLOCKi_60_Q_reg_4_inst : DFF_X1 port map( D => n5465, CK => CLK,
                           Q => n_2089, QN => 
                           DataPath_RF_bus_reg_dataout_1668_port);
   DataPath_RF_BLOCKi_60_Q_reg_3_inst : DFF_X1 port map( D => n5466, CK => CLK,
                           Q => n_2090, QN => 
                           DataPath_RF_bus_reg_dataout_1667_port);
   DataPath_RF_BLOCKi_60_Q_reg_2_inst : DFF_X1 port map( D => n5467, CK => CLK,
                           Q => n_2091, QN => 
                           DataPath_RF_bus_reg_dataout_1666_port);
   DataPath_RF_BLOCKi_60_Q_reg_1_inst : DFF_X1 port map( D => n5468, CK => CLK,
                           Q => n_2092, QN => 
                           DataPath_RF_bus_reg_dataout_1665_port);
   DataPath_RF_BLOCKi_60_Q_reg_0_inst : DFF_X1 port map( D => n5469, CK => CLK,
                           Q => n_2093, QN => 
                           DataPath_RF_bus_reg_dataout_1664_port);
   DataPath_RF_BLOCKi_76_Q_reg_31_inst : DFF_X1 port map( D => n6016, CK => CLK
                           , Q => n_2094, QN => 
                           DataPath_RF_bus_reg_dataout_2207_port);
   DataPath_RF_BLOCKi_76_Q_reg_30_inst : DFF_X1 port map( D => n6019, CK => CLK
                           , Q => n_2095, QN => 
                           DataPath_RF_bus_reg_dataout_2206_port);
   DataPath_RF_BLOCKi_76_Q_reg_29_inst : DFF_X1 port map( D => n6020, CK => CLK
                           , Q => n_2096, QN => 
                           DataPath_RF_bus_reg_dataout_2205_port);
   DataPath_RF_BLOCKi_76_Q_reg_28_inst : DFF_X1 port map( D => n6021, CK => CLK
                           , Q => n_2097, QN => 
                           DataPath_RF_bus_reg_dataout_2204_port);
   DataPath_RF_BLOCKi_76_Q_reg_27_inst : DFF_X1 port map( D => n6022, CK => CLK
                           , Q => n_2098, QN => 
                           DataPath_RF_bus_reg_dataout_2203_port);
   DataPath_RF_BLOCKi_76_Q_reg_26_inst : DFF_X1 port map( D => n6023, CK => CLK
                           , Q => n_2099, QN => 
                           DataPath_RF_bus_reg_dataout_2202_port);
   DataPath_RF_BLOCKi_76_Q_reg_25_inst : DFF_X1 port map( D => n6024, CK => CLK
                           , Q => n_2100, QN => 
                           DataPath_RF_bus_reg_dataout_2201_port);
   DataPath_RF_BLOCKi_76_Q_reg_24_inst : DFF_X1 port map( D => n6025, CK => CLK
                           , Q => n_2101, QN => 
                           DataPath_RF_bus_reg_dataout_2200_port);
   DataPath_RF_BLOCKi_76_Q_reg_23_inst : DFF_X1 port map( D => n6026, CK => CLK
                           , Q => n_2102, QN => 
                           DataPath_RF_bus_reg_dataout_2199_port);
   DataPath_RF_BLOCKi_76_Q_reg_22_inst : DFF_X1 port map( D => n6027, CK => CLK
                           , Q => n_2103, QN => 
                           DataPath_RF_bus_reg_dataout_2198_port);
   DataPath_RF_BLOCKi_76_Q_reg_21_inst : DFF_X1 port map( D => n6028, CK => CLK
                           , Q => n_2104, QN => 
                           DataPath_RF_bus_reg_dataout_2197_port);
   DataPath_RF_BLOCKi_76_Q_reg_20_inst : DFF_X1 port map( D => n6029, CK => CLK
                           , Q => n_2105, QN => 
                           DataPath_RF_bus_reg_dataout_2196_port);
   DataPath_RF_BLOCKi_76_Q_reg_19_inst : DFF_X1 port map( D => n6030, CK => CLK
                           , Q => n_2106, QN => 
                           DataPath_RF_bus_reg_dataout_2195_port);
   DataPath_RF_BLOCKi_76_Q_reg_18_inst : DFF_X1 port map( D => n6031, CK => CLK
                           , Q => n_2107, QN => 
                           DataPath_RF_bus_reg_dataout_2194_port);
   DataPath_RF_BLOCKi_76_Q_reg_17_inst : DFF_X1 port map( D => n6032, CK => CLK
                           , Q => n_2108, QN => 
                           DataPath_RF_bus_reg_dataout_2193_port);
   DataPath_RF_BLOCKi_76_Q_reg_16_inst : DFF_X1 port map( D => n6033, CK => CLK
                           , Q => n_2109, QN => 
                           DataPath_RF_bus_reg_dataout_2192_port);
   DataPath_RF_BLOCKi_76_Q_reg_15_inst : DFF_X1 port map( D => n6034, CK => CLK
                           , Q => n_2110, QN => 
                           DataPath_RF_bus_reg_dataout_2191_port);
   DataPath_RF_BLOCKi_76_Q_reg_14_inst : DFF_X1 port map( D => n6035, CK => CLK
                           , Q => n_2111, QN => 
                           DataPath_RF_bus_reg_dataout_2190_port);
   DataPath_RF_BLOCKi_76_Q_reg_13_inst : DFF_X1 port map( D => n6036, CK => CLK
                           , Q => n_2112, QN => 
                           DataPath_RF_bus_reg_dataout_2189_port);
   DataPath_RF_BLOCKi_76_Q_reg_12_inst : DFF_X1 port map( D => n6037, CK => CLK
                           , Q => n_2113, QN => 
                           DataPath_RF_bus_reg_dataout_2188_port);
   DataPath_RF_BLOCKi_76_Q_reg_11_inst : DFF_X1 port map( D => n6038, CK => CLK
                           , Q => n_2114, QN => 
                           DataPath_RF_bus_reg_dataout_2187_port);
   DataPath_RF_BLOCKi_76_Q_reg_9_inst : DFF_X1 port map( D => n6040, CK => CLK,
                           Q => n_2115, QN => 
                           DataPath_RF_bus_reg_dataout_2185_port);
   DataPath_RF_BLOCKi_76_Q_reg_8_inst : DFF_X1 port map( D => n6041, CK => CLK,
                           Q => n_2116, QN => 
                           DataPath_RF_bus_reg_dataout_2184_port);
   DataPath_RF_BLOCKi_76_Q_reg_7_inst : DFF_X1 port map( D => n6042, CK => CLK,
                           Q => n_2117, QN => 
                           DataPath_RF_bus_reg_dataout_2183_port);
   DataPath_RF_BLOCKi_76_Q_reg_6_inst : DFF_X1 port map( D => n6043, CK => CLK,
                           Q => n_2118, QN => 
                           DataPath_RF_bus_reg_dataout_2182_port);
   DataPath_RF_BLOCKi_76_Q_reg_5_inst : DFF_X1 port map( D => n6044, CK => CLK,
                           Q => n_2119, QN => 
                           DataPath_RF_bus_reg_dataout_2181_port);
   DataPath_RF_BLOCKi_76_Q_reg_4_inst : DFF_X1 port map( D => n6045, CK => CLK,
                           Q => n_2120, QN => 
                           DataPath_RF_bus_reg_dataout_2180_port);
   DataPath_RF_BLOCKi_76_Q_reg_3_inst : DFF_X1 port map( D => n6046, CK => CLK,
                           Q => n_2121, QN => 
                           DataPath_RF_bus_reg_dataout_2179_port);
   DataPath_RF_BLOCKi_76_Q_reg_2_inst : DFF_X1 port map( D => n6047, CK => CLK,
                           Q => n_2122, QN => 
                           DataPath_RF_bus_reg_dataout_2178_port);
   DataPath_RF_BLOCKi_76_Q_reg_1_inst : DFF_X1 port map( D => n6048, CK => CLK,
                           Q => n_2123, QN => 
                           DataPath_RF_bus_reg_dataout_2177_port);
   DataPath_RF_BLOCKi_76_Q_reg_0_inst : DFF_X1 port map( D => n6049, CK => CLK,
                           Q => n_2124, QN => 
                           DataPath_RF_bus_reg_dataout_2176_port);
   DataPath_RF_BLOCKi_13_Q_reg_31_inst : DFF_X1 port map( D => n3651, CK => CLK
                           , Q => n_2125, QN => 
                           DataPath_RF_bus_reg_dataout_191_port);
   DataPath_RF_BLOCKi_13_Q_reg_30_inst : DFF_X1 port map( D => n3654, CK => CLK
                           , Q => n_2126, QN => 
                           DataPath_RF_bus_reg_dataout_190_port);
   DataPath_RF_BLOCKi_13_Q_reg_29_inst : DFF_X1 port map( D => n3655, CK => CLK
                           , Q => n_2127, QN => 
                           DataPath_RF_bus_reg_dataout_189_port);
   DataPath_RF_BLOCKi_13_Q_reg_28_inst : DFF_X1 port map( D => n3656, CK => CLK
                           , Q => n_2128, QN => 
                           DataPath_RF_bus_reg_dataout_188_port);
   DataPath_RF_BLOCKi_13_Q_reg_27_inst : DFF_X1 port map( D => n3657, CK => CLK
                           , Q => n_2129, QN => 
                           DataPath_RF_bus_reg_dataout_187_port);
   DataPath_RF_BLOCKi_13_Q_reg_26_inst : DFF_X1 port map( D => n3658, CK => CLK
                           , Q => n_2130, QN => 
                           DataPath_RF_bus_reg_dataout_186_port);
   DataPath_RF_BLOCKi_13_Q_reg_25_inst : DFF_X1 port map( D => n3659, CK => CLK
                           , Q => n_2131, QN => 
                           DataPath_RF_bus_reg_dataout_185_port);
   DataPath_RF_BLOCKi_13_Q_reg_24_inst : DFF_X1 port map( D => n3660, CK => CLK
                           , Q => n_2132, QN => 
                           DataPath_RF_bus_reg_dataout_184_port);
   DataPath_RF_BLOCKi_13_Q_reg_23_inst : DFF_X1 port map( D => n3661, CK => CLK
                           , Q => n_2133, QN => 
                           DataPath_RF_bus_reg_dataout_183_port);
   DataPath_RF_BLOCKi_13_Q_reg_22_inst : DFF_X1 port map( D => n3662, CK => CLK
                           , Q => n_2134, QN => 
                           DataPath_RF_bus_reg_dataout_182_port);
   DataPath_RF_BLOCKi_13_Q_reg_21_inst : DFF_X1 port map( D => n3663, CK => CLK
                           , Q => n_2135, QN => 
                           DataPath_RF_bus_reg_dataout_181_port);
   DataPath_RF_BLOCKi_13_Q_reg_20_inst : DFF_X1 port map( D => n3664, CK => CLK
                           , Q => n_2136, QN => 
                           DataPath_RF_bus_reg_dataout_180_port);
   DataPath_RF_BLOCKi_13_Q_reg_19_inst : DFF_X1 port map( D => n3665, CK => CLK
                           , Q => n_2137, QN => 
                           DataPath_RF_bus_reg_dataout_179_port);
   DataPath_RF_BLOCKi_13_Q_reg_18_inst : DFF_X1 port map( D => n3666, CK => CLK
                           , Q => n_2138, QN => 
                           DataPath_RF_bus_reg_dataout_178_port);
   DataPath_RF_BLOCKi_13_Q_reg_17_inst : DFF_X1 port map( D => n3667, CK => CLK
                           , Q => n_2139, QN => 
                           DataPath_RF_bus_reg_dataout_177_port);
   DataPath_RF_BLOCKi_13_Q_reg_16_inst : DFF_X1 port map( D => n3668, CK => CLK
                           , Q => n_2140, QN => 
                           DataPath_RF_bus_reg_dataout_176_port);
   DataPath_RF_BLOCKi_13_Q_reg_15_inst : DFF_X1 port map( D => n3669, CK => CLK
                           , Q => n_2141, QN => 
                           DataPath_RF_bus_reg_dataout_175_port);
   DataPath_RF_BLOCKi_13_Q_reg_14_inst : DFF_X1 port map( D => n3670, CK => CLK
                           , Q => n_2142, QN => 
                           DataPath_RF_bus_reg_dataout_174_port);
   DataPath_RF_BLOCKi_13_Q_reg_13_inst : DFF_X1 port map( D => n3671, CK => CLK
                           , Q => n_2143, QN => 
                           DataPath_RF_bus_reg_dataout_173_port);
   DataPath_RF_BLOCKi_13_Q_reg_12_inst : DFF_X1 port map( D => n3672, CK => CLK
                           , Q => n_2144, QN => 
                           DataPath_RF_bus_reg_dataout_172_port);
   DataPath_RF_BLOCKi_13_Q_reg_11_inst : DFF_X1 port map( D => n3673, CK => CLK
                           , Q => n_2145, QN => 
                           DataPath_RF_bus_reg_dataout_171_port);
   DataPath_RF_BLOCKi_13_Q_reg_9_inst : DFF_X1 port map( D => n3675, CK => CLK,
                           Q => n_2146, QN => 
                           DataPath_RF_bus_reg_dataout_169_port);
   DataPath_RF_BLOCKi_13_Q_reg_8_inst : DFF_X1 port map( D => n3676, CK => CLK,
                           Q => n_2147, QN => 
                           DataPath_RF_bus_reg_dataout_168_port);
   DataPath_RF_BLOCKi_13_Q_reg_7_inst : DFF_X1 port map( D => n3677, CK => CLK,
                           Q => n_2148, QN => 
                           DataPath_RF_bus_reg_dataout_167_port);
   DataPath_RF_BLOCKi_13_Q_reg_6_inst : DFF_X1 port map( D => n3678, CK => CLK,
                           Q => n_2149, QN => 
                           DataPath_RF_bus_reg_dataout_166_port);
   DataPath_RF_BLOCKi_13_Q_reg_5_inst : DFF_X1 port map( D => n3679, CK => CLK,
                           Q => n_2150, QN => 
                           DataPath_RF_bus_reg_dataout_165_port);
   DataPath_RF_BLOCKi_13_Q_reg_4_inst : DFF_X1 port map( D => n3680, CK => CLK,
                           Q => n_2151, QN => 
                           DataPath_RF_bus_reg_dataout_164_port);
   DataPath_RF_BLOCKi_13_Q_reg_3_inst : DFF_X1 port map( D => n3681, CK => CLK,
                           Q => n_2152, QN => 
                           DataPath_RF_bus_reg_dataout_163_port);
   DataPath_RF_BLOCKi_13_Q_reg_2_inst : DFF_X1 port map( D => n3682, CK => CLK,
                           Q => n_2153, QN => 
                           DataPath_RF_bus_reg_dataout_162_port);
   DataPath_RF_BLOCKi_13_Q_reg_1_inst : DFF_X1 port map( D => n3683, CK => CLK,
                           Q => n_2154, QN => 
                           DataPath_RF_bus_reg_dataout_161_port);
   DataPath_RF_BLOCKi_13_Q_reg_0_inst : DFF_X1 port map( D => n3684, CK => CLK,
                           Q => n_2155, QN => 
                           DataPath_RF_bus_reg_dataout_160_port);
   DataPath_RF_BLOCKi_29_Q_reg_31_inst : DFF_X1 port map( D => n4285, CK => CLK
                           , Q => n_2156, QN => 
                           DataPath_RF_bus_reg_dataout_703_port);
   DataPath_RF_BLOCKi_29_Q_reg_30_inst : DFF_X1 port map( D => n4288, CK => CLK
                           , Q => n_2157, QN => 
                           DataPath_RF_bus_reg_dataout_702_port);
   DataPath_RF_BLOCKi_29_Q_reg_29_inst : DFF_X1 port map( D => n4289, CK => CLK
                           , Q => n_2158, QN => 
                           DataPath_RF_bus_reg_dataout_701_port);
   DataPath_RF_BLOCKi_29_Q_reg_28_inst : DFF_X1 port map( D => n4290, CK => CLK
                           , Q => n_2159, QN => 
                           DataPath_RF_bus_reg_dataout_700_port);
   DataPath_RF_BLOCKi_29_Q_reg_27_inst : DFF_X1 port map( D => n4291, CK => CLK
                           , Q => n_2160, QN => 
                           DataPath_RF_bus_reg_dataout_699_port);
   DataPath_RF_BLOCKi_29_Q_reg_26_inst : DFF_X1 port map( D => n4292, CK => CLK
                           , Q => n_2161, QN => 
                           DataPath_RF_bus_reg_dataout_698_port);
   DataPath_RF_BLOCKi_29_Q_reg_25_inst : DFF_X1 port map( D => n4293, CK => CLK
                           , Q => n_2162, QN => 
                           DataPath_RF_bus_reg_dataout_697_port);
   DataPath_RF_BLOCKi_29_Q_reg_24_inst : DFF_X1 port map( D => n4294, CK => CLK
                           , Q => n_2163, QN => 
                           DataPath_RF_bus_reg_dataout_696_port);
   DataPath_RF_BLOCKi_29_Q_reg_23_inst : DFF_X1 port map( D => n4295, CK => CLK
                           , Q => n_2164, QN => 
                           DataPath_RF_bus_reg_dataout_695_port);
   DataPath_RF_BLOCKi_29_Q_reg_22_inst : DFF_X1 port map( D => n4296, CK => CLK
                           , Q => n_2165, QN => 
                           DataPath_RF_bus_reg_dataout_694_port);
   DataPath_RF_BLOCKi_29_Q_reg_21_inst : DFF_X1 port map( D => n4297, CK => CLK
                           , Q => n_2166, QN => 
                           DataPath_RF_bus_reg_dataout_693_port);
   DataPath_RF_BLOCKi_29_Q_reg_20_inst : DFF_X1 port map( D => n4298, CK => CLK
                           , Q => n_2167, QN => 
                           DataPath_RF_bus_reg_dataout_692_port);
   DataPath_RF_BLOCKi_29_Q_reg_19_inst : DFF_X1 port map( D => n4299, CK => CLK
                           , Q => n_2168, QN => 
                           DataPath_RF_bus_reg_dataout_691_port);
   DataPath_RF_BLOCKi_29_Q_reg_18_inst : DFF_X1 port map( D => n4300, CK => CLK
                           , Q => n_2169, QN => 
                           DataPath_RF_bus_reg_dataout_690_port);
   DataPath_RF_BLOCKi_29_Q_reg_17_inst : DFF_X1 port map( D => n4301, CK => CLK
                           , Q => n_2170, QN => 
                           DataPath_RF_bus_reg_dataout_689_port);
   DataPath_RF_BLOCKi_29_Q_reg_16_inst : DFF_X1 port map( D => n4302, CK => CLK
                           , Q => n_2171, QN => 
                           DataPath_RF_bus_reg_dataout_688_port);
   DataPath_RF_BLOCKi_29_Q_reg_15_inst : DFF_X1 port map( D => n4303, CK => CLK
                           , Q => n_2172, QN => 
                           DataPath_RF_bus_reg_dataout_687_port);
   DataPath_RF_BLOCKi_29_Q_reg_14_inst : DFF_X1 port map( D => n4304, CK => CLK
                           , Q => n_2173, QN => 
                           DataPath_RF_bus_reg_dataout_686_port);
   DataPath_RF_BLOCKi_29_Q_reg_13_inst : DFF_X1 port map( D => n4305, CK => CLK
                           , Q => n_2174, QN => 
                           DataPath_RF_bus_reg_dataout_685_port);
   DataPath_RF_BLOCKi_29_Q_reg_12_inst : DFF_X1 port map( D => n4306, CK => CLK
                           , Q => n_2175, QN => 
                           DataPath_RF_bus_reg_dataout_684_port);
   DataPath_RF_BLOCKi_29_Q_reg_11_inst : DFF_X1 port map( D => n4307, CK => CLK
                           , Q => n_2176, QN => 
                           DataPath_RF_bus_reg_dataout_683_port);
   DataPath_RF_BLOCKi_29_Q_reg_9_inst : DFF_X1 port map( D => n4309, CK => CLK,
                           Q => n_2177, QN => 
                           DataPath_RF_bus_reg_dataout_681_port);
   DataPath_RF_BLOCKi_29_Q_reg_8_inst : DFF_X1 port map( D => n4310, CK => CLK,
                           Q => n_2178, QN => 
                           DataPath_RF_bus_reg_dataout_680_port);
   DataPath_RF_BLOCKi_29_Q_reg_7_inst : DFF_X1 port map( D => n4311, CK => CLK,
                           Q => n_2179, QN => 
                           DataPath_RF_bus_reg_dataout_679_port);
   DataPath_RF_BLOCKi_29_Q_reg_6_inst : DFF_X1 port map( D => n4312, CK => CLK,
                           Q => n_2180, QN => 
                           DataPath_RF_bus_reg_dataout_678_port);
   DataPath_RF_BLOCKi_29_Q_reg_5_inst : DFF_X1 port map( D => n4313, CK => CLK,
                           Q => n_2181, QN => 
                           DataPath_RF_bus_reg_dataout_677_port);
   DataPath_RF_BLOCKi_29_Q_reg_4_inst : DFF_X1 port map( D => n4314, CK => CLK,
                           Q => n_2182, QN => 
                           DataPath_RF_bus_reg_dataout_676_port);
   DataPath_RF_BLOCKi_29_Q_reg_3_inst : DFF_X1 port map( D => n4315, CK => CLK,
                           Q => n_2183, QN => 
                           DataPath_RF_bus_reg_dataout_675_port);
   DataPath_RF_BLOCKi_29_Q_reg_2_inst : DFF_X1 port map( D => n4316, CK => CLK,
                           Q => n_2184, QN => 
                           DataPath_RF_bus_reg_dataout_674_port);
   DataPath_RF_BLOCKi_29_Q_reg_1_inst : DFF_X1 port map( D => n4317, CK => CLK,
                           Q => n_2185, QN => 
                           DataPath_RF_bus_reg_dataout_673_port);
   DataPath_RF_BLOCKi_29_Q_reg_0_inst : DFF_X1 port map( D => n4318, CK => CLK,
                           Q => n_2186, QN => 
                           DataPath_RF_bus_reg_dataout_672_port);
   DataPath_RF_BLOCKi_45_Q_reg_31_inst : DFF_X1 port map( D => n4878, CK => CLK
                           , Q => n_2187, QN => 
                           DataPath_RF_bus_reg_dataout_1215_port);
   DataPath_RF_BLOCKi_45_Q_reg_30_inst : DFF_X1 port map( D => n4881, CK => CLK
                           , Q => n_2188, QN => 
                           DataPath_RF_bus_reg_dataout_1214_port);
   DataPath_RF_BLOCKi_45_Q_reg_29_inst : DFF_X1 port map( D => n4882, CK => CLK
                           , Q => n_2189, QN => 
                           DataPath_RF_bus_reg_dataout_1213_port);
   DataPath_RF_BLOCKi_45_Q_reg_28_inst : DFF_X1 port map( D => n4883, CK => CLK
                           , Q => n_2190, QN => 
                           DataPath_RF_bus_reg_dataout_1212_port);
   DataPath_RF_BLOCKi_45_Q_reg_27_inst : DFF_X1 port map( D => n4884, CK => CLK
                           , Q => n_2191, QN => 
                           DataPath_RF_bus_reg_dataout_1211_port);
   DataPath_RF_BLOCKi_45_Q_reg_26_inst : DFF_X1 port map( D => n4885, CK => CLK
                           , Q => n_2192, QN => 
                           DataPath_RF_bus_reg_dataout_1210_port);
   DataPath_RF_BLOCKi_45_Q_reg_25_inst : DFF_X1 port map( D => n4886, CK => CLK
                           , Q => n_2193, QN => 
                           DataPath_RF_bus_reg_dataout_1209_port);
   DataPath_RF_BLOCKi_45_Q_reg_24_inst : DFF_X1 port map( D => n4887, CK => CLK
                           , Q => n_2194, QN => 
                           DataPath_RF_bus_reg_dataout_1208_port);
   DataPath_RF_BLOCKi_45_Q_reg_23_inst : DFF_X1 port map( D => n4888, CK => CLK
                           , Q => n_2195, QN => 
                           DataPath_RF_bus_reg_dataout_1207_port);
   DataPath_RF_BLOCKi_45_Q_reg_22_inst : DFF_X1 port map( D => n4889, CK => CLK
                           , Q => n_2196, QN => 
                           DataPath_RF_bus_reg_dataout_1206_port);
   DataPath_RF_BLOCKi_45_Q_reg_21_inst : DFF_X1 port map( D => n4890, CK => CLK
                           , Q => n_2197, QN => 
                           DataPath_RF_bus_reg_dataout_1205_port);
   DataPath_RF_BLOCKi_45_Q_reg_20_inst : DFF_X1 port map( D => n4891, CK => CLK
                           , Q => n_2198, QN => 
                           DataPath_RF_bus_reg_dataout_1204_port);
   DataPath_RF_BLOCKi_45_Q_reg_19_inst : DFF_X1 port map( D => n4892, CK => CLK
                           , Q => n_2199, QN => 
                           DataPath_RF_bus_reg_dataout_1203_port);
   DataPath_RF_BLOCKi_45_Q_reg_18_inst : DFF_X1 port map( D => n4893, CK => CLK
                           , Q => n_2200, QN => 
                           DataPath_RF_bus_reg_dataout_1202_port);
   DataPath_RF_BLOCKi_45_Q_reg_17_inst : DFF_X1 port map( D => n4894, CK => CLK
                           , Q => n_2201, QN => 
                           DataPath_RF_bus_reg_dataout_1201_port);
   DataPath_RF_BLOCKi_45_Q_reg_16_inst : DFF_X1 port map( D => n4895, CK => CLK
                           , Q => n_2202, QN => 
                           DataPath_RF_bus_reg_dataout_1200_port);
   DataPath_RF_BLOCKi_45_Q_reg_15_inst : DFF_X1 port map( D => n4896, CK => CLK
                           , Q => n_2203, QN => 
                           DataPath_RF_bus_reg_dataout_1199_port);
   DataPath_RF_BLOCKi_45_Q_reg_14_inst : DFF_X1 port map( D => n4897, CK => CLK
                           , Q => n_2204, QN => 
                           DataPath_RF_bus_reg_dataout_1198_port);
   DataPath_RF_BLOCKi_45_Q_reg_13_inst : DFF_X1 port map( D => n4898, CK => CLK
                           , Q => n_2205, QN => 
                           DataPath_RF_bus_reg_dataout_1197_port);
   DataPath_RF_BLOCKi_45_Q_reg_12_inst : DFF_X1 port map( D => n4899, CK => CLK
                           , Q => n_2206, QN => 
                           DataPath_RF_bus_reg_dataout_1196_port);
   DataPath_RF_BLOCKi_45_Q_reg_11_inst : DFF_X1 port map( D => n4900, CK => CLK
                           , Q => n_2207, QN => 
                           DataPath_RF_bus_reg_dataout_1195_port);
   DataPath_RF_BLOCKi_45_Q_reg_9_inst : DFF_X1 port map( D => n4902, CK => CLK,
                           Q => n_2208, QN => 
                           DataPath_RF_bus_reg_dataout_1193_port);
   DataPath_RF_BLOCKi_45_Q_reg_8_inst : DFF_X1 port map( D => n4903, CK => CLK,
                           Q => n_2209, QN => 
                           DataPath_RF_bus_reg_dataout_1192_port);
   DataPath_RF_BLOCKi_45_Q_reg_7_inst : DFF_X1 port map( D => n4904, CK => CLK,
                           Q => n_2210, QN => 
                           DataPath_RF_bus_reg_dataout_1191_port);
   DataPath_RF_BLOCKi_45_Q_reg_6_inst : DFF_X1 port map( D => n4905, CK => CLK,
                           Q => n_2211, QN => 
                           DataPath_RF_bus_reg_dataout_1190_port);
   DataPath_RF_BLOCKi_45_Q_reg_5_inst : DFF_X1 port map( D => n4906, CK => CLK,
                           Q => n_2212, QN => 
                           DataPath_RF_bus_reg_dataout_1189_port);
   DataPath_RF_BLOCKi_45_Q_reg_4_inst : DFF_X1 port map( D => n4907, CK => CLK,
                           Q => n_2213, QN => 
                           DataPath_RF_bus_reg_dataout_1188_port);
   DataPath_RF_BLOCKi_45_Q_reg_3_inst : DFF_X1 port map( D => n4908, CK => CLK,
                           Q => n_2214, QN => 
                           DataPath_RF_bus_reg_dataout_1187_port);
   DataPath_RF_BLOCKi_45_Q_reg_2_inst : DFF_X1 port map( D => n4909, CK => CLK,
                           Q => n_2215, QN => 
                           DataPath_RF_bus_reg_dataout_1186_port);
   DataPath_RF_BLOCKi_45_Q_reg_1_inst : DFF_X1 port map( D => n4910, CK => CLK,
                           Q => n_2216, QN => 
                           DataPath_RF_bus_reg_dataout_1185_port);
   DataPath_RF_BLOCKi_45_Q_reg_0_inst : DFF_X1 port map( D => n4911, CK => CLK,
                           Q => n_2217, QN => 
                           DataPath_RF_bus_reg_dataout_1184_port);
   DataPath_RF_BLOCKi_61_Q_reg_31_inst : DFF_X1 port map( D => n5471, CK => CLK
                           , Q => n_2218, QN => 
                           DataPath_RF_bus_reg_dataout_1727_port);
   DataPath_RF_BLOCKi_61_Q_reg_30_inst : DFF_X1 port map( D => n5474, CK => CLK
                           , Q => n_2219, QN => 
                           DataPath_RF_bus_reg_dataout_1726_port);
   DataPath_RF_BLOCKi_61_Q_reg_29_inst : DFF_X1 port map( D => n5475, CK => CLK
                           , Q => n_2220, QN => 
                           DataPath_RF_bus_reg_dataout_1725_port);
   DataPath_RF_BLOCKi_61_Q_reg_28_inst : DFF_X1 port map( D => n5476, CK => CLK
                           , Q => n_2221, QN => 
                           DataPath_RF_bus_reg_dataout_1724_port);
   DataPath_RF_BLOCKi_61_Q_reg_27_inst : DFF_X1 port map( D => n5477, CK => CLK
                           , Q => n_2222, QN => 
                           DataPath_RF_bus_reg_dataout_1723_port);
   DataPath_RF_BLOCKi_61_Q_reg_26_inst : DFF_X1 port map( D => n5478, CK => CLK
                           , Q => n_2223, QN => 
                           DataPath_RF_bus_reg_dataout_1722_port);
   DataPath_RF_BLOCKi_61_Q_reg_25_inst : DFF_X1 port map( D => n5479, CK => CLK
                           , Q => n_2224, QN => 
                           DataPath_RF_bus_reg_dataout_1721_port);
   DataPath_RF_BLOCKi_61_Q_reg_24_inst : DFF_X1 port map( D => n5480, CK => CLK
                           , Q => n_2225, QN => 
                           DataPath_RF_bus_reg_dataout_1720_port);
   DataPath_RF_BLOCKi_61_Q_reg_23_inst : DFF_X1 port map( D => n5481, CK => CLK
                           , Q => n_2226, QN => 
                           DataPath_RF_bus_reg_dataout_1719_port);
   DataPath_RF_BLOCKi_61_Q_reg_22_inst : DFF_X1 port map( D => n5482, CK => CLK
                           , Q => n_2227, QN => 
                           DataPath_RF_bus_reg_dataout_1718_port);
   DataPath_RF_BLOCKi_61_Q_reg_21_inst : DFF_X1 port map( D => n5483, CK => CLK
                           , Q => n_2228, QN => 
                           DataPath_RF_bus_reg_dataout_1717_port);
   DataPath_RF_BLOCKi_61_Q_reg_20_inst : DFF_X1 port map( D => n5484, CK => CLK
                           , Q => n_2229, QN => 
                           DataPath_RF_bus_reg_dataout_1716_port);
   DataPath_RF_BLOCKi_61_Q_reg_19_inst : DFF_X1 port map( D => n5485, CK => CLK
                           , Q => n_2230, QN => 
                           DataPath_RF_bus_reg_dataout_1715_port);
   DataPath_RF_BLOCKi_61_Q_reg_18_inst : DFF_X1 port map( D => n5486, CK => CLK
                           , Q => n_2231, QN => 
                           DataPath_RF_bus_reg_dataout_1714_port);
   DataPath_RF_BLOCKi_61_Q_reg_17_inst : DFF_X1 port map( D => n5487, CK => CLK
                           , Q => n_2232, QN => 
                           DataPath_RF_bus_reg_dataout_1713_port);
   DataPath_RF_BLOCKi_61_Q_reg_16_inst : DFF_X1 port map( D => n5488, CK => CLK
                           , Q => n_2233, QN => 
                           DataPath_RF_bus_reg_dataout_1712_port);
   DataPath_RF_BLOCKi_61_Q_reg_15_inst : DFF_X1 port map( D => n5489, CK => CLK
                           , Q => n_2234, QN => 
                           DataPath_RF_bus_reg_dataout_1711_port);
   DataPath_RF_BLOCKi_61_Q_reg_14_inst : DFF_X1 port map( D => n5490, CK => CLK
                           , Q => n_2235, QN => 
                           DataPath_RF_bus_reg_dataout_1710_port);
   DataPath_RF_BLOCKi_61_Q_reg_13_inst : DFF_X1 port map( D => n5491, CK => CLK
                           , Q => n_2236, QN => 
                           DataPath_RF_bus_reg_dataout_1709_port);
   DataPath_RF_BLOCKi_61_Q_reg_12_inst : DFF_X1 port map( D => n5492, CK => CLK
                           , Q => n_2237, QN => 
                           DataPath_RF_bus_reg_dataout_1708_port);
   DataPath_RF_BLOCKi_61_Q_reg_11_inst : DFF_X1 port map( D => n5493, CK => CLK
                           , Q => n_2238, QN => 
                           DataPath_RF_bus_reg_dataout_1707_port);
   DataPath_RF_BLOCKi_61_Q_reg_9_inst : DFF_X1 port map( D => n5495, CK => CLK,
                           Q => n_2239, QN => 
                           DataPath_RF_bus_reg_dataout_1705_port);
   DataPath_RF_BLOCKi_61_Q_reg_8_inst : DFF_X1 port map( D => n5496, CK => CLK,
                           Q => n_2240, QN => 
                           DataPath_RF_bus_reg_dataout_1704_port);
   DataPath_RF_BLOCKi_61_Q_reg_7_inst : DFF_X1 port map( D => n5497, CK => CLK,
                           Q => n_2241, QN => 
                           DataPath_RF_bus_reg_dataout_1703_port);
   DataPath_RF_BLOCKi_61_Q_reg_6_inst : DFF_X1 port map( D => n5498, CK => CLK,
                           Q => n_2242, QN => 
                           DataPath_RF_bus_reg_dataout_1702_port);
   DataPath_RF_BLOCKi_61_Q_reg_5_inst : DFF_X1 port map( D => n5499, CK => CLK,
                           Q => n_2243, QN => 
                           DataPath_RF_bus_reg_dataout_1701_port);
   DataPath_RF_BLOCKi_61_Q_reg_4_inst : DFF_X1 port map( D => n5500, CK => CLK,
                           Q => n_2244, QN => 
                           DataPath_RF_bus_reg_dataout_1700_port);
   DataPath_RF_BLOCKi_61_Q_reg_3_inst : DFF_X1 port map( D => n5501, CK => CLK,
                           Q => n_2245, QN => 
                           DataPath_RF_bus_reg_dataout_1699_port);
   DataPath_RF_BLOCKi_61_Q_reg_2_inst : DFF_X1 port map( D => n5502, CK => CLK,
                           Q => n_2246, QN => 
                           DataPath_RF_bus_reg_dataout_1698_port);
   DataPath_RF_BLOCKi_61_Q_reg_1_inst : DFF_X1 port map( D => n5503, CK => CLK,
                           Q => n_2247, QN => 
                           DataPath_RF_bus_reg_dataout_1697_port);
   DataPath_RF_BLOCKi_61_Q_reg_0_inst : DFF_X1 port map( D => n5504, CK => CLK,
                           Q => n_2248, QN => 
                           DataPath_RF_bus_reg_dataout_1696_port);
   DataPath_RF_BLOCKi_77_Q_reg_31_inst : DFF_X1 port map( D => n6053, CK => CLK
                           , Q => n_2249, QN => 
                           DataPath_RF_bus_reg_dataout_2239_port);
   DataPath_RF_BLOCKi_77_Q_reg_30_inst : DFF_X1 port map( D => n6056, CK => CLK
                           , Q => n_2250, QN => 
                           DataPath_RF_bus_reg_dataout_2238_port);
   DataPath_RF_BLOCKi_77_Q_reg_29_inst : DFF_X1 port map( D => n6057, CK => CLK
                           , Q => n_2251, QN => 
                           DataPath_RF_bus_reg_dataout_2237_port);
   DataPath_RF_BLOCKi_77_Q_reg_28_inst : DFF_X1 port map( D => n6058, CK => CLK
                           , Q => n_2252, QN => 
                           DataPath_RF_bus_reg_dataout_2236_port);
   DataPath_RF_BLOCKi_77_Q_reg_27_inst : DFF_X1 port map( D => n6059, CK => CLK
                           , Q => n_2253, QN => 
                           DataPath_RF_bus_reg_dataout_2235_port);
   DataPath_RF_BLOCKi_77_Q_reg_26_inst : DFF_X1 port map( D => n6060, CK => CLK
                           , Q => n_2254, QN => 
                           DataPath_RF_bus_reg_dataout_2234_port);
   DataPath_RF_BLOCKi_77_Q_reg_25_inst : DFF_X1 port map( D => n6061, CK => CLK
                           , Q => n_2255, QN => 
                           DataPath_RF_bus_reg_dataout_2233_port);
   DataPath_RF_BLOCKi_77_Q_reg_24_inst : DFF_X1 port map( D => n6062, CK => CLK
                           , Q => n_2256, QN => 
                           DataPath_RF_bus_reg_dataout_2232_port);
   DataPath_RF_BLOCKi_77_Q_reg_23_inst : DFF_X1 port map( D => n6063, CK => CLK
                           , Q => n_2257, QN => 
                           DataPath_RF_bus_reg_dataout_2231_port);
   DataPath_RF_BLOCKi_77_Q_reg_22_inst : DFF_X1 port map( D => n6064, CK => CLK
                           , Q => n_2258, QN => 
                           DataPath_RF_bus_reg_dataout_2230_port);
   DataPath_RF_BLOCKi_77_Q_reg_21_inst : DFF_X1 port map( D => n6065, CK => CLK
                           , Q => n_2259, QN => 
                           DataPath_RF_bus_reg_dataout_2229_port);
   DataPath_RF_BLOCKi_77_Q_reg_20_inst : DFF_X1 port map( D => n6066, CK => CLK
                           , Q => n_2260, QN => 
                           DataPath_RF_bus_reg_dataout_2228_port);
   DataPath_RF_BLOCKi_77_Q_reg_19_inst : DFF_X1 port map( D => n6067, CK => CLK
                           , Q => n_2261, QN => 
                           DataPath_RF_bus_reg_dataout_2227_port);
   DataPath_RF_BLOCKi_77_Q_reg_18_inst : DFF_X1 port map( D => n6068, CK => CLK
                           , Q => n_2262, QN => 
                           DataPath_RF_bus_reg_dataout_2226_port);
   DataPath_RF_BLOCKi_77_Q_reg_17_inst : DFF_X1 port map( D => n6069, CK => CLK
                           , Q => n_2263, QN => 
                           DataPath_RF_bus_reg_dataout_2225_port);
   DataPath_RF_BLOCKi_77_Q_reg_16_inst : DFF_X1 port map( D => n6070, CK => CLK
                           , Q => n_2264, QN => 
                           DataPath_RF_bus_reg_dataout_2224_port);
   DataPath_RF_BLOCKi_77_Q_reg_15_inst : DFF_X1 port map( D => n6071, CK => CLK
                           , Q => n_2265, QN => 
                           DataPath_RF_bus_reg_dataout_2223_port);
   DataPath_RF_BLOCKi_77_Q_reg_14_inst : DFF_X1 port map( D => n6072, CK => CLK
                           , Q => n_2266, QN => 
                           DataPath_RF_bus_reg_dataout_2222_port);
   DataPath_RF_BLOCKi_77_Q_reg_13_inst : DFF_X1 port map( D => n6073, CK => CLK
                           , Q => n_2267, QN => 
                           DataPath_RF_bus_reg_dataout_2221_port);
   DataPath_RF_BLOCKi_77_Q_reg_12_inst : DFF_X1 port map( D => n6074, CK => CLK
                           , Q => n_2268, QN => 
                           DataPath_RF_bus_reg_dataout_2220_port);
   DataPath_RF_BLOCKi_77_Q_reg_11_inst : DFF_X1 port map( D => n6075, CK => CLK
                           , Q => n_2269, QN => 
                           DataPath_RF_bus_reg_dataout_2219_port);
   DataPath_RF_BLOCKi_77_Q_reg_9_inst : DFF_X1 port map( D => n6077, CK => CLK,
                           Q => n_2270, QN => 
                           DataPath_RF_bus_reg_dataout_2217_port);
   DataPath_RF_BLOCKi_77_Q_reg_8_inst : DFF_X1 port map( D => n6078, CK => CLK,
                           Q => n_2271, QN => 
                           DataPath_RF_bus_reg_dataout_2216_port);
   DataPath_RF_BLOCKi_77_Q_reg_7_inst : DFF_X1 port map( D => n6079, CK => CLK,
                           Q => n_2272, QN => 
                           DataPath_RF_bus_reg_dataout_2215_port);
   DataPath_RF_BLOCKi_77_Q_reg_6_inst : DFF_X1 port map( D => n6080, CK => CLK,
                           Q => n_2273, QN => 
                           DataPath_RF_bus_reg_dataout_2214_port);
   DataPath_RF_BLOCKi_77_Q_reg_5_inst : DFF_X1 port map( D => n6081, CK => CLK,
                           Q => n_2274, QN => 
                           DataPath_RF_bus_reg_dataout_2213_port);
   DataPath_RF_BLOCKi_77_Q_reg_4_inst : DFF_X1 port map( D => n6082, CK => CLK,
                           Q => n_2275, QN => 
                           DataPath_RF_bus_reg_dataout_2212_port);
   DataPath_RF_BLOCKi_77_Q_reg_3_inst : DFF_X1 port map( D => n6083, CK => CLK,
                           Q => n_2276, QN => 
                           DataPath_RF_bus_reg_dataout_2211_port);
   DataPath_RF_BLOCKi_77_Q_reg_2_inst : DFF_X1 port map( D => n6084, CK => CLK,
                           Q => n_2277, QN => 
                           DataPath_RF_bus_reg_dataout_2210_port);
   DataPath_RF_BLOCKi_77_Q_reg_1_inst : DFF_X1 port map( D => n6085, CK => CLK,
                           Q => n_2278, QN => 
                           DataPath_RF_bus_reg_dataout_2209_port);
   DataPath_RF_BLOCKi_77_Q_reg_0_inst : DFF_X1 port map( D => n6086, CK => CLK,
                           Q => n_2279, QN => 
                           DataPath_RF_bus_reg_dataout_2208_port);
   DataPath_RF_BLOCKi_14_Q_reg_31_inst : DFF_X1 port map( D => n3689, CK => CLK
                           , Q => n_2280, QN => 
                           DataPath_RF_bus_reg_dataout_223_port);
   DataPath_RF_BLOCKi_14_Q_reg_30_inst : DFF_X1 port map( D => n3692, CK => CLK
                           , Q => n_2281, QN => 
                           DataPath_RF_bus_reg_dataout_222_port);
   DataPath_RF_BLOCKi_14_Q_reg_29_inst : DFF_X1 port map( D => n3693, CK => CLK
                           , Q => n_2282, QN => 
                           DataPath_RF_bus_reg_dataout_221_port);
   DataPath_RF_BLOCKi_14_Q_reg_28_inst : DFF_X1 port map( D => n3694, CK => CLK
                           , Q => n_2283, QN => 
                           DataPath_RF_bus_reg_dataout_220_port);
   DataPath_RF_BLOCKi_14_Q_reg_27_inst : DFF_X1 port map( D => n3695, CK => CLK
                           , Q => n_2284, QN => 
                           DataPath_RF_bus_reg_dataout_219_port);
   DataPath_RF_BLOCKi_14_Q_reg_26_inst : DFF_X1 port map( D => n3696, CK => CLK
                           , Q => n_2285, QN => 
                           DataPath_RF_bus_reg_dataout_218_port);
   DataPath_RF_BLOCKi_14_Q_reg_25_inst : DFF_X1 port map( D => n3697, CK => CLK
                           , Q => n_2286, QN => 
                           DataPath_RF_bus_reg_dataout_217_port);
   DataPath_RF_BLOCKi_14_Q_reg_24_inst : DFF_X1 port map( D => n3698, CK => CLK
                           , Q => n_2287, QN => 
                           DataPath_RF_bus_reg_dataout_216_port);
   DataPath_RF_BLOCKi_14_Q_reg_23_inst : DFF_X1 port map( D => n3699, CK => CLK
                           , Q => n_2288, QN => 
                           DataPath_RF_bus_reg_dataout_215_port);
   DataPath_RF_BLOCKi_14_Q_reg_22_inst : DFF_X1 port map( D => n3700, CK => CLK
                           , Q => n_2289, QN => 
                           DataPath_RF_bus_reg_dataout_214_port);
   DataPath_RF_BLOCKi_14_Q_reg_21_inst : DFF_X1 port map( D => n3701, CK => CLK
                           , Q => n_2290, QN => 
                           DataPath_RF_bus_reg_dataout_213_port);
   DataPath_RF_BLOCKi_14_Q_reg_20_inst : DFF_X1 port map( D => n3702, CK => CLK
                           , Q => n_2291, QN => 
                           DataPath_RF_bus_reg_dataout_212_port);
   DataPath_RF_BLOCKi_14_Q_reg_19_inst : DFF_X1 port map( D => n3703, CK => CLK
                           , Q => n_2292, QN => 
                           DataPath_RF_bus_reg_dataout_211_port);
   DataPath_RF_BLOCKi_14_Q_reg_18_inst : DFF_X1 port map( D => n3704, CK => CLK
                           , Q => n_2293, QN => 
                           DataPath_RF_bus_reg_dataout_210_port);
   DataPath_RF_BLOCKi_14_Q_reg_17_inst : DFF_X1 port map( D => n3705, CK => CLK
                           , Q => n_2294, QN => 
                           DataPath_RF_bus_reg_dataout_209_port);
   DataPath_RF_BLOCKi_14_Q_reg_16_inst : DFF_X1 port map( D => n3706, CK => CLK
                           , Q => n_2295, QN => 
                           DataPath_RF_bus_reg_dataout_208_port);
   DataPath_RF_BLOCKi_14_Q_reg_15_inst : DFF_X1 port map( D => n3707, CK => CLK
                           , Q => n_2296, QN => 
                           DataPath_RF_bus_reg_dataout_207_port);
   DataPath_RF_BLOCKi_14_Q_reg_14_inst : DFF_X1 port map( D => n3708, CK => CLK
                           , Q => n_2297, QN => 
                           DataPath_RF_bus_reg_dataout_206_port);
   DataPath_RF_BLOCKi_14_Q_reg_13_inst : DFF_X1 port map( D => n3709, CK => CLK
                           , Q => n_2298, QN => 
                           DataPath_RF_bus_reg_dataout_205_port);
   DataPath_RF_BLOCKi_14_Q_reg_12_inst : DFF_X1 port map( D => n3710, CK => CLK
                           , Q => n_2299, QN => 
                           DataPath_RF_bus_reg_dataout_204_port);
   DataPath_RF_BLOCKi_14_Q_reg_11_inst : DFF_X1 port map( D => n3711, CK => CLK
                           , Q => n_2300, QN => 
                           DataPath_RF_bus_reg_dataout_203_port);
   DataPath_RF_BLOCKi_14_Q_reg_9_inst : DFF_X1 port map( D => n3713, CK => CLK,
                           Q => n_2301, QN => 
                           DataPath_RF_bus_reg_dataout_201_port);
   DataPath_RF_BLOCKi_14_Q_reg_8_inst : DFF_X1 port map( D => n3714, CK => CLK,
                           Q => n_2302, QN => 
                           DataPath_RF_bus_reg_dataout_200_port);
   DataPath_RF_BLOCKi_14_Q_reg_7_inst : DFF_X1 port map( D => n3715, CK => CLK,
                           Q => n_2303, QN => 
                           DataPath_RF_bus_reg_dataout_199_port);
   DataPath_RF_BLOCKi_14_Q_reg_6_inst : DFF_X1 port map( D => n3716, CK => CLK,
                           Q => n_2304, QN => 
                           DataPath_RF_bus_reg_dataout_198_port);
   DataPath_RF_BLOCKi_14_Q_reg_5_inst : DFF_X1 port map( D => n3717, CK => CLK,
                           Q => n_2305, QN => 
                           DataPath_RF_bus_reg_dataout_197_port);
   DataPath_RF_BLOCKi_14_Q_reg_4_inst : DFF_X1 port map( D => n3718, CK => CLK,
                           Q => n_2306, QN => 
                           DataPath_RF_bus_reg_dataout_196_port);
   DataPath_RF_BLOCKi_14_Q_reg_3_inst : DFF_X1 port map( D => n3719, CK => CLK,
                           Q => n_2307, QN => 
                           DataPath_RF_bus_reg_dataout_195_port);
   DataPath_RF_BLOCKi_14_Q_reg_2_inst : DFF_X1 port map( D => n3720, CK => CLK,
                           Q => n_2308, QN => 
                           DataPath_RF_bus_reg_dataout_194_port);
   DataPath_RF_BLOCKi_14_Q_reg_1_inst : DFF_X1 port map( D => n3721, CK => CLK,
                           Q => n_2309, QN => 
                           DataPath_RF_bus_reg_dataout_193_port);
   DataPath_RF_BLOCKi_14_Q_reg_0_inst : DFF_X1 port map( D => n3722, CK => CLK,
                           Q => n_2310, QN => 
                           DataPath_RF_bus_reg_dataout_192_port);
   DataPath_RF_BLOCKi_30_Q_reg_31_inst : DFF_X1 port map( D => n4320, CK => CLK
                           , Q => n_2311, QN => 
                           DataPath_RF_bus_reg_dataout_735_port);
   DataPath_RF_BLOCKi_30_Q_reg_30_inst : DFF_X1 port map( D => n4323, CK => CLK
                           , Q => n_2312, QN => 
                           DataPath_RF_bus_reg_dataout_734_port);
   DataPath_RF_BLOCKi_30_Q_reg_29_inst : DFF_X1 port map( D => n4324, CK => CLK
                           , Q => n_2313, QN => 
                           DataPath_RF_bus_reg_dataout_733_port);
   DataPath_RF_BLOCKi_30_Q_reg_28_inst : DFF_X1 port map( D => n4325, CK => CLK
                           , Q => n_2314, QN => 
                           DataPath_RF_bus_reg_dataout_732_port);
   DataPath_RF_BLOCKi_30_Q_reg_27_inst : DFF_X1 port map( D => n4326, CK => CLK
                           , Q => n_2315, QN => 
                           DataPath_RF_bus_reg_dataout_731_port);
   DataPath_RF_BLOCKi_30_Q_reg_26_inst : DFF_X1 port map( D => n4327, CK => CLK
                           , Q => n_2316, QN => 
                           DataPath_RF_bus_reg_dataout_730_port);
   DataPath_RF_BLOCKi_30_Q_reg_25_inst : DFF_X1 port map( D => n4328, CK => CLK
                           , Q => n_2317, QN => 
                           DataPath_RF_bus_reg_dataout_729_port);
   DataPath_RF_BLOCKi_30_Q_reg_24_inst : DFF_X1 port map( D => n4329, CK => CLK
                           , Q => n_2318, QN => 
                           DataPath_RF_bus_reg_dataout_728_port);
   DataPath_RF_BLOCKi_30_Q_reg_23_inst : DFF_X1 port map( D => n4330, CK => CLK
                           , Q => n_2319, QN => 
                           DataPath_RF_bus_reg_dataout_727_port);
   DataPath_RF_BLOCKi_30_Q_reg_22_inst : DFF_X1 port map( D => n4331, CK => CLK
                           , Q => n_2320, QN => 
                           DataPath_RF_bus_reg_dataout_726_port);
   DataPath_RF_BLOCKi_30_Q_reg_21_inst : DFF_X1 port map( D => n4332, CK => CLK
                           , Q => n_2321, QN => 
                           DataPath_RF_bus_reg_dataout_725_port);
   DataPath_RF_BLOCKi_30_Q_reg_20_inst : DFF_X1 port map( D => n4333, CK => CLK
                           , Q => n_2322, QN => 
                           DataPath_RF_bus_reg_dataout_724_port);
   DataPath_RF_BLOCKi_30_Q_reg_19_inst : DFF_X1 port map( D => n4334, CK => CLK
                           , Q => n_2323, QN => 
                           DataPath_RF_bus_reg_dataout_723_port);
   DataPath_RF_BLOCKi_30_Q_reg_18_inst : DFF_X1 port map( D => n4335, CK => CLK
                           , Q => n_2324, QN => 
                           DataPath_RF_bus_reg_dataout_722_port);
   DataPath_RF_BLOCKi_30_Q_reg_17_inst : DFF_X1 port map( D => n4336, CK => CLK
                           , Q => n_2325, QN => 
                           DataPath_RF_bus_reg_dataout_721_port);
   DataPath_RF_BLOCKi_30_Q_reg_16_inst : DFF_X1 port map( D => n4337, CK => CLK
                           , Q => n_2326, QN => 
                           DataPath_RF_bus_reg_dataout_720_port);
   DataPath_RF_BLOCKi_30_Q_reg_15_inst : DFF_X1 port map( D => n4338, CK => CLK
                           , Q => n_2327, QN => 
                           DataPath_RF_bus_reg_dataout_719_port);
   DataPath_RF_BLOCKi_30_Q_reg_14_inst : DFF_X1 port map( D => n4339, CK => CLK
                           , Q => n_2328, QN => 
                           DataPath_RF_bus_reg_dataout_718_port);
   DataPath_RF_BLOCKi_30_Q_reg_13_inst : DFF_X1 port map( D => n4340, CK => CLK
                           , Q => n_2329, QN => 
                           DataPath_RF_bus_reg_dataout_717_port);
   DataPath_RF_BLOCKi_30_Q_reg_12_inst : DFF_X1 port map( D => n4341, CK => CLK
                           , Q => n_2330, QN => 
                           DataPath_RF_bus_reg_dataout_716_port);
   DataPath_RF_BLOCKi_30_Q_reg_11_inst : DFF_X1 port map( D => n4342, CK => CLK
                           , Q => n_2331, QN => 
                           DataPath_RF_bus_reg_dataout_715_port);
   DataPath_RF_BLOCKi_30_Q_reg_9_inst : DFF_X1 port map( D => n4344, CK => CLK,
                           Q => n_2332, QN => 
                           DataPath_RF_bus_reg_dataout_713_port);
   DataPath_RF_BLOCKi_30_Q_reg_8_inst : DFF_X1 port map( D => n4345, CK => CLK,
                           Q => n_2333, QN => 
                           DataPath_RF_bus_reg_dataout_712_port);
   DataPath_RF_BLOCKi_30_Q_reg_7_inst : DFF_X1 port map( D => n4346, CK => CLK,
                           Q => n_2334, QN => 
                           DataPath_RF_bus_reg_dataout_711_port);
   DataPath_RF_BLOCKi_30_Q_reg_6_inst : DFF_X1 port map( D => n4347, CK => CLK,
                           Q => n_2335, QN => 
                           DataPath_RF_bus_reg_dataout_710_port);
   DataPath_RF_BLOCKi_30_Q_reg_5_inst : DFF_X1 port map( D => n4348, CK => CLK,
                           Q => n_2336, QN => 
                           DataPath_RF_bus_reg_dataout_709_port);
   DataPath_RF_BLOCKi_30_Q_reg_4_inst : DFF_X1 port map( D => n4349, CK => CLK,
                           Q => n_2337, QN => 
                           DataPath_RF_bus_reg_dataout_708_port);
   DataPath_RF_BLOCKi_30_Q_reg_3_inst : DFF_X1 port map( D => n4350, CK => CLK,
                           Q => n_2338, QN => 
                           DataPath_RF_bus_reg_dataout_707_port);
   DataPath_RF_BLOCKi_30_Q_reg_2_inst : DFF_X1 port map( D => n4351, CK => CLK,
                           Q => n_2339, QN => 
                           DataPath_RF_bus_reg_dataout_706_port);
   DataPath_RF_BLOCKi_30_Q_reg_1_inst : DFF_X1 port map( D => n4352, CK => CLK,
                           Q => n_2340, QN => 
                           DataPath_RF_bus_reg_dataout_705_port);
   DataPath_RF_BLOCKi_30_Q_reg_0_inst : DFF_X1 port map( D => n4353, CK => CLK,
                           Q => n_2341, QN => 
                           DataPath_RF_bus_reg_dataout_704_port);
   DataPath_RF_BLOCKi_46_Q_reg_31_inst : DFF_X1 port map( D => n4913, CK => CLK
                           , Q => n_2342, QN => 
                           DataPath_RF_bus_reg_dataout_1247_port);
   DataPath_RF_BLOCKi_46_Q_reg_30_inst : DFF_X1 port map( D => n4916, CK => CLK
                           , Q => n_2343, QN => 
                           DataPath_RF_bus_reg_dataout_1246_port);
   DataPath_RF_BLOCKi_46_Q_reg_29_inst : DFF_X1 port map( D => n4917, CK => CLK
                           , Q => n_2344, QN => 
                           DataPath_RF_bus_reg_dataout_1245_port);
   DataPath_RF_BLOCKi_46_Q_reg_28_inst : DFF_X1 port map( D => n4918, CK => CLK
                           , Q => n_2345, QN => 
                           DataPath_RF_bus_reg_dataout_1244_port);
   DataPath_RF_BLOCKi_46_Q_reg_27_inst : DFF_X1 port map( D => n4919, CK => CLK
                           , Q => n_2346, QN => 
                           DataPath_RF_bus_reg_dataout_1243_port);
   DataPath_RF_BLOCKi_46_Q_reg_26_inst : DFF_X1 port map( D => n4920, CK => CLK
                           , Q => n_2347, QN => 
                           DataPath_RF_bus_reg_dataout_1242_port);
   DataPath_RF_BLOCKi_46_Q_reg_25_inst : DFF_X1 port map( D => n4921, CK => CLK
                           , Q => n_2348, QN => 
                           DataPath_RF_bus_reg_dataout_1241_port);
   DataPath_RF_BLOCKi_46_Q_reg_24_inst : DFF_X1 port map( D => n4922, CK => CLK
                           , Q => n_2349, QN => 
                           DataPath_RF_bus_reg_dataout_1240_port);
   DataPath_RF_BLOCKi_46_Q_reg_23_inst : DFF_X1 port map( D => n4923, CK => CLK
                           , Q => n_2350, QN => 
                           DataPath_RF_bus_reg_dataout_1239_port);
   DataPath_RF_BLOCKi_46_Q_reg_22_inst : DFF_X1 port map( D => n4924, CK => CLK
                           , Q => n_2351, QN => 
                           DataPath_RF_bus_reg_dataout_1238_port);
   DataPath_RF_BLOCKi_46_Q_reg_21_inst : DFF_X1 port map( D => n4925, CK => CLK
                           , Q => n_2352, QN => 
                           DataPath_RF_bus_reg_dataout_1237_port);
   DataPath_RF_BLOCKi_46_Q_reg_20_inst : DFF_X1 port map( D => n4926, CK => CLK
                           , Q => n_2353, QN => 
                           DataPath_RF_bus_reg_dataout_1236_port);
   DataPath_RF_BLOCKi_46_Q_reg_19_inst : DFF_X1 port map( D => n4927, CK => CLK
                           , Q => n_2354, QN => 
                           DataPath_RF_bus_reg_dataout_1235_port);
   DataPath_RF_BLOCKi_46_Q_reg_18_inst : DFF_X1 port map( D => n4928, CK => CLK
                           , Q => n_2355, QN => 
                           DataPath_RF_bus_reg_dataout_1234_port);
   DataPath_RF_BLOCKi_46_Q_reg_17_inst : DFF_X1 port map( D => n4929, CK => CLK
                           , Q => n_2356, QN => 
                           DataPath_RF_bus_reg_dataout_1233_port);
   DataPath_RF_BLOCKi_46_Q_reg_16_inst : DFF_X1 port map( D => n4930, CK => CLK
                           , Q => n_2357, QN => 
                           DataPath_RF_bus_reg_dataout_1232_port);
   DataPath_RF_BLOCKi_46_Q_reg_15_inst : DFF_X1 port map( D => n4931, CK => CLK
                           , Q => n_2358, QN => 
                           DataPath_RF_bus_reg_dataout_1231_port);
   DataPath_RF_BLOCKi_46_Q_reg_14_inst : DFF_X1 port map( D => n4932, CK => CLK
                           , Q => n_2359, QN => 
                           DataPath_RF_bus_reg_dataout_1230_port);
   DataPath_RF_BLOCKi_46_Q_reg_13_inst : DFF_X1 port map( D => n4933, CK => CLK
                           , Q => n_2360, QN => 
                           DataPath_RF_bus_reg_dataout_1229_port);
   DataPath_RF_BLOCKi_46_Q_reg_12_inst : DFF_X1 port map( D => n4934, CK => CLK
                           , Q => n_2361, QN => 
                           DataPath_RF_bus_reg_dataout_1228_port);
   DataPath_RF_BLOCKi_46_Q_reg_11_inst : DFF_X1 port map( D => n4935, CK => CLK
                           , Q => n_2362, QN => 
                           DataPath_RF_bus_reg_dataout_1227_port);
   DataPath_RF_BLOCKi_46_Q_reg_9_inst : DFF_X1 port map( D => n4937, CK => CLK,
                           Q => n_2363, QN => 
                           DataPath_RF_bus_reg_dataout_1225_port);
   DataPath_RF_BLOCKi_46_Q_reg_8_inst : DFF_X1 port map( D => n4938, CK => CLK,
                           Q => n_2364, QN => 
                           DataPath_RF_bus_reg_dataout_1224_port);
   DataPath_RF_BLOCKi_46_Q_reg_7_inst : DFF_X1 port map( D => n4939, CK => CLK,
                           Q => n_2365, QN => 
                           DataPath_RF_bus_reg_dataout_1223_port);
   DataPath_RF_BLOCKi_46_Q_reg_6_inst : DFF_X1 port map( D => n4940, CK => CLK,
                           Q => n_2366, QN => 
                           DataPath_RF_bus_reg_dataout_1222_port);
   DataPath_RF_BLOCKi_46_Q_reg_5_inst : DFF_X1 port map( D => n4941, CK => CLK,
                           Q => n_2367, QN => 
                           DataPath_RF_bus_reg_dataout_1221_port);
   DataPath_RF_BLOCKi_46_Q_reg_4_inst : DFF_X1 port map( D => n4942, CK => CLK,
                           Q => n_2368, QN => 
                           DataPath_RF_bus_reg_dataout_1220_port);
   DataPath_RF_BLOCKi_46_Q_reg_3_inst : DFF_X1 port map( D => n4943, CK => CLK,
                           Q => n_2369, QN => 
                           DataPath_RF_bus_reg_dataout_1219_port);
   DataPath_RF_BLOCKi_46_Q_reg_2_inst : DFF_X1 port map( D => n4944, CK => CLK,
                           Q => n_2370, QN => 
                           DataPath_RF_bus_reg_dataout_1218_port);
   DataPath_RF_BLOCKi_46_Q_reg_1_inst : DFF_X1 port map( D => n4945, CK => CLK,
                           Q => n_2371, QN => 
                           DataPath_RF_bus_reg_dataout_1217_port);
   DataPath_RF_BLOCKi_46_Q_reg_0_inst : DFF_X1 port map( D => n4946, CK => CLK,
                           Q => n_2372, QN => 
                           DataPath_RF_bus_reg_dataout_1216_port);
   DataPath_RF_BLOCKi_62_Q_reg_31_inst : DFF_X1 port map( D => n5506, CK => CLK
                           , Q => n_2373, QN => 
                           DataPath_RF_bus_reg_dataout_1759_port);
   DataPath_RF_BLOCKi_62_Q_reg_30_inst : DFF_X1 port map( D => n5509, CK => CLK
                           , Q => n_2374, QN => 
                           DataPath_RF_bus_reg_dataout_1758_port);
   DataPath_RF_BLOCKi_62_Q_reg_29_inst : DFF_X1 port map( D => n5510, CK => CLK
                           , Q => n_2375, QN => 
                           DataPath_RF_bus_reg_dataout_1757_port);
   DataPath_RF_BLOCKi_62_Q_reg_28_inst : DFF_X1 port map( D => n5511, CK => CLK
                           , Q => n_2376, QN => 
                           DataPath_RF_bus_reg_dataout_1756_port);
   DataPath_RF_BLOCKi_62_Q_reg_27_inst : DFF_X1 port map( D => n5512, CK => CLK
                           , Q => n_2377, QN => 
                           DataPath_RF_bus_reg_dataout_1755_port);
   DataPath_RF_BLOCKi_62_Q_reg_26_inst : DFF_X1 port map( D => n5513, CK => CLK
                           , Q => n_2378, QN => 
                           DataPath_RF_bus_reg_dataout_1754_port);
   DataPath_RF_BLOCKi_62_Q_reg_25_inst : DFF_X1 port map( D => n5514, CK => CLK
                           , Q => n_2379, QN => 
                           DataPath_RF_bus_reg_dataout_1753_port);
   DataPath_RF_BLOCKi_62_Q_reg_24_inst : DFF_X1 port map( D => n5515, CK => CLK
                           , Q => n_2380, QN => 
                           DataPath_RF_bus_reg_dataout_1752_port);
   DataPath_RF_BLOCKi_62_Q_reg_23_inst : DFF_X1 port map( D => n5516, CK => CLK
                           , Q => n_2381, QN => 
                           DataPath_RF_bus_reg_dataout_1751_port);
   DataPath_RF_BLOCKi_62_Q_reg_22_inst : DFF_X1 port map( D => n5517, CK => CLK
                           , Q => n_2382, QN => 
                           DataPath_RF_bus_reg_dataout_1750_port);
   DataPath_RF_BLOCKi_62_Q_reg_21_inst : DFF_X1 port map( D => n5518, CK => CLK
                           , Q => n_2383, QN => 
                           DataPath_RF_bus_reg_dataout_1749_port);
   DataPath_RF_BLOCKi_62_Q_reg_20_inst : DFF_X1 port map( D => n5519, CK => CLK
                           , Q => n_2384, QN => 
                           DataPath_RF_bus_reg_dataout_1748_port);
   DataPath_RF_BLOCKi_62_Q_reg_19_inst : DFF_X1 port map( D => n5520, CK => CLK
                           , Q => n_2385, QN => 
                           DataPath_RF_bus_reg_dataout_1747_port);
   DataPath_RF_BLOCKi_62_Q_reg_18_inst : DFF_X1 port map( D => n5521, CK => CLK
                           , Q => n_2386, QN => 
                           DataPath_RF_bus_reg_dataout_1746_port);
   DataPath_RF_BLOCKi_62_Q_reg_17_inst : DFF_X1 port map( D => n5522, CK => CLK
                           , Q => n_2387, QN => 
                           DataPath_RF_bus_reg_dataout_1745_port);
   DataPath_RF_BLOCKi_62_Q_reg_16_inst : DFF_X1 port map( D => n5523, CK => CLK
                           , Q => n_2388, QN => 
                           DataPath_RF_bus_reg_dataout_1744_port);
   DataPath_RF_BLOCKi_62_Q_reg_15_inst : DFF_X1 port map( D => n5524, CK => CLK
                           , Q => n_2389, QN => 
                           DataPath_RF_bus_reg_dataout_1743_port);
   DataPath_RF_BLOCKi_62_Q_reg_14_inst : DFF_X1 port map( D => n5525, CK => CLK
                           , Q => n_2390, QN => 
                           DataPath_RF_bus_reg_dataout_1742_port);
   DataPath_RF_BLOCKi_62_Q_reg_13_inst : DFF_X1 port map( D => n5526, CK => CLK
                           , Q => n_2391, QN => 
                           DataPath_RF_bus_reg_dataout_1741_port);
   DataPath_RF_BLOCKi_62_Q_reg_12_inst : DFF_X1 port map( D => n5527, CK => CLK
                           , Q => n_2392, QN => 
                           DataPath_RF_bus_reg_dataout_1740_port);
   DataPath_RF_BLOCKi_62_Q_reg_11_inst : DFF_X1 port map( D => n5528, CK => CLK
                           , Q => n_2393, QN => 
                           DataPath_RF_bus_reg_dataout_1739_port);
   DataPath_RF_BLOCKi_62_Q_reg_9_inst : DFF_X1 port map( D => n5530, CK => CLK,
                           Q => n_2394, QN => 
                           DataPath_RF_bus_reg_dataout_1737_port);
   DataPath_RF_BLOCKi_62_Q_reg_8_inst : DFF_X1 port map( D => n5531, CK => CLK,
                           Q => n_2395, QN => 
                           DataPath_RF_bus_reg_dataout_1736_port);
   DataPath_RF_BLOCKi_62_Q_reg_7_inst : DFF_X1 port map( D => n5532, CK => CLK,
                           Q => n_2396, QN => 
                           DataPath_RF_bus_reg_dataout_1735_port);
   DataPath_RF_BLOCKi_62_Q_reg_6_inst : DFF_X1 port map( D => n5533, CK => CLK,
                           Q => n_2397, QN => 
                           DataPath_RF_bus_reg_dataout_1734_port);
   DataPath_RF_BLOCKi_62_Q_reg_5_inst : DFF_X1 port map( D => n5534, CK => CLK,
                           Q => n_2398, QN => 
                           DataPath_RF_bus_reg_dataout_1733_port);
   DataPath_RF_BLOCKi_62_Q_reg_4_inst : DFF_X1 port map( D => n5535, CK => CLK,
                           Q => n_2399, QN => 
                           DataPath_RF_bus_reg_dataout_1732_port);
   DataPath_RF_BLOCKi_62_Q_reg_3_inst : DFF_X1 port map( D => n5536, CK => CLK,
                           Q => n_2400, QN => 
                           DataPath_RF_bus_reg_dataout_1731_port);
   DataPath_RF_BLOCKi_62_Q_reg_2_inst : DFF_X1 port map( D => n5537, CK => CLK,
                           Q => n_2401, QN => 
                           DataPath_RF_bus_reg_dataout_1730_port);
   DataPath_RF_BLOCKi_62_Q_reg_1_inst : DFF_X1 port map( D => n5538, CK => CLK,
                           Q => n_2402, QN => 
                           DataPath_RF_bus_reg_dataout_1729_port);
   DataPath_RF_BLOCKi_62_Q_reg_0_inst : DFF_X1 port map( D => n5539, CK => CLK,
                           Q => n_2403, QN => 
                           DataPath_RF_bus_reg_dataout_1728_port);
   DataPath_RF_BLOCKi_78_Q_reg_31_inst : DFF_X1 port map( D => n6090, CK => CLK
                           , Q => n_2404, QN => 
                           DataPath_RF_bus_reg_dataout_2271_port);
   DataPath_RF_BLOCKi_78_Q_reg_30_inst : DFF_X1 port map( D => n6093, CK => CLK
                           , Q => n_2405, QN => 
                           DataPath_RF_bus_reg_dataout_2270_port);
   DataPath_RF_BLOCKi_78_Q_reg_29_inst : DFF_X1 port map( D => n6094, CK => CLK
                           , Q => n_2406, QN => 
                           DataPath_RF_bus_reg_dataout_2269_port);
   DataPath_RF_BLOCKi_78_Q_reg_28_inst : DFF_X1 port map( D => n6095, CK => CLK
                           , Q => n_2407, QN => 
                           DataPath_RF_bus_reg_dataout_2268_port);
   DataPath_RF_BLOCKi_78_Q_reg_27_inst : DFF_X1 port map( D => n6096, CK => CLK
                           , Q => n_2408, QN => 
                           DataPath_RF_bus_reg_dataout_2267_port);
   DataPath_RF_BLOCKi_78_Q_reg_26_inst : DFF_X1 port map( D => n6097, CK => CLK
                           , Q => n_2409, QN => 
                           DataPath_RF_bus_reg_dataout_2266_port);
   DataPath_RF_BLOCKi_78_Q_reg_25_inst : DFF_X1 port map( D => n6098, CK => CLK
                           , Q => n_2410, QN => 
                           DataPath_RF_bus_reg_dataout_2265_port);
   DataPath_RF_BLOCKi_78_Q_reg_24_inst : DFF_X1 port map( D => n6099, CK => CLK
                           , Q => n_2411, QN => 
                           DataPath_RF_bus_reg_dataout_2264_port);
   DataPath_RF_BLOCKi_78_Q_reg_23_inst : DFF_X1 port map( D => n6100, CK => CLK
                           , Q => n_2412, QN => 
                           DataPath_RF_bus_reg_dataout_2263_port);
   DataPath_RF_BLOCKi_78_Q_reg_22_inst : DFF_X1 port map( D => n6101, CK => CLK
                           , Q => n_2413, QN => 
                           DataPath_RF_bus_reg_dataout_2262_port);
   DataPath_RF_BLOCKi_78_Q_reg_21_inst : DFF_X1 port map( D => n6102, CK => CLK
                           , Q => n_2414, QN => 
                           DataPath_RF_bus_reg_dataout_2261_port);
   DataPath_RF_BLOCKi_78_Q_reg_20_inst : DFF_X1 port map( D => n6103, CK => CLK
                           , Q => n_2415, QN => 
                           DataPath_RF_bus_reg_dataout_2260_port);
   DataPath_RF_BLOCKi_78_Q_reg_19_inst : DFF_X1 port map( D => n6104, CK => CLK
                           , Q => n_2416, QN => 
                           DataPath_RF_bus_reg_dataout_2259_port);
   DataPath_RF_BLOCKi_78_Q_reg_18_inst : DFF_X1 port map( D => n6105, CK => CLK
                           , Q => n_2417, QN => 
                           DataPath_RF_bus_reg_dataout_2258_port);
   DataPath_RF_BLOCKi_78_Q_reg_17_inst : DFF_X1 port map( D => n6106, CK => CLK
                           , Q => n_2418, QN => 
                           DataPath_RF_bus_reg_dataout_2257_port);
   DataPath_RF_BLOCKi_78_Q_reg_16_inst : DFF_X1 port map( D => n6107, CK => CLK
                           , Q => n_2419, QN => 
                           DataPath_RF_bus_reg_dataout_2256_port);
   DataPath_RF_BLOCKi_78_Q_reg_15_inst : DFF_X1 port map( D => n6108, CK => CLK
                           , Q => n_2420, QN => 
                           DataPath_RF_bus_reg_dataout_2255_port);
   DataPath_RF_BLOCKi_78_Q_reg_14_inst : DFF_X1 port map( D => n6109, CK => CLK
                           , Q => n_2421, QN => 
                           DataPath_RF_bus_reg_dataout_2254_port);
   DataPath_RF_BLOCKi_78_Q_reg_13_inst : DFF_X1 port map( D => n6110, CK => CLK
                           , Q => n_2422, QN => 
                           DataPath_RF_bus_reg_dataout_2253_port);
   DataPath_RF_BLOCKi_78_Q_reg_12_inst : DFF_X1 port map( D => n6111, CK => CLK
                           , Q => n_2423, QN => 
                           DataPath_RF_bus_reg_dataout_2252_port);
   DataPath_RF_BLOCKi_78_Q_reg_11_inst : DFF_X1 port map( D => n6112, CK => CLK
                           , Q => n_2424, QN => 
                           DataPath_RF_bus_reg_dataout_2251_port);
   DataPath_RF_BLOCKi_78_Q_reg_9_inst : DFF_X1 port map( D => n6114, CK => CLK,
                           Q => n_2425, QN => 
                           DataPath_RF_bus_reg_dataout_2249_port);
   DataPath_RF_BLOCKi_78_Q_reg_8_inst : DFF_X1 port map( D => n6115, CK => CLK,
                           Q => n_2426, QN => 
                           DataPath_RF_bus_reg_dataout_2248_port);
   DataPath_RF_BLOCKi_78_Q_reg_7_inst : DFF_X1 port map( D => n6116, CK => CLK,
                           Q => n_2427, QN => 
                           DataPath_RF_bus_reg_dataout_2247_port);
   DataPath_RF_BLOCKi_78_Q_reg_6_inst : DFF_X1 port map( D => n6117, CK => CLK,
                           Q => n_2428, QN => 
                           DataPath_RF_bus_reg_dataout_2246_port);
   DataPath_RF_BLOCKi_78_Q_reg_5_inst : DFF_X1 port map( D => n6118, CK => CLK,
                           Q => n_2429, QN => 
                           DataPath_RF_bus_reg_dataout_2245_port);
   DataPath_RF_BLOCKi_78_Q_reg_4_inst : DFF_X1 port map( D => n6119, CK => CLK,
                           Q => n_2430, QN => 
                           DataPath_RF_bus_reg_dataout_2244_port);
   DataPath_RF_BLOCKi_78_Q_reg_3_inst : DFF_X1 port map( D => n6120, CK => CLK,
                           Q => n_2431, QN => 
                           DataPath_RF_bus_reg_dataout_2243_port);
   DataPath_RF_BLOCKi_78_Q_reg_2_inst : DFF_X1 port map( D => n6121, CK => CLK,
                           Q => n_2432, QN => 
                           DataPath_RF_bus_reg_dataout_2242_port);
   DataPath_RF_BLOCKi_78_Q_reg_1_inst : DFF_X1 port map( D => n6122, CK => CLK,
                           Q => n_2433, QN => 
                           DataPath_RF_bus_reg_dataout_2241_port);
   DataPath_RF_BLOCKi_78_Q_reg_0_inst : DFF_X1 port map( D => n6123, CK => CLK,
                           Q => n_2434, QN => 
                           DataPath_RF_bus_reg_dataout_2240_port);
   DataPath_RF_BLOCKi_15_Q_reg_31_inst : DFF_X1 port map( D => n3727, CK => CLK
                           , Q => n_2435, QN => 
                           DataPath_RF_bus_reg_dataout_255_port);
   DataPath_RF_BLOCKi_15_Q_reg_30_inst : DFF_X1 port map( D => n3730, CK => CLK
                           , Q => n_2436, QN => 
                           DataPath_RF_bus_reg_dataout_254_port);
   DataPath_RF_BLOCKi_15_Q_reg_29_inst : DFF_X1 port map( D => n3731, CK => CLK
                           , Q => n_2437, QN => 
                           DataPath_RF_bus_reg_dataout_253_port);
   DataPath_RF_BLOCKi_15_Q_reg_28_inst : DFF_X1 port map( D => n3732, CK => CLK
                           , Q => n_2438, QN => 
                           DataPath_RF_bus_reg_dataout_252_port);
   DataPath_RF_BLOCKi_15_Q_reg_27_inst : DFF_X1 port map( D => n3733, CK => CLK
                           , Q => n_2439, QN => 
                           DataPath_RF_bus_reg_dataout_251_port);
   DataPath_RF_BLOCKi_15_Q_reg_26_inst : DFF_X1 port map( D => n3734, CK => CLK
                           , Q => n_2440, QN => 
                           DataPath_RF_bus_reg_dataout_250_port);
   DataPath_RF_BLOCKi_15_Q_reg_25_inst : DFF_X1 port map( D => n3735, CK => CLK
                           , Q => n_2441, QN => 
                           DataPath_RF_bus_reg_dataout_249_port);
   DataPath_RF_BLOCKi_15_Q_reg_24_inst : DFF_X1 port map( D => n3736, CK => CLK
                           , Q => n_2442, QN => 
                           DataPath_RF_bus_reg_dataout_248_port);
   DataPath_RF_BLOCKi_15_Q_reg_23_inst : DFF_X1 port map( D => n3737, CK => CLK
                           , Q => n_2443, QN => 
                           DataPath_RF_bus_reg_dataout_247_port);
   DataPath_RF_BLOCKi_15_Q_reg_22_inst : DFF_X1 port map( D => n3738, CK => CLK
                           , Q => n_2444, QN => 
                           DataPath_RF_bus_reg_dataout_246_port);
   DataPath_RF_BLOCKi_15_Q_reg_21_inst : DFF_X1 port map( D => n3739, CK => CLK
                           , Q => n_2445, QN => 
                           DataPath_RF_bus_reg_dataout_245_port);
   DataPath_RF_BLOCKi_15_Q_reg_20_inst : DFF_X1 port map( D => n3740, CK => CLK
                           , Q => n_2446, QN => 
                           DataPath_RF_bus_reg_dataout_244_port);
   DataPath_RF_BLOCKi_15_Q_reg_19_inst : DFF_X1 port map( D => n3741, CK => CLK
                           , Q => n_2447, QN => 
                           DataPath_RF_bus_reg_dataout_243_port);
   DataPath_RF_BLOCKi_15_Q_reg_18_inst : DFF_X1 port map( D => n3742, CK => CLK
                           , Q => n_2448, QN => 
                           DataPath_RF_bus_reg_dataout_242_port);
   DataPath_RF_BLOCKi_15_Q_reg_17_inst : DFF_X1 port map( D => n3743, CK => CLK
                           , Q => n_2449, QN => 
                           DataPath_RF_bus_reg_dataout_241_port);
   DataPath_RF_BLOCKi_15_Q_reg_16_inst : DFF_X1 port map( D => n3744, CK => CLK
                           , Q => n_2450, QN => 
                           DataPath_RF_bus_reg_dataout_240_port);
   DataPath_RF_BLOCKi_15_Q_reg_15_inst : DFF_X1 port map( D => n3745, CK => CLK
                           , Q => n_2451, QN => 
                           DataPath_RF_bus_reg_dataout_239_port);
   DataPath_RF_BLOCKi_15_Q_reg_14_inst : DFF_X1 port map( D => n3746, CK => CLK
                           , Q => n_2452, QN => 
                           DataPath_RF_bus_reg_dataout_238_port);
   DataPath_RF_BLOCKi_15_Q_reg_13_inst : DFF_X1 port map( D => n3747, CK => CLK
                           , Q => n_2453, QN => 
                           DataPath_RF_bus_reg_dataout_237_port);
   DataPath_RF_BLOCKi_15_Q_reg_12_inst : DFF_X1 port map( D => n3748, CK => CLK
                           , Q => n_2454, QN => 
                           DataPath_RF_bus_reg_dataout_236_port);
   DataPath_RF_BLOCKi_15_Q_reg_11_inst : DFF_X1 port map( D => n3749, CK => CLK
                           , Q => n_2455, QN => 
                           DataPath_RF_bus_reg_dataout_235_port);
   DataPath_RF_BLOCKi_15_Q_reg_9_inst : DFF_X1 port map( D => n3751, CK => CLK,
                           Q => n_2456, QN => 
                           DataPath_RF_bus_reg_dataout_233_port);
   DataPath_RF_BLOCKi_15_Q_reg_8_inst : DFF_X1 port map( D => n3752, CK => CLK,
                           Q => n_2457, QN => 
                           DataPath_RF_bus_reg_dataout_232_port);
   DataPath_RF_BLOCKi_15_Q_reg_7_inst : DFF_X1 port map( D => n3753, CK => CLK,
                           Q => n_2458, QN => 
                           DataPath_RF_bus_reg_dataout_231_port);
   DataPath_RF_BLOCKi_15_Q_reg_6_inst : DFF_X1 port map( D => n3754, CK => CLK,
                           Q => n_2459, QN => 
                           DataPath_RF_bus_reg_dataout_230_port);
   DataPath_RF_BLOCKi_15_Q_reg_5_inst : DFF_X1 port map( D => n3755, CK => CLK,
                           Q => n_2460, QN => 
                           DataPath_RF_bus_reg_dataout_229_port);
   DataPath_RF_BLOCKi_15_Q_reg_4_inst : DFF_X1 port map( D => n3756, CK => CLK,
                           Q => n_2461, QN => 
                           DataPath_RF_bus_reg_dataout_228_port);
   DataPath_RF_BLOCKi_15_Q_reg_3_inst : DFF_X1 port map( D => n3757, CK => CLK,
                           Q => n_2462, QN => 
                           DataPath_RF_bus_reg_dataout_227_port);
   DataPath_RF_BLOCKi_15_Q_reg_2_inst : DFF_X1 port map( D => n3758, CK => CLK,
                           Q => n_2463, QN => 
                           DataPath_RF_bus_reg_dataout_226_port);
   DataPath_RF_BLOCKi_15_Q_reg_1_inst : DFF_X1 port map( D => n3759, CK => CLK,
                           Q => n_2464, QN => 
                           DataPath_RF_bus_reg_dataout_225_port);
   DataPath_RF_BLOCKi_15_Q_reg_0_inst : DFF_X1 port map( D => n3760, CK => CLK,
                           Q => n_2465, QN => 
                           DataPath_RF_bus_reg_dataout_224_port);
   DataPath_RF_BLOCKi_31_Q_reg_31_inst : DFF_X1 port map( D => n4355, CK => CLK
                           , Q => n_2466, QN => 
                           DataPath_RF_bus_reg_dataout_767_port);
   DataPath_RF_BLOCKi_31_Q_reg_30_inst : DFF_X1 port map( D => n4358, CK => CLK
                           , Q => n_2467, QN => 
                           DataPath_RF_bus_reg_dataout_766_port);
   DataPath_RF_BLOCKi_31_Q_reg_29_inst : DFF_X1 port map( D => n4359, CK => CLK
                           , Q => n_2468, QN => 
                           DataPath_RF_bus_reg_dataout_765_port);
   DataPath_RF_BLOCKi_31_Q_reg_28_inst : DFF_X1 port map( D => n4360, CK => CLK
                           , Q => n_2469, QN => 
                           DataPath_RF_bus_reg_dataout_764_port);
   DataPath_RF_BLOCKi_31_Q_reg_27_inst : DFF_X1 port map( D => n4361, CK => CLK
                           , Q => n_2470, QN => 
                           DataPath_RF_bus_reg_dataout_763_port);
   DataPath_RF_BLOCKi_31_Q_reg_26_inst : DFF_X1 port map( D => n4362, CK => CLK
                           , Q => n_2471, QN => 
                           DataPath_RF_bus_reg_dataout_762_port);
   DataPath_RF_BLOCKi_31_Q_reg_25_inst : DFF_X1 port map( D => n4363, CK => CLK
                           , Q => n_2472, QN => 
                           DataPath_RF_bus_reg_dataout_761_port);
   DataPath_RF_BLOCKi_31_Q_reg_24_inst : DFF_X1 port map( D => n4364, CK => CLK
                           , Q => n_2473, QN => 
                           DataPath_RF_bus_reg_dataout_760_port);
   DataPath_RF_BLOCKi_31_Q_reg_23_inst : DFF_X1 port map( D => n4365, CK => CLK
                           , Q => n_2474, QN => 
                           DataPath_RF_bus_reg_dataout_759_port);
   DataPath_RF_BLOCKi_31_Q_reg_22_inst : DFF_X1 port map( D => n4366, CK => CLK
                           , Q => n_2475, QN => 
                           DataPath_RF_bus_reg_dataout_758_port);
   DataPath_RF_BLOCKi_31_Q_reg_21_inst : DFF_X1 port map( D => n4367, CK => CLK
                           , Q => n_2476, QN => 
                           DataPath_RF_bus_reg_dataout_757_port);
   DataPath_RF_BLOCKi_31_Q_reg_20_inst : DFF_X1 port map( D => n4368, CK => CLK
                           , Q => n_2477, QN => 
                           DataPath_RF_bus_reg_dataout_756_port);
   DataPath_RF_BLOCKi_31_Q_reg_19_inst : DFF_X1 port map( D => n4369, CK => CLK
                           , Q => n_2478, QN => 
                           DataPath_RF_bus_reg_dataout_755_port);
   DataPath_RF_BLOCKi_31_Q_reg_18_inst : DFF_X1 port map( D => n4370, CK => CLK
                           , Q => n_2479, QN => 
                           DataPath_RF_bus_reg_dataout_754_port);
   DataPath_RF_BLOCKi_31_Q_reg_17_inst : DFF_X1 port map( D => n4371, CK => CLK
                           , Q => n_2480, QN => 
                           DataPath_RF_bus_reg_dataout_753_port);
   DataPath_RF_BLOCKi_31_Q_reg_16_inst : DFF_X1 port map( D => n4372, CK => CLK
                           , Q => n_2481, QN => 
                           DataPath_RF_bus_reg_dataout_752_port);
   DataPath_RF_BLOCKi_31_Q_reg_15_inst : DFF_X1 port map( D => n4373, CK => CLK
                           , Q => n_2482, QN => 
                           DataPath_RF_bus_reg_dataout_751_port);
   DataPath_RF_BLOCKi_31_Q_reg_14_inst : DFF_X1 port map( D => n4374, CK => CLK
                           , Q => n_2483, QN => 
                           DataPath_RF_bus_reg_dataout_750_port);
   DataPath_RF_BLOCKi_31_Q_reg_13_inst : DFF_X1 port map( D => n4375, CK => CLK
                           , Q => n_2484, QN => 
                           DataPath_RF_bus_reg_dataout_749_port);
   DataPath_RF_BLOCKi_31_Q_reg_12_inst : DFF_X1 port map( D => n4376, CK => CLK
                           , Q => n_2485, QN => 
                           DataPath_RF_bus_reg_dataout_748_port);
   DataPath_RF_BLOCKi_31_Q_reg_11_inst : DFF_X1 port map( D => n4377, CK => CLK
                           , Q => n_2486, QN => 
                           DataPath_RF_bus_reg_dataout_747_port);
   DataPath_RF_BLOCKi_31_Q_reg_9_inst : DFF_X1 port map( D => n4379, CK => CLK,
                           Q => n_2487, QN => 
                           DataPath_RF_bus_reg_dataout_745_port);
   DataPath_RF_BLOCKi_31_Q_reg_8_inst : DFF_X1 port map( D => n4380, CK => CLK,
                           Q => n_2488, QN => 
                           DataPath_RF_bus_reg_dataout_744_port);
   DataPath_RF_BLOCKi_31_Q_reg_7_inst : DFF_X1 port map( D => n4381, CK => CLK,
                           Q => n_2489, QN => 
                           DataPath_RF_bus_reg_dataout_743_port);
   DataPath_RF_BLOCKi_31_Q_reg_6_inst : DFF_X1 port map( D => n4382, CK => CLK,
                           Q => n_2490, QN => 
                           DataPath_RF_bus_reg_dataout_742_port);
   DataPath_RF_BLOCKi_31_Q_reg_5_inst : DFF_X1 port map( D => n4383, CK => CLK,
                           Q => n_2491, QN => 
                           DataPath_RF_bus_reg_dataout_741_port);
   DataPath_RF_BLOCKi_31_Q_reg_4_inst : DFF_X1 port map( D => n4384, CK => CLK,
                           Q => n_2492, QN => 
                           DataPath_RF_bus_reg_dataout_740_port);
   DataPath_RF_BLOCKi_31_Q_reg_3_inst : DFF_X1 port map( D => n4385, CK => CLK,
                           Q => n_2493, QN => 
                           DataPath_RF_bus_reg_dataout_739_port);
   DataPath_RF_BLOCKi_31_Q_reg_2_inst : DFF_X1 port map( D => n4386, CK => CLK,
                           Q => n_2494, QN => 
                           DataPath_RF_bus_reg_dataout_738_port);
   DataPath_RF_BLOCKi_31_Q_reg_1_inst : DFF_X1 port map( D => n4387, CK => CLK,
                           Q => n_2495, QN => 
                           DataPath_RF_bus_reg_dataout_737_port);
   DataPath_RF_BLOCKi_31_Q_reg_0_inst : DFF_X1 port map( D => n4388, CK => CLK,
                           Q => n_2496, QN => 
                           DataPath_RF_bus_reg_dataout_736_port);
   DataPath_RF_BLOCKi_47_Q_reg_31_inst : DFF_X1 port map( D => n4948, CK => CLK
                           , Q => n_2497, QN => 
                           DataPath_RF_bus_reg_dataout_1279_port);
   DataPath_RF_BLOCKi_47_Q_reg_30_inst : DFF_X1 port map( D => n4951, CK => CLK
                           , Q => n_2498, QN => 
                           DataPath_RF_bus_reg_dataout_1278_port);
   DataPath_RF_BLOCKi_47_Q_reg_29_inst : DFF_X1 port map( D => n4952, CK => CLK
                           , Q => n_2499, QN => 
                           DataPath_RF_bus_reg_dataout_1277_port);
   DataPath_RF_BLOCKi_47_Q_reg_28_inst : DFF_X1 port map( D => n4953, CK => CLK
                           , Q => n_2500, QN => 
                           DataPath_RF_bus_reg_dataout_1276_port);
   DataPath_RF_BLOCKi_47_Q_reg_27_inst : DFF_X1 port map( D => n4954, CK => CLK
                           , Q => n_2501, QN => 
                           DataPath_RF_bus_reg_dataout_1275_port);
   DataPath_RF_BLOCKi_47_Q_reg_26_inst : DFF_X1 port map( D => n4955, CK => CLK
                           , Q => n_2502, QN => 
                           DataPath_RF_bus_reg_dataout_1274_port);
   DataPath_RF_BLOCKi_47_Q_reg_25_inst : DFF_X1 port map( D => n4956, CK => CLK
                           , Q => n_2503, QN => 
                           DataPath_RF_bus_reg_dataout_1273_port);
   DataPath_RF_BLOCKi_47_Q_reg_24_inst : DFF_X1 port map( D => n4957, CK => CLK
                           , Q => n_2504, QN => 
                           DataPath_RF_bus_reg_dataout_1272_port);
   DataPath_RF_BLOCKi_47_Q_reg_23_inst : DFF_X1 port map( D => n4958, CK => CLK
                           , Q => n_2505, QN => 
                           DataPath_RF_bus_reg_dataout_1271_port);
   DataPath_RF_BLOCKi_47_Q_reg_22_inst : DFF_X1 port map( D => n4959, CK => CLK
                           , Q => n_2506, QN => 
                           DataPath_RF_bus_reg_dataout_1270_port);
   DataPath_RF_BLOCKi_47_Q_reg_21_inst : DFF_X1 port map( D => n4960, CK => CLK
                           , Q => n_2507, QN => 
                           DataPath_RF_bus_reg_dataout_1269_port);
   DataPath_RF_BLOCKi_47_Q_reg_20_inst : DFF_X1 port map( D => n4961, CK => CLK
                           , Q => n_2508, QN => 
                           DataPath_RF_bus_reg_dataout_1268_port);
   DataPath_RF_BLOCKi_47_Q_reg_19_inst : DFF_X1 port map( D => n4962, CK => CLK
                           , Q => n_2509, QN => 
                           DataPath_RF_bus_reg_dataout_1267_port);
   DataPath_RF_BLOCKi_47_Q_reg_18_inst : DFF_X1 port map( D => n4963, CK => CLK
                           , Q => n_2510, QN => 
                           DataPath_RF_bus_reg_dataout_1266_port);
   DataPath_RF_BLOCKi_47_Q_reg_17_inst : DFF_X1 port map( D => n4964, CK => CLK
                           , Q => n_2511, QN => 
                           DataPath_RF_bus_reg_dataout_1265_port);
   DataPath_RF_BLOCKi_47_Q_reg_16_inst : DFF_X1 port map( D => n4965, CK => CLK
                           , Q => n_2512, QN => 
                           DataPath_RF_bus_reg_dataout_1264_port);
   DataPath_RF_BLOCKi_47_Q_reg_15_inst : DFF_X1 port map( D => n4966, CK => CLK
                           , Q => n_2513, QN => 
                           DataPath_RF_bus_reg_dataout_1263_port);
   DataPath_RF_BLOCKi_47_Q_reg_14_inst : DFF_X1 port map( D => n4967, CK => CLK
                           , Q => n_2514, QN => 
                           DataPath_RF_bus_reg_dataout_1262_port);
   DataPath_RF_BLOCKi_47_Q_reg_13_inst : DFF_X1 port map( D => n4968, CK => CLK
                           , Q => n_2515, QN => 
                           DataPath_RF_bus_reg_dataout_1261_port);
   DataPath_RF_BLOCKi_47_Q_reg_12_inst : DFF_X1 port map( D => n4969, CK => CLK
                           , Q => n_2516, QN => 
                           DataPath_RF_bus_reg_dataout_1260_port);
   DataPath_RF_BLOCKi_47_Q_reg_11_inst : DFF_X1 port map( D => n4970, CK => CLK
                           , Q => n_2517, QN => 
                           DataPath_RF_bus_reg_dataout_1259_port);
   DataPath_RF_BLOCKi_47_Q_reg_9_inst : DFF_X1 port map( D => n4972, CK => CLK,
                           Q => n_2518, QN => 
                           DataPath_RF_bus_reg_dataout_1257_port);
   DataPath_RF_BLOCKi_47_Q_reg_8_inst : DFF_X1 port map( D => n4973, CK => CLK,
                           Q => n_2519, QN => 
                           DataPath_RF_bus_reg_dataout_1256_port);
   DataPath_RF_BLOCKi_47_Q_reg_7_inst : DFF_X1 port map( D => n4974, CK => CLK,
                           Q => n_2520, QN => 
                           DataPath_RF_bus_reg_dataout_1255_port);
   DataPath_RF_BLOCKi_47_Q_reg_6_inst : DFF_X1 port map( D => n4975, CK => CLK,
                           Q => n_2521, QN => 
                           DataPath_RF_bus_reg_dataout_1254_port);
   DataPath_RF_BLOCKi_47_Q_reg_5_inst : DFF_X1 port map( D => n4976, CK => CLK,
                           Q => n_2522, QN => 
                           DataPath_RF_bus_reg_dataout_1253_port);
   DataPath_RF_BLOCKi_47_Q_reg_4_inst : DFF_X1 port map( D => n4977, CK => CLK,
                           Q => n_2523, QN => 
                           DataPath_RF_bus_reg_dataout_1252_port);
   DataPath_RF_BLOCKi_47_Q_reg_3_inst : DFF_X1 port map( D => n4978, CK => CLK,
                           Q => n_2524, QN => 
                           DataPath_RF_bus_reg_dataout_1251_port);
   DataPath_RF_BLOCKi_47_Q_reg_2_inst : DFF_X1 port map( D => n4979, CK => CLK,
                           Q => n_2525, QN => 
                           DataPath_RF_bus_reg_dataout_1250_port);
   DataPath_RF_BLOCKi_47_Q_reg_1_inst : DFF_X1 port map( D => n4980, CK => CLK,
                           Q => n_2526, QN => 
                           DataPath_RF_bus_reg_dataout_1249_port);
   DataPath_RF_BLOCKi_47_Q_reg_0_inst : DFF_X1 port map( D => n4981, CK => CLK,
                           Q => n_2527, QN => 
                           DataPath_RF_bus_reg_dataout_1248_port);
   DataPath_RF_BLOCKi_63_Q_reg_31_inst : DFF_X1 port map( D => n5541, CK => CLK
                           , Q => n_2528, QN => 
                           DataPath_RF_bus_reg_dataout_1791_port);
   DataPath_RF_BLOCKi_63_Q_reg_30_inst : DFF_X1 port map( D => n5544, CK => CLK
                           , Q => n_2529, QN => 
                           DataPath_RF_bus_reg_dataout_1790_port);
   DataPath_RF_BLOCKi_63_Q_reg_29_inst : DFF_X1 port map( D => n5545, CK => CLK
                           , Q => n_2530, QN => 
                           DataPath_RF_bus_reg_dataout_1789_port);
   DataPath_RF_BLOCKi_63_Q_reg_28_inst : DFF_X1 port map( D => n5546, CK => CLK
                           , Q => n_2531, QN => 
                           DataPath_RF_bus_reg_dataout_1788_port);
   DataPath_RF_BLOCKi_63_Q_reg_27_inst : DFF_X1 port map( D => n5547, CK => CLK
                           , Q => n_2532, QN => 
                           DataPath_RF_bus_reg_dataout_1787_port);
   DataPath_RF_BLOCKi_63_Q_reg_26_inst : DFF_X1 port map( D => n5548, CK => CLK
                           , Q => n_2533, QN => 
                           DataPath_RF_bus_reg_dataout_1786_port);
   DataPath_RF_BLOCKi_63_Q_reg_25_inst : DFF_X1 port map( D => n5549, CK => CLK
                           , Q => n_2534, QN => 
                           DataPath_RF_bus_reg_dataout_1785_port);
   DataPath_RF_BLOCKi_63_Q_reg_24_inst : DFF_X1 port map( D => n5550, CK => CLK
                           , Q => n_2535, QN => 
                           DataPath_RF_bus_reg_dataout_1784_port);
   DataPath_RF_BLOCKi_63_Q_reg_23_inst : DFF_X1 port map( D => n5551, CK => CLK
                           , Q => n_2536, QN => 
                           DataPath_RF_bus_reg_dataout_1783_port);
   DataPath_RF_BLOCKi_63_Q_reg_22_inst : DFF_X1 port map( D => n5552, CK => CLK
                           , Q => n_2537, QN => 
                           DataPath_RF_bus_reg_dataout_1782_port);
   DataPath_RF_BLOCKi_63_Q_reg_21_inst : DFF_X1 port map( D => n5553, CK => CLK
                           , Q => n_2538, QN => 
                           DataPath_RF_bus_reg_dataout_1781_port);
   DataPath_RF_BLOCKi_63_Q_reg_20_inst : DFF_X1 port map( D => n5554, CK => CLK
                           , Q => n_2539, QN => 
                           DataPath_RF_bus_reg_dataout_1780_port);
   DataPath_RF_BLOCKi_63_Q_reg_19_inst : DFF_X1 port map( D => n5555, CK => CLK
                           , Q => n_2540, QN => 
                           DataPath_RF_bus_reg_dataout_1779_port);
   DataPath_RF_BLOCKi_63_Q_reg_18_inst : DFF_X1 port map( D => n5556, CK => CLK
                           , Q => n_2541, QN => 
                           DataPath_RF_bus_reg_dataout_1778_port);
   DataPath_RF_BLOCKi_63_Q_reg_17_inst : DFF_X1 port map( D => n5557, CK => CLK
                           , Q => n_2542, QN => 
                           DataPath_RF_bus_reg_dataout_1777_port);
   DataPath_RF_BLOCKi_63_Q_reg_16_inst : DFF_X1 port map( D => n5558, CK => CLK
                           , Q => n_2543, QN => 
                           DataPath_RF_bus_reg_dataout_1776_port);
   DataPath_RF_BLOCKi_63_Q_reg_15_inst : DFF_X1 port map( D => n5559, CK => CLK
                           , Q => n_2544, QN => 
                           DataPath_RF_bus_reg_dataout_1775_port);
   DataPath_RF_BLOCKi_63_Q_reg_14_inst : DFF_X1 port map( D => n5560, CK => CLK
                           , Q => n_2545, QN => 
                           DataPath_RF_bus_reg_dataout_1774_port);
   DataPath_RF_BLOCKi_63_Q_reg_13_inst : DFF_X1 port map( D => n5561, CK => CLK
                           , Q => n_2546, QN => 
                           DataPath_RF_bus_reg_dataout_1773_port);
   DataPath_RF_BLOCKi_63_Q_reg_12_inst : DFF_X1 port map( D => n5562, CK => CLK
                           , Q => n_2547, QN => 
                           DataPath_RF_bus_reg_dataout_1772_port);
   DataPath_RF_BLOCKi_63_Q_reg_11_inst : DFF_X1 port map( D => n5563, CK => CLK
                           , Q => n_2548, QN => 
                           DataPath_RF_bus_reg_dataout_1771_port);
   DataPath_RF_BLOCKi_63_Q_reg_9_inst : DFF_X1 port map( D => n5565, CK => CLK,
                           Q => n_2549, QN => 
                           DataPath_RF_bus_reg_dataout_1769_port);
   DataPath_RF_BLOCKi_63_Q_reg_8_inst : DFF_X1 port map( D => n5566, CK => CLK,
                           Q => n_2550, QN => 
                           DataPath_RF_bus_reg_dataout_1768_port);
   DataPath_RF_BLOCKi_63_Q_reg_7_inst : DFF_X1 port map( D => n5567, CK => CLK,
                           Q => n_2551, QN => 
                           DataPath_RF_bus_reg_dataout_1767_port);
   DataPath_RF_BLOCKi_63_Q_reg_6_inst : DFF_X1 port map( D => n5568, CK => CLK,
                           Q => n_2552, QN => 
                           DataPath_RF_bus_reg_dataout_1766_port);
   DataPath_RF_BLOCKi_63_Q_reg_5_inst : DFF_X1 port map( D => n5569, CK => CLK,
                           Q => n_2553, QN => 
                           DataPath_RF_bus_reg_dataout_1765_port);
   DataPath_RF_BLOCKi_63_Q_reg_4_inst : DFF_X1 port map( D => n5570, CK => CLK,
                           Q => n_2554, QN => 
                           DataPath_RF_bus_reg_dataout_1764_port);
   DataPath_RF_BLOCKi_63_Q_reg_3_inst : DFF_X1 port map( D => n5571, CK => CLK,
                           Q => n_2555, QN => 
                           DataPath_RF_bus_reg_dataout_1763_port);
   DataPath_RF_BLOCKi_63_Q_reg_2_inst : DFF_X1 port map( D => n5572, CK => CLK,
                           Q => n_2556, QN => 
                           DataPath_RF_bus_reg_dataout_1762_port);
   DataPath_RF_BLOCKi_63_Q_reg_1_inst : DFF_X1 port map( D => n5573, CK => CLK,
                           Q => n_2557, QN => 
                           DataPath_RF_bus_reg_dataout_1761_port);
   DataPath_RF_BLOCKi_63_Q_reg_0_inst : DFF_X1 port map( D => n5574, CK => CLK,
                           Q => n_2558, QN => 
                           DataPath_RF_bus_reg_dataout_1760_port);
   DataPath_RF_BLOCKi_79_Q_reg_15_inst : DFF_X1 port map( D => n879, CK => CLK,
                           Q => n_2559, QN => 
                           DataPath_RF_bus_reg_dataout_2287_port);
   DataPath_RF_BLOCKi_79_Q_reg_14_inst : DFF_X1 port map( D => n883, CK => CLK,
                           Q => n_2560, QN => 
                           DataPath_RF_bus_reg_dataout_2286_port);
   DataPath_RF_BLOCKi_79_Q_reg_13_inst : DFF_X1 port map( D => n885, CK => CLK,
                           Q => n_2561, QN => 
                           DataPath_RF_bus_reg_dataout_2285_port);
   DataPath_RF_BLOCKi_79_Q_reg_12_inst : DFF_X1 port map( D => n887, CK => CLK,
                           Q => n_2562, QN => 
                           DataPath_RF_bus_reg_dataout_2284_port);
   DataPath_RF_BLOCKi_79_Q_reg_11_inst : DFF_X1 port map( D => n889, CK => CLK,
                           Q => n_2563, QN => 
                           DataPath_RF_bus_reg_dataout_2283_port);
   DataPath_RF_BLOCKi_79_Q_reg_9_inst : DFF_X1 port map( D => n893, CK => CLK, 
                           Q => n_2564, QN => 
                           DataPath_RF_bus_reg_dataout_2281_port);
   DataPath_RF_BLOCKi_79_Q_reg_8_inst : DFF_X1 port map( D => n895, CK => CLK, 
                           Q => n_2565, QN => 
                           DataPath_RF_bus_reg_dataout_2280_port);
   DataPath_RF_BLOCKi_79_Q_reg_7_inst : DFF_X1 port map( D => n897, CK => CLK, 
                           Q => n_2566, QN => 
                           DataPath_RF_bus_reg_dataout_2279_port);
   DataPath_RF_BLOCKi_79_Q_reg_6_inst : DFF_X1 port map( D => n899, CK => CLK, 
                           Q => n_2567, QN => 
                           DataPath_RF_bus_reg_dataout_2278_port);
   DataPath_RF_BLOCKi_79_Q_reg_5_inst : DFF_X1 port map( D => n901, CK => CLK, 
                           Q => n_2568, QN => 
                           DataPath_RF_bus_reg_dataout_2277_port);
   DataPath_RF_BLOCKi_79_Q_reg_4_inst : DFF_X1 port map( D => n903, CK => CLK, 
                           Q => n_2569, QN => 
                           DataPath_RF_bus_reg_dataout_2276_port);
   DataPath_RF_BLOCKi_79_Q_reg_3_inst : DFF_X1 port map( D => n905, CK => CLK, 
                           Q => n_2570, QN => 
                           DataPath_RF_bus_reg_dataout_2275_port);
   DataPath_RF_BLOCKi_79_Q_reg_2_inst : DFF_X1 port map( D => n907, CK => CLK, 
                           Q => n_2571, QN => 
                           DataPath_RF_bus_reg_dataout_2274_port);
   DataPath_RF_BLOCKi_79_Q_reg_1_inst : DFF_X1 port map( D => n909, CK => CLK, 
                           Q => n_2572, QN => 
                           DataPath_RF_bus_reg_dataout_2273_port);
   DataPath_RF_BLOCKi_79_Q_reg_0_inst : DFF_X1 port map( D => n911, CK => CLK, 
                           Q => n_2573, QN => 
                           DataPath_RF_bus_reg_dataout_2272_port);
   DataPath_RF_BLOCKi_79_Q_reg_31_inst : DFF_X1 port map( D => n6127, CK => CLK
                           , Q => n_2574, QN => 
                           DataPath_RF_bus_reg_dataout_2303_port);
   DataPath_RF_BLOCKi_79_Q_reg_30_inst : DFF_X1 port map( D => n6128, CK => CLK
                           , Q => n_2575, QN => 
                           DataPath_RF_bus_reg_dataout_2302_port);
   DataPath_RF_BLOCKi_79_Q_reg_29_inst : DFF_X1 port map( D => n6129, CK => CLK
                           , Q => n_2576, QN => 
                           DataPath_RF_bus_reg_dataout_2301_port);
   DataPath_RF_BLOCKi_79_Q_reg_28_inst : DFF_X1 port map( D => n6130, CK => CLK
                           , Q => n_2577, QN => 
                           DataPath_RF_bus_reg_dataout_2300_port);
   DataPath_RF_BLOCKi_79_Q_reg_27_inst : DFF_X1 port map( D => n6131, CK => CLK
                           , Q => n_2578, QN => 
                           DataPath_RF_bus_reg_dataout_2299_port);
   DataPath_RF_BLOCKi_79_Q_reg_26_inst : DFF_X1 port map( D => n6132, CK => CLK
                           , Q => n_2579, QN => 
                           DataPath_RF_bus_reg_dataout_2298_port);
   DataPath_RF_BLOCKi_79_Q_reg_25_inst : DFF_X1 port map( D => n6133, CK => CLK
                           , Q => n_2580, QN => 
                           DataPath_RF_bus_reg_dataout_2297_port);
   DataPath_RF_BLOCKi_79_Q_reg_24_inst : DFF_X1 port map( D => n6134, CK => CLK
                           , Q => n_2581, QN => 
                           DataPath_RF_bus_reg_dataout_2296_port);
   DataPath_RF_BLOCKi_79_Q_reg_23_inst : DFF_X1 port map( D => n6135, CK => CLK
                           , Q => n_2582, QN => 
                           DataPath_RF_bus_reg_dataout_2295_port);
   DataPath_RF_BLOCKi_79_Q_reg_22_inst : DFF_X1 port map( D => n6136, CK => CLK
                           , Q => n_2583, QN => 
                           DataPath_RF_bus_reg_dataout_2294_port);
   DataPath_RF_BLOCKi_79_Q_reg_21_inst : DFF_X1 port map( D => n6137, CK => CLK
                           , Q => n_2584, QN => 
                           DataPath_RF_bus_reg_dataout_2293_port);
   DataPath_RF_BLOCKi_79_Q_reg_20_inst : DFF_X1 port map( D => n6138, CK => CLK
                           , Q => n_2585, QN => 
                           DataPath_RF_bus_reg_dataout_2292_port);
   DataPath_RF_BLOCKi_79_Q_reg_19_inst : DFF_X1 port map( D => n6139, CK => CLK
                           , Q => n_2586, QN => 
                           DataPath_RF_bus_reg_dataout_2291_port);
   DataPath_RF_BLOCKi_79_Q_reg_18_inst : DFF_X1 port map( D => n6140, CK => CLK
                           , Q => n_2587, QN => 
                           DataPath_RF_bus_reg_dataout_2290_port);
   DataPath_RF_BLOCKi_79_Q_reg_17_inst : DFF_X1 port map( D => n6141, CK => CLK
                           , Q => n_2588, QN => 
                           DataPath_RF_bus_reg_dataout_2289_port);
   DataPath_RF_BLOCKi_79_Q_reg_16_inst : DFF_X1 port map( D => n6142, CK => CLK
                           , Q => n_2589, QN => 
                           DataPath_RF_bus_reg_dataout_2288_port);
   DataPath_RF_BLOCKi_81_Q_reg_31_inst : DFF_X1 port map( D => n966, CK => CLK,
                           Q => n_2590, QN => 
                           DataPath_RF_bus_reg_dataout_2367_port);
   DataPath_RF_BLOCKi_81_Q_reg_30_inst : DFF_X1 port map( D => n969, CK => CLK,
                           Q => n_2591, QN => 
                           DataPath_RF_bus_reg_dataout_2366_port);
   DataPath_RF_BLOCKi_81_Q_reg_29_inst : DFF_X1 port map( D => n970, CK => CLK,
                           Q => n_2592, QN => 
                           DataPath_RF_bus_reg_dataout_2365_port);
   DataPath_RF_BLOCKi_81_Q_reg_28_inst : DFF_X1 port map( D => n971, CK => CLK,
                           Q => n_2593, QN => 
                           DataPath_RF_bus_reg_dataout_2364_port);
   DataPath_RF_BLOCKi_81_Q_reg_27_inst : DFF_X1 port map( D => n972, CK => CLK,
                           Q => n_2594, QN => 
                           DataPath_RF_bus_reg_dataout_2363_port);
   DataPath_RF_BLOCKi_81_Q_reg_26_inst : DFF_X1 port map( D => n973, CK => CLK,
                           Q => n_2595, QN => 
                           DataPath_RF_bus_reg_dataout_2362_port);
   DataPath_RF_BLOCKi_81_Q_reg_25_inst : DFF_X1 port map( D => n974, CK => CLK,
                           Q => n_2596, QN => 
                           DataPath_RF_bus_reg_dataout_2361_port);
   DataPath_RF_BLOCKi_81_Q_reg_24_inst : DFF_X1 port map( D => n975, CK => CLK,
                           Q => n_2597, QN => 
                           DataPath_RF_bus_reg_dataout_2360_port);
   DataPath_RF_BLOCKi_81_Q_reg_23_inst : DFF_X1 port map( D => n976, CK => CLK,
                           Q => n_2598, QN => 
                           DataPath_RF_bus_reg_dataout_2359_port);
   DataPath_RF_BLOCKi_81_Q_reg_22_inst : DFF_X1 port map( D => n977, CK => CLK,
                           Q => n_2599, QN => 
                           DataPath_RF_bus_reg_dataout_2358_port);
   DataPath_RF_BLOCKi_81_Q_reg_21_inst : DFF_X1 port map( D => n978, CK => CLK,
                           Q => n_2600, QN => 
                           DataPath_RF_bus_reg_dataout_2357_port);
   DataPath_RF_BLOCKi_81_Q_reg_20_inst : DFF_X1 port map( D => n979, CK => CLK,
                           Q => n_2601, QN => 
                           DataPath_RF_bus_reg_dataout_2356_port);
   DataPath_RF_BLOCKi_81_Q_reg_19_inst : DFF_X1 port map( D => n980, CK => CLK,
                           Q => n_2602, QN => 
                           DataPath_RF_bus_reg_dataout_2355_port);
   DataPath_RF_BLOCKi_81_Q_reg_18_inst : DFF_X1 port map( D => n981, CK => CLK,
                           Q => n_2603, QN => 
                           DataPath_RF_bus_reg_dataout_2354_port);
   DataPath_RF_BLOCKi_81_Q_reg_17_inst : DFF_X1 port map( D => n982, CK => CLK,
                           Q => n_2604, QN => 
                           DataPath_RF_bus_reg_dataout_2353_port);
   DataPath_RF_BLOCKi_81_Q_reg_16_inst : DFF_X1 port map( D => n983, CK => CLK,
                           Q => n_2605, QN => 
                           DataPath_RF_bus_reg_dataout_2352_port);
   DataPath_RF_BLOCKi_81_Q_reg_15_inst : DFF_X1 port map( D => n984, CK => CLK,
                           Q => n_2606, QN => 
                           DataPath_RF_bus_reg_dataout_2351_port);
   DataPath_RF_BLOCKi_81_Q_reg_14_inst : DFF_X1 port map( D => n985, CK => CLK,
                           Q => n_2607, QN => 
                           DataPath_RF_bus_reg_dataout_2350_port);
   DataPath_RF_BLOCKi_81_Q_reg_13_inst : DFF_X1 port map( D => n986, CK => CLK,
                           Q => n_2608, QN => 
                           DataPath_RF_bus_reg_dataout_2349_port);
   DataPath_RF_BLOCKi_81_Q_reg_12_inst : DFF_X1 port map( D => n987, CK => CLK,
                           Q => n_2609, QN => 
                           DataPath_RF_bus_reg_dataout_2348_port);
   DataPath_RF_BLOCKi_81_Q_reg_11_inst : DFF_X1 port map( D => n988, CK => CLK,
                           Q => n_2610, QN => 
                           DataPath_RF_bus_reg_dataout_2347_port);
   DataPath_RF_BLOCKi_81_Q_reg_9_inst : DFF_X1 port map( D => n990, CK => CLK, 
                           Q => n_2611, QN => 
                           DataPath_RF_bus_reg_dataout_2345_port);
   DataPath_RF_BLOCKi_81_Q_reg_8_inst : DFF_X1 port map( D => n991, CK => CLK, 
                           Q => n_2612, QN => 
                           DataPath_RF_bus_reg_dataout_2344_port);
   DataPath_RF_BLOCKi_81_Q_reg_7_inst : DFF_X1 port map( D => n992, CK => CLK, 
                           Q => n_2613, QN => 
                           DataPath_RF_bus_reg_dataout_2343_port);
   DataPath_RF_BLOCKi_81_Q_reg_6_inst : DFF_X1 port map( D => n993, CK => CLK, 
                           Q => n_2614, QN => 
                           DataPath_RF_bus_reg_dataout_2342_port);
   DataPath_RF_BLOCKi_81_Q_reg_5_inst : DFF_X1 port map( D => n994, CK => CLK, 
                           Q => n_2615, QN => 
                           DataPath_RF_bus_reg_dataout_2341_port);
   DataPath_RF_BLOCKi_81_Q_reg_4_inst : DFF_X1 port map( D => n995, CK => CLK, 
                           Q => n_2616, QN => 
                           DataPath_RF_bus_reg_dataout_2340_port);
   DataPath_RF_BLOCKi_81_Q_reg_3_inst : DFF_X1 port map( D => n996, CK => CLK, 
                           Q => n_2617, QN => 
                           DataPath_RF_bus_reg_dataout_2339_port);
   DataPath_RF_BLOCKi_81_Q_reg_2_inst : DFF_X1 port map( D => n997, CK => CLK, 
                           Q => n_2618, QN => 
                           DataPath_RF_bus_reg_dataout_2338_port);
   DataPath_RF_BLOCKi_81_Q_reg_1_inst : DFF_X1 port map( D => n998, CK => CLK, 
                           Q => n_2619, QN => 
                           DataPath_RF_bus_reg_dataout_2337_port);
   DataPath_RF_BLOCKi_81_Q_reg_0_inst : DFF_X1 port map( D => n999, CK => CLK, 
                           Q => n_2620, QN => 
                           DataPath_RF_bus_reg_dataout_2336_port);
   DataPath_RF_BLOCKi_17_Q_reg_31_inst : DFF_X1 port map( D => n3800, CK => CLK
                           , Q => n_2621, QN => 
                           DataPath_RF_bus_reg_dataout_319_port);
   DataPath_RF_BLOCKi_17_Q_reg_30_inst : DFF_X1 port map( D => n3803, CK => CLK
                           , Q => n_2622, QN => 
                           DataPath_RF_bus_reg_dataout_318_port);
   DataPath_RF_BLOCKi_17_Q_reg_29_inst : DFF_X1 port map( D => n3804, CK => CLK
                           , Q => n_2623, QN => 
                           DataPath_RF_bus_reg_dataout_317_port);
   DataPath_RF_BLOCKi_17_Q_reg_28_inst : DFF_X1 port map( D => n3805, CK => CLK
                           , Q => n_2624, QN => 
                           DataPath_RF_bus_reg_dataout_316_port);
   DataPath_RF_BLOCKi_17_Q_reg_27_inst : DFF_X1 port map( D => n3806, CK => CLK
                           , Q => n_2625, QN => 
                           DataPath_RF_bus_reg_dataout_315_port);
   DataPath_RF_BLOCKi_17_Q_reg_26_inst : DFF_X1 port map( D => n3807, CK => CLK
                           , Q => n_2626, QN => 
                           DataPath_RF_bus_reg_dataout_314_port);
   DataPath_RF_BLOCKi_17_Q_reg_25_inst : DFF_X1 port map( D => n3808, CK => CLK
                           , Q => n_2627, QN => 
                           DataPath_RF_bus_reg_dataout_313_port);
   DataPath_RF_BLOCKi_17_Q_reg_24_inst : DFF_X1 port map( D => n3809, CK => CLK
                           , Q => n_2628, QN => 
                           DataPath_RF_bus_reg_dataout_312_port);
   DataPath_RF_BLOCKi_17_Q_reg_23_inst : DFF_X1 port map( D => n3810, CK => CLK
                           , Q => n_2629, QN => 
                           DataPath_RF_bus_reg_dataout_311_port);
   DataPath_RF_BLOCKi_17_Q_reg_22_inst : DFF_X1 port map( D => n3811, CK => CLK
                           , Q => n_2630, QN => 
                           DataPath_RF_bus_reg_dataout_310_port);
   DataPath_RF_BLOCKi_17_Q_reg_21_inst : DFF_X1 port map( D => n3812, CK => CLK
                           , Q => n_2631, QN => 
                           DataPath_RF_bus_reg_dataout_309_port);
   DataPath_RF_BLOCKi_17_Q_reg_20_inst : DFF_X1 port map( D => n3813, CK => CLK
                           , Q => n_2632, QN => 
                           DataPath_RF_bus_reg_dataout_308_port);
   DataPath_RF_BLOCKi_17_Q_reg_19_inst : DFF_X1 port map( D => n3814, CK => CLK
                           , Q => n_2633, QN => 
                           DataPath_RF_bus_reg_dataout_307_port);
   DataPath_RF_BLOCKi_17_Q_reg_18_inst : DFF_X1 port map( D => n3815, CK => CLK
                           , Q => n_2634, QN => 
                           DataPath_RF_bus_reg_dataout_306_port);
   DataPath_RF_BLOCKi_17_Q_reg_17_inst : DFF_X1 port map( D => n3816, CK => CLK
                           , Q => n_2635, QN => 
                           DataPath_RF_bus_reg_dataout_305_port);
   DataPath_RF_BLOCKi_17_Q_reg_16_inst : DFF_X1 port map( D => n3817, CK => CLK
                           , Q => n_2636, QN => 
                           DataPath_RF_bus_reg_dataout_304_port);
   DataPath_RF_BLOCKi_17_Q_reg_15_inst : DFF_X1 port map( D => n3818, CK => CLK
                           , Q => n_2637, QN => 
                           DataPath_RF_bus_reg_dataout_303_port);
   DataPath_RF_BLOCKi_17_Q_reg_14_inst : DFF_X1 port map( D => n3819, CK => CLK
                           , Q => n_2638, QN => 
                           DataPath_RF_bus_reg_dataout_302_port);
   DataPath_RF_BLOCKi_17_Q_reg_13_inst : DFF_X1 port map( D => n3820, CK => CLK
                           , Q => n_2639, QN => 
                           DataPath_RF_bus_reg_dataout_301_port);
   DataPath_RF_BLOCKi_17_Q_reg_12_inst : DFF_X1 port map( D => n3821, CK => CLK
                           , Q => n_2640, QN => 
                           DataPath_RF_bus_reg_dataout_300_port);
   DataPath_RF_BLOCKi_17_Q_reg_11_inst : DFF_X1 port map( D => n3822, CK => CLK
                           , Q => n_2641, QN => 
                           DataPath_RF_bus_reg_dataout_299_port);
   DataPath_RF_BLOCKi_17_Q_reg_9_inst : DFF_X1 port map( D => n3824, CK => CLK,
                           Q => n_2642, QN => 
                           DataPath_RF_bus_reg_dataout_297_port);
   DataPath_RF_BLOCKi_17_Q_reg_8_inst : DFF_X1 port map( D => n3825, CK => CLK,
                           Q => n_2643, QN => 
                           DataPath_RF_bus_reg_dataout_296_port);
   DataPath_RF_BLOCKi_17_Q_reg_7_inst : DFF_X1 port map( D => n3826, CK => CLK,
                           Q => n_2644, QN => 
                           DataPath_RF_bus_reg_dataout_295_port);
   DataPath_RF_BLOCKi_17_Q_reg_6_inst : DFF_X1 port map( D => n3827, CK => CLK,
                           Q => n_2645, QN => 
                           DataPath_RF_bus_reg_dataout_294_port);
   DataPath_RF_BLOCKi_17_Q_reg_5_inst : DFF_X1 port map( D => n3828, CK => CLK,
                           Q => n_2646, QN => 
                           DataPath_RF_bus_reg_dataout_293_port);
   DataPath_RF_BLOCKi_17_Q_reg_4_inst : DFF_X1 port map( D => n3829, CK => CLK,
                           Q => n_2647, QN => 
                           DataPath_RF_bus_reg_dataout_292_port);
   DataPath_RF_BLOCKi_17_Q_reg_3_inst : DFF_X1 port map( D => n3830, CK => CLK,
                           Q => n_2648, QN => 
                           DataPath_RF_bus_reg_dataout_291_port);
   DataPath_RF_BLOCKi_17_Q_reg_2_inst : DFF_X1 port map( D => n3831, CK => CLK,
                           Q => n_2649, QN => 
                           DataPath_RF_bus_reg_dataout_290_port);
   DataPath_RF_BLOCKi_17_Q_reg_1_inst : DFF_X1 port map( D => n3832, CK => CLK,
                           Q => n_2650, QN => 
                           DataPath_RF_bus_reg_dataout_289_port);
   DataPath_RF_BLOCKi_17_Q_reg_0_inst : DFF_X1 port map( D => n3833, CK => CLK,
                           Q => n_2651, QN => 
                           DataPath_RF_bus_reg_dataout_288_port);
   DataPath_RF_BLOCKi_33_Q_reg_31_inst : DFF_X1 port map( D => n4425, CK => CLK
                           , Q => n_2652, QN => 
                           DataPath_RF_bus_reg_dataout_831_port);
   DataPath_RF_BLOCKi_33_Q_reg_30_inst : DFF_X1 port map( D => n4428, CK => CLK
                           , Q => n_2653, QN => 
                           DataPath_RF_bus_reg_dataout_830_port);
   DataPath_RF_BLOCKi_33_Q_reg_29_inst : DFF_X1 port map( D => n4429, CK => CLK
                           , Q => n_2654, QN => 
                           DataPath_RF_bus_reg_dataout_829_port);
   DataPath_RF_BLOCKi_33_Q_reg_28_inst : DFF_X1 port map( D => n4430, CK => CLK
                           , Q => n_2655, QN => 
                           DataPath_RF_bus_reg_dataout_828_port);
   DataPath_RF_BLOCKi_33_Q_reg_27_inst : DFF_X1 port map( D => n4431, CK => CLK
                           , Q => n_2656, QN => 
                           DataPath_RF_bus_reg_dataout_827_port);
   DataPath_RF_BLOCKi_33_Q_reg_26_inst : DFF_X1 port map( D => n4432, CK => CLK
                           , Q => n_2657, QN => 
                           DataPath_RF_bus_reg_dataout_826_port);
   DataPath_RF_BLOCKi_33_Q_reg_25_inst : DFF_X1 port map( D => n4433, CK => CLK
                           , Q => n_2658, QN => 
                           DataPath_RF_bus_reg_dataout_825_port);
   DataPath_RF_BLOCKi_33_Q_reg_24_inst : DFF_X1 port map( D => n4434, CK => CLK
                           , Q => n_2659, QN => 
                           DataPath_RF_bus_reg_dataout_824_port);
   DataPath_RF_BLOCKi_33_Q_reg_23_inst : DFF_X1 port map( D => n4435, CK => CLK
                           , Q => n_2660, QN => 
                           DataPath_RF_bus_reg_dataout_823_port);
   DataPath_RF_BLOCKi_33_Q_reg_22_inst : DFF_X1 port map( D => n4436, CK => CLK
                           , Q => n_2661, QN => 
                           DataPath_RF_bus_reg_dataout_822_port);
   DataPath_RF_BLOCKi_33_Q_reg_21_inst : DFF_X1 port map( D => n4437, CK => CLK
                           , Q => n_2662, QN => 
                           DataPath_RF_bus_reg_dataout_821_port);
   DataPath_RF_BLOCKi_33_Q_reg_20_inst : DFF_X1 port map( D => n4438, CK => CLK
                           , Q => n_2663, QN => 
                           DataPath_RF_bus_reg_dataout_820_port);
   DataPath_RF_BLOCKi_33_Q_reg_19_inst : DFF_X1 port map( D => n4439, CK => CLK
                           , Q => n_2664, QN => 
                           DataPath_RF_bus_reg_dataout_819_port);
   DataPath_RF_BLOCKi_33_Q_reg_18_inst : DFF_X1 port map( D => n4440, CK => CLK
                           , Q => n_2665, QN => 
                           DataPath_RF_bus_reg_dataout_818_port);
   DataPath_RF_BLOCKi_33_Q_reg_17_inst : DFF_X1 port map( D => n4441, CK => CLK
                           , Q => n_2666, QN => 
                           DataPath_RF_bus_reg_dataout_817_port);
   DataPath_RF_BLOCKi_33_Q_reg_16_inst : DFF_X1 port map( D => n4442, CK => CLK
                           , Q => n_2667, QN => 
                           DataPath_RF_bus_reg_dataout_816_port);
   DataPath_RF_BLOCKi_33_Q_reg_15_inst : DFF_X1 port map( D => n4443, CK => CLK
                           , Q => n_2668, QN => 
                           DataPath_RF_bus_reg_dataout_815_port);
   DataPath_RF_BLOCKi_33_Q_reg_14_inst : DFF_X1 port map( D => n4444, CK => CLK
                           , Q => n_2669, QN => 
                           DataPath_RF_bus_reg_dataout_814_port);
   DataPath_RF_BLOCKi_33_Q_reg_13_inst : DFF_X1 port map( D => n4445, CK => CLK
                           , Q => n_2670, QN => 
                           DataPath_RF_bus_reg_dataout_813_port);
   DataPath_RF_BLOCKi_33_Q_reg_12_inst : DFF_X1 port map( D => n4446, CK => CLK
                           , Q => n_2671, QN => 
                           DataPath_RF_bus_reg_dataout_812_port);
   DataPath_RF_BLOCKi_33_Q_reg_11_inst : DFF_X1 port map( D => n4447, CK => CLK
                           , Q => n_2672, QN => 
                           DataPath_RF_bus_reg_dataout_811_port);
   DataPath_RF_BLOCKi_33_Q_reg_9_inst : DFF_X1 port map( D => n4449, CK => CLK,
                           Q => n_2673, QN => 
                           DataPath_RF_bus_reg_dataout_809_port);
   DataPath_RF_BLOCKi_33_Q_reg_8_inst : DFF_X1 port map( D => n4450, CK => CLK,
                           Q => n_2674, QN => 
                           DataPath_RF_bus_reg_dataout_808_port);
   DataPath_RF_BLOCKi_33_Q_reg_7_inst : DFF_X1 port map( D => n4451, CK => CLK,
                           Q => n_2675, QN => 
                           DataPath_RF_bus_reg_dataout_807_port);
   DataPath_RF_BLOCKi_33_Q_reg_6_inst : DFF_X1 port map( D => n4452, CK => CLK,
                           Q => n_2676, QN => 
                           DataPath_RF_bus_reg_dataout_806_port);
   DataPath_RF_BLOCKi_33_Q_reg_5_inst : DFF_X1 port map( D => n4453, CK => CLK,
                           Q => n_2677, QN => 
                           DataPath_RF_bus_reg_dataout_805_port);
   DataPath_RF_BLOCKi_33_Q_reg_4_inst : DFF_X1 port map( D => n4454, CK => CLK,
                           Q => n_2678, QN => 
                           DataPath_RF_bus_reg_dataout_804_port);
   DataPath_RF_BLOCKi_33_Q_reg_3_inst : DFF_X1 port map( D => n4455, CK => CLK,
                           Q => n_2679, QN => 
                           DataPath_RF_bus_reg_dataout_803_port);
   DataPath_RF_BLOCKi_33_Q_reg_2_inst : DFF_X1 port map( D => n4456, CK => CLK,
                           Q => n_2680, QN => 
                           DataPath_RF_bus_reg_dataout_802_port);
   DataPath_RF_BLOCKi_33_Q_reg_1_inst : DFF_X1 port map( D => n4457, CK => CLK,
                           Q => n_2681, QN => 
                           DataPath_RF_bus_reg_dataout_801_port);
   DataPath_RF_BLOCKi_33_Q_reg_0_inst : DFF_X1 port map( D => n4458, CK => CLK,
                           Q => n_2682, QN => 
                           DataPath_RF_bus_reg_dataout_800_port);
   DataPath_RF_BLOCKi_49_Q_reg_31_inst : DFF_X1 port map( D => n5018, CK => CLK
                           , Q => n_2683, QN => 
                           DataPath_RF_bus_reg_dataout_1343_port);
   DataPath_RF_BLOCKi_49_Q_reg_30_inst : DFF_X1 port map( D => n5021, CK => CLK
                           , Q => n_2684, QN => 
                           DataPath_RF_bus_reg_dataout_1342_port);
   DataPath_RF_BLOCKi_49_Q_reg_29_inst : DFF_X1 port map( D => n5022, CK => CLK
                           , Q => n_2685, QN => 
                           DataPath_RF_bus_reg_dataout_1341_port);
   DataPath_RF_BLOCKi_49_Q_reg_28_inst : DFF_X1 port map( D => n5023, CK => CLK
                           , Q => n_2686, QN => 
                           DataPath_RF_bus_reg_dataout_1340_port);
   DataPath_RF_BLOCKi_49_Q_reg_27_inst : DFF_X1 port map( D => n5024, CK => CLK
                           , Q => n_2687, QN => 
                           DataPath_RF_bus_reg_dataout_1339_port);
   DataPath_RF_BLOCKi_49_Q_reg_26_inst : DFF_X1 port map( D => n5025, CK => CLK
                           , Q => n_2688, QN => 
                           DataPath_RF_bus_reg_dataout_1338_port);
   DataPath_RF_BLOCKi_49_Q_reg_25_inst : DFF_X1 port map( D => n5026, CK => CLK
                           , Q => n_2689, QN => 
                           DataPath_RF_bus_reg_dataout_1337_port);
   DataPath_RF_BLOCKi_49_Q_reg_24_inst : DFF_X1 port map( D => n5027, CK => CLK
                           , Q => n_2690, QN => 
                           DataPath_RF_bus_reg_dataout_1336_port);
   DataPath_RF_BLOCKi_49_Q_reg_23_inst : DFF_X1 port map( D => n5028, CK => CLK
                           , Q => n_2691, QN => 
                           DataPath_RF_bus_reg_dataout_1335_port);
   DataPath_RF_BLOCKi_49_Q_reg_22_inst : DFF_X1 port map( D => n5029, CK => CLK
                           , Q => n_2692, QN => 
                           DataPath_RF_bus_reg_dataout_1334_port);
   DataPath_RF_BLOCKi_49_Q_reg_21_inst : DFF_X1 port map( D => n5030, CK => CLK
                           , Q => n_2693, QN => 
                           DataPath_RF_bus_reg_dataout_1333_port);
   DataPath_RF_BLOCKi_49_Q_reg_20_inst : DFF_X1 port map( D => n5031, CK => CLK
                           , Q => n_2694, QN => 
                           DataPath_RF_bus_reg_dataout_1332_port);
   DataPath_RF_BLOCKi_49_Q_reg_19_inst : DFF_X1 port map( D => n5032, CK => CLK
                           , Q => n_2695, QN => 
                           DataPath_RF_bus_reg_dataout_1331_port);
   DataPath_RF_BLOCKi_49_Q_reg_18_inst : DFF_X1 port map( D => n5033, CK => CLK
                           , Q => n_2696, QN => 
                           DataPath_RF_bus_reg_dataout_1330_port);
   DataPath_RF_BLOCKi_49_Q_reg_17_inst : DFF_X1 port map( D => n5034, CK => CLK
                           , Q => n_2697, QN => 
                           DataPath_RF_bus_reg_dataout_1329_port);
   DataPath_RF_BLOCKi_49_Q_reg_16_inst : DFF_X1 port map( D => n5035, CK => CLK
                           , Q => n_2698, QN => 
                           DataPath_RF_bus_reg_dataout_1328_port);
   DataPath_RF_BLOCKi_49_Q_reg_15_inst : DFF_X1 port map( D => n5036, CK => CLK
                           , Q => n_2699, QN => 
                           DataPath_RF_bus_reg_dataout_1327_port);
   DataPath_RF_BLOCKi_49_Q_reg_14_inst : DFF_X1 port map( D => n5037, CK => CLK
                           , Q => n_2700, QN => 
                           DataPath_RF_bus_reg_dataout_1326_port);
   DataPath_RF_BLOCKi_49_Q_reg_13_inst : DFF_X1 port map( D => n5038, CK => CLK
                           , Q => n_2701, QN => 
                           DataPath_RF_bus_reg_dataout_1325_port);
   DataPath_RF_BLOCKi_49_Q_reg_12_inst : DFF_X1 port map( D => n5039, CK => CLK
                           , Q => n_2702, QN => 
                           DataPath_RF_bus_reg_dataout_1324_port);
   DataPath_RF_BLOCKi_49_Q_reg_11_inst : DFF_X1 port map( D => n5040, CK => CLK
                           , Q => n_2703, QN => 
                           DataPath_RF_bus_reg_dataout_1323_port);
   DataPath_RF_BLOCKi_49_Q_reg_9_inst : DFF_X1 port map( D => n5042, CK => CLK,
                           Q => n_2704, QN => 
                           DataPath_RF_bus_reg_dataout_1321_port);
   DataPath_RF_BLOCKi_49_Q_reg_8_inst : DFF_X1 port map( D => n5043, CK => CLK,
                           Q => n_2705, QN => 
                           DataPath_RF_bus_reg_dataout_1320_port);
   DataPath_RF_BLOCKi_49_Q_reg_7_inst : DFF_X1 port map( D => n5044, CK => CLK,
                           Q => n_2706, QN => 
                           DataPath_RF_bus_reg_dataout_1319_port);
   DataPath_RF_BLOCKi_49_Q_reg_6_inst : DFF_X1 port map( D => n5045, CK => CLK,
                           Q => n_2707, QN => 
                           DataPath_RF_bus_reg_dataout_1318_port);
   DataPath_RF_BLOCKi_49_Q_reg_5_inst : DFF_X1 port map( D => n5046, CK => CLK,
                           Q => n_2708, QN => 
                           DataPath_RF_bus_reg_dataout_1317_port);
   DataPath_RF_BLOCKi_49_Q_reg_4_inst : DFF_X1 port map( D => n5047, CK => CLK,
                           Q => n_2709, QN => 
                           DataPath_RF_bus_reg_dataout_1316_port);
   DataPath_RF_BLOCKi_49_Q_reg_3_inst : DFF_X1 port map( D => n5048, CK => CLK,
                           Q => n_2710, QN => 
                           DataPath_RF_bus_reg_dataout_1315_port);
   DataPath_RF_BLOCKi_49_Q_reg_2_inst : DFF_X1 port map( D => n5049, CK => CLK,
                           Q => n_2711, QN => 
                           DataPath_RF_bus_reg_dataout_1314_port);
   DataPath_RF_BLOCKi_49_Q_reg_1_inst : DFF_X1 port map( D => n5050, CK => CLK,
                           Q => n_2712, QN => 
                           DataPath_RF_bus_reg_dataout_1313_port);
   DataPath_RF_BLOCKi_49_Q_reg_0_inst : DFF_X1 port map( D => n5051, CK => CLK,
                           Q => n_2713, QN => 
                           DataPath_RF_bus_reg_dataout_1312_port);
   DataPath_RF_BLOCKi_65_Q_reg_31_inst : DFF_X1 port map( D => n5615, CK => CLK
                           , Q => n_2714, QN => 
                           DataPath_RF_bus_reg_dataout_1855_port);
   DataPath_RF_BLOCKi_65_Q_reg_30_inst : DFF_X1 port map( D => n5618, CK => CLK
                           , Q => n_2715, QN => 
                           DataPath_RF_bus_reg_dataout_1854_port);
   DataPath_RF_BLOCKi_65_Q_reg_29_inst : DFF_X1 port map( D => n5619, CK => CLK
                           , Q => n_2716, QN => 
                           DataPath_RF_bus_reg_dataout_1853_port);
   DataPath_RF_BLOCKi_65_Q_reg_28_inst : DFF_X1 port map( D => n5620, CK => CLK
                           , Q => n_2717, QN => 
                           DataPath_RF_bus_reg_dataout_1852_port);
   DataPath_RF_BLOCKi_65_Q_reg_27_inst : DFF_X1 port map( D => n5621, CK => CLK
                           , Q => n_2718, QN => 
                           DataPath_RF_bus_reg_dataout_1851_port);
   DataPath_RF_BLOCKi_65_Q_reg_26_inst : DFF_X1 port map( D => n5622, CK => CLK
                           , Q => n_2719, QN => 
                           DataPath_RF_bus_reg_dataout_1850_port);
   DataPath_RF_BLOCKi_65_Q_reg_25_inst : DFF_X1 port map( D => n5623, CK => CLK
                           , Q => n_2720, QN => 
                           DataPath_RF_bus_reg_dataout_1849_port);
   DataPath_RF_BLOCKi_65_Q_reg_24_inst : DFF_X1 port map( D => n5624, CK => CLK
                           , Q => n_2721, QN => 
                           DataPath_RF_bus_reg_dataout_1848_port);
   DataPath_RF_BLOCKi_65_Q_reg_23_inst : DFF_X1 port map( D => n5625, CK => CLK
                           , Q => n_2722, QN => 
                           DataPath_RF_bus_reg_dataout_1847_port);
   DataPath_RF_BLOCKi_65_Q_reg_22_inst : DFF_X1 port map( D => n5626, CK => CLK
                           , Q => n_2723, QN => 
                           DataPath_RF_bus_reg_dataout_1846_port);
   DataPath_RF_BLOCKi_65_Q_reg_21_inst : DFF_X1 port map( D => n5627, CK => CLK
                           , Q => n_2724, QN => 
                           DataPath_RF_bus_reg_dataout_1845_port);
   DataPath_RF_BLOCKi_65_Q_reg_20_inst : DFF_X1 port map( D => n5628, CK => CLK
                           , Q => n_2725, QN => 
                           DataPath_RF_bus_reg_dataout_1844_port);
   DataPath_RF_BLOCKi_65_Q_reg_19_inst : DFF_X1 port map( D => n5629, CK => CLK
                           , Q => n_2726, QN => 
                           DataPath_RF_bus_reg_dataout_1843_port);
   DataPath_RF_BLOCKi_65_Q_reg_18_inst : DFF_X1 port map( D => n5630, CK => CLK
                           , Q => n_2727, QN => 
                           DataPath_RF_bus_reg_dataout_1842_port);
   DataPath_RF_BLOCKi_65_Q_reg_17_inst : DFF_X1 port map( D => n5631, CK => CLK
                           , Q => n_2728, QN => 
                           DataPath_RF_bus_reg_dataout_1841_port);
   DataPath_RF_BLOCKi_65_Q_reg_16_inst : DFF_X1 port map( D => n5632, CK => CLK
                           , Q => n_2729, QN => 
                           DataPath_RF_bus_reg_dataout_1840_port);
   DataPath_RF_BLOCKi_65_Q_reg_15_inst : DFF_X1 port map( D => n5633, CK => CLK
                           , Q => n_2730, QN => 
                           DataPath_RF_bus_reg_dataout_1839_port);
   DataPath_RF_BLOCKi_65_Q_reg_14_inst : DFF_X1 port map( D => n5634, CK => CLK
                           , Q => n_2731, QN => 
                           DataPath_RF_bus_reg_dataout_1838_port);
   DataPath_RF_BLOCKi_65_Q_reg_13_inst : DFF_X1 port map( D => n5635, CK => CLK
                           , Q => n_2732, QN => 
                           DataPath_RF_bus_reg_dataout_1837_port);
   DataPath_RF_BLOCKi_65_Q_reg_12_inst : DFF_X1 port map( D => n5636, CK => CLK
                           , Q => n_2733, QN => 
                           DataPath_RF_bus_reg_dataout_1836_port);
   DataPath_RF_BLOCKi_65_Q_reg_11_inst : DFF_X1 port map( D => n5637, CK => CLK
                           , Q => n_2734, QN => 
                           DataPath_RF_bus_reg_dataout_1835_port);
   DataPath_RF_BLOCKi_65_Q_reg_9_inst : DFF_X1 port map( D => n5639, CK => CLK,
                           Q => n_2735, QN => 
                           DataPath_RF_bus_reg_dataout_1833_port);
   DataPath_RF_BLOCKi_65_Q_reg_8_inst : DFF_X1 port map( D => n5640, CK => CLK,
                           Q => n_2736, QN => 
                           DataPath_RF_bus_reg_dataout_1832_port);
   DataPath_RF_BLOCKi_65_Q_reg_7_inst : DFF_X1 port map( D => n5641, CK => CLK,
                           Q => n_2737, QN => 
                           DataPath_RF_bus_reg_dataout_1831_port);
   DataPath_RF_BLOCKi_65_Q_reg_6_inst : DFF_X1 port map( D => n5642, CK => CLK,
                           Q => n_2738, QN => 
                           DataPath_RF_bus_reg_dataout_1830_port);
   DataPath_RF_BLOCKi_65_Q_reg_5_inst : DFF_X1 port map( D => n5643, CK => CLK,
                           Q => n_2739, QN => 
                           DataPath_RF_bus_reg_dataout_1829_port);
   DataPath_RF_BLOCKi_65_Q_reg_4_inst : DFF_X1 port map( D => n5644, CK => CLK,
                           Q => n_2740, QN => 
                           DataPath_RF_bus_reg_dataout_1828_port);
   DataPath_RF_BLOCKi_65_Q_reg_3_inst : DFF_X1 port map( D => n5645, CK => CLK,
                           Q => n_2741, QN => 
                           DataPath_RF_bus_reg_dataout_1827_port);
   DataPath_RF_BLOCKi_65_Q_reg_2_inst : DFF_X1 port map( D => n5646, CK => CLK,
                           Q => n_2742, QN => 
                           DataPath_RF_bus_reg_dataout_1826_port);
   DataPath_RF_BLOCKi_65_Q_reg_1_inst : DFF_X1 port map( D => n5647, CK => CLK,
                           Q => n_2743, QN => 
                           DataPath_RF_bus_reg_dataout_1825_port);
   DataPath_RF_BLOCKi_65_Q_reg_0_inst : DFF_X1 port map( D => n5648, CK => CLK,
                           Q => n_2744, QN => 
                           DataPath_RF_bus_reg_dataout_1824_port);
   DataPath_RF_BLOCKi_82_Q_reg_31_inst : DFF_X1 port map( D => n1003, CK => CLK
                           , Q => n_2745, QN => 
                           DataPath_RF_bus_reg_dataout_2399_port);
   DataPath_RF_BLOCKi_82_Q_reg_30_inst : DFF_X1 port map( D => n1006, CK => CLK
                           , Q => n_2746, QN => 
                           DataPath_RF_bus_reg_dataout_2398_port);
   DataPath_RF_BLOCKi_82_Q_reg_29_inst : DFF_X1 port map( D => n1007, CK => CLK
                           , Q => n_2747, QN => 
                           DataPath_RF_bus_reg_dataout_2397_port);
   DataPath_RF_BLOCKi_82_Q_reg_28_inst : DFF_X1 port map( D => n1008, CK => CLK
                           , Q => n_2748, QN => 
                           DataPath_RF_bus_reg_dataout_2396_port);
   DataPath_RF_BLOCKi_82_Q_reg_27_inst : DFF_X1 port map( D => n1009, CK => CLK
                           , Q => n_2749, QN => 
                           DataPath_RF_bus_reg_dataout_2395_port);
   DataPath_RF_BLOCKi_82_Q_reg_26_inst : DFF_X1 port map( D => n1010, CK => CLK
                           , Q => n_2750, QN => 
                           DataPath_RF_bus_reg_dataout_2394_port);
   DataPath_RF_BLOCKi_82_Q_reg_25_inst : DFF_X1 port map( D => n1011, CK => CLK
                           , Q => n_2751, QN => 
                           DataPath_RF_bus_reg_dataout_2393_port);
   DataPath_RF_BLOCKi_82_Q_reg_24_inst : DFF_X1 port map( D => n1012, CK => CLK
                           , Q => n_2752, QN => 
                           DataPath_RF_bus_reg_dataout_2392_port);
   DataPath_RF_BLOCKi_82_Q_reg_23_inst : DFF_X1 port map( D => n1013, CK => CLK
                           , Q => n_2753, QN => 
                           DataPath_RF_bus_reg_dataout_2391_port);
   DataPath_RF_BLOCKi_82_Q_reg_22_inst : DFF_X1 port map( D => n1014, CK => CLK
                           , Q => n_2754, QN => 
                           DataPath_RF_bus_reg_dataout_2390_port);
   DataPath_RF_BLOCKi_82_Q_reg_21_inst : DFF_X1 port map( D => n1015, CK => CLK
                           , Q => n_2755, QN => 
                           DataPath_RF_bus_reg_dataout_2389_port);
   DataPath_RF_BLOCKi_82_Q_reg_20_inst : DFF_X1 port map( D => n1016, CK => CLK
                           , Q => n_2756, QN => 
                           DataPath_RF_bus_reg_dataout_2388_port);
   DataPath_RF_BLOCKi_82_Q_reg_19_inst : DFF_X1 port map( D => n1017, CK => CLK
                           , Q => n_2757, QN => 
                           DataPath_RF_bus_reg_dataout_2387_port);
   DataPath_RF_BLOCKi_82_Q_reg_18_inst : DFF_X1 port map( D => n1018, CK => CLK
                           , Q => n_2758, QN => 
                           DataPath_RF_bus_reg_dataout_2386_port);
   DataPath_RF_BLOCKi_82_Q_reg_17_inst : DFF_X1 port map( D => n1019, CK => CLK
                           , Q => n_2759, QN => 
                           DataPath_RF_bus_reg_dataout_2385_port);
   DataPath_RF_BLOCKi_82_Q_reg_16_inst : DFF_X1 port map( D => n1020, CK => CLK
                           , Q => n_2760, QN => 
                           DataPath_RF_bus_reg_dataout_2384_port);
   DataPath_RF_BLOCKi_82_Q_reg_15_inst : DFF_X1 port map( D => n1021, CK => CLK
                           , Q => n_2761, QN => 
                           DataPath_RF_bus_reg_dataout_2383_port);
   DataPath_RF_BLOCKi_82_Q_reg_14_inst : DFF_X1 port map( D => n1022, CK => CLK
                           , Q => n_2762, QN => 
                           DataPath_RF_bus_reg_dataout_2382_port);
   DataPath_RF_BLOCKi_82_Q_reg_13_inst : DFF_X1 port map( D => n1023, CK => CLK
                           , Q => n_2763, QN => 
                           DataPath_RF_bus_reg_dataout_2381_port);
   DataPath_RF_BLOCKi_82_Q_reg_12_inst : DFF_X1 port map( D => n1024, CK => CLK
                           , Q => n_2764, QN => 
                           DataPath_RF_bus_reg_dataout_2380_port);
   DataPath_RF_BLOCKi_82_Q_reg_11_inst : DFF_X1 port map( D => n1025, CK => CLK
                           , Q => n_2765, QN => 
                           DataPath_RF_bus_reg_dataout_2379_port);
   DataPath_RF_BLOCKi_82_Q_reg_9_inst : DFF_X1 port map( D => n1027, CK => CLK,
                           Q => n_2766, QN => 
                           DataPath_RF_bus_reg_dataout_2377_port);
   DataPath_RF_BLOCKi_82_Q_reg_8_inst : DFF_X1 port map( D => n1028, CK => CLK,
                           Q => n_2767, QN => 
                           DataPath_RF_bus_reg_dataout_2376_port);
   DataPath_RF_BLOCKi_82_Q_reg_7_inst : DFF_X1 port map( D => n1029, CK => CLK,
                           Q => n_2768, QN => 
                           DataPath_RF_bus_reg_dataout_2375_port);
   DataPath_RF_BLOCKi_82_Q_reg_6_inst : DFF_X1 port map( D => n1030, CK => CLK,
                           Q => n_2769, QN => 
                           DataPath_RF_bus_reg_dataout_2374_port);
   DataPath_RF_BLOCKi_82_Q_reg_5_inst : DFF_X1 port map( D => n1031, CK => CLK,
                           Q => n_2770, QN => 
                           DataPath_RF_bus_reg_dataout_2373_port);
   DataPath_RF_BLOCKi_82_Q_reg_4_inst : DFF_X1 port map( D => n1032, CK => CLK,
                           Q => n_2771, QN => 
                           DataPath_RF_bus_reg_dataout_2372_port);
   DataPath_RF_BLOCKi_82_Q_reg_3_inst : DFF_X1 port map( D => n1033, CK => CLK,
                           Q => n_2772, QN => 
                           DataPath_RF_bus_reg_dataout_2371_port);
   DataPath_RF_BLOCKi_82_Q_reg_2_inst : DFF_X1 port map( D => n1034, CK => CLK,
                           Q => n_2773, QN => 
                           DataPath_RF_bus_reg_dataout_2370_port);
   DataPath_RF_BLOCKi_82_Q_reg_1_inst : DFF_X1 port map( D => n1035, CK => CLK,
                           Q => n_2774, QN => 
                           DataPath_RF_bus_reg_dataout_2369_port);
   DataPath_RF_BLOCKi_82_Q_reg_0_inst : DFF_X1 port map( D => n1036, CK => CLK,
                           Q => n_2775, QN => 
                           DataPath_RF_bus_reg_dataout_2368_port);
   DataPath_RF_BLOCKi_18_Q_reg_31_inst : DFF_X1 port map( D => n3835, CK => CLK
                           , Q => n_2776, QN => 
                           DataPath_RF_bus_reg_dataout_351_port);
   DataPath_RF_BLOCKi_18_Q_reg_30_inst : DFF_X1 port map( D => n3838, CK => CLK
                           , Q => n_2777, QN => 
                           DataPath_RF_bus_reg_dataout_350_port);
   DataPath_RF_BLOCKi_18_Q_reg_29_inst : DFF_X1 port map( D => n3839, CK => CLK
                           , Q => n_2778, QN => 
                           DataPath_RF_bus_reg_dataout_349_port);
   DataPath_RF_BLOCKi_18_Q_reg_28_inst : DFF_X1 port map( D => n3840, CK => CLK
                           , Q => n_2779, QN => 
                           DataPath_RF_bus_reg_dataout_348_port);
   DataPath_RF_BLOCKi_18_Q_reg_27_inst : DFF_X1 port map( D => n3841, CK => CLK
                           , Q => n_2780, QN => 
                           DataPath_RF_bus_reg_dataout_347_port);
   DataPath_RF_BLOCKi_18_Q_reg_26_inst : DFF_X1 port map( D => n3842, CK => CLK
                           , Q => n_2781, QN => 
                           DataPath_RF_bus_reg_dataout_346_port);
   DataPath_RF_BLOCKi_18_Q_reg_25_inst : DFF_X1 port map( D => n3843, CK => CLK
                           , Q => n_2782, QN => 
                           DataPath_RF_bus_reg_dataout_345_port);
   DataPath_RF_BLOCKi_18_Q_reg_24_inst : DFF_X1 port map( D => n3844, CK => CLK
                           , Q => n_2783, QN => 
                           DataPath_RF_bus_reg_dataout_344_port);
   DataPath_RF_BLOCKi_18_Q_reg_23_inst : DFF_X1 port map( D => n3845, CK => CLK
                           , Q => n_2784, QN => 
                           DataPath_RF_bus_reg_dataout_343_port);
   DataPath_RF_BLOCKi_18_Q_reg_22_inst : DFF_X1 port map( D => n3846, CK => CLK
                           , Q => n_2785, QN => 
                           DataPath_RF_bus_reg_dataout_342_port);
   DataPath_RF_BLOCKi_18_Q_reg_21_inst : DFF_X1 port map( D => n3847, CK => CLK
                           , Q => n_2786, QN => 
                           DataPath_RF_bus_reg_dataout_341_port);
   DataPath_RF_BLOCKi_18_Q_reg_20_inst : DFF_X1 port map( D => n3848, CK => CLK
                           , Q => n_2787, QN => 
                           DataPath_RF_bus_reg_dataout_340_port);
   DataPath_RF_BLOCKi_18_Q_reg_19_inst : DFF_X1 port map( D => n3849, CK => CLK
                           , Q => n_2788, QN => 
                           DataPath_RF_bus_reg_dataout_339_port);
   DataPath_RF_BLOCKi_18_Q_reg_18_inst : DFF_X1 port map( D => n3850, CK => CLK
                           , Q => n_2789, QN => 
                           DataPath_RF_bus_reg_dataout_338_port);
   DataPath_RF_BLOCKi_18_Q_reg_17_inst : DFF_X1 port map( D => n3851, CK => CLK
                           , Q => n_2790, QN => 
                           DataPath_RF_bus_reg_dataout_337_port);
   DataPath_RF_BLOCKi_18_Q_reg_16_inst : DFF_X1 port map( D => n3852, CK => CLK
                           , Q => n_2791, QN => 
                           DataPath_RF_bus_reg_dataout_336_port);
   DataPath_RF_BLOCKi_18_Q_reg_15_inst : DFF_X1 port map( D => n3853, CK => CLK
                           , Q => n_2792, QN => 
                           DataPath_RF_bus_reg_dataout_335_port);
   DataPath_RF_BLOCKi_18_Q_reg_14_inst : DFF_X1 port map( D => n3854, CK => CLK
                           , Q => n_2793, QN => 
                           DataPath_RF_bus_reg_dataout_334_port);
   DataPath_RF_BLOCKi_18_Q_reg_13_inst : DFF_X1 port map( D => n3855, CK => CLK
                           , Q => n_2794, QN => 
                           DataPath_RF_bus_reg_dataout_333_port);
   DataPath_RF_BLOCKi_18_Q_reg_12_inst : DFF_X1 port map( D => n3856, CK => CLK
                           , Q => n_2795, QN => 
                           DataPath_RF_bus_reg_dataout_332_port);
   DataPath_RF_BLOCKi_18_Q_reg_11_inst : DFF_X1 port map( D => n3857, CK => CLK
                           , Q => n_2796, QN => 
                           DataPath_RF_bus_reg_dataout_331_port);
   DataPath_RF_BLOCKi_18_Q_reg_9_inst : DFF_X1 port map( D => n3859, CK => CLK,
                           Q => n_2797, QN => 
                           DataPath_RF_bus_reg_dataout_329_port);
   DataPath_RF_BLOCKi_18_Q_reg_8_inst : DFF_X1 port map( D => n3860, CK => CLK,
                           Q => n_2798, QN => 
                           DataPath_RF_bus_reg_dataout_328_port);
   DataPath_RF_BLOCKi_18_Q_reg_7_inst : DFF_X1 port map( D => n3861, CK => CLK,
                           Q => n_2799, QN => 
                           DataPath_RF_bus_reg_dataout_327_port);
   DataPath_RF_BLOCKi_18_Q_reg_6_inst : DFF_X1 port map( D => n3862, CK => CLK,
                           Q => n_2800, QN => 
                           DataPath_RF_bus_reg_dataout_326_port);
   DataPath_RF_BLOCKi_18_Q_reg_5_inst : DFF_X1 port map( D => n3863, CK => CLK,
                           Q => n_2801, QN => 
                           DataPath_RF_bus_reg_dataout_325_port);
   DataPath_RF_BLOCKi_18_Q_reg_4_inst : DFF_X1 port map( D => n3864, CK => CLK,
                           Q => n_2802, QN => 
                           DataPath_RF_bus_reg_dataout_324_port);
   DataPath_RF_BLOCKi_18_Q_reg_3_inst : DFF_X1 port map( D => n3865, CK => CLK,
                           Q => n_2803, QN => 
                           DataPath_RF_bus_reg_dataout_323_port);
   DataPath_RF_BLOCKi_18_Q_reg_2_inst : DFF_X1 port map( D => n3866, CK => CLK,
                           Q => n_2804, QN => 
                           DataPath_RF_bus_reg_dataout_322_port);
   DataPath_RF_BLOCKi_18_Q_reg_1_inst : DFF_X1 port map( D => n3867, CK => CLK,
                           Q => n_2805, QN => 
                           DataPath_RF_bus_reg_dataout_321_port);
   DataPath_RF_BLOCKi_18_Q_reg_0_inst : DFF_X1 port map( D => n3868, CK => CLK,
                           Q => n_2806, QN => 
                           DataPath_RF_bus_reg_dataout_320_port);
   DataPath_RF_BLOCKi_34_Q_reg_31_inst : DFF_X1 port map( D => n4460, CK => CLK
                           , Q => n_2807, QN => 
                           DataPath_RF_bus_reg_dataout_863_port);
   DataPath_RF_BLOCKi_34_Q_reg_30_inst : DFF_X1 port map( D => n4463, CK => CLK
                           , Q => n_2808, QN => 
                           DataPath_RF_bus_reg_dataout_862_port);
   DataPath_RF_BLOCKi_34_Q_reg_29_inst : DFF_X1 port map( D => n4464, CK => CLK
                           , Q => n_2809, QN => 
                           DataPath_RF_bus_reg_dataout_861_port);
   DataPath_RF_BLOCKi_34_Q_reg_28_inst : DFF_X1 port map( D => n4465, CK => CLK
                           , Q => n_2810, QN => 
                           DataPath_RF_bus_reg_dataout_860_port);
   DataPath_RF_BLOCKi_34_Q_reg_27_inst : DFF_X1 port map( D => n4466, CK => CLK
                           , Q => n_2811, QN => 
                           DataPath_RF_bus_reg_dataout_859_port);
   DataPath_RF_BLOCKi_34_Q_reg_26_inst : DFF_X1 port map( D => n4467, CK => CLK
                           , Q => n_2812, QN => 
                           DataPath_RF_bus_reg_dataout_858_port);
   DataPath_RF_BLOCKi_34_Q_reg_25_inst : DFF_X1 port map( D => n4468, CK => CLK
                           , Q => n_2813, QN => 
                           DataPath_RF_bus_reg_dataout_857_port);
   DataPath_RF_BLOCKi_34_Q_reg_24_inst : DFF_X1 port map( D => n4469, CK => CLK
                           , Q => n_2814, QN => 
                           DataPath_RF_bus_reg_dataout_856_port);
   DataPath_RF_BLOCKi_34_Q_reg_23_inst : DFF_X1 port map( D => n4470, CK => CLK
                           , Q => n_2815, QN => 
                           DataPath_RF_bus_reg_dataout_855_port);
   DataPath_RF_BLOCKi_34_Q_reg_22_inst : DFF_X1 port map( D => n4471, CK => CLK
                           , Q => n_2816, QN => 
                           DataPath_RF_bus_reg_dataout_854_port);
   DataPath_RF_BLOCKi_34_Q_reg_21_inst : DFF_X1 port map( D => n4472, CK => CLK
                           , Q => n_2817, QN => 
                           DataPath_RF_bus_reg_dataout_853_port);
   DataPath_RF_BLOCKi_34_Q_reg_20_inst : DFF_X1 port map( D => n4473, CK => CLK
                           , Q => n_2818, QN => 
                           DataPath_RF_bus_reg_dataout_852_port);
   DataPath_RF_BLOCKi_34_Q_reg_19_inst : DFF_X1 port map( D => n4474, CK => CLK
                           , Q => n_2819, QN => 
                           DataPath_RF_bus_reg_dataout_851_port);
   DataPath_RF_BLOCKi_34_Q_reg_18_inst : DFF_X1 port map( D => n4475, CK => CLK
                           , Q => n_2820, QN => 
                           DataPath_RF_bus_reg_dataout_850_port);
   DataPath_RF_BLOCKi_34_Q_reg_17_inst : DFF_X1 port map( D => n4476, CK => CLK
                           , Q => n_2821, QN => 
                           DataPath_RF_bus_reg_dataout_849_port);
   DataPath_RF_BLOCKi_34_Q_reg_16_inst : DFF_X1 port map( D => n4477, CK => CLK
                           , Q => n_2822, QN => 
                           DataPath_RF_bus_reg_dataout_848_port);
   DataPath_RF_BLOCKi_34_Q_reg_15_inst : DFF_X1 port map( D => n4478, CK => CLK
                           , Q => n_2823, QN => 
                           DataPath_RF_bus_reg_dataout_847_port);
   DataPath_RF_BLOCKi_34_Q_reg_14_inst : DFF_X1 port map( D => n4479, CK => CLK
                           , Q => n_2824, QN => 
                           DataPath_RF_bus_reg_dataout_846_port);
   DataPath_RF_BLOCKi_34_Q_reg_13_inst : DFF_X1 port map( D => n4480, CK => CLK
                           , Q => n_2825, QN => 
                           DataPath_RF_bus_reg_dataout_845_port);
   DataPath_RF_BLOCKi_34_Q_reg_12_inst : DFF_X1 port map( D => n4481, CK => CLK
                           , Q => n_2826, QN => 
                           DataPath_RF_bus_reg_dataout_844_port);
   DataPath_RF_BLOCKi_34_Q_reg_11_inst : DFF_X1 port map( D => n4482, CK => CLK
                           , Q => n_2827, QN => 
                           DataPath_RF_bus_reg_dataout_843_port);
   DataPath_RF_BLOCKi_34_Q_reg_9_inst : DFF_X1 port map( D => n4484, CK => CLK,
                           Q => n_2828, QN => 
                           DataPath_RF_bus_reg_dataout_841_port);
   DataPath_RF_BLOCKi_34_Q_reg_8_inst : DFF_X1 port map( D => n4485, CK => CLK,
                           Q => n_2829, QN => 
                           DataPath_RF_bus_reg_dataout_840_port);
   DataPath_RF_BLOCKi_34_Q_reg_7_inst : DFF_X1 port map( D => n4486, CK => CLK,
                           Q => n_2830, QN => 
                           DataPath_RF_bus_reg_dataout_839_port);
   DataPath_RF_BLOCKi_34_Q_reg_6_inst : DFF_X1 port map( D => n4487, CK => CLK,
                           Q => n_2831, QN => 
                           DataPath_RF_bus_reg_dataout_838_port);
   DataPath_RF_BLOCKi_34_Q_reg_5_inst : DFF_X1 port map( D => n4488, CK => CLK,
                           Q => n_2832, QN => 
                           DataPath_RF_bus_reg_dataout_837_port);
   DataPath_RF_BLOCKi_34_Q_reg_4_inst : DFF_X1 port map( D => n4489, CK => CLK,
                           Q => n_2833, QN => 
                           DataPath_RF_bus_reg_dataout_836_port);
   DataPath_RF_BLOCKi_34_Q_reg_3_inst : DFF_X1 port map( D => n4490, CK => CLK,
                           Q => n_2834, QN => 
                           DataPath_RF_bus_reg_dataout_835_port);
   DataPath_RF_BLOCKi_34_Q_reg_2_inst : DFF_X1 port map( D => n4491, CK => CLK,
                           Q => n_2835, QN => 
                           DataPath_RF_bus_reg_dataout_834_port);
   DataPath_RF_BLOCKi_34_Q_reg_1_inst : DFF_X1 port map( D => n4492, CK => CLK,
                           Q => n_2836, QN => 
                           DataPath_RF_bus_reg_dataout_833_port);
   DataPath_RF_BLOCKi_34_Q_reg_0_inst : DFF_X1 port map( D => n4493, CK => CLK,
                           Q => n_2837, QN => 
                           DataPath_RF_bus_reg_dataout_832_port);
   DataPath_RF_BLOCKi_50_Q_reg_31_inst : DFF_X1 port map( D => n5053, CK => CLK
                           , Q => n_2838, QN => 
                           DataPath_RF_bus_reg_dataout_1375_port);
   DataPath_RF_BLOCKi_50_Q_reg_30_inst : DFF_X1 port map( D => n5056, CK => CLK
                           , Q => n_2839, QN => 
                           DataPath_RF_bus_reg_dataout_1374_port);
   DataPath_RF_BLOCKi_50_Q_reg_29_inst : DFF_X1 port map( D => n5057, CK => CLK
                           , Q => n_2840, QN => 
                           DataPath_RF_bus_reg_dataout_1373_port);
   DataPath_RF_BLOCKi_50_Q_reg_28_inst : DFF_X1 port map( D => n5058, CK => CLK
                           , Q => n_2841, QN => 
                           DataPath_RF_bus_reg_dataout_1372_port);
   DataPath_RF_BLOCKi_50_Q_reg_27_inst : DFF_X1 port map( D => n5059, CK => CLK
                           , Q => n_2842, QN => 
                           DataPath_RF_bus_reg_dataout_1371_port);
   DataPath_RF_BLOCKi_50_Q_reg_26_inst : DFF_X1 port map( D => n5060, CK => CLK
                           , Q => n_2843, QN => 
                           DataPath_RF_bus_reg_dataout_1370_port);
   DataPath_RF_BLOCKi_50_Q_reg_25_inst : DFF_X1 port map( D => n5061, CK => CLK
                           , Q => n_2844, QN => 
                           DataPath_RF_bus_reg_dataout_1369_port);
   DataPath_RF_BLOCKi_50_Q_reg_24_inst : DFF_X1 port map( D => n5062, CK => CLK
                           , Q => n_2845, QN => 
                           DataPath_RF_bus_reg_dataout_1368_port);
   DataPath_RF_BLOCKi_50_Q_reg_23_inst : DFF_X1 port map( D => n5063, CK => CLK
                           , Q => n_2846, QN => 
                           DataPath_RF_bus_reg_dataout_1367_port);
   DataPath_RF_BLOCKi_50_Q_reg_22_inst : DFF_X1 port map( D => n5064, CK => CLK
                           , Q => n_2847, QN => 
                           DataPath_RF_bus_reg_dataout_1366_port);
   DataPath_RF_BLOCKi_50_Q_reg_21_inst : DFF_X1 port map( D => n5065, CK => CLK
                           , Q => n_2848, QN => 
                           DataPath_RF_bus_reg_dataout_1365_port);
   DataPath_RF_BLOCKi_50_Q_reg_20_inst : DFF_X1 port map( D => n5066, CK => CLK
                           , Q => n_2849, QN => 
                           DataPath_RF_bus_reg_dataout_1364_port);
   DataPath_RF_BLOCKi_50_Q_reg_19_inst : DFF_X1 port map( D => n5067, CK => CLK
                           , Q => n_2850, QN => 
                           DataPath_RF_bus_reg_dataout_1363_port);
   DataPath_RF_BLOCKi_50_Q_reg_18_inst : DFF_X1 port map( D => n5068, CK => CLK
                           , Q => n_2851, QN => 
                           DataPath_RF_bus_reg_dataout_1362_port);
   DataPath_RF_BLOCKi_50_Q_reg_17_inst : DFF_X1 port map( D => n5069, CK => CLK
                           , Q => n_2852, QN => 
                           DataPath_RF_bus_reg_dataout_1361_port);
   DataPath_RF_BLOCKi_50_Q_reg_16_inst : DFF_X1 port map( D => n5070, CK => CLK
                           , Q => n_2853, QN => 
                           DataPath_RF_bus_reg_dataout_1360_port);
   DataPath_RF_BLOCKi_50_Q_reg_15_inst : DFF_X1 port map( D => n5071, CK => CLK
                           , Q => n_2854, QN => 
                           DataPath_RF_bus_reg_dataout_1359_port);
   DataPath_RF_BLOCKi_50_Q_reg_14_inst : DFF_X1 port map( D => n5072, CK => CLK
                           , Q => n_2855, QN => 
                           DataPath_RF_bus_reg_dataout_1358_port);
   DataPath_RF_BLOCKi_50_Q_reg_13_inst : DFF_X1 port map( D => n5073, CK => CLK
                           , Q => n_2856, QN => 
                           DataPath_RF_bus_reg_dataout_1357_port);
   DataPath_RF_BLOCKi_50_Q_reg_12_inst : DFF_X1 port map( D => n5074, CK => CLK
                           , Q => n_2857, QN => 
                           DataPath_RF_bus_reg_dataout_1356_port);
   DataPath_RF_BLOCKi_50_Q_reg_11_inst : DFF_X1 port map( D => n5075, CK => CLK
                           , Q => n_2858, QN => 
                           DataPath_RF_bus_reg_dataout_1355_port);
   DataPath_RF_BLOCKi_50_Q_reg_9_inst : DFF_X1 port map( D => n5077, CK => CLK,
                           Q => n_2859, QN => 
                           DataPath_RF_bus_reg_dataout_1353_port);
   DataPath_RF_BLOCKi_50_Q_reg_8_inst : DFF_X1 port map( D => n5078, CK => CLK,
                           Q => n_2860, QN => 
                           DataPath_RF_bus_reg_dataout_1352_port);
   DataPath_RF_BLOCKi_50_Q_reg_7_inst : DFF_X1 port map( D => n5079, CK => CLK,
                           Q => n_2861, QN => 
                           DataPath_RF_bus_reg_dataout_1351_port);
   DataPath_RF_BLOCKi_50_Q_reg_6_inst : DFF_X1 port map( D => n5080, CK => CLK,
                           Q => n_2862, QN => 
                           DataPath_RF_bus_reg_dataout_1350_port);
   DataPath_RF_BLOCKi_50_Q_reg_5_inst : DFF_X1 port map( D => n5081, CK => CLK,
                           Q => n_2863, QN => 
                           DataPath_RF_bus_reg_dataout_1349_port);
   DataPath_RF_BLOCKi_50_Q_reg_4_inst : DFF_X1 port map( D => n5082, CK => CLK,
                           Q => n_2864, QN => 
                           DataPath_RF_bus_reg_dataout_1348_port);
   DataPath_RF_BLOCKi_50_Q_reg_3_inst : DFF_X1 port map( D => n5083, CK => CLK,
                           Q => n_2865, QN => 
                           DataPath_RF_bus_reg_dataout_1347_port);
   DataPath_RF_BLOCKi_50_Q_reg_2_inst : DFF_X1 port map( D => n5084, CK => CLK,
                           Q => n_2866, QN => 
                           DataPath_RF_bus_reg_dataout_1346_port);
   DataPath_RF_BLOCKi_50_Q_reg_1_inst : DFF_X1 port map( D => n5085, CK => CLK,
                           Q => n_2867, QN => 
                           DataPath_RF_bus_reg_dataout_1345_port);
   DataPath_RF_BLOCKi_50_Q_reg_0_inst : DFF_X1 port map( D => n5086, CK => CLK,
                           Q => n_2868, QN => 
                           DataPath_RF_bus_reg_dataout_1344_port);
   DataPath_RF_BLOCKi_66_Q_reg_31_inst : DFF_X1 port map( D => n5651, CK => CLK
                           , Q => n_2869, QN => 
                           DataPath_RF_bus_reg_dataout_1887_port);
   DataPath_RF_BLOCKi_66_Q_reg_30_inst : DFF_X1 port map( D => n5654, CK => CLK
                           , Q => n_2870, QN => 
                           DataPath_RF_bus_reg_dataout_1886_port);
   DataPath_RF_BLOCKi_66_Q_reg_29_inst : DFF_X1 port map( D => n5655, CK => CLK
                           , Q => n_2871, QN => 
                           DataPath_RF_bus_reg_dataout_1885_port);
   DataPath_RF_BLOCKi_66_Q_reg_28_inst : DFF_X1 port map( D => n5656, CK => CLK
                           , Q => n_2872, QN => 
                           DataPath_RF_bus_reg_dataout_1884_port);
   DataPath_RF_BLOCKi_66_Q_reg_27_inst : DFF_X1 port map( D => n5657, CK => CLK
                           , Q => n_2873, QN => 
                           DataPath_RF_bus_reg_dataout_1883_port);
   DataPath_RF_BLOCKi_66_Q_reg_26_inst : DFF_X1 port map( D => n5658, CK => CLK
                           , Q => n_2874, QN => 
                           DataPath_RF_bus_reg_dataout_1882_port);
   DataPath_RF_BLOCKi_66_Q_reg_25_inst : DFF_X1 port map( D => n5659, CK => CLK
                           , Q => n_2875, QN => 
                           DataPath_RF_bus_reg_dataout_1881_port);
   DataPath_RF_BLOCKi_66_Q_reg_24_inst : DFF_X1 port map( D => n5660, CK => CLK
                           , Q => n_2876, QN => 
                           DataPath_RF_bus_reg_dataout_1880_port);
   DataPath_RF_BLOCKi_66_Q_reg_23_inst : DFF_X1 port map( D => n5661, CK => CLK
                           , Q => n_2877, QN => 
                           DataPath_RF_bus_reg_dataout_1879_port);
   DataPath_RF_BLOCKi_66_Q_reg_22_inst : DFF_X1 port map( D => n5662, CK => CLK
                           , Q => n_2878, QN => 
                           DataPath_RF_bus_reg_dataout_1878_port);
   DataPath_RF_BLOCKi_66_Q_reg_21_inst : DFF_X1 port map( D => n5663, CK => CLK
                           , Q => n_2879, QN => 
                           DataPath_RF_bus_reg_dataout_1877_port);
   DataPath_RF_BLOCKi_66_Q_reg_20_inst : DFF_X1 port map( D => n5664, CK => CLK
                           , Q => n_2880, QN => 
                           DataPath_RF_bus_reg_dataout_1876_port);
   DataPath_RF_BLOCKi_66_Q_reg_19_inst : DFF_X1 port map( D => n5665, CK => CLK
                           , Q => n_2881, QN => 
                           DataPath_RF_bus_reg_dataout_1875_port);
   DataPath_RF_BLOCKi_66_Q_reg_18_inst : DFF_X1 port map( D => n5666, CK => CLK
                           , Q => n_2882, QN => 
                           DataPath_RF_bus_reg_dataout_1874_port);
   DataPath_RF_BLOCKi_66_Q_reg_17_inst : DFF_X1 port map( D => n5667, CK => CLK
                           , Q => n_2883, QN => 
                           DataPath_RF_bus_reg_dataout_1873_port);
   DataPath_RF_BLOCKi_66_Q_reg_16_inst : DFF_X1 port map( D => n5668, CK => CLK
                           , Q => n_2884, QN => 
                           DataPath_RF_bus_reg_dataout_1872_port);
   DataPath_RF_BLOCKi_66_Q_reg_15_inst : DFF_X1 port map( D => n5669, CK => CLK
                           , Q => n_2885, QN => 
                           DataPath_RF_bus_reg_dataout_1871_port);
   DataPath_RF_BLOCKi_66_Q_reg_14_inst : DFF_X1 port map( D => n5670, CK => CLK
                           , Q => n_2886, QN => 
                           DataPath_RF_bus_reg_dataout_1870_port);
   DataPath_RF_BLOCKi_66_Q_reg_13_inst : DFF_X1 port map( D => n5671, CK => CLK
                           , Q => n_2887, QN => 
                           DataPath_RF_bus_reg_dataout_1869_port);
   DataPath_RF_BLOCKi_66_Q_reg_12_inst : DFF_X1 port map( D => n5672, CK => CLK
                           , Q => n_2888, QN => 
                           DataPath_RF_bus_reg_dataout_1868_port);
   DataPath_RF_BLOCKi_66_Q_reg_11_inst : DFF_X1 port map( D => n5673, CK => CLK
                           , Q => n_2889, QN => 
                           DataPath_RF_bus_reg_dataout_1867_port);
   DataPath_RF_BLOCKi_66_Q_reg_9_inst : DFF_X1 port map( D => n5675, CK => CLK,
                           Q => n_2890, QN => 
                           DataPath_RF_bus_reg_dataout_1865_port);
   DataPath_RF_BLOCKi_66_Q_reg_8_inst : DFF_X1 port map( D => n5676, CK => CLK,
                           Q => n_2891, QN => 
                           DataPath_RF_bus_reg_dataout_1864_port);
   DataPath_RF_BLOCKi_66_Q_reg_7_inst : DFF_X1 port map( D => n5677, CK => CLK,
                           Q => n_2892, QN => 
                           DataPath_RF_bus_reg_dataout_1863_port);
   DataPath_RF_BLOCKi_66_Q_reg_6_inst : DFF_X1 port map( D => n5678, CK => CLK,
                           Q => n_2893, QN => 
                           DataPath_RF_bus_reg_dataout_1862_port);
   DataPath_RF_BLOCKi_66_Q_reg_5_inst : DFF_X1 port map( D => n5679, CK => CLK,
                           Q => n_2894, QN => 
                           DataPath_RF_bus_reg_dataout_1861_port);
   DataPath_RF_BLOCKi_66_Q_reg_4_inst : DFF_X1 port map( D => n5680, CK => CLK,
                           Q => n_2895, QN => 
                           DataPath_RF_bus_reg_dataout_1860_port);
   DataPath_RF_BLOCKi_66_Q_reg_3_inst : DFF_X1 port map( D => n5681, CK => CLK,
                           Q => n_2896, QN => 
                           DataPath_RF_bus_reg_dataout_1859_port);
   DataPath_RF_BLOCKi_66_Q_reg_2_inst : DFF_X1 port map( D => n5682, CK => CLK,
                           Q => n_2897, QN => 
                           DataPath_RF_bus_reg_dataout_1858_port);
   DataPath_RF_BLOCKi_66_Q_reg_1_inst : DFF_X1 port map( D => n5683, CK => CLK,
                           Q => n_2898, QN => 
                           DataPath_RF_bus_reg_dataout_1857_port);
   DataPath_RF_BLOCKi_66_Q_reg_0_inst : DFF_X1 port map( D => n5684, CK => CLK,
                           Q => n_2899, QN => 
                           DataPath_RF_bus_reg_dataout_1856_port);
   DataPath_RF_BLOCKi_83_Q_reg_31_inst : DFF_X1 port map( D => n1040, CK => CLK
                           , Q => n_2900, QN => 
                           DataPath_RF_bus_reg_dataout_2431_port);
   DataPath_RF_BLOCKi_83_Q_reg_30_inst : DFF_X1 port map( D => n1043, CK => CLK
                           , Q => n_2901, QN => 
                           DataPath_RF_bus_reg_dataout_2430_port);
   DataPath_RF_BLOCKi_83_Q_reg_29_inst : DFF_X1 port map( D => n1044, CK => CLK
                           , Q => n_2902, QN => 
                           DataPath_RF_bus_reg_dataout_2429_port);
   DataPath_RF_BLOCKi_83_Q_reg_28_inst : DFF_X1 port map( D => n1045, CK => CLK
                           , Q => n_2903, QN => 
                           DataPath_RF_bus_reg_dataout_2428_port);
   DataPath_RF_BLOCKi_83_Q_reg_27_inst : DFF_X1 port map( D => n1046, CK => CLK
                           , Q => n_2904, QN => 
                           DataPath_RF_bus_reg_dataout_2427_port);
   DataPath_RF_BLOCKi_83_Q_reg_26_inst : DFF_X1 port map( D => n1047, CK => CLK
                           , Q => n_2905, QN => 
                           DataPath_RF_bus_reg_dataout_2426_port);
   DataPath_RF_BLOCKi_83_Q_reg_25_inst : DFF_X1 port map( D => n1048, CK => CLK
                           , Q => n_2906, QN => 
                           DataPath_RF_bus_reg_dataout_2425_port);
   DataPath_RF_BLOCKi_83_Q_reg_24_inst : DFF_X1 port map( D => n1049, CK => CLK
                           , Q => n_2907, QN => 
                           DataPath_RF_bus_reg_dataout_2424_port);
   DataPath_RF_BLOCKi_83_Q_reg_23_inst : DFF_X1 port map( D => n1050, CK => CLK
                           , Q => n_2908, QN => 
                           DataPath_RF_bus_reg_dataout_2423_port);
   DataPath_RF_BLOCKi_83_Q_reg_22_inst : DFF_X1 port map( D => n1051, CK => CLK
                           , Q => n_2909, QN => 
                           DataPath_RF_bus_reg_dataout_2422_port);
   DataPath_RF_BLOCKi_83_Q_reg_21_inst : DFF_X1 port map( D => n1052, CK => CLK
                           , Q => n_2910, QN => 
                           DataPath_RF_bus_reg_dataout_2421_port);
   DataPath_RF_BLOCKi_83_Q_reg_20_inst : DFF_X1 port map( D => n1053, CK => CLK
                           , Q => n_2911, QN => 
                           DataPath_RF_bus_reg_dataout_2420_port);
   DataPath_RF_BLOCKi_83_Q_reg_19_inst : DFF_X1 port map( D => n1054, CK => CLK
                           , Q => n_2912, QN => 
                           DataPath_RF_bus_reg_dataout_2419_port);
   DataPath_RF_BLOCKi_83_Q_reg_18_inst : DFF_X1 port map( D => n1055, CK => CLK
                           , Q => n_2913, QN => 
                           DataPath_RF_bus_reg_dataout_2418_port);
   DataPath_RF_BLOCKi_83_Q_reg_17_inst : DFF_X1 port map( D => n1056, CK => CLK
                           , Q => n_2914, QN => 
                           DataPath_RF_bus_reg_dataout_2417_port);
   DataPath_RF_BLOCKi_83_Q_reg_16_inst : DFF_X1 port map( D => n1057, CK => CLK
                           , Q => n_2915, QN => 
                           DataPath_RF_bus_reg_dataout_2416_port);
   DataPath_RF_BLOCKi_83_Q_reg_15_inst : DFF_X1 port map( D => n1058, CK => CLK
                           , Q => n_2916, QN => 
                           DataPath_RF_bus_reg_dataout_2415_port);
   DataPath_RF_BLOCKi_83_Q_reg_14_inst : DFF_X1 port map( D => n1059, CK => CLK
                           , Q => n_2917, QN => 
                           DataPath_RF_bus_reg_dataout_2414_port);
   DataPath_RF_BLOCKi_83_Q_reg_13_inst : DFF_X1 port map( D => n1060, CK => CLK
                           , Q => n_2918, QN => 
                           DataPath_RF_bus_reg_dataout_2413_port);
   DataPath_RF_BLOCKi_83_Q_reg_12_inst : DFF_X1 port map( D => n1061, CK => CLK
                           , Q => n_2919, QN => 
                           DataPath_RF_bus_reg_dataout_2412_port);
   DataPath_RF_BLOCKi_83_Q_reg_11_inst : DFF_X1 port map( D => n1062, CK => CLK
                           , Q => n_2920, QN => 
                           DataPath_RF_bus_reg_dataout_2411_port);
   DataPath_RF_BLOCKi_83_Q_reg_9_inst : DFF_X1 port map( D => n1064, CK => CLK,
                           Q => n_2921, QN => 
                           DataPath_RF_bus_reg_dataout_2409_port);
   DataPath_RF_BLOCKi_83_Q_reg_8_inst : DFF_X1 port map( D => n1065, CK => CLK,
                           Q => n_2922, QN => 
                           DataPath_RF_bus_reg_dataout_2408_port);
   DataPath_RF_BLOCKi_83_Q_reg_7_inst : DFF_X1 port map( D => n1066, CK => CLK,
                           Q => n_2923, QN => 
                           DataPath_RF_bus_reg_dataout_2407_port);
   DataPath_RF_BLOCKi_83_Q_reg_6_inst : DFF_X1 port map( D => n1067, CK => CLK,
                           Q => n_2924, QN => 
                           DataPath_RF_bus_reg_dataout_2406_port);
   DataPath_RF_BLOCKi_83_Q_reg_5_inst : DFF_X1 port map( D => n1068, CK => CLK,
                           Q => n_2925, QN => 
                           DataPath_RF_bus_reg_dataout_2405_port);
   DataPath_RF_BLOCKi_83_Q_reg_4_inst : DFF_X1 port map( D => n1069, CK => CLK,
                           Q => n_2926, QN => 
                           DataPath_RF_bus_reg_dataout_2404_port);
   DataPath_RF_BLOCKi_83_Q_reg_3_inst : DFF_X1 port map( D => n1070, CK => CLK,
                           Q => n_2927, QN => 
                           DataPath_RF_bus_reg_dataout_2403_port);
   DataPath_RF_BLOCKi_83_Q_reg_2_inst : DFF_X1 port map( D => n1071, CK => CLK,
                           Q => n_2928, QN => 
                           DataPath_RF_bus_reg_dataout_2402_port);
   DataPath_RF_BLOCKi_83_Q_reg_1_inst : DFF_X1 port map( D => n1072, CK => CLK,
                           Q => n_2929, QN => 
                           DataPath_RF_bus_reg_dataout_2401_port);
   DataPath_RF_BLOCKi_83_Q_reg_0_inst : DFF_X1 port map( D => n1073, CK => CLK,
                           Q => n_2930, QN => 
                           DataPath_RF_bus_reg_dataout_2400_port);
   DataPath_RF_BLOCKi_19_Q_reg_31_inst : DFF_X1 port map( D => n3870, CK => CLK
                           , Q => n_2931, QN => 
                           DataPath_RF_bus_reg_dataout_383_port);
   DataPath_RF_BLOCKi_19_Q_reg_30_inst : DFF_X1 port map( D => n3873, CK => CLK
                           , Q => n_2932, QN => 
                           DataPath_RF_bus_reg_dataout_382_port);
   DataPath_RF_BLOCKi_19_Q_reg_29_inst : DFF_X1 port map( D => n3874, CK => CLK
                           , Q => n_2933, QN => 
                           DataPath_RF_bus_reg_dataout_381_port);
   DataPath_RF_BLOCKi_19_Q_reg_28_inst : DFF_X1 port map( D => n3875, CK => CLK
                           , Q => n_2934, QN => 
                           DataPath_RF_bus_reg_dataout_380_port);
   DataPath_RF_BLOCKi_19_Q_reg_27_inst : DFF_X1 port map( D => n3876, CK => CLK
                           , Q => n_2935, QN => 
                           DataPath_RF_bus_reg_dataout_379_port);
   DataPath_RF_BLOCKi_19_Q_reg_26_inst : DFF_X1 port map( D => n3877, CK => CLK
                           , Q => n_2936, QN => 
                           DataPath_RF_bus_reg_dataout_378_port);
   DataPath_RF_BLOCKi_19_Q_reg_25_inst : DFF_X1 port map( D => n3878, CK => CLK
                           , Q => n_2937, QN => 
                           DataPath_RF_bus_reg_dataout_377_port);
   DataPath_RF_BLOCKi_19_Q_reg_24_inst : DFF_X1 port map( D => n3879, CK => CLK
                           , Q => n_2938, QN => 
                           DataPath_RF_bus_reg_dataout_376_port);
   DataPath_RF_BLOCKi_19_Q_reg_23_inst : DFF_X1 port map( D => n3880, CK => CLK
                           , Q => n_2939, QN => 
                           DataPath_RF_bus_reg_dataout_375_port);
   DataPath_RF_BLOCKi_19_Q_reg_22_inst : DFF_X1 port map( D => n3881, CK => CLK
                           , Q => n_2940, QN => 
                           DataPath_RF_bus_reg_dataout_374_port);
   DataPath_RF_BLOCKi_19_Q_reg_21_inst : DFF_X1 port map( D => n3882, CK => CLK
                           , Q => n_2941, QN => 
                           DataPath_RF_bus_reg_dataout_373_port);
   DataPath_RF_BLOCKi_19_Q_reg_20_inst : DFF_X1 port map( D => n3883, CK => CLK
                           , Q => n_2942, QN => 
                           DataPath_RF_bus_reg_dataout_372_port);
   DataPath_RF_BLOCKi_19_Q_reg_19_inst : DFF_X1 port map( D => n3884, CK => CLK
                           , Q => n_2943, QN => 
                           DataPath_RF_bus_reg_dataout_371_port);
   DataPath_RF_BLOCKi_19_Q_reg_18_inst : DFF_X1 port map( D => n3885, CK => CLK
                           , Q => n_2944, QN => 
                           DataPath_RF_bus_reg_dataout_370_port);
   DataPath_RF_BLOCKi_19_Q_reg_17_inst : DFF_X1 port map( D => n3886, CK => CLK
                           , Q => n_2945, QN => 
                           DataPath_RF_bus_reg_dataout_369_port);
   DataPath_RF_BLOCKi_19_Q_reg_16_inst : DFF_X1 port map( D => n3887, CK => CLK
                           , Q => n_2946, QN => 
                           DataPath_RF_bus_reg_dataout_368_port);
   DataPath_RF_BLOCKi_19_Q_reg_15_inst : DFF_X1 port map( D => n3888, CK => CLK
                           , Q => n_2947, QN => 
                           DataPath_RF_bus_reg_dataout_367_port);
   DataPath_RF_BLOCKi_19_Q_reg_14_inst : DFF_X1 port map( D => n3889, CK => CLK
                           , Q => n_2948, QN => 
                           DataPath_RF_bus_reg_dataout_366_port);
   DataPath_RF_BLOCKi_19_Q_reg_13_inst : DFF_X1 port map( D => n3890, CK => CLK
                           , Q => n_2949, QN => 
                           DataPath_RF_bus_reg_dataout_365_port);
   DataPath_RF_BLOCKi_19_Q_reg_12_inst : DFF_X1 port map( D => n3891, CK => CLK
                           , Q => n_2950, QN => 
                           DataPath_RF_bus_reg_dataout_364_port);
   DataPath_RF_BLOCKi_19_Q_reg_11_inst : DFF_X1 port map( D => n3892, CK => CLK
                           , Q => n_2951, QN => 
                           DataPath_RF_bus_reg_dataout_363_port);
   DataPath_RF_BLOCKi_19_Q_reg_9_inst : DFF_X1 port map( D => n3894, CK => CLK,
                           Q => n_2952, QN => 
                           DataPath_RF_bus_reg_dataout_361_port);
   DataPath_RF_BLOCKi_19_Q_reg_8_inst : DFF_X1 port map( D => n3895, CK => CLK,
                           Q => n_2953, QN => 
                           DataPath_RF_bus_reg_dataout_360_port);
   DataPath_RF_BLOCKi_19_Q_reg_7_inst : DFF_X1 port map( D => n3896, CK => CLK,
                           Q => n_2954, QN => 
                           DataPath_RF_bus_reg_dataout_359_port);
   DataPath_RF_BLOCKi_19_Q_reg_6_inst : DFF_X1 port map( D => n3897, CK => CLK,
                           Q => n_2955, QN => 
                           DataPath_RF_bus_reg_dataout_358_port);
   DataPath_RF_BLOCKi_19_Q_reg_5_inst : DFF_X1 port map( D => n3898, CK => CLK,
                           Q => n_2956, QN => 
                           DataPath_RF_bus_reg_dataout_357_port);
   DataPath_RF_BLOCKi_19_Q_reg_4_inst : DFF_X1 port map( D => n3899, CK => CLK,
                           Q => n_2957, QN => 
                           DataPath_RF_bus_reg_dataout_356_port);
   DataPath_RF_BLOCKi_19_Q_reg_3_inst : DFF_X1 port map( D => n3900, CK => CLK,
                           Q => n_2958, QN => 
                           DataPath_RF_bus_reg_dataout_355_port);
   DataPath_RF_BLOCKi_19_Q_reg_2_inst : DFF_X1 port map( D => n3901, CK => CLK,
                           Q => n_2959, QN => 
                           DataPath_RF_bus_reg_dataout_354_port);
   DataPath_RF_BLOCKi_19_Q_reg_1_inst : DFF_X1 port map( D => n3902, CK => CLK,
                           Q => n_2960, QN => 
                           DataPath_RF_bus_reg_dataout_353_port);
   DataPath_RF_BLOCKi_19_Q_reg_0_inst : DFF_X1 port map( D => n3903, CK => CLK,
                           Q => n_2961, QN => 
                           DataPath_RF_bus_reg_dataout_352_port);
   DataPath_RF_BLOCKi_35_Q_reg_31_inst : DFF_X1 port map( D => n4495, CK => CLK
                           , Q => n_2962, QN => 
                           DataPath_RF_bus_reg_dataout_895_port);
   DataPath_RF_BLOCKi_35_Q_reg_30_inst : DFF_X1 port map( D => n4498, CK => CLK
                           , Q => n_2963, QN => 
                           DataPath_RF_bus_reg_dataout_894_port);
   DataPath_RF_BLOCKi_35_Q_reg_29_inst : DFF_X1 port map( D => n4499, CK => CLK
                           , Q => n_2964, QN => 
                           DataPath_RF_bus_reg_dataout_893_port);
   DataPath_RF_BLOCKi_35_Q_reg_28_inst : DFF_X1 port map( D => n4500, CK => CLK
                           , Q => n_2965, QN => 
                           DataPath_RF_bus_reg_dataout_892_port);
   DataPath_RF_BLOCKi_35_Q_reg_27_inst : DFF_X1 port map( D => n4501, CK => CLK
                           , Q => n_2966, QN => 
                           DataPath_RF_bus_reg_dataout_891_port);
   DataPath_RF_BLOCKi_35_Q_reg_26_inst : DFF_X1 port map( D => n4502, CK => CLK
                           , Q => n_2967, QN => 
                           DataPath_RF_bus_reg_dataout_890_port);
   DataPath_RF_BLOCKi_35_Q_reg_25_inst : DFF_X1 port map( D => n4503, CK => CLK
                           , Q => n_2968, QN => 
                           DataPath_RF_bus_reg_dataout_889_port);
   DataPath_RF_BLOCKi_35_Q_reg_24_inst : DFF_X1 port map( D => n4504, CK => CLK
                           , Q => n_2969, QN => 
                           DataPath_RF_bus_reg_dataout_888_port);
   DataPath_RF_BLOCKi_35_Q_reg_23_inst : DFF_X1 port map( D => n4505, CK => CLK
                           , Q => n_2970, QN => 
                           DataPath_RF_bus_reg_dataout_887_port);
   DataPath_RF_BLOCKi_35_Q_reg_22_inst : DFF_X1 port map( D => n4506, CK => CLK
                           , Q => n_2971, QN => 
                           DataPath_RF_bus_reg_dataout_886_port);
   DataPath_RF_BLOCKi_35_Q_reg_21_inst : DFF_X1 port map( D => n4507, CK => CLK
                           , Q => n_2972, QN => 
                           DataPath_RF_bus_reg_dataout_885_port);
   DataPath_RF_BLOCKi_35_Q_reg_20_inst : DFF_X1 port map( D => n4508, CK => CLK
                           , Q => n_2973, QN => 
                           DataPath_RF_bus_reg_dataout_884_port);
   DataPath_RF_BLOCKi_35_Q_reg_19_inst : DFF_X1 port map( D => n4509, CK => CLK
                           , Q => n_2974, QN => 
                           DataPath_RF_bus_reg_dataout_883_port);
   DataPath_RF_BLOCKi_35_Q_reg_18_inst : DFF_X1 port map( D => n4510, CK => CLK
                           , Q => n_2975, QN => 
                           DataPath_RF_bus_reg_dataout_882_port);
   DataPath_RF_BLOCKi_35_Q_reg_17_inst : DFF_X1 port map( D => n4511, CK => CLK
                           , Q => n_2976, QN => 
                           DataPath_RF_bus_reg_dataout_881_port);
   DataPath_RF_BLOCKi_35_Q_reg_16_inst : DFF_X1 port map( D => n4512, CK => CLK
                           , Q => n_2977, QN => 
                           DataPath_RF_bus_reg_dataout_880_port);
   DataPath_RF_BLOCKi_35_Q_reg_15_inst : DFF_X1 port map( D => n4513, CK => CLK
                           , Q => n_2978, QN => 
                           DataPath_RF_bus_reg_dataout_879_port);
   DataPath_RF_BLOCKi_35_Q_reg_14_inst : DFF_X1 port map( D => n4514, CK => CLK
                           , Q => n_2979, QN => 
                           DataPath_RF_bus_reg_dataout_878_port);
   DataPath_RF_BLOCKi_35_Q_reg_13_inst : DFF_X1 port map( D => n4515, CK => CLK
                           , Q => n_2980, QN => 
                           DataPath_RF_bus_reg_dataout_877_port);
   DataPath_RF_BLOCKi_35_Q_reg_12_inst : DFF_X1 port map( D => n4516, CK => CLK
                           , Q => n_2981, QN => 
                           DataPath_RF_bus_reg_dataout_876_port);
   DataPath_RF_BLOCKi_35_Q_reg_11_inst : DFF_X1 port map( D => n4517, CK => CLK
                           , Q => n_2982, QN => 
                           DataPath_RF_bus_reg_dataout_875_port);
   DataPath_RF_BLOCKi_35_Q_reg_9_inst : DFF_X1 port map( D => n4519, CK => CLK,
                           Q => n_2983, QN => 
                           DataPath_RF_bus_reg_dataout_873_port);
   DataPath_RF_BLOCKi_35_Q_reg_8_inst : DFF_X1 port map( D => n4520, CK => CLK,
                           Q => n_2984, QN => 
                           DataPath_RF_bus_reg_dataout_872_port);
   DataPath_RF_BLOCKi_35_Q_reg_7_inst : DFF_X1 port map( D => n4521, CK => CLK,
                           Q => n_2985, QN => 
                           DataPath_RF_bus_reg_dataout_871_port);
   DataPath_RF_BLOCKi_35_Q_reg_6_inst : DFF_X1 port map( D => n4522, CK => CLK,
                           Q => n_2986, QN => 
                           DataPath_RF_bus_reg_dataout_870_port);
   DataPath_RF_BLOCKi_35_Q_reg_5_inst : DFF_X1 port map( D => n4523, CK => CLK,
                           Q => n_2987, QN => 
                           DataPath_RF_bus_reg_dataout_869_port);
   DataPath_RF_BLOCKi_35_Q_reg_4_inst : DFF_X1 port map( D => n4524, CK => CLK,
                           Q => n_2988, QN => 
                           DataPath_RF_bus_reg_dataout_868_port);
   DataPath_RF_BLOCKi_35_Q_reg_3_inst : DFF_X1 port map( D => n4525, CK => CLK,
                           Q => n_2989, QN => 
                           DataPath_RF_bus_reg_dataout_867_port);
   DataPath_RF_BLOCKi_35_Q_reg_2_inst : DFF_X1 port map( D => n4526, CK => CLK,
                           Q => n_2990, QN => 
                           DataPath_RF_bus_reg_dataout_866_port);
   DataPath_RF_BLOCKi_35_Q_reg_1_inst : DFF_X1 port map( D => n4527, CK => CLK,
                           Q => n_2991, QN => 
                           DataPath_RF_bus_reg_dataout_865_port);
   DataPath_RF_BLOCKi_35_Q_reg_0_inst : DFF_X1 port map( D => n4528, CK => CLK,
                           Q => n_2992, QN => 
                           DataPath_RF_bus_reg_dataout_864_port);
   DataPath_RF_BLOCKi_51_Q_reg_31_inst : DFF_X1 port map( D => n5088, CK => CLK
                           , Q => n_2993, QN => 
                           DataPath_RF_bus_reg_dataout_1407_port);
   DataPath_RF_BLOCKi_51_Q_reg_30_inst : DFF_X1 port map( D => n5091, CK => CLK
                           , Q => n_2994, QN => 
                           DataPath_RF_bus_reg_dataout_1406_port);
   DataPath_RF_BLOCKi_51_Q_reg_29_inst : DFF_X1 port map( D => n5092, CK => CLK
                           , Q => n_2995, QN => 
                           DataPath_RF_bus_reg_dataout_1405_port);
   DataPath_RF_BLOCKi_51_Q_reg_28_inst : DFF_X1 port map( D => n5093, CK => CLK
                           , Q => n_2996, QN => 
                           DataPath_RF_bus_reg_dataout_1404_port);
   DataPath_RF_BLOCKi_51_Q_reg_27_inst : DFF_X1 port map( D => n5094, CK => CLK
                           , Q => n_2997, QN => 
                           DataPath_RF_bus_reg_dataout_1403_port);
   DataPath_RF_BLOCKi_51_Q_reg_26_inst : DFF_X1 port map( D => n5095, CK => CLK
                           , Q => n_2998, QN => 
                           DataPath_RF_bus_reg_dataout_1402_port);
   DataPath_RF_BLOCKi_51_Q_reg_25_inst : DFF_X1 port map( D => n5096, CK => CLK
                           , Q => n_2999, QN => 
                           DataPath_RF_bus_reg_dataout_1401_port);
   DataPath_RF_BLOCKi_51_Q_reg_24_inst : DFF_X1 port map( D => n5097, CK => CLK
                           , Q => n_3000, QN => 
                           DataPath_RF_bus_reg_dataout_1400_port);
   DataPath_RF_BLOCKi_51_Q_reg_23_inst : DFF_X1 port map( D => n5098, CK => CLK
                           , Q => n_3001, QN => 
                           DataPath_RF_bus_reg_dataout_1399_port);
   DataPath_RF_BLOCKi_51_Q_reg_22_inst : DFF_X1 port map( D => n5099, CK => CLK
                           , Q => n_3002, QN => 
                           DataPath_RF_bus_reg_dataout_1398_port);
   DataPath_RF_BLOCKi_51_Q_reg_21_inst : DFF_X1 port map( D => n5100, CK => CLK
                           , Q => n_3003, QN => 
                           DataPath_RF_bus_reg_dataout_1397_port);
   DataPath_RF_BLOCKi_51_Q_reg_20_inst : DFF_X1 port map( D => n5101, CK => CLK
                           , Q => n_3004, QN => 
                           DataPath_RF_bus_reg_dataout_1396_port);
   DataPath_RF_BLOCKi_51_Q_reg_19_inst : DFF_X1 port map( D => n5102, CK => CLK
                           , Q => n_3005, QN => 
                           DataPath_RF_bus_reg_dataout_1395_port);
   DataPath_RF_BLOCKi_51_Q_reg_18_inst : DFF_X1 port map( D => n5103, CK => CLK
                           , Q => n_3006, QN => 
                           DataPath_RF_bus_reg_dataout_1394_port);
   DataPath_RF_BLOCKi_51_Q_reg_17_inst : DFF_X1 port map( D => n5104, CK => CLK
                           , Q => n_3007, QN => 
                           DataPath_RF_bus_reg_dataout_1393_port);
   DataPath_RF_BLOCKi_51_Q_reg_16_inst : DFF_X1 port map( D => n5105, CK => CLK
                           , Q => n_3008, QN => 
                           DataPath_RF_bus_reg_dataout_1392_port);
   DataPath_RF_BLOCKi_51_Q_reg_15_inst : DFF_X1 port map( D => n5106, CK => CLK
                           , Q => n_3009, QN => 
                           DataPath_RF_bus_reg_dataout_1391_port);
   DataPath_RF_BLOCKi_51_Q_reg_14_inst : DFF_X1 port map( D => n5107, CK => CLK
                           , Q => n_3010, QN => 
                           DataPath_RF_bus_reg_dataout_1390_port);
   DataPath_RF_BLOCKi_51_Q_reg_13_inst : DFF_X1 port map( D => n5108, CK => CLK
                           , Q => n_3011, QN => 
                           DataPath_RF_bus_reg_dataout_1389_port);
   DataPath_RF_BLOCKi_51_Q_reg_12_inst : DFF_X1 port map( D => n5109, CK => CLK
                           , Q => n_3012, QN => 
                           DataPath_RF_bus_reg_dataout_1388_port);
   DataPath_RF_BLOCKi_51_Q_reg_11_inst : DFF_X1 port map( D => n5110, CK => CLK
                           , Q => n_3013, QN => 
                           DataPath_RF_bus_reg_dataout_1387_port);
   DataPath_RF_BLOCKi_51_Q_reg_9_inst : DFF_X1 port map( D => n5112, CK => CLK,
                           Q => n_3014, QN => 
                           DataPath_RF_bus_reg_dataout_1385_port);
   DataPath_RF_BLOCKi_51_Q_reg_8_inst : DFF_X1 port map( D => n5113, CK => CLK,
                           Q => n_3015, QN => 
                           DataPath_RF_bus_reg_dataout_1384_port);
   DataPath_RF_BLOCKi_51_Q_reg_7_inst : DFF_X1 port map( D => n5114, CK => CLK,
                           Q => n_3016, QN => 
                           DataPath_RF_bus_reg_dataout_1383_port);
   DataPath_RF_BLOCKi_51_Q_reg_6_inst : DFF_X1 port map( D => n5115, CK => CLK,
                           Q => n_3017, QN => 
                           DataPath_RF_bus_reg_dataout_1382_port);
   DataPath_RF_BLOCKi_51_Q_reg_5_inst : DFF_X1 port map( D => n5116, CK => CLK,
                           Q => n_3018, QN => 
                           DataPath_RF_bus_reg_dataout_1381_port);
   DataPath_RF_BLOCKi_51_Q_reg_4_inst : DFF_X1 port map( D => n5117, CK => CLK,
                           Q => n_3019, QN => 
                           DataPath_RF_bus_reg_dataout_1380_port);
   DataPath_RF_BLOCKi_51_Q_reg_3_inst : DFF_X1 port map( D => n5118, CK => CLK,
                           Q => n_3020, QN => 
                           DataPath_RF_bus_reg_dataout_1379_port);
   DataPath_RF_BLOCKi_51_Q_reg_2_inst : DFF_X1 port map( D => n5119, CK => CLK,
                           Q => n_3021, QN => 
                           DataPath_RF_bus_reg_dataout_1378_port);
   DataPath_RF_BLOCKi_51_Q_reg_1_inst : DFF_X1 port map( D => n5120, CK => CLK,
                           Q => n_3022, QN => 
                           DataPath_RF_bus_reg_dataout_1377_port);
   DataPath_RF_BLOCKi_51_Q_reg_0_inst : DFF_X1 port map( D => n5121, CK => CLK,
                           Q => n_3023, QN => 
                           DataPath_RF_bus_reg_dataout_1376_port);
   DataPath_RF_BLOCKi_67_Q_reg_31_inst : DFF_X1 port map( D => n5687, CK => CLK
                           , Q => n_3024, QN => 
                           DataPath_RF_bus_reg_dataout_1919_port);
   DataPath_RF_BLOCKi_67_Q_reg_30_inst : DFF_X1 port map( D => n5690, CK => CLK
                           , Q => n_3025, QN => 
                           DataPath_RF_bus_reg_dataout_1918_port);
   DataPath_RF_BLOCKi_67_Q_reg_29_inst : DFF_X1 port map( D => n5691, CK => CLK
                           , Q => n_3026, QN => 
                           DataPath_RF_bus_reg_dataout_1917_port);
   DataPath_RF_BLOCKi_67_Q_reg_28_inst : DFF_X1 port map( D => n5692, CK => CLK
                           , Q => n_3027, QN => 
                           DataPath_RF_bus_reg_dataout_1916_port);
   DataPath_RF_BLOCKi_67_Q_reg_27_inst : DFF_X1 port map( D => n5693, CK => CLK
                           , Q => n_3028, QN => 
                           DataPath_RF_bus_reg_dataout_1915_port);
   DataPath_RF_BLOCKi_67_Q_reg_26_inst : DFF_X1 port map( D => n5694, CK => CLK
                           , Q => n_3029, QN => 
                           DataPath_RF_bus_reg_dataout_1914_port);
   DataPath_RF_BLOCKi_67_Q_reg_25_inst : DFF_X1 port map( D => n5695, CK => CLK
                           , Q => n_3030, QN => 
                           DataPath_RF_bus_reg_dataout_1913_port);
   DataPath_RF_BLOCKi_67_Q_reg_24_inst : DFF_X1 port map( D => n5696, CK => CLK
                           , Q => n_3031, QN => 
                           DataPath_RF_bus_reg_dataout_1912_port);
   DataPath_RF_BLOCKi_67_Q_reg_23_inst : DFF_X1 port map( D => n5697, CK => CLK
                           , Q => n_3032, QN => 
                           DataPath_RF_bus_reg_dataout_1911_port);
   DataPath_RF_BLOCKi_67_Q_reg_22_inst : DFF_X1 port map( D => n5698, CK => CLK
                           , Q => n_3033, QN => 
                           DataPath_RF_bus_reg_dataout_1910_port);
   DataPath_RF_BLOCKi_67_Q_reg_21_inst : DFF_X1 port map( D => n5699, CK => CLK
                           , Q => n_3034, QN => 
                           DataPath_RF_bus_reg_dataout_1909_port);
   DataPath_RF_BLOCKi_67_Q_reg_20_inst : DFF_X1 port map( D => n5700, CK => CLK
                           , Q => n_3035, QN => 
                           DataPath_RF_bus_reg_dataout_1908_port);
   DataPath_RF_BLOCKi_67_Q_reg_19_inst : DFF_X1 port map( D => n5701, CK => CLK
                           , Q => n_3036, QN => 
                           DataPath_RF_bus_reg_dataout_1907_port);
   DataPath_RF_BLOCKi_67_Q_reg_18_inst : DFF_X1 port map( D => n5702, CK => CLK
                           , Q => n_3037, QN => 
                           DataPath_RF_bus_reg_dataout_1906_port);
   DataPath_RF_BLOCKi_67_Q_reg_17_inst : DFF_X1 port map( D => n5703, CK => CLK
                           , Q => n_3038, QN => 
                           DataPath_RF_bus_reg_dataout_1905_port);
   DataPath_RF_BLOCKi_67_Q_reg_16_inst : DFF_X1 port map( D => n5704, CK => CLK
                           , Q => n_3039, QN => 
                           DataPath_RF_bus_reg_dataout_1904_port);
   DataPath_RF_BLOCKi_67_Q_reg_15_inst : DFF_X1 port map( D => n5705, CK => CLK
                           , Q => n_3040, QN => 
                           DataPath_RF_bus_reg_dataout_1903_port);
   DataPath_RF_BLOCKi_67_Q_reg_14_inst : DFF_X1 port map( D => n5706, CK => CLK
                           , Q => n_3041, QN => 
                           DataPath_RF_bus_reg_dataout_1902_port);
   DataPath_RF_BLOCKi_67_Q_reg_13_inst : DFF_X1 port map( D => n5707, CK => CLK
                           , Q => n_3042, QN => 
                           DataPath_RF_bus_reg_dataout_1901_port);
   DataPath_RF_BLOCKi_67_Q_reg_12_inst : DFF_X1 port map( D => n5708, CK => CLK
                           , Q => n_3043, QN => 
                           DataPath_RF_bus_reg_dataout_1900_port);
   DataPath_RF_BLOCKi_67_Q_reg_11_inst : DFF_X1 port map( D => n5709, CK => CLK
                           , Q => n_3044, QN => 
                           DataPath_RF_bus_reg_dataout_1899_port);
   DataPath_RF_BLOCKi_67_Q_reg_9_inst : DFF_X1 port map( D => n5711, CK => CLK,
                           Q => n_3045, QN => 
                           DataPath_RF_bus_reg_dataout_1897_port);
   DataPath_RF_BLOCKi_67_Q_reg_8_inst : DFF_X1 port map( D => n5712, CK => CLK,
                           Q => n_3046, QN => 
                           DataPath_RF_bus_reg_dataout_1896_port);
   DataPath_RF_BLOCKi_67_Q_reg_7_inst : DFF_X1 port map( D => n5713, CK => CLK,
                           Q => n_3047, QN => 
                           DataPath_RF_bus_reg_dataout_1895_port);
   DataPath_RF_BLOCKi_67_Q_reg_6_inst : DFF_X1 port map( D => n5714, CK => CLK,
                           Q => n_3048, QN => 
                           DataPath_RF_bus_reg_dataout_1894_port);
   DataPath_RF_BLOCKi_67_Q_reg_5_inst : DFF_X1 port map( D => n5715, CK => CLK,
                           Q => n_3049, QN => 
                           DataPath_RF_bus_reg_dataout_1893_port);
   DataPath_RF_BLOCKi_67_Q_reg_4_inst : DFF_X1 port map( D => n5716, CK => CLK,
                           Q => n_3050, QN => 
                           DataPath_RF_bus_reg_dataout_1892_port);
   DataPath_RF_BLOCKi_67_Q_reg_3_inst : DFF_X1 port map( D => n5717, CK => CLK,
                           Q => n_3051, QN => 
                           DataPath_RF_bus_reg_dataout_1891_port);
   DataPath_RF_BLOCKi_67_Q_reg_2_inst : DFF_X1 port map( D => n5718, CK => CLK,
                           Q => n_3052, QN => 
                           DataPath_RF_bus_reg_dataout_1890_port);
   DataPath_RF_BLOCKi_67_Q_reg_1_inst : DFF_X1 port map( D => n5719, CK => CLK,
                           Q => n_3053, QN => 
                           DataPath_RF_bus_reg_dataout_1889_port);
   DataPath_RF_BLOCKi_67_Q_reg_0_inst : DFF_X1 port map( D => n5720, CK => CLK,
                           Q => n_3054, QN => 
                           DataPath_RF_bus_reg_dataout_1888_port);
   DataPath_RF_BLOCKi_84_Q_reg_31_inst : DFF_X1 port map( D => n1077, CK => CLK
                           , Q => n_3055, QN => 
                           DataPath_RF_bus_reg_dataout_2463_port);
   DataPath_RF_BLOCKi_84_Q_reg_30_inst : DFF_X1 port map( D => n1080, CK => CLK
                           , Q => n_3056, QN => 
                           DataPath_RF_bus_reg_dataout_2462_port);
   DataPath_RF_BLOCKi_84_Q_reg_29_inst : DFF_X1 port map( D => n1081, CK => CLK
                           , Q => n_3057, QN => 
                           DataPath_RF_bus_reg_dataout_2461_port);
   DataPath_RF_BLOCKi_84_Q_reg_28_inst : DFF_X1 port map( D => n1082, CK => CLK
                           , Q => n_3058, QN => 
                           DataPath_RF_bus_reg_dataout_2460_port);
   DataPath_RF_BLOCKi_84_Q_reg_27_inst : DFF_X1 port map( D => n1083, CK => CLK
                           , Q => n_3059, QN => 
                           DataPath_RF_bus_reg_dataout_2459_port);
   DataPath_RF_BLOCKi_84_Q_reg_26_inst : DFF_X1 port map( D => n1084, CK => CLK
                           , Q => n_3060, QN => 
                           DataPath_RF_bus_reg_dataout_2458_port);
   DataPath_RF_BLOCKi_84_Q_reg_25_inst : DFF_X1 port map( D => n1085, CK => CLK
                           , Q => n_3061, QN => 
                           DataPath_RF_bus_reg_dataout_2457_port);
   DataPath_RF_BLOCKi_84_Q_reg_24_inst : DFF_X1 port map( D => n1086, CK => CLK
                           , Q => n_3062, QN => 
                           DataPath_RF_bus_reg_dataout_2456_port);
   DataPath_RF_BLOCKi_84_Q_reg_23_inst : DFF_X1 port map( D => n1087, CK => CLK
                           , Q => n_3063, QN => 
                           DataPath_RF_bus_reg_dataout_2455_port);
   DataPath_RF_BLOCKi_84_Q_reg_22_inst : DFF_X1 port map( D => n1088, CK => CLK
                           , Q => n_3064, QN => 
                           DataPath_RF_bus_reg_dataout_2454_port);
   DataPath_RF_BLOCKi_84_Q_reg_21_inst : DFF_X1 port map( D => n1089, CK => CLK
                           , Q => n_3065, QN => 
                           DataPath_RF_bus_reg_dataout_2453_port);
   DataPath_RF_BLOCKi_84_Q_reg_20_inst : DFF_X1 port map( D => n1090, CK => CLK
                           , Q => n_3066, QN => 
                           DataPath_RF_bus_reg_dataout_2452_port);
   DataPath_RF_BLOCKi_84_Q_reg_19_inst : DFF_X1 port map( D => n1091, CK => CLK
                           , Q => n_3067, QN => 
                           DataPath_RF_bus_reg_dataout_2451_port);
   DataPath_RF_BLOCKi_84_Q_reg_18_inst : DFF_X1 port map( D => n1092, CK => CLK
                           , Q => n_3068, QN => 
                           DataPath_RF_bus_reg_dataout_2450_port);
   DataPath_RF_BLOCKi_84_Q_reg_17_inst : DFF_X1 port map( D => n1093, CK => CLK
                           , Q => n_3069, QN => 
                           DataPath_RF_bus_reg_dataout_2449_port);
   DataPath_RF_BLOCKi_84_Q_reg_16_inst : DFF_X1 port map( D => n1094, CK => CLK
                           , Q => n_3070, QN => 
                           DataPath_RF_bus_reg_dataout_2448_port);
   DataPath_RF_BLOCKi_84_Q_reg_15_inst : DFF_X1 port map( D => n1095, CK => CLK
                           , Q => n_3071, QN => 
                           DataPath_RF_bus_reg_dataout_2447_port);
   DataPath_RF_BLOCKi_84_Q_reg_14_inst : DFF_X1 port map( D => n1096, CK => CLK
                           , Q => n_3072, QN => 
                           DataPath_RF_bus_reg_dataout_2446_port);
   DataPath_RF_BLOCKi_84_Q_reg_13_inst : DFF_X1 port map( D => n1097, CK => CLK
                           , Q => n_3073, QN => 
                           DataPath_RF_bus_reg_dataout_2445_port);
   DataPath_RF_BLOCKi_84_Q_reg_12_inst : DFF_X1 port map( D => n1098, CK => CLK
                           , Q => n_3074, QN => 
                           DataPath_RF_bus_reg_dataout_2444_port);
   DataPath_RF_BLOCKi_84_Q_reg_11_inst : DFF_X1 port map( D => n1099, CK => CLK
                           , Q => n_3075, QN => 
                           DataPath_RF_bus_reg_dataout_2443_port);
   DataPath_RF_BLOCKi_84_Q_reg_9_inst : DFF_X1 port map( D => n1101, CK => CLK,
                           Q => n_3076, QN => 
                           DataPath_RF_bus_reg_dataout_2441_port);
   DataPath_RF_BLOCKi_84_Q_reg_8_inst : DFF_X1 port map( D => n1102, CK => CLK,
                           Q => n_3077, QN => 
                           DataPath_RF_bus_reg_dataout_2440_port);
   DataPath_RF_BLOCKi_84_Q_reg_7_inst : DFF_X1 port map( D => n1103, CK => CLK,
                           Q => n_3078, QN => 
                           DataPath_RF_bus_reg_dataout_2439_port);
   DataPath_RF_BLOCKi_84_Q_reg_6_inst : DFF_X1 port map( D => n1104, CK => CLK,
                           Q => n_3079, QN => 
                           DataPath_RF_bus_reg_dataout_2438_port);
   DataPath_RF_BLOCKi_84_Q_reg_5_inst : DFF_X1 port map( D => n1105, CK => CLK,
                           Q => n_3080, QN => 
                           DataPath_RF_bus_reg_dataout_2437_port);
   DataPath_RF_BLOCKi_84_Q_reg_4_inst : DFF_X1 port map( D => n1106, CK => CLK,
                           Q => n_3081, QN => 
                           DataPath_RF_bus_reg_dataout_2436_port);
   DataPath_RF_BLOCKi_84_Q_reg_3_inst : DFF_X1 port map( D => n1107, CK => CLK,
                           Q => n_3082, QN => 
                           DataPath_RF_bus_reg_dataout_2435_port);
   DataPath_RF_BLOCKi_84_Q_reg_2_inst : DFF_X1 port map( D => n1108, CK => CLK,
                           Q => n_3083, QN => 
                           DataPath_RF_bus_reg_dataout_2434_port);
   DataPath_RF_BLOCKi_84_Q_reg_1_inst : DFF_X1 port map( D => n1109, CK => CLK,
                           Q => n_3084, QN => 
                           DataPath_RF_bus_reg_dataout_2433_port);
   DataPath_RF_BLOCKi_84_Q_reg_0_inst : DFF_X1 port map( D => n1110, CK => CLK,
                           Q => n_3085, QN => 
                           DataPath_RF_bus_reg_dataout_2432_port);
   DataPath_RF_BLOCKi_20_Q_reg_31_inst : DFF_X1 port map( D => n3905, CK => CLK
                           , Q => n_3086, QN => 
                           DataPath_RF_bus_reg_dataout_415_port);
   DataPath_RF_BLOCKi_20_Q_reg_30_inst : DFF_X1 port map( D => n3908, CK => CLK
                           , Q => n_3087, QN => 
                           DataPath_RF_bus_reg_dataout_414_port);
   DataPath_RF_BLOCKi_20_Q_reg_29_inst : DFF_X1 port map( D => n3909, CK => CLK
                           , Q => n_3088, QN => 
                           DataPath_RF_bus_reg_dataout_413_port);
   DataPath_RF_BLOCKi_20_Q_reg_28_inst : DFF_X1 port map( D => n3910, CK => CLK
                           , Q => n_3089, QN => 
                           DataPath_RF_bus_reg_dataout_412_port);
   DataPath_RF_BLOCKi_20_Q_reg_27_inst : DFF_X1 port map( D => n3911, CK => CLK
                           , Q => n_3090, QN => 
                           DataPath_RF_bus_reg_dataout_411_port);
   DataPath_RF_BLOCKi_20_Q_reg_26_inst : DFF_X1 port map( D => n3912, CK => CLK
                           , Q => n_3091, QN => 
                           DataPath_RF_bus_reg_dataout_410_port);
   DataPath_RF_BLOCKi_20_Q_reg_25_inst : DFF_X1 port map( D => n3913, CK => CLK
                           , Q => n_3092, QN => 
                           DataPath_RF_bus_reg_dataout_409_port);
   DataPath_RF_BLOCKi_20_Q_reg_24_inst : DFF_X1 port map( D => n3914, CK => CLK
                           , Q => n_3093, QN => 
                           DataPath_RF_bus_reg_dataout_408_port);
   DataPath_RF_BLOCKi_20_Q_reg_23_inst : DFF_X1 port map( D => n3915, CK => CLK
                           , Q => n_3094, QN => 
                           DataPath_RF_bus_reg_dataout_407_port);
   DataPath_RF_BLOCKi_20_Q_reg_22_inst : DFF_X1 port map( D => n3916, CK => CLK
                           , Q => n_3095, QN => 
                           DataPath_RF_bus_reg_dataout_406_port);
   DataPath_RF_BLOCKi_20_Q_reg_21_inst : DFF_X1 port map( D => n3917, CK => CLK
                           , Q => n_3096, QN => 
                           DataPath_RF_bus_reg_dataout_405_port);
   DataPath_RF_BLOCKi_20_Q_reg_20_inst : DFF_X1 port map( D => n3918, CK => CLK
                           , Q => n_3097, QN => 
                           DataPath_RF_bus_reg_dataout_404_port);
   DataPath_RF_BLOCKi_20_Q_reg_19_inst : DFF_X1 port map( D => n3919, CK => CLK
                           , Q => n_3098, QN => 
                           DataPath_RF_bus_reg_dataout_403_port);
   DataPath_RF_BLOCKi_20_Q_reg_18_inst : DFF_X1 port map( D => n3920, CK => CLK
                           , Q => n_3099, QN => 
                           DataPath_RF_bus_reg_dataout_402_port);
   DataPath_RF_BLOCKi_20_Q_reg_17_inst : DFF_X1 port map( D => n3921, CK => CLK
                           , Q => n_3100, QN => 
                           DataPath_RF_bus_reg_dataout_401_port);
   DataPath_RF_BLOCKi_20_Q_reg_16_inst : DFF_X1 port map( D => n3922, CK => CLK
                           , Q => n_3101, QN => 
                           DataPath_RF_bus_reg_dataout_400_port);
   DataPath_RF_BLOCKi_20_Q_reg_15_inst : DFF_X1 port map( D => n3923, CK => CLK
                           , Q => n_3102, QN => 
                           DataPath_RF_bus_reg_dataout_399_port);
   DataPath_RF_BLOCKi_20_Q_reg_14_inst : DFF_X1 port map( D => n3924, CK => CLK
                           , Q => n_3103, QN => 
                           DataPath_RF_bus_reg_dataout_398_port);
   DataPath_RF_BLOCKi_20_Q_reg_13_inst : DFF_X1 port map( D => n3925, CK => CLK
                           , Q => n_3104, QN => 
                           DataPath_RF_bus_reg_dataout_397_port);
   DataPath_RF_BLOCKi_20_Q_reg_12_inst : DFF_X1 port map( D => n3926, CK => CLK
                           , Q => n_3105, QN => 
                           DataPath_RF_bus_reg_dataout_396_port);
   DataPath_RF_BLOCKi_20_Q_reg_11_inst : DFF_X1 port map( D => n3927, CK => CLK
                           , Q => n_3106, QN => 
                           DataPath_RF_bus_reg_dataout_395_port);
   DataPath_RF_BLOCKi_20_Q_reg_9_inst : DFF_X1 port map( D => n3929, CK => CLK,
                           Q => n_3107, QN => 
                           DataPath_RF_bus_reg_dataout_393_port);
   DataPath_RF_BLOCKi_20_Q_reg_8_inst : DFF_X1 port map( D => n3930, CK => CLK,
                           Q => n_3108, QN => 
                           DataPath_RF_bus_reg_dataout_392_port);
   DataPath_RF_BLOCKi_20_Q_reg_7_inst : DFF_X1 port map( D => n3931, CK => CLK,
                           Q => n_3109, QN => 
                           DataPath_RF_bus_reg_dataout_391_port);
   DataPath_RF_BLOCKi_20_Q_reg_6_inst : DFF_X1 port map( D => n3932, CK => CLK,
                           Q => n_3110, QN => 
                           DataPath_RF_bus_reg_dataout_390_port);
   DataPath_RF_BLOCKi_20_Q_reg_5_inst : DFF_X1 port map( D => n3933, CK => CLK,
                           Q => n_3111, QN => 
                           DataPath_RF_bus_reg_dataout_389_port);
   DataPath_RF_BLOCKi_20_Q_reg_4_inst : DFF_X1 port map( D => n3934, CK => CLK,
                           Q => n_3112, QN => 
                           DataPath_RF_bus_reg_dataout_388_port);
   DataPath_RF_BLOCKi_20_Q_reg_3_inst : DFF_X1 port map( D => n3935, CK => CLK,
                           Q => n_3113, QN => 
                           DataPath_RF_bus_reg_dataout_387_port);
   DataPath_RF_BLOCKi_20_Q_reg_2_inst : DFF_X1 port map( D => n3936, CK => CLK,
                           Q => n_3114, QN => 
                           DataPath_RF_bus_reg_dataout_386_port);
   DataPath_RF_BLOCKi_20_Q_reg_1_inst : DFF_X1 port map( D => n3937, CK => CLK,
                           Q => n_3115, QN => 
                           DataPath_RF_bus_reg_dataout_385_port);
   DataPath_RF_BLOCKi_20_Q_reg_0_inst : DFF_X1 port map( D => n3938, CK => CLK,
                           Q => n_3116, QN => 
                           DataPath_RF_bus_reg_dataout_384_port);
   DataPath_RF_BLOCKi_36_Q_reg_31_inst : DFF_X1 port map( D => n4530, CK => CLK
                           , Q => n_3117, QN => 
                           DataPath_RF_bus_reg_dataout_927_port);
   DataPath_RF_BLOCKi_36_Q_reg_30_inst : DFF_X1 port map( D => n4533, CK => CLK
                           , Q => n_3118, QN => 
                           DataPath_RF_bus_reg_dataout_926_port);
   DataPath_RF_BLOCKi_36_Q_reg_29_inst : DFF_X1 port map( D => n4534, CK => CLK
                           , Q => n_3119, QN => 
                           DataPath_RF_bus_reg_dataout_925_port);
   DataPath_RF_BLOCKi_36_Q_reg_28_inst : DFF_X1 port map( D => n4535, CK => CLK
                           , Q => n_3120, QN => 
                           DataPath_RF_bus_reg_dataout_924_port);
   DataPath_RF_BLOCKi_36_Q_reg_27_inst : DFF_X1 port map( D => n4536, CK => CLK
                           , Q => n_3121, QN => 
                           DataPath_RF_bus_reg_dataout_923_port);
   DataPath_RF_BLOCKi_36_Q_reg_26_inst : DFF_X1 port map( D => n4537, CK => CLK
                           , Q => n_3122, QN => 
                           DataPath_RF_bus_reg_dataout_922_port);
   DataPath_RF_BLOCKi_36_Q_reg_25_inst : DFF_X1 port map( D => n4538, CK => CLK
                           , Q => n_3123, QN => 
                           DataPath_RF_bus_reg_dataout_921_port);
   DataPath_RF_BLOCKi_36_Q_reg_24_inst : DFF_X1 port map( D => n4539, CK => CLK
                           , Q => n_3124, QN => 
                           DataPath_RF_bus_reg_dataout_920_port);
   DataPath_RF_BLOCKi_36_Q_reg_23_inst : DFF_X1 port map( D => n4540, CK => CLK
                           , Q => n_3125, QN => 
                           DataPath_RF_bus_reg_dataout_919_port);
   DataPath_RF_BLOCKi_36_Q_reg_22_inst : DFF_X1 port map( D => n4541, CK => CLK
                           , Q => n_3126, QN => 
                           DataPath_RF_bus_reg_dataout_918_port);
   DataPath_RF_BLOCKi_36_Q_reg_21_inst : DFF_X1 port map( D => n4542, CK => CLK
                           , Q => n_3127, QN => 
                           DataPath_RF_bus_reg_dataout_917_port);
   DataPath_RF_BLOCKi_36_Q_reg_20_inst : DFF_X1 port map( D => n4543, CK => CLK
                           , Q => n_3128, QN => 
                           DataPath_RF_bus_reg_dataout_916_port);
   DataPath_RF_BLOCKi_36_Q_reg_19_inst : DFF_X1 port map( D => n4544, CK => CLK
                           , Q => n_3129, QN => 
                           DataPath_RF_bus_reg_dataout_915_port);
   DataPath_RF_BLOCKi_36_Q_reg_18_inst : DFF_X1 port map( D => n4545, CK => CLK
                           , Q => n_3130, QN => 
                           DataPath_RF_bus_reg_dataout_914_port);
   DataPath_RF_BLOCKi_36_Q_reg_17_inst : DFF_X1 port map( D => n4546, CK => CLK
                           , Q => n_3131, QN => 
                           DataPath_RF_bus_reg_dataout_913_port);
   DataPath_RF_BLOCKi_36_Q_reg_16_inst : DFF_X1 port map( D => n4547, CK => CLK
                           , Q => n_3132, QN => 
                           DataPath_RF_bus_reg_dataout_912_port);
   DataPath_RF_BLOCKi_36_Q_reg_15_inst : DFF_X1 port map( D => n4548, CK => CLK
                           , Q => n_3133, QN => 
                           DataPath_RF_bus_reg_dataout_911_port);
   DataPath_RF_BLOCKi_36_Q_reg_14_inst : DFF_X1 port map( D => n4549, CK => CLK
                           , Q => n_3134, QN => 
                           DataPath_RF_bus_reg_dataout_910_port);
   DataPath_RF_BLOCKi_36_Q_reg_13_inst : DFF_X1 port map( D => n4550, CK => CLK
                           , Q => n_3135, QN => 
                           DataPath_RF_bus_reg_dataout_909_port);
   DataPath_RF_BLOCKi_36_Q_reg_12_inst : DFF_X1 port map( D => n4551, CK => CLK
                           , Q => n_3136, QN => 
                           DataPath_RF_bus_reg_dataout_908_port);
   DataPath_RF_BLOCKi_36_Q_reg_11_inst : DFF_X1 port map( D => n4552, CK => CLK
                           , Q => n_3137, QN => 
                           DataPath_RF_bus_reg_dataout_907_port);
   DataPath_RF_BLOCKi_36_Q_reg_9_inst : DFF_X1 port map( D => n4554, CK => CLK,
                           Q => n_3138, QN => 
                           DataPath_RF_bus_reg_dataout_905_port);
   DataPath_RF_BLOCKi_36_Q_reg_8_inst : DFF_X1 port map( D => n4555, CK => CLK,
                           Q => n_3139, QN => 
                           DataPath_RF_bus_reg_dataout_904_port);
   DataPath_RF_BLOCKi_36_Q_reg_7_inst : DFF_X1 port map( D => n4556, CK => CLK,
                           Q => n_3140, QN => 
                           DataPath_RF_bus_reg_dataout_903_port);
   DataPath_RF_BLOCKi_36_Q_reg_6_inst : DFF_X1 port map( D => n4557, CK => CLK,
                           Q => n_3141, QN => 
                           DataPath_RF_bus_reg_dataout_902_port);
   DataPath_RF_BLOCKi_36_Q_reg_5_inst : DFF_X1 port map( D => n4558, CK => CLK,
                           Q => n_3142, QN => 
                           DataPath_RF_bus_reg_dataout_901_port);
   DataPath_RF_BLOCKi_36_Q_reg_4_inst : DFF_X1 port map( D => n4559, CK => CLK,
                           Q => n_3143, QN => 
                           DataPath_RF_bus_reg_dataout_900_port);
   DataPath_RF_BLOCKi_36_Q_reg_3_inst : DFF_X1 port map( D => n4560, CK => CLK,
                           Q => n_3144, QN => 
                           DataPath_RF_bus_reg_dataout_899_port);
   DataPath_RF_BLOCKi_36_Q_reg_2_inst : DFF_X1 port map( D => n4561, CK => CLK,
                           Q => n_3145, QN => 
                           DataPath_RF_bus_reg_dataout_898_port);
   DataPath_RF_BLOCKi_36_Q_reg_1_inst : DFF_X1 port map( D => n4562, CK => CLK,
                           Q => n_3146, QN => 
                           DataPath_RF_bus_reg_dataout_897_port);
   DataPath_RF_BLOCKi_36_Q_reg_0_inst : DFF_X1 port map( D => n4563, CK => CLK,
                           Q => n_3147, QN => 
                           DataPath_RF_bus_reg_dataout_896_port);
   DataPath_RF_BLOCKi_52_Q_reg_31_inst : DFF_X1 port map( D => n5123, CK => CLK
                           , Q => n_3148, QN => 
                           DataPath_RF_bus_reg_dataout_1439_port);
   DataPath_RF_BLOCKi_52_Q_reg_30_inst : DFF_X1 port map( D => n5126, CK => CLK
                           , Q => n_3149, QN => 
                           DataPath_RF_bus_reg_dataout_1438_port);
   DataPath_RF_BLOCKi_52_Q_reg_29_inst : DFF_X1 port map( D => n5127, CK => CLK
                           , Q => n_3150, QN => 
                           DataPath_RF_bus_reg_dataout_1437_port);
   DataPath_RF_BLOCKi_52_Q_reg_28_inst : DFF_X1 port map( D => n5128, CK => CLK
                           , Q => n_3151, QN => 
                           DataPath_RF_bus_reg_dataout_1436_port);
   DataPath_RF_BLOCKi_52_Q_reg_27_inst : DFF_X1 port map( D => n5129, CK => CLK
                           , Q => n_3152, QN => 
                           DataPath_RF_bus_reg_dataout_1435_port);
   DataPath_RF_BLOCKi_52_Q_reg_26_inst : DFF_X1 port map( D => n5130, CK => CLK
                           , Q => n_3153, QN => 
                           DataPath_RF_bus_reg_dataout_1434_port);
   DataPath_RF_BLOCKi_52_Q_reg_25_inst : DFF_X1 port map( D => n5131, CK => CLK
                           , Q => n_3154, QN => 
                           DataPath_RF_bus_reg_dataout_1433_port);
   DataPath_RF_BLOCKi_52_Q_reg_24_inst : DFF_X1 port map( D => n5132, CK => CLK
                           , Q => n_3155, QN => 
                           DataPath_RF_bus_reg_dataout_1432_port);
   DataPath_RF_BLOCKi_52_Q_reg_23_inst : DFF_X1 port map( D => n5133, CK => CLK
                           , Q => n_3156, QN => 
                           DataPath_RF_bus_reg_dataout_1431_port);
   DataPath_RF_BLOCKi_52_Q_reg_22_inst : DFF_X1 port map( D => n5134, CK => CLK
                           , Q => n_3157, QN => 
                           DataPath_RF_bus_reg_dataout_1430_port);
   DataPath_RF_BLOCKi_52_Q_reg_21_inst : DFF_X1 port map( D => n5135, CK => CLK
                           , Q => n_3158, QN => 
                           DataPath_RF_bus_reg_dataout_1429_port);
   DataPath_RF_BLOCKi_52_Q_reg_20_inst : DFF_X1 port map( D => n5136, CK => CLK
                           , Q => n_3159, QN => 
                           DataPath_RF_bus_reg_dataout_1428_port);
   DataPath_RF_BLOCKi_52_Q_reg_19_inst : DFF_X1 port map( D => n5137, CK => CLK
                           , Q => n_3160, QN => 
                           DataPath_RF_bus_reg_dataout_1427_port);
   DataPath_RF_BLOCKi_52_Q_reg_18_inst : DFF_X1 port map( D => n5138, CK => CLK
                           , Q => n_3161, QN => 
                           DataPath_RF_bus_reg_dataout_1426_port);
   DataPath_RF_BLOCKi_52_Q_reg_17_inst : DFF_X1 port map( D => n5139, CK => CLK
                           , Q => n_3162, QN => 
                           DataPath_RF_bus_reg_dataout_1425_port);
   DataPath_RF_BLOCKi_52_Q_reg_16_inst : DFF_X1 port map( D => n5140, CK => CLK
                           , Q => n_3163, QN => 
                           DataPath_RF_bus_reg_dataout_1424_port);
   DataPath_RF_BLOCKi_52_Q_reg_15_inst : DFF_X1 port map( D => n5141, CK => CLK
                           , Q => n_3164, QN => 
                           DataPath_RF_bus_reg_dataout_1423_port);
   DataPath_RF_BLOCKi_52_Q_reg_14_inst : DFF_X1 port map( D => n5142, CK => CLK
                           , Q => n_3165, QN => 
                           DataPath_RF_bus_reg_dataout_1422_port);
   DataPath_RF_BLOCKi_52_Q_reg_13_inst : DFF_X1 port map( D => n5143, CK => CLK
                           , Q => n_3166, QN => 
                           DataPath_RF_bus_reg_dataout_1421_port);
   DataPath_RF_BLOCKi_52_Q_reg_12_inst : DFF_X1 port map( D => n5144, CK => CLK
                           , Q => n_3167, QN => 
                           DataPath_RF_bus_reg_dataout_1420_port);
   DataPath_RF_BLOCKi_52_Q_reg_11_inst : DFF_X1 port map( D => n5145, CK => CLK
                           , Q => n_3168, QN => 
                           DataPath_RF_bus_reg_dataout_1419_port);
   DataPath_RF_BLOCKi_52_Q_reg_9_inst : DFF_X1 port map( D => n5147, CK => CLK,
                           Q => n_3169, QN => 
                           DataPath_RF_bus_reg_dataout_1417_port);
   DataPath_RF_BLOCKi_52_Q_reg_8_inst : DFF_X1 port map( D => n5148, CK => CLK,
                           Q => n_3170, QN => 
                           DataPath_RF_bus_reg_dataout_1416_port);
   DataPath_RF_BLOCKi_52_Q_reg_7_inst : DFF_X1 port map( D => n5149, CK => CLK,
                           Q => n_3171, QN => 
                           DataPath_RF_bus_reg_dataout_1415_port);
   DataPath_RF_BLOCKi_52_Q_reg_6_inst : DFF_X1 port map( D => n5150, CK => CLK,
                           Q => n_3172, QN => 
                           DataPath_RF_bus_reg_dataout_1414_port);
   DataPath_RF_BLOCKi_52_Q_reg_5_inst : DFF_X1 port map( D => n5151, CK => CLK,
                           Q => n_3173, QN => 
                           DataPath_RF_bus_reg_dataout_1413_port);
   DataPath_RF_BLOCKi_52_Q_reg_4_inst : DFF_X1 port map( D => n5152, CK => CLK,
                           Q => n_3174, QN => 
                           DataPath_RF_bus_reg_dataout_1412_port);
   DataPath_RF_BLOCKi_52_Q_reg_3_inst : DFF_X1 port map( D => n5153, CK => CLK,
                           Q => n_3175, QN => 
                           DataPath_RF_bus_reg_dataout_1411_port);
   DataPath_RF_BLOCKi_52_Q_reg_2_inst : DFF_X1 port map( D => n5154, CK => CLK,
                           Q => n_3176, QN => 
                           DataPath_RF_bus_reg_dataout_1410_port);
   DataPath_RF_BLOCKi_52_Q_reg_1_inst : DFF_X1 port map( D => n5155, CK => CLK,
                           Q => n_3177, QN => 
                           DataPath_RF_bus_reg_dataout_1409_port);
   DataPath_RF_BLOCKi_52_Q_reg_0_inst : DFF_X1 port map( D => n5156, CK => CLK,
                           Q => n_3178, QN => 
                           DataPath_RF_bus_reg_dataout_1408_port);
   DataPath_RF_BLOCKi_68_Q_reg_31_inst : DFF_X1 port map( D => n5723, CK => CLK
                           , Q => n_3179, QN => 
                           DataPath_RF_bus_reg_dataout_1951_port);
   DataPath_RF_BLOCKi_68_Q_reg_30_inst : DFF_X1 port map( D => n5726, CK => CLK
                           , Q => n_3180, QN => 
                           DataPath_RF_bus_reg_dataout_1950_port);
   DataPath_RF_BLOCKi_68_Q_reg_29_inst : DFF_X1 port map( D => n5727, CK => CLK
                           , Q => n_3181, QN => 
                           DataPath_RF_bus_reg_dataout_1949_port);
   DataPath_RF_BLOCKi_68_Q_reg_28_inst : DFF_X1 port map( D => n5728, CK => CLK
                           , Q => n_3182, QN => 
                           DataPath_RF_bus_reg_dataout_1948_port);
   DataPath_RF_BLOCKi_68_Q_reg_27_inst : DFF_X1 port map( D => n5729, CK => CLK
                           , Q => n_3183, QN => 
                           DataPath_RF_bus_reg_dataout_1947_port);
   DataPath_RF_BLOCKi_68_Q_reg_26_inst : DFF_X1 port map( D => n5730, CK => CLK
                           , Q => n_3184, QN => 
                           DataPath_RF_bus_reg_dataout_1946_port);
   DataPath_RF_BLOCKi_68_Q_reg_25_inst : DFF_X1 port map( D => n5731, CK => CLK
                           , Q => n_3185, QN => 
                           DataPath_RF_bus_reg_dataout_1945_port);
   DataPath_RF_BLOCKi_68_Q_reg_24_inst : DFF_X1 port map( D => n5732, CK => CLK
                           , Q => n_3186, QN => 
                           DataPath_RF_bus_reg_dataout_1944_port);
   DataPath_RF_BLOCKi_68_Q_reg_23_inst : DFF_X1 port map( D => n5733, CK => CLK
                           , Q => n_3187, QN => 
                           DataPath_RF_bus_reg_dataout_1943_port);
   DataPath_RF_BLOCKi_68_Q_reg_22_inst : DFF_X1 port map( D => n5734, CK => CLK
                           , Q => n_3188, QN => 
                           DataPath_RF_bus_reg_dataout_1942_port);
   DataPath_RF_BLOCKi_68_Q_reg_21_inst : DFF_X1 port map( D => n5735, CK => CLK
                           , Q => n_3189, QN => 
                           DataPath_RF_bus_reg_dataout_1941_port);
   DataPath_RF_BLOCKi_68_Q_reg_20_inst : DFF_X1 port map( D => n5736, CK => CLK
                           , Q => n_3190, QN => 
                           DataPath_RF_bus_reg_dataout_1940_port);
   DataPath_RF_BLOCKi_68_Q_reg_19_inst : DFF_X1 port map( D => n5737, CK => CLK
                           , Q => n_3191, QN => 
                           DataPath_RF_bus_reg_dataout_1939_port);
   DataPath_RF_BLOCKi_68_Q_reg_18_inst : DFF_X1 port map( D => n5738, CK => CLK
                           , Q => n_3192, QN => 
                           DataPath_RF_bus_reg_dataout_1938_port);
   DataPath_RF_BLOCKi_68_Q_reg_17_inst : DFF_X1 port map( D => n5739, CK => CLK
                           , Q => n_3193, QN => 
                           DataPath_RF_bus_reg_dataout_1937_port);
   DataPath_RF_BLOCKi_68_Q_reg_16_inst : DFF_X1 port map( D => n5740, CK => CLK
                           , Q => n_3194, QN => 
                           DataPath_RF_bus_reg_dataout_1936_port);
   DataPath_RF_BLOCKi_68_Q_reg_15_inst : DFF_X1 port map( D => n5741, CK => CLK
                           , Q => n_3195, QN => 
                           DataPath_RF_bus_reg_dataout_1935_port);
   DataPath_RF_BLOCKi_68_Q_reg_14_inst : DFF_X1 port map( D => n5742, CK => CLK
                           , Q => n_3196, QN => 
                           DataPath_RF_bus_reg_dataout_1934_port);
   DataPath_RF_BLOCKi_68_Q_reg_13_inst : DFF_X1 port map( D => n5743, CK => CLK
                           , Q => n_3197, QN => 
                           DataPath_RF_bus_reg_dataout_1933_port);
   DataPath_RF_BLOCKi_68_Q_reg_12_inst : DFF_X1 port map( D => n5744, CK => CLK
                           , Q => n_3198, QN => 
                           DataPath_RF_bus_reg_dataout_1932_port);
   DataPath_RF_BLOCKi_68_Q_reg_11_inst : DFF_X1 port map( D => n5745, CK => CLK
                           , Q => n_3199, QN => 
                           DataPath_RF_bus_reg_dataout_1931_port);
   DataPath_RF_BLOCKi_68_Q_reg_9_inst : DFF_X1 port map( D => n5747, CK => CLK,
                           Q => n_3200, QN => 
                           DataPath_RF_bus_reg_dataout_1929_port);
   DataPath_RF_BLOCKi_68_Q_reg_8_inst : DFF_X1 port map( D => n5748, CK => CLK,
                           Q => n_3201, QN => 
                           DataPath_RF_bus_reg_dataout_1928_port);
   DataPath_RF_BLOCKi_68_Q_reg_7_inst : DFF_X1 port map( D => n5749, CK => CLK,
                           Q => n_3202, QN => 
                           DataPath_RF_bus_reg_dataout_1927_port);
   DataPath_RF_BLOCKi_68_Q_reg_6_inst : DFF_X1 port map( D => n5750, CK => CLK,
                           Q => n_3203, QN => 
                           DataPath_RF_bus_reg_dataout_1926_port);
   DataPath_RF_BLOCKi_68_Q_reg_5_inst : DFF_X1 port map( D => n5751, CK => CLK,
                           Q => n_3204, QN => 
                           DataPath_RF_bus_reg_dataout_1925_port);
   DataPath_RF_BLOCKi_68_Q_reg_4_inst : DFF_X1 port map( D => n5752, CK => CLK,
                           Q => n_3205, QN => 
                           DataPath_RF_bus_reg_dataout_1924_port);
   DataPath_RF_BLOCKi_68_Q_reg_3_inst : DFF_X1 port map( D => n5753, CK => CLK,
                           Q => n_3206, QN => 
                           DataPath_RF_bus_reg_dataout_1923_port);
   DataPath_RF_BLOCKi_68_Q_reg_2_inst : DFF_X1 port map( D => n5754, CK => CLK,
                           Q => n_3207, QN => 
                           DataPath_RF_bus_reg_dataout_1922_port);
   DataPath_RF_BLOCKi_68_Q_reg_1_inst : DFF_X1 port map( D => n5755, CK => CLK,
                           Q => n_3208, QN => 
                           DataPath_RF_bus_reg_dataout_1921_port);
   DataPath_RF_BLOCKi_68_Q_reg_0_inst : DFF_X1 port map( D => n5756, CK => CLK,
                           Q => n_3209, QN => 
                           DataPath_RF_bus_reg_dataout_1920_port);
   DataPath_RF_BLOCKi_85_Q_reg_31_inst : DFF_X1 port map( D => n1114, CK => CLK
                           , Q => n_3210, QN => 
                           DataPath_RF_bus_reg_dataout_2495_port);
   DataPath_RF_BLOCKi_85_Q_reg_30_inst : DFF_X1 port map( D => n1117, CK => CLK
                           , Q => n_3211, QN => 
                           DataPath_RF_bus_reg_dataout_2494_port);
   DataPath_RF_BLOCKi_85_Q_reg_29_inst : DFF_X1 port map( D => n1118, CK => CLK
                           , Q => n_3212, QN => 
                           DataPath_RF_bus_reg_dataout_2493_port);
   DataPath_RF_BLOCKi_85_Q_reg_28_inst : DFF_X1 port map( D => n1119, CK => CLK
                           , Q => n_3213, QN => 
                           DataPath_RF_bus_reg_dataout_2492_port);
   DataPath_RF_BLOCKi_85_Q_reg_27_inst : DFF_X1 port map( D => n1120, CK => CLK
                           , Q => n_3214, QN => 
                           DataPath_RF_bus_reg_dataout_2491_port);
   DataPath_RF_BLOCKi_85_Q_reg_26_inst : DFF_X1 port map( D => n1121, CK => CLK
                           , Q => n_3215, QN => 
                           DataPath_RF_bus_reg_dataout_2490_port);
   DataPath_RF_BLOCKi_85_Q_reg_25_inst : DFF_X1 port map( D => n1122, CK => CLK
                           , Q => n_3216, QN => 
                           DataPath_RF_bus_reg_dataout_2489_port);
   DataPath_RF_BLOCKi_85_Q_reg_24_inst : DFF_X1 port map( D => n1123, CK => CLK
                           , Q => n_3217, QN => 
                           DataPath_RF_bus_reg_dataout_2488_port);
   DataPath_RF_BLOCKi_85_Q_reg_23_inst : DFF_X1 port map( D => n1124, CK => CLK
                           , Q => n_3218, QN => 
                           DataPath_RF_bus_reg_dataout_2487_port);
   DataPath_RF_BLOCKi_85_Q_reg_22_inst : DFF_X1 port map( D => n1125, CK => CLK
                           , Q => n_3219, QN => 
                           DataPath_RF_bus_reg_dataout_2486_port);
   DataPath_RF_BLOCKi_85_Q_reg_21_inst : DFF_X1 port map( D => n1126, CK => CLK
                           , Q => n_3220, QN => 
                           DataPath_RF_bus_reg_dataout_2485_port);
   DataPath_RF_BLOCKi_85_Q_reg_20_inst : DFF_X1 port map( D => n1127, CK => CLK
                           , Q => n_3221, QN => 
                           DataPath_RF_bus_reg_dataout_2484_port);
   DataPath_RF_BLOCKi_85_Q_reg_19_inst : DFF_X1 port map( D => n1128, CK => CLK
                           , Q => n_3222, QN => 
                           DataPath_RF_bus_reg_dataout_2483_port);
   DataPath_RF_BLOCKi_85_Q_reg_18_inst : DFF_X1 port map( D => n1129, CK => CLK
                           , Q => n_3223, QN => 
                           DataPath_RF_bus_reg_dataout_2482_port);
   DataPath_RF_BLOCKi_85_Q_reg_17_inst : DFF_X1 port map( D => n1130, CK => CLK
                           , Q => n_3224, QN => 
                           DataPath_RF_bus_reg_dataout_2481_port);
   DataPath_RF_BLOCKi_85_Q_reg_16_inst : DFF_X1 port map( D => n1131, CK => CLK
                           , Q => n_3225, QN => 
                           DataPath_RF_bus_reg_dataout_2480_port);
   DataPath_RF_BLOCKi_85_Q_reg_15_inst : DFF_X1 port map( D => n1132, CK => CLK
                           , Q => n_3226, QN => 
                           DataPath_RF_bus_reg_dataout_2479_port);
   DataPath_RF_BLOCKi_85_Q_reg_14_inst : DFF_X1 port map( D => n1133, CK => CLK
                           , Q => n_3227, QN => 
                           DataPath_RF_bus_reg_dataout_2478_port);
   DataPath_RF_BLOCKi_85_Q_reg_13_inst : DFF_X1 port map( D => n1134, CK => CLK
                           , Q => n_3228, QN => 
                           DataPath_RF_bus_reg_dataout_2477_port);
   DataPath_RF_BLOCKi_85_Q_reg_12_inst : DFF_X1 port map( D => n1135, CK => CLK
                           , Q => n_3229, QN => 
                           DataPath_RF_bus_reg_dataout_2476_port);
   DataPath_RF_BLOCKi_85_Q_reg_11_inst : DFF_X1 port map( D => n1136, CK => CLK
                           , Q => n_3230, QN => 
                           DataPath_RF_bus_reg_dataout_2475_port);
   DataPath_RF_BLOCKi_85_Q_reg_9_inst : DFF_X1 port map( D => n1138, CK => CLK,
                           Q => n_3231, QN => 
                           DataPath_RF_bus_reg_dataout_2473_port);
   DataPath_RF_BLOCKi_85_Q_reg_8_inst : DFF_X1 port map( D => n1139, CK => CLK,
                           Q => n_3232, QN => 
                           DataPath_RF_bus_reg_dataout_2472_port);
   DataPath_RF_BLOCKi_85_Q_reg_7_inst : DFF_X1 port map( D => n1140, CK => CLK,
                           Q => n_3233, QN => 
                           DataPath_RF_bus_reg_dataout_2471_port);
   DataPath_RF_BLOCKi_85_Q_reg_6_inst : DFF_X1 port map( D => n1141, CK => CLK,
                           Q => n_3234, QN => 
                           DataPath_RF_bus_reg_dataout_2470_port);
   DataPath_RF_BLOCKi_85_Q_reg_5_inst : DFF_X1 port map( D => n1142, CK => CLK,
                           Q => n_3235, QN => 
                           DataPath_RF_bus_reg_dataout_2469_port);
   DataPath_RF_BLOCKi_85_Q_reg_4_inst : DFF_X1 port map( D => n1143, CK => CLK,
                           Q => n_3236, QN => 
                           DataPath_RF_bus_reg_dataout_2468_port);
   DataPath_RF_BLOCKi_85_Q_reg_3_inst : DFF_X1 port map( D => n1144, CK => CLK,
                           Q => n_3237, QN => 
                           DataPath_RF_bus_reg_dataout_2467_port);
   DataPath_RF_BLOCKi_85_Q_reg_2_inst : DFF_X1 port map( D => n1145, CK => CLK,
                           Q => n_3238, QN => 
                           DataPath_RF_bus_reg_dataout_2466_port);
   DataPath_RF_BLOCKi_85_Q_reg_1_inst : DFF_X1 port map( D => n1146, CK => CLK,
                           Q => n_3239, QN => 
                           DataPath_RF_bus_reg_dataout_2465_port);
   DataPath_RF_BLOCKi_85_Q_reg_0_inst : DFF_X1 port map( D => n1147, CK => CLK,
                           Q => n_3240, QN => 
                           DataPath_RF_bus_reg_dataout_2464_port);
   DataPath_RF_BLOCKi_21_Q_reg_31_inst : DFF_X1 port map( D => n3940, CK => CLK
                           , Q => n_3241, QN => 
                           DataPath_RF_bus_reg_dataout_447_port);
   DataPath_RF_BLOCKi_21_Q_reg_30_inst : DFF_X1 port map( D => n3943, CK => CLK
                           , Q => n_3242, QN => 
                           DataPath_RF_bus_reg_dataout_446_port);
   DataPath_RF_BLOCKi_21_Q_reg_29_inst : DFF_X1 port map( D => n3944, CK => CLK
                           , Q => n_3243, QN => 
                           DataPath_RF_bus_reg_dataout_445_port);
   DataPath_RF_BLOCKi_21_Q_reg_28_inst : DFF_X1 port map( D => n3945, CK => CLK
                           , Q => n_3244, QN => 
                           DataPath_RF_bus_reg_dataout_444_port);
   DataPath_RF_BLOCKi_21_Q_reg_27_inst : DFF_X1 port map( D => n3946, CK => CLK
                           , Q => n_3245, QN => 
                           DataPath_RF_bus_reg_dataout_443_port);
   DataPath_RF_BLOCKi_21_Q_reg_26_inst : DFF_X1 port map( D => n3947, CK => CLK
                           , Q => n_3246, QN => 
                           DataPath_RF_bus_reg_dataout_442_port);
   DataPath_RF_BLOCKi_21_Q_reg_25_inst : DFF_X1 port map( D => n3948, CK => CLK
                           , Q => n_3247, QN => 
                           DataPath_RF_bus_reg_dataout_441_port);
   DataPath_RF_BLOCKi_21_Q_reg_24_inst : DFF_X1 port map( D => n3949, CK => CLK
                           , Q => n_3248, QN => 
                           DataPath_RF_bus_reg_dataout_440_port);
   DataPath_RF_BLOCKi_21_Q_reg_23_inst : DFF_X1 port map( D => n3950, CK => CLK
                           , Q => n_3249, QN => 
                           DataPath_RF_bus_reg_dataout_439_port);
   DataPath_RF_BLOCKi_21_Q_reg_22_inst : DFF_X1 port map( D => n3951, CK => CLK
                           , Q => n_3250, QN => 
                           DataPath_RF_bus_reg_dataout_438_port);
   DataPath_RF_BLOCKi_21_Q_reg_21_inst : DFF_X1 port map( D => n3952, CK => CLK
                           , Q => n_3251, QN => 
                           DataPath_RF_bus_reg_dataout_437_port);
   DataPath_RF_BLOCKi_21_Q_reg_20_inst : DFF_X1 port map( D => n3953, CK => CLK
                           , Q => n_3252, QN => 
                           DataPath_RF_bus_reg_dataout_436_port);
   DataPath_RF_BLOCKi_21_Q_reg_19_inst : DFF_X1 port map( D => n3954, CK => CLK
                           , Q => n_3253, QN => 
                           DataPath_RF_bus_reg_dataout_435_port);
   DataPath_RF_BLOCKi_21_Q_reg_18_inst : DFF_X1 port map( D => n3955, CK => CLK
                           , Q => n_3254, QN => 
                           DataPath_RF_bus_reg_dataout_434_port);
   DataPath_RF_BLOCKi_21_Q_reg_17_inst : DFF_X1 port map( D => n3956, CK => CLK
                           , Q => n_3255, QN => 
                           DataPath_RF_bus_reg_dataout_433_port);
   DataPath_RF_BLOCKi_21_Q_reg_16_inst : DFF_X1 port map( D => n3957, CK => CLK
                           , Q => n_3256, QN => 
                           DataPath_RF_bus_reg_dataout_432_port);
   DataPath_RF_BLOCKi_21_Q_reg_15_inst : DFF_X1 port map( D => n3958, CK => CLK
                           , Q => n_3257, QN => 
                           DataPath_RF_bus_reg_dataout_431_port);
   DataPath_RF_BLOCKi_21_Q_reg_14_inst : DFF_X1 port map( D => n3959, CK => CLK
                           , Q => n_3258, QN => 
                           DataPath_RF_bus_reg_dataout_430_port);
   DataPath_RF_BLOCKi_21_Q_reg_13_inst : DFF_X1 port map( D => n3960, CK => CLK
                           , Q => n_3259, QN => 
                           DataPath_RF_bus_reg_dataout_429_port);
   DataPath_RF_BLOCKi_21_Q_reg_12_inst : DFF_X1 port map( D => n3961, CK => CLK
                           , Q => n_3260, QN => 
                           DataPath_RF_bus_reg_dataout_428_port);
   DataPath_RF_BLOCKi_21_Q_reg_11_inst : DFF_X1 port map( D => n3962, CK => CLK
                           , Q => n_3261, QN => 
                           DataPath_RF_bus_reg_dataout_427_port);
   DataPath_RF_BLOCKi_21_Q_reg_9_inst : DFF_X1 port map( D => n3964, CK => CLK,
                           Q => n_3262, QN => 
                           DataPath_RF_bus_reg_dataout_425_port);
   DataPath_RF_BLOCKi_21_Q_reg_8_inst : DFF_X1 port map( D => n3965, CK => CLK,
                           Q => n_3263, QN => 
                           DataPath_RF_bus_reg_dataout_424_port);
   DataPath_RF_BLOCKi_21_Q_reg_7_inst : DFF_X1 port map( D => n3966, CK => CLK,
                           Q => n_3264, QN => 
                           DataPath_RF_bus_reg_dataout_423_port);
   DataPath_RF_BLOCKi_21_Q_reg_6_inst : DFF_X1 port map( D => n3967, CK => CLK,
                           Q => n_3265, QN => 
                           DataPath_RF_bus_reg_dataout_422_port);
   DataPath_RF_BLOCKi_21_Q_reg_5_inst : DFF_X1 port map( D => n3968, CK => CLK,
                           Q => n_3266, QN => 
                           DataPath_RF_bus_reg_dataout_421_port);
   DataPath_RF_BLOCKi_21_Q_reg_4_inst : DFF_X1 port map( D => n3969, CK => CLK,
                           Q => n_3267, QN => 
                           DataPath_RF_bus_reg_dataout_420_port);
   DataPath_RF_BLOCKi_21_Q_reg_3_inst : DFF_X1 port map( D => n3970, CK => CLK,
                           Q => n_3268, QN => 
                           DataPath_RF_bus_reg_dataout_419_port);
   DataPath_RF_BLOCKi_21_Q_reg_2_inst : DFF_X1 port map( D => n3971, CK => CLK,
                           Q => n_3269, QN => 
                           DataPath_RF_bus_reg_dataout_418_port);
   DataPath_RF_BLOCKi_21_Q_reg_1_inst : DFF_X1 port map( D => n3972, CK => CLK,
                           Q => n_3270, QN => 
                           DataPath_RF_bus_reg_dataout_417_port);
   DataPath_RF_BLOCKi_21_Q_reg_0_inst : DFF_X1 port map( D => n3973, CK => CLK,
                           Q => n_3271, QN => 
                           DataPath_RF_bus_reg_dataout_416_port);
   DataPath_RF_BLOCKi_37_Q_reg_31_inst : DFF_X1 port map( D => n4565, CK => CLK
                           , Q => n_3272, QN => 
                           DataPath_RF_bus_reg_dataout_959_port);
   DataPath_RF_BLOCKi_37_Q_reg_30_inst : DFF_X1 port map( D => n4568, CK => CLK
                           , Q => n_3273, QN => 
                           DataPath_RF_bus_reg_dataout_958_port);
   DataPath_RF_BLOCKi_37_Q_reg_29_inst : DFF_X1 port map( D => n4569, CK => CLK
                           , Q => n_3274, QN => 
                           DataPath_RF_bus_reg_dataout_957_port);
   DataPath_RF_BLOCKi_37_Q_reg_28_inst : DFF_X1 port map( D => n4570, CK => CLK
                           , Q => n_3275, QN => 
                           DataPath_RF_bus_reg_dataout_956_port);
   DataPath_RF_BLOCKi_37_Q_reg_27_inst : DFF_X1 port map( D => n4571, CK => CLK
                           , Q => n_3276, QN => 
                           DataPath_RF_bus_reg_dataout_955_port);
   DataPath_RF_BLOCKi_37_Q_reg_26_inst : DFF_X1 port map( D => n4572, CK => CLK
                           , Q => n_3277, QN => 
                           DataPath_RF_bus_reg_dataout_954_port);
   DataPath_RF_BLOCKi_37_Q_reg_25_inst : DFF_X1 port map( D => n4573, CK => CLK
                           , Q => n_3278, QN => 
                           DataPath_RF_bus_reg_dataout_953_port);
   DataPath_RF_BLOCKi_37_Q_reg_24_inst : DFF_X1 port map( D => n4574, CK => CLK
                           , Q => n_3279, QN => 
                           DataPath_RF_bus_reg_dataout_952_port);
   DataPath_RF_BLOCKi_37_Q_reg_23_inst : DFF_X1 port map( D => n4575, CK => CLK
                           , Q => n_3280, QN => 
                           DataPath_RF_bus_reg_dataout_951_port);
   DataPath_RF_BLOCKi_37_Q_reg_22_inst : DFF_X1 port map( D => n4576, CK => CLK
                           , Q => n_3281, QN => 
                           DataPath_RF_bus_reg_dataout_950_port);
   DataPath_RF_BLOCKi_37_Q_reg_21_inst : DFF_X1 port map( D => n4577, CK => CLK
                           , Q => n_3282, QN => 
                           DataPath_RF_bus_reg_dataout_949_port);
   DataPath_RF_BLOCKi_37_Q_reg_20_inst : DFF_X1 port map( D => n4578, CK => CLK
                           , Q => n_3283, QN => 
                           DataPath_RF_bus_reg_dataout_948_port);
   DataPath_RF_BLOCKi_37_Q_reg_19_inst : DFF_X1 port map( D => n4579, CK => CLK
                           , Q => n_3284, QN => 
                           DataPath_RF_bus_reg_dataout_947_port);
   DataPath_RF_BLOCKi_37_Q_reg_18_inst : DFF_X1 port map( D => n4580, CK => CLK
                           , Q => n_3285, QN => 
                           DataPath_RF_bus_reg_dataout_946_port);
   DataPath_RF_BLOCKi_37_Q_reg_17_inst : DFF_X1 port map( D => n4581, CK => CLK
                           , Q => n_3286, QN => 
                           DataPath_RF_bus_reg_dataout_945_port);
   DataPath_RF_BLOCKi_37_Q_reg_16_inst : DFF_X1 port map( D => n4582, CK => CLK
                           , Q => n_3287, QN => 
                           DataPath_RF_bus_reg_dataout_944_port);
   DataPath_RF_BLOCKi_37_Q_reg_15_inst : DFF_X1 port map( D => n4583, CK => CLK
                           , Q => n_3288, QN => 
                           DataPath_RF_bus_reg_dataout_943_port);
   DataPath_RF_BLOCKi_37_Q_reg_14_inst : DFF_X1 port map( D => n4584, CK => CLK
                           , Q => n_3289, QN => 
                           DataPath_RF_bus_reg_dataout_942_port);
   DataPath_RF_BLOCKi_37_Q_reg_13_inst : DFF_X1 port map( D => n4585, CK => CLK
                           , Q => n_3290, QN => 
                           DataPath_RF_bus_reg_dataout_941_port);
   DataPath_RF_BLOCKi_37_Q_reg_12_inst : DFF_X1 port map( D => n4586, CK => CLK
                           , Q => n_3291, QN => 
                           DataPath_RF_bus_reg_dataout_940_port);
   DataPath_RF_BLOCKi_37_Q_reg_11_inst : DFF_X1 port map( D => n4587, CK => CLK
                           , Q => n_3292, QN => 
                           DataPath_RF_bus_reg_dataout_939_port);
   DataPath_RF_BLOCKi_37_Q_reg_9_inst : DFF_X1 port map( D => n4589, CK => CLK,
                           Q => n_3293, QN => 
                           DataPath_RF_bus_reg_dataout_937_port);
   DataPath_RF_BLOCKi_37_Q_reg_8_inst : DFF_X1 port map( D => n4590, CK => CLK,
                           Q => n_3294, QN => 
                           DataPath_RF_bus_reg_dataout_936_port);
   DataPath_RF_BLOCKi_37_Q_reg_7_inst : DFF_X1 port map( D => n4591, CK => CLK,
                           Q => n_3295, QN => 
                           DataPath_RF_bus_reg_dataout_935_port);
   DataPath_RF_BLOCKi_37_Q_reg_6_inst : DFF_X1 port map( D => n4592, CK => CLK,
                           Q => n_3296, QN => 
                           DataPath_RF_bus_reg_dataout_934_port);
   DataPath_RF_BLOCKi_37_Q_reg_5_inst : DFF_X1 port map( D => n4593, CK => CLK,
                           Q => n_3297, QN => 
                           DataPath_RF_bus_reg_dataout_933_port);
   DataPath_RF_BLOCKi_37_Q_reg_4_inst : DFF_X1 port map( D => n4594, CK => CLK,
                           Q => n_3298, QN => 
                           DataPath_RF_bus_reg_dataout_932_port);
   DataPath_RF_BLOCKi_37_Q_reg_3_inst : DFF_X1 port map( D => n4595, CK => CLK,
                           Q => n_3299, QN => 
                           DataPath_RF_bus_reg_dataout_931_port);
   DataPath_RF_BLOCKi_37_Q_reg_2_inst : DFF_X1 port map( D => n4596, CK => CLK,
                           Q => n_3300, QN => 
                           DataPath_RF_bus_reg_dataout_930_port);
   DataPath_RF_BLOCKi_37_Q_reg_1_inst : DFF_X1 port map( D => n4597, CK => CLK,
                           Q => n_3301, QN => 
                           DataPath_RF_bus_reg_dataout_929_port);
   DataPath_RF_BLOCKi_37_Q_reg_0_inst : DFF_X1 port map( D => n4598, CK => CLK,
                           Q => n_3302, QN => 
                           DataPath_RF_bus_reg_dataout_928_port);
   DataPath_RF_BLOCKi_53_Q_reg_31_inst : DFF_X1 port map( D => n5158, CK => CLK
                           , Q => n_3303, QN => 
                           DataPath_RF_bus_reg_dataout_1471_port);
   DataPath_RF_BLOCKi_53_Q_reg_30_inst : DFF_X1 port map( D => n5161, CK => CLK
                           , Q => n_3304, QN => 
                           DataPath_RF_bus_reg_dataout_1470_port);
   DataPath_RF_BLOCKi_53_Q_reg_29_inst : DFF_X1 port map( D => n5162, CK => CLK
                           , Q => n_3305, QN => 
                           DataPath_RF_bus_reg_dataout_1469_port);
   DataPath_RF_BLOCKi_53_Q_reg_28_inst : DFF_X1 port map( D => n5163, CK => CLK
                           , Q => n_3306, QN => 
                           DataPath_RF_bus_reg_dataout_1468_port);
   DataPath_RF_BLOCKi_53_Q_reg_27_inst : DFF_X1 port map( D => n5164, CK => CLK
                           , Q => n_3307, QN => 
                           DataPath_RF_bus_reg_dataout_1467_port);
   DataPath_RF_BLOCKi_53_Q_reg_26_inst : DFF_X1 port map( D => n5165, CK => CLK
                           , Q => n_3308, QN => 
                           DataPath_RF_bus_reg_dataout_1466_port);
   DataPath_RF_BLOCKi_53_Q_reg_25_inst : DFF_X1 port map( D => n5166, CK => CLK
                           , Q => n_3309, QN => 
                           DataPath_RF_bus_reg_dataout_1465_port);
   DataPath_RF_BLOCKi_53_Q_reg_24_inst : DFF_X1 port map( D => n5167, CK => CLK
                           , Q => n_3310, QN => 
                           DataPath_RF_bus_reg_dataout_1464_port);
   DataPath_RF_BLOCKi_53_Q_reg_23_inst : DFF_X1 port map( D => n5168, CK => CLK
                           , Q => n_3311, QN => 
                           DataPath_RF_bus_reg_dataout_1463_port);
   DataPath_RF_BLOCKi_53_Q_reg_22_inst : DFF_X1 port map( D => n5169, CK => CLK
                           , Q => n_3312, QN => 
                           DataPath_RF_bus_reg_dataout_1462_port);
   DataPath_RF_BLOCKi_53_Q_reg_21_inst : DFF_X1 port map( D => n5170, CK => CLK
                           , Q => n_3313, QN => 
                           DataPath_RF_bus_reg_dataout_1461_port);
   DataPath_RF_BLOCKi_53_Q_reg_20_inst : DFF_X1 port map( D => n5171, CK => CLK
                           , Q => n_3314, QN => 
                           DataPath_RF_bus_reg_dataout_1460_port);
   DataPath_RF_BLOCKi_53_Q_reg_19_inst : DFF_X1 port map( D => n5172, CK => CLK
                           , Q => n_3315, QN => 
                           DataPath_RF_bus_reg_dataout_1459_port);
   DataPath_RF_BLOCKi_53_Q_reg_18_inst : DFF_X1 port map( D => n5173, CK => CLK
                           , Q => n_3316, QN => 
                           DataPath_RF_bus_reg_dataout_1458_port);
   DataPath_RF_BLOCKi_53_Q_reg_17_inst : DFF_X1 port map( D => n5174, CK => CLK
                           , Q => n_3317, QN => 
                           DataPath_RF_bus_reg_dataout_1457_port);
   DataPath_RF_BLOCKi_53_Q_reg_16_inst : DFF_X1 port map( D => n5175, CK => CLK
                           , Q => n_3318, QN => 
                           DataPath_RF_bus_reg_dataout_1456_port);
   DataPath_RF_BLOCKi_53_Q_reg_15_inst : DFF_X1 port map( D => n5176, CK => CLK
                           , Q => n_3319, QN => 
                           DataPath_RF_bus_reg_dataout_1455_port);
   DataPath_RF_BLOCKi_53_Q_reg_14_inst : DFF_X1 port map( D => n5177, CK => CLK
                           , Q => n_3320, QN => 
                           DataPath_RF_bus_reg_dataout_1454_port);
   DataPath_RF_BLOCKi_53_Q_reg_13_inst : DFF_X1 port map( D => n5178, CK => CLK
                           , Q => n_3321, QN => 
                           DataPath_RF_bus_reg_dataout_1453_port);
   DataPath_RF_BLOCKi_53_Q_reg_12_inst : DFF_X1 port map( D => n5179, CK => CLK
                           , Q => n_3322, QN => 
                           DataPath_RF_bus_reg_dataout_1452_port);
   DataPath_RF_BLOCKi_53_Q_reg_11_inst : DFF_X1 port map( D => n5180, CK => CLK
                           , Q => n_3323, QN => 
                           DataPath_RF_bus_reg_dataout_1451_port);
   DataPath_RF_BLOCKi_53_Q_reg_9_inst : DFF_X1 port map( D => n5182, CK => CLK,
                           Q => n_3324, QN => 
                           DataPath_RF_bus_reg_dataout_1449_port);
   DataPath_RF_BLOCKi_53_Q_reg_8_inst : DFF_X1 port map( D => n5183, CK => CLK,
                           Q => n_3325, QN => 
                           DataPath_RF_bus_reg_dataout_1448_port);
   DataPath_RF_BLOCKi_53_Q_reg_7_inst : DFF_X1 port map( D => n5184, CK => CLK,
                           Q => n_3326, QN => 
                           DataPath_RF_bus_reg_dataout_1447_port);
   DataPath_RF_BLOCKi_53_Q_reg_6_inst : DFF_X1 port map( D => n5185, CK => CLK,
                           Q => n_3327, QN => 
                           DataPath_RF_bus_reg_dataout_1446_port);
   DataPath_RF_BLOCKi_53_Q_reg_5_inst : DFF_X1 port map( D => n5186, CK => CLK,
                           Q => n_3328, QN => 
                           DataPath_RF_bus_reg_dataout_1445_port);
   DataPath_RF_BLOCKi_53_Q_reg_4_inst : DFF_X1 port map( D => n5187, CK => CLK,
                           Q => n_3329, QN => 
                           DataPath_RF_bus_reg_dataout_1444_port);
   DataPath_RF_BLOCKi_53_Q_reg_3_inst : DFF_X1 port map( D => n5188, CK => CLK,
                           Q => n_3330, QN => 
                           DataPath_RF_bus_reg_dataout_1443_port);
   DataPath_RF_BLOCKi_53_Q_reg_2_inst : DFF_X1 port map( D => n5189, CK => CLK,
                           Q => n_3331, QN => 
                           DataPath_RF_bus_reg_dataout_1442_port);
   DataPath_RF_BLOCKi_53_Q_reg_1_inst : DFF_X1 port map( D => n5190, CK => CLK,
                           Q => n_3332, QN => 
                           DataPath_RF_bus_reg_dataout_1441_port);
   DataPath_RF_BLOCKi_53_Q_reg_0_inst : DFF_X1 port map( D => n5191, CK => CLK,
                           Q => n_3333, QN => 
                           DataPath_RF_bus_reg_dataout_1440_port);
   DataPath_RF_BLOCKi_69_Q_reg_31_inst : DFF_X1 port map( D => n5759, CK => CLK
                           , Q => n_3334, QN => 
                           DataPath_RF_bus_reg_dataout_1983_port);
   DataPath_RF_BLOCKi_69_Q_reg_30_inst : DFF_X1 port map( D => n5762, CK => CLK
                           , Q => n_3335, QN => 
                           DataPath_RF_bus_reg_dataout_1982_port);
   DataPath_RF_BLOCKi_69_Q_reg_29_inst : DFF_X1 port map( D => n5763, CK => CLK
                           , Q => n_3336, QN => 
                           DataPath_RF_bus_reg_dataout_1981_port);
   DataPath_RF_BLOCKi_69_Q_reg_28_inst : DFF_X1 port map( D => n5764, CK => CLK
                           , Q => n_3337, QN => 
                           DataPath_RF_bus_reg_dataout_1980_port);
   DataPath_RF_BLOCKi_69_Q_reg_27_inst : DFF_X1 port map( D => n5765, CK => CLK
                           , Q => n_3338, QN => 
                           DataPath_RF_bus_reg_dataout_1979_port);
   DataPath_RF_BLOCKi_69_Q_reg_26_inst : DFF_X1 port map( D => n5766, CK => CLK
                           , Q => n_3339, QN => 
                           DataPath_RF_bus_reg_dataout_1978_port);
   DataPath_RF_BLOCKi_69_Q_reg_25_inst : DFF_X1 port map( D => n5767, CK => CLK
                           , Q => n_3340, QN => 
                           DataPath_RF_bus_reg_dataout_1977_port);
   DataPath_RF_BLOCKi_69_Q_reg_24_inst : DFF_X1 port map( D => n5768, CK => CLK
                           , Q => n_3341, QN => 
                           DataPath_RF_bus_reg_dataout_1976_port);
   DataPath_RF_BLOCKi_69_Q_reg_23_inst : DFF_X1 port map( D => n5769, CK => CLK
                           , Q => n_3342, QN => 
                           DataPath_RF_bus_reg_dataout_1975_port);
   DataPath_RF_BLOCKi_69_Q_reg_22_inst : DFF_X1 port map( D => n5770, CK => CLK
                           , Q => n_3343, QN => 
                           DataPath_RF_bus_reg_dataout_1974_port);
   DataPath_RF_BLOCKi_69_Q_reg_21_inst : DFF_X1 port map( D => n5771, CK => CLK
                           , Q => n_3344, QN => 
                           DataPath_RF_bus_reg_dataout_1973_port);
   DataPath_RF_BLOCKi_69_Q_reg_20_inst : DFF_X1 port map( D => n5772, CK => CLK
                           , Q => n_3345, QN => 
                           DataPath_RF_bus_reg_dataout_1972_port);
   DataPath_RF_BLOCKi_69_Q_reg_19_inst : DFF_X1 port map( D => n5773, CK => CLK
                           , Q => n_3346, QN => 
                           DataPath_RF_bus_reg_dataout_1971_port);
   DataPath_RF_BLOCKi_69_Q_reg_18_inst : DFF_X1 port map( D => n5774, CK => CLK
                           , Q => n_3347, QN => 
                           DataPath_RF_bus_reg_dataout_1970_port);
   DataPath_RF_BLOCKi_69_Q_reg_17_inst : DFF_X1 port map( D => n5775, CK => CLK
                           , Q => n_3348, QN => 
                           DataPath_RF_bus_reg_dataout_1969_port);
   DataPath_RF_BLOCKi_69_Q_reg_16_inst : DFF_X1 port map( D => n5776, CK => CLK
                           , Q => n_3349, QN => 
                           DataPath_RF_bus_reg_dataout_1968_port);
   DataPath_RF_BLOCKi_69_Q_reg_15_inst : DFF_X1 port map( D => n5777, CK => CLK
                           , Q => n_3350, QN => 
                           DataPath_RF_bus_reg_dataout_1967_port);
   DataPath_RF_BLOCKi_69_Q_reg_14_inst : DFF_X1 port map( D => n5778, CK => CLK
                           , Q => n_3351, QN => 
                           DataPath_RF_bus_reg_dataout_1966_port);
   DataPath_RF_BLOCKi_69_Q_reg_13_inst : DFF_X1 port map( D => n5779, CK => CLK
                           , Q => n_3352, QN => 
                           DataPath_RF_bus_reg_dataout_1965_port);
   DataPath_RF_BLOCKi_69_Q_reg_12_inst : DFF_X1 port map( D => n5780, CK => CLK
                           , Q => n_3353, QN => 
                           DataPath_RF_bus_reg_dataout_1964_port);
   DataPath_RF_BLOCKi_69_Q_reg_11_inst : DFF_X1 port map( D => n5781, CK => CLK
                           , Q => n_3354, QN => 
                           DataPath_RF_bus_reg_dataout_1963_port);
   DataPath_RF_BLOCKi_69_Q_reg_9_inst : DFF_X1 port map( D => n5783, CK => CLK,
                           Q => n_3355, QN => 
                           DataPath_RF_bus_reg_dataout_1961_port);
   DataPath_RF_BLOCKi_69_Q_reg_8_inst : DFF_X1 port map( D => n5784, CK => CLK,
                           Q => n_3356, QN => 
                           DataPath_RF_bus_reg_dataout_1960_port);
   DataPath_RF_BLOCKi_69_Q_reg_7_inst : DFF_X1 port map( D => n5785, CK => CLK,
                           Q => n_3357, QN => 
                           DataPath_RF_bus_reg_dataout_1959_port);
   DataPath_RF_BLOCKi_69_Q_reg_6_inst : DFF_X1 port map( D => n5786, CK => CLK,
                           Q => n_3358, QN => 
                           DataPath_RF_bus_reg_dataout_1958_port);
   DataPath_RF_BLOCKi_69_Q_reg_5_inst : DFF_X1 port map( D => n5787, CK => CLK,
                           Q => n_3359, QN => 
                           DataPath_RF_bus_reg_dataout_1957_port);
   DataPath_RF_BLOCKi_69_Q_reg_4_inst : DFF_X1 port map( D => n5788, CK => CLK,
                           Q => n_3360, QN => 
                           DataPath_RF_bus_reg_dataout_1956_port);
   DataPath_RF_BLOCKi_69_Q_reg_3_inst : DFF_X1 port map( D => n5789, CK => CLK,
                           Q => n_3361, QN => 
                           DataPath_RF_bus_reg_dataout_1955_port);
   DataPath_RF_BLOCKi_69_Q_reg_2_inst : DFF_X1 port map( D => n5790, CK => CLK,
                           Q => n_3362, QN => 
                           DataPath_RF_bus_reg_dataout_1954_port);
   DataPath_RF_BLOCKi_69_Q_reg_1_inst : DFF_X1 port map( D => n5791, CK => CLK,
                           Q => n_3363, QN => 
                           DataPath_RF_bus_reg_dataout_1953_port);
   DataPath_RF_BLOCKi_69_Q_reg_0_inst : DFF_X1 port map( D => n5792, CK => CLK,
                           Q => n_3364, QN => 
                           DataPath_RF_bus_reg_dataout_1952_port);
   DataPath_RF_BLOCKi_86_Q_reg_31_inst : DFF_X1 port map( D => n1151, CK => CLK
                           , Q => n_3365, QN => 
                           DataPath_RF_bus_reg_dataout_2527_port);
   DataPath_RF_BLOCKi_86_Q_reg_30_inst : DFF_X1 port map( D => n1154, CK => CLK
                           , Q => n_3366, QN => 
                           DataPath_RF_bus_reg_dataout_2526_port);
   DataPath_RF_BLOCKi_86_Q_reg_29_inst : DFF_X1 port map( D => n1155, CK => CLK
                           , Q => n_3367, QN => 
                           DataPath_RF_bus_reg_dataout_2525_port);
   DataPath_RF_BLOCKi_86_Q_reg_28_inst : DFF_X1 port map( D => n1156, CK => CLK
                           , Q => n_3368, QN => 
                           DataPath_RF_bus_reg_dataout_2524_port);
   DataPath_RF_BLOCKi_86_Q_reg_27_inst : DFF_X1 port map( D => n1157, CK => CLK
                           , Q => n_3369, QN => 
                           DataPath_RF_bus_reg_dataout_2523_port);
   DataPath_RF_BLOCKi_86_Q_reg_26_inst : DFF_X1 port map( D => n1158, CK => CLK
                           , Q => n_3370, QN => 
                           DataPath_RF_bus_reg_dataout_2522_port);
   DataPath_RF_BLOCKi_86_Q_reg_25_inst : DFF_X1 port map( D => n1159, CK => CLK
                           , Q => n_3371, QN => 
                           DataPath_RF_bus_reg_dataout_2521_port);
   DataPath_RF_BLOCKi_86_Q_reg_24_inst : DFF_X1 port map( D => n1160, CK => CLK
                           , Q => n_3372, QN => 
                           DataPath_RF_bus_reg_dataout_2520_port);
   DataPath_RF_BLOCKi_86_Q_reg_23_inst : DFF_X1 port map( D => n1161, CK => CLK
                           , Q => n_3373, QN => 
                           DataPath_RF_bus_reg_dataout_2519_port);
   DataPath_RF_BLOCKi_86_Q_reg_22_inst : DFF_X1 port map( D => n1162, CK => CLK
                           , Q => n_3374, QN => 
                           DataPath_RF_bus_reg_dataout_2518_port);
   DataPath_RF_BLOCKi_86_Q_reg_21_inst : DFF_X1 port map( D => n1163, CK => CLK
                           , Q => n_3375, QN => 
                           DataPath_RF_bus_reg_dataout_2517_port);
   DataPath_RF_BLOCKi_86_Q_reg_20_inst : DFF_X1 port map( D => n1164, CK => CLK
                           , Q => n_3376, QN => 
                           DataPath_RF_bus_reg_dataout_2516_port);
   DataPath_RF_BLOCKi_86_Q_reg_19_inst : DFF_X1 port map( D => n1165, CK => CLK
                           , Q => n_3377, QN => 
                           DataPath_RF_bus_reg_dataout_2515_port);
   DataPath_RF_BLOCKi_86_Q_reg_18_inst : DFF_X1 port map( D => n1166, CK => CLK
                           , Q => n_3378, QN => 
                           DataPath_RF_bus_reg_dataout_2514_port);
   DataPath_RF_BLOCKi_86_Q_reg_17_inst : DFF_X1 port map( D => n1167, CK => CLK
                           , Q => n_3379, QN => 
                           DataPath_RF_bus_reg_dataout_2513_port);
   DataPath_RF_BLOCKi_86_Q_reg_16_inst : DFF_X1 port map( D => n1168, CK => CLK
                           , Q => n_3380, QN => 
                           DataPath_RF_bus_reg_dataout_2512_port);
   DataPath_RF_BLOCKi_86_Q_reg_15_inst : DFF_X1 port map( D => n1169, CK => CLK
                           , Q => n_3381, QN => 
                           DataPath_RF_bus_reg_dataout_2511_port);
   DataPath_RF_BLOCKi_86_Q_reg_14_inst : DFF_X1 port map( D => n1170, CK => CLK
                           , Q => n_3382, QN => 
                           DataPath_RF_bus_reg_dataout_2510_port);
   DataPath_RF_BLOCKi_86_Q_reg_13_inst : DFF_X1 port map( D => n1171, CK => CLK
                           , Q => n_3383, QN => 
                           DataPath_RF_bus_reg_dataout_2509_port);
   DataPath_RF_BLOCKi_86_Q_reg_12_inst : DFF_X1 port map( D => n1172, CK => CLK
                           , Q => n_3384, QN => 
                           DataPath_RF_bus_reg_dataout_2508_port);
   DataPath_RF_BLOCKi_86_Q_reg_11_inst : DFF_X1 port map( D => n1173, CK => CLK
                           , Q => n_3385, QN => 
                           DataPath_RF_bus_reg_dataout_2507_port);
   DataPath_RF_BLOCKi_86_Q_reg_9_inst : DFF_X1 port map( D => n1175, CK => CLK,
                           Q => n_3386, QN => 
                           DataPath_RF_bus_reg_dataout_2505_port);
   DataPath_RF_BLOCKi_86_Q_reg_8_inst : DFF_X1 port map( D => n1176, CK => CLK,
                           Q => n_3387, QN => 
                           DataPath_RF_bus_reg_dataout_2504_port);
   DataPath_RF_BLOCKi_86_Q_reg_7_inst : DFF_X1 port map( D => n1177, CK => CLK,
                           Q => n_3388, QN => 
                           DataPath_RF_bus_reg_dataout_2503_port);
   DataPath_RF_BLOCKi_86_Q_reg_6_inst : DFF_X1 port map( D => n1178, CK => CLK,
                           Q => n_3389, QN => 
                           DataPath_RF_bus_reg_dataout_2502_port);
   DataPath_RF_BLOCKi_86_Q_reg_5_inst : DFF_X1 port map( D => n1179, CK => CLK,
                           Q => n_3390, QN => 
                           DataPath_RF_bus_reg_dataout_2501_port);
   DataPath_RF_BLOCKi_86_Q_reg_4_inst : DFF_X1 port map( D => n1180, CK => CLK,
                           Q => n_3391, QN => 
                           DataPath_RF_bus_reg_dataout_2500_port);
   DataPath_RF_BLOCKi_86_Q_reg_3_inst : DFF_X1 port map( D => n1181, CK => CLK,
                           Q => n_3392, QN => 
                           DataPath_RF_bus_reg_dataout_2499_port);
   DataPath_RF_BLOCKi_86_Q_reg_2_inst : DFF_X1 port map( D => n1182, CK => CLK,
                           Q => n_3393, QN => 
                           DataPath_RF_bus_reg_dataout_2498_port);
   DataPath_RF_BLOCKi_86_Q_reg_1_inst : DFF_X1 port map( D => n1183, CK => CLK,
                           Q => n_3394, QN => 
                           DataPath_RF_bus_reg_dataout_2497_port);
   DataPath_RF_BLOCKi_86_Q_reg_0_inst : DFF_X1 port map( D => n1184, CK => CLK,
                           Q => n_3395, QN => 
                           DataPath_RF_bus_reg_dataout_2496_port);
   DataPath_RF_BLOCKi_22_Q_reg_31_inst : DFF_X1 port map( D => n3975, CK => CLK
                           , Q => n_3396, QN => 
                           DataPath_RF_bus_reg_dataout_479_port);
   DataPath_RF_BLOCKi_22_Q_reg_30_inst : DFF_X1 port map( D => n3978, CK => CLK
                           , Q => n_3397, QN => 
                           DataPath_RF_bus_reg_dataout_478_port);
   DataPath_RF_BLOCKi_22_Q_reg_29_inst : DFF_X1 port map( D => n3979, CK => CLK
                           , Q => n_3398, QN => 
                           DataPath_RF_bus_reg_dataout_477_port);
   DataPath_RF_BLOCKi_22_Q_reg_28_inst : DFF_X1 port map( D => n3980, CK => CLK
                           , Q => n_3399, QN => 
                           DataPath_RF_bus_reg_dataout_476_port);
   DataPath_RF_BLOCKi_22_Q_reg_27_inst : DFF_X1 port map( D => n3981, CK => CLK
                           , Q => n_3400, QN => 
                           DataPath_RF_bus_reg_dataout_475_port);
   DataPath_RF_BLOCKi_22_Q_reg_26_inst : DFF_X1 port map( D => n3982, CK => CLK
                           , Q => n_3401, QN => 
                           DataPath_RF_bus_reg_dataout_474_port);
   DataPath_RF_BLOCKi_22_Q_reg_25_inst : DFF_X1 port map( D => n3983, CK => CLK
                           , Q => n_3402, QN => 
                           DataPath_RF_bus_reg_dataout_473_port);
   DataPath_RF_BLOCKi_22_Q_reg_24_inst : DFF_X1 port map( D => n3984, CK => CLK
                           , Q => n_3403, QN => 
                           DataPath_RF_bus_reg_dataout_472_port);
   DataPath_RF_BLOCKi_22_Q_reg_23_inst : DFF_X1 port map( D => n3985, CK => CLK
                           , Q => n_3404, QN => 
                           DataPath_RF_bus_reg_dataout_471_port);
   DataPath_RF_BLOCKi_22_Q_reg_22_inst : DFF_X1 port map( D => n3986, CK => CLK
                           , Q => n_3405, QN => 
                           DataPath_RF_bus_reg_dataout_470_port);
   DataPath_RF_BLOCKi_22_Q_reg_21_inst : DFF_X1 port map( D => n3987, CK => CLK
                           , Q => n_3406, QN => 
                           DataPath_RF_bus_reg_dataout_469_port);
   DataPath_RF_BLOCKi_22_Q_reg_20_inst : DFF_X1 port map( D => n3988, CK => CLK
                           , Q => n_3407, QN => 
                           DataPath_RF_bus_reg_dataout_468_port);
   DataPath_RF_BLOCKi_22_Q_reg_19_inst : DFF_X1 port map( D => n3989, CK => CLK
                           , Q => n_3408, QN => 
                           DataPath_RF_bus_reg_dataout_467_port);
   DataPath_RF_BLOCKi_22_Q_reg_18_inst : DFF_X1 port map( D => n3990, CK => CLK
                           , Q => n_3409, QN => 
                           DataPath_RF_bus_reg_dataout_466_port);
   DataPath_RF_BLOCKi_22_Q_reg_17_inst : DFF_X1 port map( D => n3991, CK => CLK
                           , Q => n_3410, QN => 
                           DataPath_RF_bus_reg_dataout_465_port);
   DataPath_RF_BLOCKi_22_Q_reg_16_inst : DFF_X1 port map( D => n3992, CK => CLK
                           , Q => n_3411, QN => 
                           DataPath_RF_bus_reg_dataout_464_port);
   DataPath_RF_BLOCKi_22_Q_reg_15_inst : DFF_X1 port map( D => n3993, CK => CLK
                           , Q => n_3412, QN => 
                           DataPath_RF_bus_reg_dataout_463_port);
   DataPath_RF_BLOCKi_22_Q_reg_14_inst : DFF_X1 port map( D => n3994, CK => CLK
                           , Q => n_3413, QN => 
                           DataPath_RF_bus_reg_dataout_462_port);
   DataPath_RF_BLOCKi_22_Q_reg_13_inst : DFF_X1 port map( D => n3995, CK => CLK
                           , Q => n_3414, QN => 
                           DataPath_RF_bus_reg_dataout_461_port);
   DataPath_RF_BLOCKi_22_Q_reg_12_inst : DFF_X1 port map( D => n3996, CK => CLK
                           , Q => n_3415, QN => 
                           DataPath_RF_bus_reg_dataout_460_port);
   DataPath_RF_BLOCKi_22_Q_reg_11_inst : DFF_X1 port map( D => n3997, CK => CLK
                           , Q => n_3416, QN => 
                           DataPath_RF_bus_reg_dataout_459_port);
   DataPath_RF_BLOCKi_22_Q_reg_9_inst : DFF_X1 port map( D => n3999, CK => CLK,
                           Q => n_3417, QN => 
                           DataPath_RF_bus_reg_dataout_457_port);
   DataPath_RF_BLOCKi_22_Q_reg_8_inst : DFF_X1 port map( D => n4000, CK => CLK,
                           Q => n_3418, QN => 
                           DataPath_RF_bus_reg_dataout_456_port);
   DataPath_RF_BLOCKi_22_Q_reg_7_inst : DFF_X1 port map( D => n4001, CK => CLK,
                           Q => n_3419, QN => 
                           DataPath_RF_bus_reg_dataout_455_port);
   DataPath_RF_BLOCKi_22_Q_reg_6_inst : DFF_X1 port map( D => n4002, CK => CLK,
                           Q => n_3420, QN => 
                           DataPath_RF_bus_reg_dataout_454_port);
   DataPath_RF_BLOCKi_22_Q_reg_5_inst : DFF_X1 port map( D => n4003, CK => CLK,
                           Q => n_3421, QN => 
                           DataPath_RF_bus_reg_dataout_453_port);
   DataPath_RF_BLOCKi_22_Q_reg_4_inst : DFF_X1 port map( D => n4004, CK => CLK,
                           Q => n_3422, QN => 
                           DataPath_RF_bus_reg_dataout_452_port);
   DataPath_RF_BLOCKi_22_Q_reg_3_inst : DFF_X1 port map( D => n4005, CK => CLK,
                           Q => n_3423, QN => 
                           DataPath_RF_bus_reg_dataout_451_port);
   DataPath_RF_BLOCKi_22_Q_reg_2_inst : DFF_X1 port map( D => n4006, CK => CLK,
                           Q => n_3424, QN => 
                           DataPath_RF_bus_reg_dataout_450_port);
   DataPath_RF_BLOCKi_22_Q_reg_1_inst : DFF_X1 port map( D => n4007, CK => CLK,
                           Q => n_3425, QN => 
                           DataPath_RF_bus_reg_dataout_449_port);
   DataPath_RF_BLOCKi_22_Q_reg_0_inst : DFF_X1 port map( D => n4008, CK => CLK,
                           Q => n_3426, QN => 
                           DataPath_RF_bus_reg_dataout_448_port);
   DataPath_RF_BLOCKi_38_Q_reg_31_inst : DFF_X1 port map( D => n4600, CK => CLK
                           , Q => n_3427, QN => 
                           DataPath_RF_bus_reg_dataout_991_port);
   DataPath_RF_BLOCKi_38_Q_reg_30_inst : DFF_X1 port map( D => n4603, CK => CLK
                           , Q => n_3428, QN => 
                           DataPath_RF_bus_reg_dataout_990_port);
   DataPath_RF_BLOCKi_38_Q_reg_29_inst : DFF_X1 port map( D => n4604, CK => CLK
                           , Q => n_3429, QN => 
                           DataPath_RF_bus_reg_dataout_989_port);
   DataPath_RF_BLOCKi_38_Q_reg_28_inst : DFF_X1 port map( D => n4605, CK => CLK
                           , Q => n_3430, QN => 
                           DataPath_RF_bus_reg_dataout_988_port);
   DataPath_RF_BLOCKi_38_Q_reg_27_inst : DFF_X1 port map( D => n4606, CK => CLK
                           , Q => n_3431, QN => 
                           DataPath_RF_bus_reg_dataout_987_port);
   DataPath_RF_BLOCKi_38_Q_reg_26_inst : DFF_X1 port map( D => n4607, CK => CLK
                           , Q => n_3432, QN => 
                           DataPath_RF_bus_reg_dataout_986_port);
   DataPath_RF_BLOCKi_38_Q_reg_25_inst : DFF_X1 port map( D => n4608, CK => CLK
                           , Q => n_3433, QN => 
                           DataPath_RF_bus_reg_dataout_985_port);
   DataPath_RF_BLOCKi_38_Q_reg_24_inst : DFF_X1 port map( D => n4609, CK => CLK
                           , Q => n_3434, QN => 
                           DataPath_RF_bus_reg_dataout_984_port);
   DataPath_RF_BLOCKi_38_Q_reg_23_inst : DFF_X1 port map( D => n4610, CK => CLK
                           , Q => n_3435, QN => 
                           DataPath_RF_bus_reg_dataout_983_port);
   DataPath_RF_BLOCKi_38_Q_reg_22_inst : DFF_X1 port map( D => n4611, CK => CLK
                           , Q => n_3436, QN => 
                           DataPath_RF_bus_reg_dataout_982_port);
   DataPath_RF_BLOCKi_38_Q_reg_21_inst : DFF_X1 port map( D => n4612, CK => CLK
                           , Q => n_3437, QN => 
                           DataPath_RF_bus_reg_dataout_981_port);
   DataPath_RF_BLOCKi_38_Q_reg_20_inst : DFF_X1 port map( D => n4613, CK => CLK
                           , Q => n_3438, QN => 
                           DataPath_RF_bus_reg_dataout_980_port);
   DataPath_RF_BLOCKi_38_Q_reg_19_inst : DFF_X1 port map( D => n4614, CK => CLK
                           , Q => n_3439, QN => 
                           DataPath_RF_bus_reg_dataout_979_port);
   DataPath_RF_BLOCKi_38_Q_reg_18_inst : DFF_X1 port map( D => n4615, CK => CLK
                           , Q => n_3440, QN => 
                           DataPath_RF_bus_reg_dataout_978_port);
   DataPath_RF_BLOCKi_38_Q_reg_17_inst : DFF_X1 port map( D => n4616, CK => CLK
                           , Q => n_3441, QN => 
                           DataPath_RF_bus_reg_dataout_977_port);
   DataPath_RF_BLOCKi_38_Q_reg_16_inst : DFF_X1 port map( D => n4617, CK => CLK
                           , Q => n_3442, QN => 
                           DataPath_RF_bus_reg_dataout_976_port);
   DataPath_RF_BLOCKi_38_Q_reg_15_inst : DFF_X1 port map( D => n4618, CK => CLK
                           , Q => n_3443, QN => 
                           DataPath_RF_bus_reg_dataout_975_port);
   DataPath_RF_BLOCKi_38_Q_reg_14_inst : DFF_X1 port map( D => n4619, CK => CLK
                           , Q => n_3444, QN => 
                           DataPath_RF_bus_reg_dataout_974_port);
   DataPath_RF_BLOCKi_38_Q_reg_13_inst : DFF_X1 port map( D => n4620, CK => CLK
                           , Q => n_3445, QN => 
                           DataPath_RF_bus_reg_dataout_973_port);
   DataPath_RF_BLOCKi_38_Q_reg_12_inst : DFF_X1 port map( D => n4621, CK => CLK
                           , Q => n_3446, QN => 
                           DataPath_RF_bus_reg_dataout_972_port);
   DataPath_RF_BLOCKi_38_Q_reg_11_inst : DFF_X1 port map( D => n4622, CK => CLK
                           , Q => n_3447, QN => 
                           DataPath_RF_bus_reg_dataout_971_port);
   DataPath_RF_BLOCKi_38_Q_reg_9_inst : DFF_X1 port map( D => n4624, CK => CLK,
                           Q => n_3448, QN => 
                           DataPath_RF_bus_reg_dataout_969_port);
   DataPath_RF_BLOCKi_38_Q_reg_8_inst : DFF_X1 port map( D => n4625, CK => CLK,
                           Q => n_3449, QN => 
                           DataPath_RF_bus_reg_dataout_968_port);
   DataPath_RF_BLOCKi_38_Q_reg_7_inst : DFF_X1 port map( D => n4626, CK => CLK,
                           Q => n_3450, QN => 
                           DataPath_RF_bus_reg_dataout_967_port);
   DataPath_RF_BLOCKi_38_Q_reg_6_inst : DFF_X1 port map( D => n4627, CK => CLK,
                           Q => n_3451, QN => 
                           DataPath_RF_bus_reg_dataout_966_port);
   DataPath_RF_BLOCKi_38_Q_reg_5_inst : DFF_X1 port map( D => n4628, CK => CLK,
                           Q => n_3452, QN => 
                           DataPath_RF_bus_reg_dataout_965_port);
   DataPath_RF_BLOCKi_38_Q_reg_4_inst : DFF_X1 port map( D => n4629, CK => CLK,
                           Q => n_3453, QN => 
                           DataPath_RF_bus_reg_dataout_964_port);
   DataPath_RF_BLOCKi_38_Q_reg_3_inst : DFF_X1 port map( D => n4630, CK => CLK,
                           Q => n_3454, QN => 
                           DataPath_RF_bus_reg_dataout_963_port);
   DataPath_RF_BLOCKi_38_Q_reg_2_inst : DFF_X1 port map( D => n4631, CK => CLK,
                           Q => n_3455, QN => 
                           DataPath_RF_bus_reg_dataout_962_port);
   DataPath_RF_BLOCKi_38_Q_reg_1_inst : DFF_X1 port map( D => n4632, CK => CLK,
                           Q => n_3456, QN => 
                           DataPath_RF_bus_reg_dataout_961_port);
   DataPath_RF_BLOCKi_38_Q_reg_0_inst : DFF_X1 port map( D => n4633, CK => CLK,
                           Q => n_3457, QN => 
                           DataPath_RF_bus_reg_dataout_960_port);
   DataPath_RF_BLOCKi_54_Q_reg_31_inst : DFF_X1 port map( D => n5193, CK => CLK
                           , Q => n_3458, QN => 
                           DataPath_RF_bus_reg_dataout_1503_port);
   DataPath_RF_BLOCKi_54_Q_reg_30_inst : DFF_X1 port map( D => n5196, CK => CLK
                           , Q => n_3459, QN => 
                           DataPath_RF_bus_reg_dataout_1502_port);
   DataPath_RF_BLOCKi_54_Q_reg_29_inst : DFF_X1 port map( D => n5197, CK => CLK
                           , Q => n_3460, QN => 
                           DataPath_RF_bus_reg_dataout_1501_port);
   DataPath_RF_BLOCKi_54_Q_reg_28_inst : DFF_X1 port map( D => n5198, CK => CLK
                           , Q => n_3461, QN => 
                           DataPath_RF_bus_reg_dataout_1500_port);
   DataPath_RF_BLOCKi_54_Q_reg_27_inst : DFF_X1 port map( D => n5199, CK => CLK
                           , Q => n_3462, QN => 
                           DataPath_RF_bus_reg_dataout_1499_port);
   DataPath_RF_BLOCKi_54_Q_reg_26_inst : DFF_X1 port map( D => n5200, CK => CLK
                           , Q => n_3463, QN => 
                           DataPath_RF_bus_reg_dataout_1498_port);
   DataPath_RF_BLOCKi_54_Q_reg_25_inst : DFF_X1 port map( D => n5201, CK => CLK
                           , Q => n_3464, QN => 
                           DataPath_RF_bus_reg_dataout_1497_port);
   DataPath_RF_BLOCKi_54_Q_reg_24_inst : DFF_X1 port map( D => n5202, CK => CLK
                           , Q => n_3465, QN => 
                           DataPath_RF_bus_reg_dataout_1496_port);
   DataPath_RF_BLOCKi_54_Q_reg_23_inst : DFF_X1 port map( D => n5203, CK => CLK
                           , Q => n_3466, QN => 
                           DataPath_RF_bus_reg_dataout_1495_port);
   DataPath_RF_BLOCKi_54_Q_reg_22_inst : DFF_X1 port map( D => n5204, CK => CLK
                           , Q => n_3467, QN => 
                           DataPath_RF_bus_reg_dataout_1494_port);
   DataPath_RF_BLOCKi_54_Q_reg_21_inst : DFF_X1 port map( D => n5205, CK => CLK
                           , Q => n_3468, QN => 
                           DataPath_RF_bus_reg_dataout_1493_port);
   DataPath_RF_BLOCKi_54_Q_reg_20_inst : DFF_X1 port map( D => n5206, CK => CLK
                           , Q => n_3469, QN => 
                           DataPath_RF_bus_reg_dataout_1492_port);
   DataPath_RF_BLOCKi_54_Q_reg_19_inst : DFF_X1 port map( D => n5207, CK => CLK
                           , Q => n_3470, QN => 
                           DataPath_RF_bus_reg_dataout_1491_port);
   DataPath_RF_BLOCKi_54_Q_reg_18_inst : DFF_X1 port map( D => n5208, CK => CLK
                           , Q => n_3471, QN => 
                           DataPath_RF_bus_reg_dataout_1490_port);
   DataPath_RF_BLOCKi_54_Q_reg_17_inst : DFF_X1 port map( D => n5209, CK => CLK
                           , Q => n_3472, QN => 
                           DataPath_RF_bus_reg_dataout_1489_port);
   DataPath_RF_BLOCKi_54_Q_reg_16_inst : DFF_X1 port map( D => n5210, CK => CLK
                           , Q => n_3473, QN => 
                           DataPath_RF_bus_reg_dataout_1488_port);
   DataPath_RF_BLOCKi_54_Q_reg_15_inst : DFF_X1 port map( D => n5211, CK => CLK
                           , Q => n_3474, QN => 
                           DataPath_RF_bus_reg_dataout_1487_port);
   DataPath_RF_BLOCKi_54_Q_reg_14_inst : DFF_X1 port map( D => n5212, CK => CLK
                           , Q => n_3475, QN => 
                           DataPath_RF_bus_reg_dataout_1486_port);
   DataPath_RF_BLOCKi_54_Q_reg_13_inst : DFF_X1 port map( D => n5213, CK => CLK
                           , Q => n_3476, QN => 
                           DataPath_RF_bus_reg_dataout_1485_port);
   DataPath_RF_BLOCKi_54_Q_reg_12_inst : DFF_X1 port map( D => n5214, CK => CLK
                           , Q => n_3477, QN => 
                           DataPath_RF_bus_reg_dataout_1484_port);
   DataPath_RF_BLOCKi_54_Q_reg_11_inst : DFF_X1 port map( D => n5215, CK => CLK
                           , Q => n_3478, QN => 
                           DataPath_RF_bus_reg_dataout_1483_port);
   DataPath_RF_BLOCKi_54_Q_reg_9_inst : DFF_X1 port map( D => n5217, CK => CLK,
                           Q => n_3479, QN => 
                           DataPath_RF_bus_reg_dataout_1481_port);
   DataPath_RF_BLOCKi_54_Q_reg_8_inst : DFF_X1 port map( D => n5218, CK => CLK,
                           Q => n_3480, QN => 
                           DataPath_RF_bus_reg_dataout_1480_port);
   DataPath_RF_BLOCKi_54_Q_reg_7_inst : DFF_X1 port map( D => n5219, CK => CLK,
                           Q => n_3481, QN => 
                           DataPath_RF_bus_reg_dataout_1479_port);
   DataPath_RF_BLOCKi_54_Q_reg_6_inst : DFF_X1 port map( D => n5220, CK => CLK,
                           Q => n_3482, QN => 
                           DataPath_RF_bus_reg_dataout_1478_port);
   DataPath_RF_BLOCKi_54_Q_reg_5_inst : DFF_X1 port map( D => n5221, CK => CLK,
                           Q => n_3483, QN => 
                           DataPath_RF_bus_reg_dataout_1477_port);
   DataPath_RF_BLOCKi_54_Q_reg_4_inst : DFF_X1 port map( D => n5222, CK => CLK,
                           Q => n_3484, QN => 
                           DataPath_RF_bus_reg_dataout_1476_port);
   DataPath_RF_BLOCKi_54_Q_reg_3_inst : DFF_X1 port map( D => n5223, CK => CLK,
                           Q => n_3485, QN => 
                           DataPath_RF_bus_reg_dataout_1475_port);
   DataPath_RF_BLOCKi_54_Q_reg_2_inst : DFF_X1 port map( D => n5224, CK => CLK,
                           Q => n_3486, QN => 
                           DataPath_RF_bus_reg_dataout_1474_port);
   DataPath_RF_BLOCKi_54_Q_reg_1_inst : DFF_X1 port map( D => n5225, CK => CLK,
                           Q => n_3487, QN => 
                           DataPath_RF_bus_reg_dataout_1473_port);
   DataPath_RF_BLOCKi_54_Q_reg_0_inst : DFF_X1 port map( D => n5226, CK => CLK,
                           Q => n_3488, QN => 
                           DataPath_RF_bus_reg_dataout_1472_port);
   DataPath_RF_BLOCKi_70_Q_reg_31_inst : DFF_X1 port map( D => n5795, CK => CLK
                           , Q => n_3489, QN => 
                           DataPath_RF_bus_reg_dataout_2015_port);
   DataPath_RF_BLOCKi_70_Q_reg_30_inst : DFF_X1 port map( D => n5798, CK => CLK
                           , Q => n_3490, QN => 
                           DataPath_RF_bus_reg_dataout_2014_port);
   DataPath_RF_BLOCKi_70_Q_reg_29_inst : DFF_X1 port map( D => n5799, CK => CLK
                           , Q => n_3491, QN => 
                           DataPath_RF_bus_reg_dataout_2013_port);
   DataPath_RF_BLOCKi_70_Q_reg_28_inst : DFF_X1 port map( D => n5800, CK => CLK
                           , Q => n_3492, QN => 
                           DataPath_RF_bus_reg_dataout_2012_port);
   DataPath_RF_BLOCKi_70_Q_reg_27_inst : DFF_X1 port map( D => n5801, CK => CLK
                           , Q => n_3493, QN => 
                           DataPath_RF_bus_reg_dataout_2011_port);
   DataPath_RF_BLOCKi_70_Q_reg_26_inst : DFF_X1 port map( D => n5802, CK => CLK
                           , Q => n_3494, QN => 
                           DataPath_RF_bus_reg_dataout_2010_port);
   DataPath_RF_BLOCKi_70_Q_reg_25_inst : DFF_X1 port map( D => n5803, CK => CLK
                           , Q => n_3495, QN => 
                           DataPath_RF_bus_reg_dataout_2009_port);
   DataPath_RF_BLOCKi_70_Q_reg_24_inst : DFF_X1 port map( D => n5804, CK => CLK
                           , Q => n_3496, QN => 
                           DataPath_RF_bus_reg_dataout_2008_port);
   DataPath_RF_BLOCKi_70_Q_reg_23_inst : DFF_X1 port map( D => n5805, CK => CLK
                           , Q => n_3497, QN => 
                           DataPath_RF_bus_reg_dataout_2007_port);
   DataPath_RF_BLOCKi_70_Q_reg_22_inst : DFF_X1 port map( D => n5806, CK => CLK
                           , Q => n_3498, QN => 
                           DataPath_RF_bus_reg_dataout_2006_port);
   DataPath_RF_BLOCKi_70_Q_reg_21_inst : DFF_X1 port map( D => n5807, CK => CLK
                           , Q => n_3499, QN => 
                           DataPath_RF_bus_reg_dataout_2005_port);
   DataPath_RF_BLOCKi_70_Q_reg_20_inst : DFF_X1 port map( D => n5808, CK => CLK
                           , Q => n_3500, QN => 
                           DataPath_RF_bus_reg_dataout_2004_port);
   DataPath_RF_BLOCKi_70_Q_reg_19_inst : DFF_X1 port map( D => n5809, CK => CLK
                           , Q => n_3501, QN => 
                           DataPath_RF_bus_reg_dataout_2003_port);
   DataPath_RF_BLOCKi_70_Q_reg_18_inst : DFF_X1 port map( D => n5810, CK => CLK
                           , Q => n_3502, QN => 
                           DataPath_RF_bus_reg_dataout_2002_port);
   DataPath_RF_BLOCKi_70_Q_reg_17_inst : DFF_X1 port map( D => n5811, CK => CLK
                           , Q => n_3503, QN => 
                           DataPath_RF_bus_reg_dataout_2001_port);
   DataPath_RF_BLOCKi_70_Q_reg_16_inst : DFF_X1 port map( D => n5812, CK => CLK
                           , Q => n_3504, QN => 
                           DataPath_RF_bus_reg_dataout_2000_port);
   DataPath_RF_BLOCKi_70_Q_reg_15_inst : DFF_X1 port map( D => n5813, CK => CLK
                           , Q => n_3505, QN => 
                           DataPath_RF_bus_reg_dataout_1999_port);
   DataPath_RF_BLOCKi_70_Q_reg_14_inst : DFF_X1 port map( D => n5814, CK => CLK
                           , Q => n_3506, QN => 
                           DataPath_RF_bus_reg_dataout_1998_port);
   DataPath_RF_BLOCKi_70_Q_reg_13_inst : DFF_X1 port map( D => n5815, CK => CLK
                           , Q => n_3507, QN => 
                           DataPath_RF_bus_reg_dataout_1997_port);
   DataPath_RF_BLOCKi_70_Q_reg_12_inst : DFF_X1 port map( D => n5816, CK => CLK
                           , Q => n_3508, QN => 
                           DataPath_RF_bus_reg_dataout_1996_port);
   DataPath_RF_BLOCKi_70_Q_reg_11_inst : DFF_X1 port map( D => n5817, CK => CLK
                           , Q => n_3509, QN => 
                           DataPath_RF_bus_reg_dataout_1995_port);
   DataPath_RF_BLOCKi_70_Q_reg_9_inst : DFF_X1 port map( D => n5819, CK => CLK,
                           Q => n_3510, QN => 
                           DataPath_RF_bus_reg_dataout_1993_port);
   DataPath_RF_BLOCKi_70_Q_reg_8_inst : DFF_X1 port map( D => n5820, CK => CLK,
                           Q => n_3511, QN => 
                           DataPath_RF_bus_reg_dataout_1992_port);
   DataPath_RF_BLOCKi_70_Q_reg_7_inst : DFF_X1 port map( D => n5821, CK => CLK,
                           Q => n_3512, QN => 
                           DataPath_RF_bus_reg_dataout_1991_port);
   DataPath_RF_BLOCKi_70_Q_reg_6_inst : DFF_X1 port map( D => n5822, CK => CLK,
                           Q => n_3513, QN => 
                           DataPath_RF_bus_reg_dataout_1990_port);
   DataPath_RF_BLOCKi_70_Q_reg_5_inst : DFF_X1 port map( D => n5823, CK => CLK,
                           Q => n_3514, QN => 
                           DataPath_RF_bus_reg_dataout_1989_port);
   DataPath_RF_BLOCKi_70_Q_reg_4_inst : DFF_X1 port map( D => n5824, CK => CLK,
                           Q => n_3515, QN => 
                           DataPath_RF_bus_reg_dataout_1988_port);
   DataPath_RF_BLOCKi_70_Q_reg_3_inst : DFF_X1 port map( D => n5825, CK => CLK,
                           Q => n_3516, QN => 
                           DataPath_RF_bus_reg_dataout_1987_port);
   DataPath_RF_BLOCKi_70_Q_reg_2_inst : DFF_X1 port map( D => n5826, CK => CLK,
                           Q => n_3517, QN => 
                           DataPath_RF_bus_reg_dataout_1986_port);
   DataPath_RF_BLOCKi_70_Q_reg_1_inst : DFF_X1 port map( D => n5827, CK => CLK,
                           Q => n_3518, QN => 
                           DataPath_RF_bus_reg_dataout_1985_port);
   DataPath_RF_BLOCKi_70_Q_reg_0_inst : DFF_X1 port map( D => n5828, CK => CLK,
                           Q => n_3519, QN => 
                           DataPath_RF_bus_reg_dataout_1984_port);
   DataPath_RF_BLOCKi_87_Q_reg_31_inst : DFF_X1 port map( D => n1188, CK => CLK
                           , Q => n_3520, QN => 
                           DataPath_RF_bus_reg_dataout_2559_port);
   DataPath_RF_BLOCKi_87_Q_reg_30_inst : DFF_X1 port map( D => n1191, CK => CLK
                           , Q => n_3521, QN => 
                           DataPath_RF_bus_reg_dataout_2558_port);
   DataPath_RF_BLOCKi_87_Q_reg_29_inst : DFF_X1 port map( D => n1192, CK => CLK
                           , Q => n_3522, QN => 
                           DataPath_RF_bus_reg_dataout_2557_port);
   DataPath_RF_BLOCKi_87_Q_reg_28_inst : DFF_X1 port map( D => n1193, CK => CLK
                           , Q => n_3523, QN => 
                           DataPath_RF_bus_reg_dataout_2556_port);
   DataPath_RF_BLOCKi_87_Q_reg_27_inst : DFF_X1 port map( D => n1194, CK => CLK
                           , Q => n_3524, QN => 
                           DataPath_RF_bus_reg_dataout_2555_port);
   DataPath_RF_BLOCKi_87_Q_reg_26_inst : DFF_X1 port map( D => n1195, CK => CLK
                           , Q => n_3525, QN => 
                           DataPath_RF_bus_reg_dataout_2554_port);
   DataPath_RF_BLOCKi_87_Q_reg_25_inst : DFF_X1 port map( D => n1196, CK => CLK
                           , Q => n_3526, QN => 
                           DataPath_RF_bus_reg_dataout_2553_port);
   DataPath_RF_BLOCKi_87_Q_reg_24_inst : DFF_X1 port map( D => n1197, CK => CLK
                           , Q => n_3527, QN => 
                           DataPath_RF_bus_reg_dataout_2552_port);
   DataPath_RF_BLOCKi_87_Q_reg_23_inst : DFF_X1 port map( D => n1198, CK => CLK
                           , Q => n_3528, QN => 
                           DataPath_RF_bus_reg_dataout_2551_port);
   DataPath_RF_BLOCKi_87_Q_reg_22_inst : DFF_X1 port map( D => n1199, CK => CLK
                           , Q => n_3529, QN => 
                           DataPath_RF_bus_reg_dataout_2550_port);
   DataPath_RF_BLOCKi_87_Q_reg_21_inst : DFF_X1 port map( D => n1200, CK => CLK
                           , Q => n_3530, QN => 
                           DataPath_RF_bus_reg_dataout_2549_port);
   DataPath_RF_BLOCKi_87_Q_reg_20_inst : DFF_X1 port map( D => n1201, CK => CLK
                           , Q => n_3531, QN => 
                           DataPath_RF_bus_reg_dataout_2548_port);
   DataPath_RF_BLOCKi_87_Q_reg_19_inst : DFF_X1 port map( D => n1202, CK => CLK
                           , Q => n_3532, QN => 
                           DataPath_RF_bus_reg_dataout_2547_port);
   DataPath_RF_BLOCKi_87_Q_reg_18_inst : DFF_X1 port map( D => n1203, CK => CLK
                           , Q => n_3533, QN => 
                           DataPath_RF_bus_reg_dataout_2546_port);
   DataPath_RF_BLOCKi_87_Q_reg_17_inst : DFF_X1 port map( D => n1204, CK => CLK
                           , Q => n_3534, QN => 
                           DataPath_RF_bus_reg_dataout_2545_port);
   DataPath_RF_BLOCKi_87_Q_reg_16_inst : DFF_X1 port map( D => n1205, CK => CLK
                           , Q => n_3535, QN => 
                           DataPath_RF_bus_reg_dataout_2544_port);
   DataPath_RF_BLOCKi_87_Q_reg_15_inst : DFF_X1 port map( D => n1206, CK => CLK
                           , Q => n_3536, QN => 
                           DataPath_RF_bus_reg_dataout_2543_port);
   DataPath_RF_BLOCKi_87_Q_reg_14_inst : DFF_X1 port map( D => n1207, CK => CLK
                           , Q => n_3537, QN => 
                           DataPath_RF_bus_reg_dataout_2542_port);
   DataPath_RF_BLOCKi_87_Q_reg_13_inst : DFF_X1 port map( D => n1208, CK => CLK
                           , Q => n_3538, QN => 
                           DataPath_RF_bus_reg_dataout_2541_port);
   DataPath_RF_BLOCKi_87_Q_reg_12_inst : DFF_X1 port map( D => n1209, CK => CLK
                           , Q => n_3539, QN => 
                           DataPath_RF_bus_reg_dataout_2540_port);
   DataPath_RF_BLOCKi_87_Q_reg_11_inst : DFF_X1 port map( D => n1210, CK => CLK
                           , Q => n_3540, QN => 
                           DataPath_RF_bus_reg_dataout_2539_port);
   DataPath_RF_BLOCKi_87_Q_reg_9_inst : DFF_X1 port map( D => n1212, CK => CLK,
                           Q => n_3541, QN => 
                           DataPath_RF_bus_reg_dataout_2537_port);
   DataPath_RF_BLOCKi_87_Q_reg_8_inst : DFF_X1 port map( D => n1213, CK => CLK,
                           Q => n_3542, QN => 
                           DataPath_RF_bus_reg_dataout_2536_port);
   DataPath_RF_BLOCKi_87_Q_reg_7_inst : DFF_X1 port map( D => n1214, CK => CLK,
                           Q => n_3543, QN => 
                           DataPath_RF_bus_reg_dataout_2535_port);
   DataPath_RF_BLOCKi_87_Q_reg_6_inst : DFF_X1 port map( D => n1215, CK => CLK,
                           Q => n_3544, QN => 
                           DataPath_RF_bus_reg_dataout_2534_port);
   DataPath_RF_BLOCKi_87_Q_reg_5_inst : DFF_X1 port map( D => n1216, CK => CLK,
                           Q => n_3545, QN => 
                           DataPath_RF_bus_reg_dataout_2533_port);
   DataPath_RF_BLOCKi_87_Q_reg_4_inst : DFF_X1 port map( D => n1217, CK => CLK,
                           Q => n_3546, QN => 
                           DataPath_RF_bus_reg_dataout_2532_port);
   DataPath_RF_BLOCKi_87_Q_reg_3_inst : DFF_X1 port map( D => n1218, CK => CLK,
                           Q => n_3547, QN => 
                           DataPath_RF_bus_reg_dataout_2531_port);
   DataPath_RF_BLOCKi_87_Q_reg_2_inst : DFF_X1 port map( D => n1219, CK => CLK,
                           Q => n_3548, QN => 
                           DataPath_RF_bus_reg_dataout_2530_port);
   DataPath_RF_BLOCKi_87_Q_reg_1_inst : DFF_X1 port map( D => n1220, CK => CLK,
                           Q => n_3549, QN => 
                           DataPath_RF_bus_reg_dataout_2529_port);
   DataPath_RF_BLOCKi_87_Q_reg_0_inst : DFF_X1 port map( D => n1221, CK => CLK,
                           Q => n_3550, QN => 
                           DataPath_RF_bus_reg_dataout_2528_port);
   DataPath_RF_BLOCKi_23_Q_reg_31_inst : DFF_X1 port map( D => n4010, CK => CLK
                           , Q => n_3551, QN => 
                           DataPath_RF_bus_reg_dataout_511_port);
   DataPath_RF_BLOCKi_23_Q_reg_30_inst : DFF_X1 port map( D => n4014, CK => CLK
                           , Q => n_3552, QN => 
                           DataPath_RF_bus_reg_dataout_510_port);
   DataPath_RF_BLOCKi_23_Q_reg_29_inst : DFF_X1 port map( D => n4016, CK => CLK
                           , Q => n_3553, QN => 
                           DataPath_RF_bus_reg_dataout_509_port);
   DataPath_RF_BLOCKi_23_Q_reg_28_inst : DFF_X1 port map( D => n4018, CK => CLK
                           , Q => n_3554, QN => 
                           DataPath_RF_bus_reg_dataout_508_port);
   DataPath_RF_BLOCKi_23_Q_reg_27_inst : DFF_X1 port map( D => n4020, CK => CLK
                           , Q => n_3555, QN => 
                           DataPath_RF_bus_reg_dataout_507_port);
   DataPath_RF_BLOCKi_23_Q_reg_26_inst : DFF_X1 port map( D => n4022, CK => CLK
                           , Q => n_3556, QN => 
                           DataPath_RF_bus_reg_dataout_506_port);
   DataPath_RF_BLOCKi_23_Q_reg_25_inst : DFF_X1 port map( D => n4024, CK => CLK
                           , Q => n_3557, QN => 
                           DataPath_RF_bus_reg_dataout_505_port);
   DataPath_RF_BLOCKi_23_Q_reg_24_inst : DFF_X1 port map( D => n4026, CK => CLK
                           , Q => n_3558, QN => 
                           DataPath_RF_bus_reg_dataout_504_port);
   DataPath_RF_BLOCKi_23_Q_reg_23_inst : DFF_X1 port map( D => n4028, CK => CLK
                           , Q => n_3559, QN => 
                           DataPath_RF_bus_reg_dataout_503_port);
   DataPath_RF_BLOCKi_23_Q_reg_22_inst : DFF_X1 port map( D => n4030, CK => CLK
                           , Q => n_3560, QN => 
                           DataPath_RF_bus_reg_dataout_502_port);
   DataPath_RF_BLOCKi_23_Q_reg_21_inst : DFF_X1 port map( D => n4032, CK => CLK
                           , Q => n_3561, QN => 
                           DataPath_RF_bus_reg_dataout_501_port);
   DataPath_RF_BLOCKi_23_Q_reg_20_inst : DFF_X1 port map( D => n4034, CK => CLK
                           , Q => n_3562, QN => 
                           DataPath_RF_bus_reg_dataout_500_port);
   DataPath_RF_BLOCKi_23_Q_reg_19_inst : DFF_X1 port map( D => n4036, CK => CLK
                           , Q => n_3563, QN => 
                           DataPath_RF_bus_reg_dataout_499_port);
   DataPath_RF_BLOCKi_23_Q_reg_18_inst : DFF_X1 port map( D => n4038, CK => CLK
                           , Q => n_3564, QN => 
                           DataPath_RF_bus_reg_dataout_498_port);
   DataPath_RF_BLOCKi_23_Q_reg_17_inst : DFF_X1 port map( D => n4040, CK => CLK
                           , Q => n_3565, QN => 
                           DataPath_RF_bus_reg_dataout_497_port);
   DataPath_RF_BLOCKi_23_Q_reg_16_inst : DFF_X1 port map( D => n4042, CK => CLK
                           , Q => n_3566, QN => 
                           DataPath_RF_bus_reg_dataout_496_port);
   DataPath_RF_BLOCKi_23_Q_reg_15_inst : DFF_X1 port map( D => n4044, CK => CLK
                           , Q => n_3567, QN => 
                           DataPath_RF_bus_reg_dataout_495_port);
   DataPath_RF_BLOCKi_23_Q_reg_14_inst : DFF_X1 port map( D => n4046, CK => CLK
                           , Q => n_3568, QN => 
                           DataPath_RF_bus_reg_dataout_494_port);
   DataPath_RF_BLOCKi_23_Q_reg_13_inst : DFF_X1 port map( D => n4048, CK => CLK
                           , Q => n_3569, QN => 
                           DataPath_RF_bus_reg_dataout_493_port);
   DataPath_RF_BLOCKi_23_Q_reg_12_inst : DFF_X1 port map( D => n4050, CK => CLK
                           , Q => n_3570, QN => 
                           DataPath_RF_bus_reg_dataout_492_port);
   DataPath_RF_BLOCKi_23_Q_reg_11_inst : DFF_X1 port map( D => n4052, CK => CLK
                           , Q => n_3571, QN => 
                           DataPath_RF_bus_reg_dataout_491_port);
   DataPath_RF_BLOCKi_23_Q_reg_9_inst : DFF_X1 port map( D => n4056, CK => CLK,
                           Q => n_3572, QN => 
                           DataPath_RF_bus_reg_dataout_489_port);
   DataPath_RF_BLOCKi_23_Q_reg_8_inst : DFF_X1 port map( D => n4058, CK => CLK,
                           Q => n_3573, QN => 
                           DataPath_RF_bus_reg_dataout_488_port);
   DataPath_RF_BLOCKi_23_Q_reg_7_inst : DFF_X1 port map( D => n4060, CK => CLK,
                           Q => n_3574, QN => 
                           DataPath_RF_bus_reg_dataout_487_port);
   DataPath_RF_BLOCKi_23_Q_reg_6_inst : DFF_X1 port map( D => n4062, CK => CLK,
                           Q => n_3575, QN => 
                           DataPath_RF_bus_reg_dataout_486_port);
   DataPath_RF_BLOCKi_23_Q_reg_5_inst : DFF_X1 port map( D => n4064, CK => CLK,
                           Q => n_3576, QN => 
                           DataPath_RF_bus_reg_dataout_485_port);
   DataPath_RF_BLOCKi_23_Q_reg_4_inst : DFF_X1 port map( D => n4066, CK => CLK,
                           Q => n_3577, QN => 
                           DataPath_RF_bus_reg_dataout_484_port);
   DataPath_RF_BLOCKi_23_Q_reg_3_inst : DFF_X1 port map( D => n4068, CK => CLK,
                           Q => n_3578, QN => 
                           DataPath_RF_bus_reg_dataout_483_port);
   DataPath_RF_BLOCKi_23_Q_reg_2_inst : DFF_X1 port map( D => n4070, CK => CLK,
                           Q => n_3579, QN => 
                           DataPath_RF_bus_reg_dataout_482_port);
   DataPath_RF_BLOCKi_23_Q_reg_1_inst : DFF_X1 port map( D => n4072, CK => CLK,
                           Q => n_3580, QN => 
                           DataPath_RF_bus_reg_dataout_481_port);
   DataPath_RF_BLOCKi_23_Q_reg_0_inst : DFF_X1 port map( D => n4074, CK => CLK,
                           Q => n_3581, QN => 
                           DataPath_RF_bus_reg_dataout_480_port);
   DataPath_RF_BLOCKi_39_Q_reg_31_inst : DFF_X1 port map( D => n4635, CK => CLK
                           , Q => n_3582, QN => 
                           DataPath_RF_bus_reg_dataout_1023_port);
   DataPath_RF_BLOCKi_39_Q_reg_30_inst : DFF_X1 port map( D => n4638, CK => CLK
                           , Q => n_3583, QN => 
                           DataPath_RF_bus_reg_dataout_1022_port);
   DataPath_RF_BLOCKi_39_Q_reg_29_inst : DFF_X1 port map( D => n4639, CK => CLK
                           , Q => n_3584, QN => 
                           DataPath_RF_bus_reg_dataout_1021_port);
   DataPath_RF_BLOCKi_39_Q_reg_28_inst : DFF_X1 port map( D => n4640, CK => CLK
                           , Q => n_3585, QN => 
                           DataPath_RF_bus_reg_dataout_1020_port);
   DataPath_RF_BLOCKi_39_Q_reg_27_inst : DFF_X1 port map( D => n4641, CK => CLK
                           , Q => n_3586, QN => 
                           DataPath_RF_bus_reg_dataout_1019_port);
   DataPath_RF_BLOCKi_39_Q_reg_26_inst : DFF_X1 port map( D => n4642, CK => CLK
                           , Q => n_3587, QN => 
                           DataPath_RF_bus_reg_dataout_1018_port);
   DataPath_RF_BLOCKi_39_Q_reg_25_inst : DFF_X1 port map( D => n4643, CK => CLK
                           , Q => n_3588, QN => 
                           DataPath_RF_bus_reg_dataout_1017_port);
   DataPath_RF_BLOCKi_39_Q_reg_24_inst : DFF_X1 port map( D => n4644, CK => CLK
                           , Q => n_3589, QN => 
                           DataPath_RF_bus_reg_dataout_1016_port);
   DataPath_RF_BLOCKi_39_Q_reg_23_inst : DFF_X1 port map( D => n4645, CK => CLK
                           , Q => n_3590, QN => 
                           DataPath_RF_bus_reg_dataout_1015_port);
   DataPath_RF_BLOCKi_39_Q_reg_22_inst : DFF_X1 port map( D => n4646, CK => CLK
                           , Q => n_3591, QN => 
                           DataPath_RF_bus_reg_dataout_1014_port);
   DataPath_RF_BLOCKi_39_Q_reg_21_inst : DFF_X1 port map( D => n4647, CK => CLK
                           , Q => n_3592, QN => 
                           DataPath_RF_bus_reg_dataout_1013_port);
   DataPath_RF_BLOCKi_39_Q_reg_20_inst : DFF_X1 port map( D => n4648, CK => CLK
                           , Q => n_3593, QN => 
                           DataPath_RF_bus_reg_dataout_1012_port);
   DataPath_RF_BLOCKi_39_Q_reg_19_inst : DFF_X1 port map( D => n4649, CK => CLK
                           , Q => n_3594, QN => 
                           DataPath_RF_bus_reg_dataout_1011_port);
   DataPath_RF_BLOCKi_39_Q_reg_18_inst : DFF_X1 port map( D => n4650, CK => CLK
                           , Q => n_3595, QN => 
                           DataPath_RF_bus_reg_dataout_1010_port);
   DataPath_RF_BLOCKi_39_Q_reg_17_inst : DFF_X1 port map( D => n4651, CK => CLK
                           , Q => n_3596, QN => 
                           DataPath_RF_bus_reg_dataout_1009_port);
   DataPath_RF_BLOCKi_39_Q_reg_16_inst : DFF_X1 port map( D => n4652, CK => CLK
                           , Q => n_3597, QN => 
                           DataPath_RF_bus_reg_dataout_1008_port);
   DataPath_RF_BLOCKi_39_Q_reg_15_inst : DFF_X1 port map( D => n4653, CK => CLK
                           , Q => n_3598, QN => 
                           DataPath_RF_bus_reg_dataout_1007_port);
   DataPath_RF_BLOCKi_39_Q_reg_14_inst : DFF_X1 port map( D => n4654, CK => CLK
                           , Q => n_3599, QN => 
                           DataPath_RF_bus_reg_dataout_1006_port);
   DataPath_RF_BLOCKi_39_Q_reg_13_inst : DFF_X1 port map( D => n4655, CK => CLK
                           , Q => n_3600, QN => 
                           DataPath_RF_bus_reg_dataout_1005_port);
   DataPath_RF_BLOCKi_39_Q_reg_12_inst : DFF_X1 port map( D => n4656, CK => CLK
                           , Q => n_3601, QN => 
                           DataPath_RF_bus_reg_dataout_1004_port);
   DataPath_RF_BLOCKi_39_Q_reg_11_inst : DFF_X1 port map( D => n4657, CK => CLK
                           , Q => n_3602, QN => 
                           DataPath_RF_bus_reg_dataout_1003_port);
   DataPath_RF_BLOCKi_39_Q_reg_9_inst : DFF_X1 port map( D => n4659, CK => CLK,
                           Q => n_3603, QN => 
                           DataPath_RF_bus_reg_dataout_1001_port);
   DataPath_RF_BLOCKi_39_Q_reg_8_inst : DFF_X1 port map( D => n4660, CK => CLK,
                           Q => n_3604, QN => 
                           DataPath_RF_bus_reg_dataout_1000_port);
   DataPath_RF_BLOCKi_39_Q_reg_7_inst : DFF_X1 port map( D => n4661, CK => CLK,
                           Q => n_3605, QN => 
                           DataPath_RF_bus_reg_dataout_999_port);
   DataPath_RF_BLOCKi_39_Q_reg_6_inst : DFF_X1 port map( D => n4662, CK => CLK,
                           Q => n_3606, QN => 
                           DataPath_RF_bus_reg_dataout_998_port);
   DataPath_RF_BLOCKi_39_Q_reg_5_inst : DFF_X1 port map( D => n4663, CK => CLK,
                           Q => n_3607, QN => 
                           DataPath_RF_bus_reg_dataout_997_port);
   DataPath_RF_BLOCKi_39_Q_reg_4_inst : DFF_X1 port map( D => n4664, CK => CLK,
                           Q => n_3608, QN => 
                           DataPath_RF_bus_reg_dataout_996_port);
   DataPath_RF_BLOCKi_39_Q_reg_3_inst : DFF_X1 port map( D => n4665, CK => CLK,
                           Q => n_3609, QN => 
                           DataPath_RF_bus_reg_dataout_995_port);
   DataPath_RF_BLOCKi_39_Q_reg_2_inst : DFF_X1 port map( D => n4666, CK => CLK,
                           Q => n_3610, QN => 
                           DataPath_RF_bus_reg_dataout_994_port);
   DataPath_RF_BLOCKi_39_Q_reg_1_inst : DFF_X1 port map( D => n4667, CK => CLK,
                           Q => n_3611, QN => 
                           DataPath_RF_bus_reg_dataout_993_port);
   DataPath_RF_BLOCKi_39_Q_reg_0_inst : DFF_X1 port map( D => n4668, CK => CLK,
                           Q => n_3612, QN => 
                           DataPath_RF_bus_reg_dataout_992_port);
   DataPath_RF_BLOCKi_55_Q_reg_31_inst : DFF_X1 port map( D => n5228, CK => CLK
                           , Q => n_3613, QN => 
                           DataPath_RF_bus_reg_dataout_1535_port);
   DataPath_RF_BLOCKi_55_Q_reg_30_inst : DFF_X1 port map( D => n5231, CK => CLK
                           , Q => n_3614, QN => 
                           DataPath_RF_bus_reg_dataout_1534_port);
   DataPath_RF_BLOCKi_55_Q_reg_29_inst : DFF_X1 port map( D => n5232, CK => CLK
                           , Q => n_3615, QN => 
                           DataPath_RF_bus_reg_dataout_1533_port);
   DataPath_RF_BLOCKi_55_Q_reg_28_inst : DFF_X1 port map( D => n5233, CK => CLK
                           , Q => n_3616, QN => 
                           DataPath_RF_bus_reg_dataout_1532_port);
   DataPath_RF_BLOCKi_55_Q_reg_27_inst : DFF_X1 port map( D => n5234, CK => CLK
                           , Q => n_3617, QN => 
                           DataPath_RF_bus_reg_dataout_1531_port);
   DataPath_RF_BLOCKi_55_Q_reg_26_inst : DFF_X1 port map( D => n5235, CK => CLK
                           , Q => n_3618, QN => 
                           DataPath_RF_bus_reg_dataout_1530_port);
   DataPath_RF_BLOCKi_55_Q_reg_25_inst : DFF_X1 port map( D => n5236, CK => CLK
                           , Q => n_3619, QN => 
                           DataPath_RF_bus_reg_dataout_1529_port);
   DataPath_RF_BLOCKi_55_Q_reg_24_inst : DFF_X1 port map( D => n5237, CK => CLK
                           , Q => n_3620, QN => 
                           DataPath_RF_bus_reg_dataout_1528_port);
   DataPath_RF_BLOCKi_55_Q_reg_23_inst : DFF_X1 port map( D => n5238, CK => CLK
                           , Q => n_3621, QN => 
                           DataPath_RF_bus_reg_dataout_1527_port);
   DataPath_RF_BLOCKi_55_Q_reg_22_inst : DFF_X1 port map( D => n5239, CK => CLK
                           , Q => n_3622, QN => 
                           DataPath_RF_bus_reg_dataout_1526_port);
   DataPath_RF_BLOCKi_55_Q_reg_21_inst : DFF_X1 port map( D => n5240, CK => CLK
                           , Q => n_3623, QN => 
                           DataPath_RF_bus_reg_dataout_1525_port);
   DataPath_RF_BLOCKi_55_Q_reg_20_inst : DFF_X1 port map( D => n5241, CK => CLK
                           , Q => n_3624, QN => 
                           DataPath_RF_bus_reg_dataout_1524_port);
   DataPath_RF_BLOCKi_55_Q_reg_19_inst : DFF_X1 port map( D => n5242, CK => CLK
                           , Q => n_3625, QN => 
                           DataPath_RF_bus_reg_dataout_1523_port);
   DataPath_RF_BLOCKi_55_Q_reg_18_inst : DFF_X1 port map( D => n5243, CK => CLK
                           , Q => n_3626, QN => 
                           DataPath_RF_bus_reg_dataout_1522_port);
   DataPath_RF_BLOCKi_55_Q_reg_17_inst : DFF_X1 port map( D => n5244, CK => CLK
                           , Q => n_3627, QN => 
                           DataPath_RF_bus_reg_dataout_1521_port);
   DataPath_RF_BLOCKi_55_Q_reg_16_inst : DFF_X1 port map( D => n5245, CK => CLK
                           , Q => n_3628, QN => 
                           DataPath_RF_bus_reg_dataout_1520_port);
   DataPath_RF_BLOCKi_55_Q_reg_15_inst : DFF_X1 port map( D => n5246, CK => CLK
                           , Q => n_3629, QN => 
                           DataPath_RF_bus_reg_dataout_1519_port);
   DataPath_RF_BLOCKi_55_Q_reg_14_inst : DFF_X1 port map( D => n5247, CK => CLK
                           , Q => n_3630, QN => 
                           DataPath_RF_bus_reg_dataout_1518_port);
   DataPath_RF_BLOCKi_55_Q_reg_13_inst : DFF_X1 port map( D => n5248, CK => CLK
                           , Q => n_3631, QN => 
                           DataPath_RF_bus_reg_dataout_1517_port);
   DataPath_RF_BLOCKi_55_Q_reg_12_inst : DFF_X1 port map( D => n5249, CK => CLK
                           , Q => n_3632, QN => 
                           DataPath_RF_bus_reg_dataout_1516_port);
   DataPath_RF_BLOCKi_55_Q_reg_11_inst : DFF_X1 port map( D => n5250, CK => CLK
                           , Q => n_3633, QN => 
                           DataPath_RF_bus_reg_dataout_1515_port);
   DataPath_RF_BLOCKi_55_Q_reg_9_inst : DFF_X1 port map( D => n5252, CK => CLK,
                           Q => n_3634, QN => 
                           DataPath_RF_bus_reg_dataout_1513_port);
   DataPath_RF_BLOCKi_55_Q_reg_8_inst : DFF_X1 port map( D => n5253, CK => CLK,
                           Q => n_3635, QN => 
                           DataPath_RF_bus_reg_dataout_1512_port);
   DataPath_RF_BLOCKi_55_Q_reg_7_inst : DFF_X1 port map( D => n5254, CK => CLK,
                           Q => n_3636, QN => 
                           DataPath_RF_bus_reg_dataout_1511_port);
   DataPath_RF_BLOCKi_55_Q_reg_6_inst : DFF_X1 port map( D => n5255, CK => CLK,
                           Q => n_3637, QN => 
                           DataPath_RF_bus_reg_dataout_1510_port);
   DataPath_RF_BLOCKi_55_Q_reg_5_inst : DFF_X1 port map( D => n5256, CK => CLK,
                           Q => n_3638, QN => 
                           DataPath_RF_bus_reg_dataout_1509_port);
   DataPath_RF_BLOCKi_55_Q_reg_4_inst : DFF_X1 port map( D => n5257, CK => CLK,
                           Q => n_3639, QN => 
                           DataPath_RF_bus_reg_dataout_1508_port);
   DataPath_RF_BLOCKi_55_Q_reg_3_inst : DFF_X1 port map( D => n5258, CK => CLK,
                           Q => n_3640, QN => 
                           DataPath_RF_bus_reg_dataout_1507_port);
   DataPath_RF_BLOCKi_55_Q_reg_2_inst : DFF_X1 port map( D => n5259, CK => CLK,
                           Q => n_3641, QN => 
                           DataPath_RF_bus_reg_dataout_1506_port);
   DataPath_RF_BLOCKi_55_Q_reg_1_inst : DFF_X1 port map( D => n5260, CK => CLK,
                           Q => n_3642, QN => 
                           DataPath_RF_bus_reg_dataout_1505_port);
   DataPath_RF_BLOCKi_55_Q_reg_0_inst : DFF_X1 port map( D => n5261, CK => CLK,
                           Q => n_3643, QN => 
                           DataPath_RF_bus_reg_dataout_1504_port);
   DataPath_RF_BLOCKi_71_Q_reg_31_inst : DFF_X1 port map( D => n5831, CK => CLK
                           , Q => n_3644, QN => 
                           DataPath_RF_bus_reg_dataout_2047_port);
   DataPath_RF_BLOCKi_71_Q_reg_30_inst : DFF_X1 port map( D => n5834, CK => CLK
                           , Q => n_3645, QN => 
                           DataPath_RF_bus_reg_dataout_2046_port);
   DataPath_RF_BLOCKi_71_Q_reg_29_inst : DFF_X1 port map( D => n5835, CK => CLK
                           , Q => n_3646, QN => 
                           DataPath_RF_bus_reg_dataout_2045_port);
   DataPath_RF_BLOCKi_71_Q_reg_28_inst : DFF_X1 port map( D => n5836, CK => CLK
                           , Q => n_3647, QN => 
                           DataPath_RF_bus_reg_dataout_2044_port);
   DataPath_RF_BLOCKi_71_Q_reg_27_inst : DFF_X1 port map( D => n5837, CK => CLK
                           , Q => n_3648, QN => 
                           DataPath_RF_bus_reg_dataout_2043_port);
   DataPath_RF_BLOCKi_71_Q_reg_26_inst : DFF_X1 port map( D => n5838, CK => CLK
                           , Q => n_3649, QN => 
                           DataPath_RF_bus_reg_dataout_2042_port);
   DataPath_RF_BLOCKi_71_Q_reg_25_inst : DFF_X1 port map( D => n5839, CK => CLK
                           , Q => n_3650, QN => 
                           DataPath_RF_bus_reg_dataout_2041_port);
   DataPath_RF_BLOCKi_71_Q_reg_24_inst : DFF_X1 port map( D => n5840, CK => CLK
                           , Q => n_3651, QN => 
                           DataPath_RF_bus_reg_dataout_2040_port);
   DataPath_RF_BLOCKi_71_Q_reg_23_inst : DFF_X1 port map( D => n5841, CK => CLK
                           , Q => n_3652, QN => 
                           DataPath_RF_bus_reg_dataout_2039_port);
   DataPath_RF_BLOCKi_71_Q_reg_22_inst : DFF_X1 port map( D => n5842, CK => CLK
                           , Q => n_3653, QN => 
                           DataPath_RF_bus_reg_dataout_2038_port);
   DataPath_RF_BLOCKi_71_Q_reg_21_inst : DFF_X1 port map( D => n5843, CK => CLK
                           , Q => n_3654, QN => 
                           DataPath_RF_bus_reg_dataout_2037_port);
   DataPath_RF_BLOCKi_71_Q_reg_20_inst : DFF_X1 port map( D => n5844, CK => CLK
                           , Q => n_3655, QN => 
                           DataPath_RF_bus_reg_dataout_2036_port);
   DataPath_RF_BLOCKi_71_Q_reg_19_inst : DFF_X1 port map( D => n5845, CK => CLK
                           , Q => n_3656, QN => 
                           DataPath_RF_bus_reg_dataout_2035_port);
   DataPath_RF_BLOCKi_71_Q_reg_18_inst : DFF_X1 port map( D => n5846, CK => CLK
                           , Q => n_3657, QN => 
                           DataPath_RF_bus_reg_dataout_2034_port);
   DataPath_RF_BLOCKi_71_Q_reg_17_inst : DFF_X1 port map( D => n5847, CK => CLK
                           , Q => n_3658, QN => 
                           DataPath_RF_bus_reg_dataout_2033_port);
   DataPath_RF_BLOCKi_71_Q_reg_16_inst : DFF_X1 port map( D => n5848, CK => CLK
                           , Q => n_3659, QN => 
                           DataPath_RF_bus_reg_dataout_2032_port);
   DataPath_RF_BLOCKi_71_Q_reg_15_inst : DFF_X1 port map( D => n5849, CK => CLK
                           , Q => n_3660, QN => 
                           DataPath_RF_bus_reg_dataout_2031_port);
   DataPath_RF_BLOCKi_71_Q_reg_14_inst : DFF_X1 port map( D => n5850, CK => CLK
                           , Q => n_3661, QN => 
                           DataPath_RF_bus_reg_dataout_2030_port);
   DataPath_RF_BLOCKi_71_Q_reg_13_inst : DFF_X1 port map( D => n5851, CK => CLK
                           , Q => n_3662, QN => 
                           DataPath_RF_bus_reg_dataout_2029_port);
   DataPath_RF_BLOCKi_71_Q_reg_12_inst : DFF_X1 port map( D => n5852, CK => CLK
                           , Q => n_3663, QN => 
                           DataPath_RF_bus_reg_dataout_2028_port);
   DataPath_RF_BLOCKi_71_Q_reg_11_inst : DFF_X1 port map( D => n5853, CK => CLK
                           , Q => n_3664, QN => 
                           DataPath_RF_bus_reg_dataout_2027_port);
   DataPath_RF_BLOCKi_71_Q_reg_9_inst : DFF_X1 port map( D => n5855, CK => CLK,
                           Q => n_3665, QN => 
                           DataPath_RF_bus_reg_dataout_2025_port);
   DataPath_RF_BLOCKi_71_Q_reg_8_inst : DFF_X1 port map( D => n5856, CK => CLK,
                           Q => n_3666, QN => 
                           DataPath_RF_bus_reg_dataout_2024_port);
   DataPath_RF_BLOCKi_71_Q_reg_7_inst : DFF_X1 port map( D => n5857, CK => CLK,
                           Q => n_3667, QN => 
                           DataPath_RF_bus_reg_dataout_2023_port);
   DataPath_RF_BLOCKi_71_Q_reg_6_inst : DFF_X1 port map( D => n5858, CK => CLK,
                           Q => n_3668, QN => 
                           DataPath_RF_bus_reg_dataout_2022_port);
   DataPath_RF_BLOCKi_71_Q_reg_5_inst : DFF_X1 port map( D => n5859, CK => CLK,
                           Q => n_3669, QN => 
                           DataPath_RF_bus_reg_dataout_2021_port);
   DataPath_RF_BLOCKi_71_Q_reg_4_inst : DFF_X1 port map( D => n5860, CK => CLK,
                           Q => n_3670, QN => 
                           DataPath_RF_bus_reg_dataout_2020_port);
   DataPath_RF_BLOCKi_71_Q_reg_3_inst : DFF_X1 port map( D => n5861, CK => CLK,
                           Q => n_3671, QN => 
                           DataPath_RF_bus_reg_dataout_2019_port);
   DataPath_RF_BLOCKi_71_Q_reg_2_inst : DFF_X1 port map( D => n5862, CK => CLK,
                           Q => n_3672, QN => 
                           DataPath_RF_bus_reg_dataout_2018_port);
   DataPath_RF_BLOCKi_71_Q_reg_1_inst : DFF_X1 port map( D => n5863, CK => CLK,
                           Q => n_3673, QN => 
                           DataPath_RF_bus_reg_dataout_2017_port);
   DataPath_RF_BLOCKi_71_Q_reg_0_inst : DFF_X1 port map( D => n5864, CK => CLK,
                           Q => n_3674, QN => 
                           DataPath_RF_bus_reg_dataout_2016_port);
   DataPath_RF_BLOCKi_80_Q_reg_31_inst : DFF_X1 port map( D => n913, CK => CLK,
                           Q => n_3675, QN => 
                           DataPath_RF_bus_reg_dataout_2335_port);
   DataPath_RF_BLOCKi_80_Q_reg_30_inst : DFF_X1 port map( D => n917, CK => CLK,
                           Q => n_3676, QN => 
                           DataPath_RF_bus_reg_dataout_2334_port);
   DataPath_RF_BLOCKi_80_Q_reg_29_inst : DFF_X1 port map( D => n919, CK => CLK,
                           Q => n_3677, QN => 
                           DataPath_RF_bus_reg_dataout_2333_port);
   DataPath_RF_BLOCKi_80_Q_reg_28_inst : DFF_X1 port map( D => n921, CK => CLK,
                           Q => n_3678, QN => 
                           DataPath_RF_bus_reg_dataout_2332_port);
   DataPath_RF_BLOCKi_80_Q_reg_27_inst : DFF_X1 port map( D => n923, CK => CLK,
                           Q => n_3679, QN => 
                           DataPath_RF_bus_reg_dataout_2331_port);
   DataPath_RF_BLOCKi_80_Q_reg_26_inst : DFF_X1 port map( D => n925, CK => CLK,
                           Q => n_3680, QN => 
                           DataPath_RF_bus_reg_dataout_2330_port);
   DataPath_RF_BLOCKi_80_Q_reg_25_inst : DFF_X1 port map( D => n927, CK => CLK,
                           Q => n_3681, QN => 
                           DataPath_RF_bus_reg_dataout_2329_port);
   DataPath_RF_BLOCKi_80_Q_reg_24_inst : DFF_X1 port map( D => n929, CK => CLK,
                           Q => n_3682, QN => 
                           DataPath_RF_bus_reg_dataout_2328_port);
   DataPath_RF_BLOCKi_80_Q_reg_23_inst : DFF_X1 port map( D => n931, CK => CLK,
                           Q => n_3683, QN => 
                           DataPath_RF_bus_reg_dataout_2327_port);
   DataPath_RF_BLOCKi_80_Q_reg_22_inst : DFF_X1 port map( D => n933, CK => CLK,
                           Q => n_3684, QN => 
                           DataPath_RF_bus_reg_dataout_2326_port);
   DataPath_RF_BLOCKi_80_Q_reg_21_inst : DFF_X1 port map( D => n935, CK => CLK,
                           Q => n_3685, QN => 
                           DataPath_RF_bus_reg_dataout_2325_port);
   DataPath_RF_BLOCKi_80_Q_reg_20_inst : DFF_X1 port map( D => n937, CK => CLK,
                           Q => n_3686, QN => 
                           DataPath_RF_bus_reg_dataout_2324_port);
   DataPath_RF_BLOCKi_80_Q_reg_19_inst : DFF_X1 port map( D => n939, CK => CLK,
                           Q => n_3687, QN => 
                           DataPath_RF_bus_reg_dataout_2323_port);
   DataPath_RF_BLOCKi_80_Q_reg_18_inst : DFF_X1 port map( D => n941, CK => CLK,
                           Q => n_3688, QN => 
                           DataPath_RF_bus_reg_dataout_2322_port);
   DataPath_RF_BLOCKi_80_Q_reg_17_inst : DFF_X1 port map( D => n943, CK => CLK,
                           Q => n_3689, QN => 
                           DataPath_RF_bus_reg_dataout_2321_port);
   DataPath_RF_BLOCKi_80_Q_reg_16_inst : DFF_X1 port map( D => n945, CK => CLK,
                           Q => n_3690, QN => 
                           DataPath_RF_bus_reg_dataout_2320_port);
   DataPath_RF_BLOCKi_80_Q_reg_15_inst : DFF_X1 port map( D => n947, CK => CLK,
                           Q => n_3691, QN => 
                           DataPath_RF_bus_reg_dataout_2319_port);
   DataPath_RF_BLOCKi_80_Q_reg_14_inst : DFF_X1 port map( D => n948, CK => CLK,
                           Q => n_3692, QN => 
                           DataPath_RF_bus_reg_dataout_2318_port);
   DataPath_RF_BLOCKi_80_Q_reg_13_inst : DFF_X1 port map( D => n949, CK => CLK,
                           Q => n_3693, QN => 
                           DataPath_RF_bus_reg_dataout_2317_port);
   DataPath_RF_BLOCKi_80_Q_reg_12_inst : DFF_X1 port map( D => n950, CK => CLK,
                           Q => n_3694, QN => 
                           DataPath_RF_bus_reg_dataout_2316_port);
   DataPath_RF_BLOCKi_80_Q_reg_11_inst : DFF_X1 port map( D => n951, CK => CLK,
                           Q => n_3695, QN => 
                           DataPath_RF_bus_reg_dataout_2315_port);
   DataPath_RF_BLOCKi_80_Q_reg_9_inst : DFF_X1 port map( D => n953, CK => CLK, 
                           Q => n_3696, QN => 
                           DataPath_RF_bus_reg_dataout_2313_port);
   DataPath_RF_BLOCKi_80_Q_reg_8_inst : DFF_X1 port map( D => n954, CK => CLK, 
                           Q => n_3697, QN => 
                           DataPath_RF_bus_reg_dataout_2312_port);
   DataPath_RF_BLOCKi_80_Q_reg_7_inst : DFF_X1 port map( D => n955, CK => CLK, 
                           Q => n_3698, QN => 
                           DataPath_RF_bus_reg_dataout_2311_port);
   DataPath_RF_BLOCKi_80_Q_reg_6_inst : DFF_X1 port map( D => n956, CK => CLK, 
                           Q => n_3699, QN => 
                           DataPath_RF_bus_reg_dataout_2310_port);
   DataPath_RF_BLOCKi_80_Q_reg_5_inst : DFF_X1 port map( D => n957, CK => CLK, 
                           Q => n_3700, QN => 
                           DataPath_RF_bus_reg_dataout_2309_port);
   DataPath_RF_BLOCKi_80_Q_reg_4_inst : DFF_X1 port map( D => n958, CK => CLK, 
                           Q => n_3701, QN => 
                           DataPath_RF_bus_reg_dataout_2308_port);
   DataPath_RF_BLOCKi_80_Q_reg_3_inst : DFF_X1 port map( D => n959, CK => CLK, 
                           Q => n_3702, QN => 
                           DataPath_RF_bus_reg_dataout_2307_port);
   DataPath_RF_BLOCKi_80_Q_reg_2_inst : DFF_X1 port map( D => n960, CK => CLK, 
                           Q => n_3703, QN => 
                           DataPath_RF_bus_reg_dataout_2306_port);
   DataPath_RF_BLOCKi_80_Q_reg_1_inst : DFF_X1 port map( D => n961, CK => CLK, 
                           Q => n_3704, QN => 
                           DataPath_RF_bus_reg_dataout_2305_port);
   DataPath_RF_BLOCKi_80_Q_reg_0_inst : DFF_X1 port map( D => n962, CK => CLK, 
                           Q => n_3705, QN => 
                           DataPath_RF_bus_reg_dataout_2304_port);
   DataPath_RF_BLOCKi_16_Q_reg_31_inst : DFF_X1 port map( D => n3765, CK => CLK
                           , Q => n_3706, QN => 
                           DataPath_RF_bus_reg_dataout_287_port);
   DataPath_RF_BLOCKi_16_Q_reg_30_inst : DFF_X1 port map( D => n3768, CK => CLK
                           , Q => n_3707, QN => 
                           DataPath_RF_bus_reg_dataout_286_port);
   DataPath_RF_BLOCKi_16_Q_reg_29_inst : DFF_X1 port map( D => n3769, CK => CLK
                           , Q => n_3708, QN => 
                           DataPath_RF_bus_reg_dataout_285_port);
   DataPath_RF_BLOCKi_16_Q_reg_28_inst : DFF_X1 port map( D => n3770, CK => CLK
                           , Q => n_3709, QN => 
                           DataPath_RF_bus_reg_dataout_284_port);
   DataPath_RF_BLOCKi_16_Q_reg_27_inst : DFF_X1 port map( D => n3771, CK => CLK
                           , Q => n_3710, QN => 
                           DataPath_RF_bus_reg_dataout_283_port);
   DataPath_RF_BLOCKi_16_Q_reg_26_inst : DFF_X1 port map( D => n3772, CK => CLK
                           , Q => n_3711, QN => 
                           DataPath_RF_bus_reg_dataout_282_port);
   DataPath_RF_BLOCKi_16_Q_reg_25_inst : DFF_X1 port map( D => n3773, CK => CLK
                           , Q => n_3712, QN => 
                           DataPath_RF_bus_reg_dataout_281_port);
   DataPath_RF_BLOCKi_16_Q_reg_24_inst : DFF_X1 port map( D => n3774, CK => CLK
                           , Q => n_3713, QN => 
                           DataPath_RF_bus_reg_dataout_280_port);
   DataPath_RF_BLOCKi_16_Q_reg_23_inst : DFF_X1 port map( D => n3775, CK => CLK
                           , Q => n_3714, QN => 
                           DataPath_RF_bus_reg_dataout_279_port);
   DataPath_RF_BLOCKi_16_Q_reg_22_inst : DFF_X1 port map( D => n3776, CK => CLK
                           , Q => n_3715, QN => 
                           DataPath_RF_bus_reg_dataout_278_port);
   DataPath_RF_BLOCKi_16_Q_reg_21_inst : DFF_X1 port map( D => n3777, CK => CLK
                           , Q => n_3716, QN => 
                           DataPath_RF_bus_reg_dataout_277_port);
   DataPath_RF_BLOCKi_16_Q_reg_20_inst : DFF_X1 port map( D => n3778, CK => CLK
                           , Q => n_3717, QN => 
                           DataPath_RF_bus_reg_dataout_276_port);
   DataPath_RF_BLOCKi_16_Q_reg_19_inst : DFF_X1 port map( D => n3779, CK => CLK
                           , Q => n_3718, QN => 
                           DataPath_RF_bus_reg_dataout_275_port);
   DataPath_RF_BLOCKi_16_Q_reg_18_inst : DFF_X1 port map( D => n3780, CK => CLK
                           , Q => n_3719, QN => 
                           DataPath_RF_bus_reg_dataout_274_port);
   DataPath_RF_BLOCKi_16_Q_reg_17_inst : DFF_X1 port map( D => n3781, CK => CLK
                           , Q => n_3720, QN => 
                           DataPath_RF_bus_reg_dataout_273_port);
   DataPath_RF_BLOCKi_16_Q_reg_16_inst : DFF_X1 port map( D => n3782, CK => CLK
                           , Q => n_3721, QN => 
                           DataPath_RF_bus_reg_dataout_272_port);
   DataPath_RF_BLOCKi_16_Q_reg_15_inst : DFF_X1 port map( D => n3783, CK => CLK
                           , Q => n_3722, QN => 
                           DataPath_RF_bus_reg_dataout_271_port);
   DataPath_RF_BLOCKi_16_Q_reg_14_inst : DFF_X1 port map( D => n3784, CK => CLK
                           , Q => n_3723, QN => 
                           DataPath_RF_bus_reg_dataout_270_port);
   DataPath_RF_BLOCKi_16_Q_reg_13_inst : DFF_X1 port map( D => n3785, CK => CLK
                           , Q => n_3724, QN => 
                           DataPath_RF_bus_reg_dataout_269_port);
   DataPath_RF_BLOCKi_16_Q_reg_12_inst : DFF_X1 port map( D => n3786, CK => CLK
                           , Q => n_3725, QN => 
                           DataPath_RF_bus_reg_dataout_268_port);
   DataPath_RF_BLOCKi_16_Q_reg_11_inst : DFF_X1 port map( D => n3787, CK => CLK
                           , Q => n_3726, QN => 
                           DataPath_RF_bus_reg_dataout_267_port);
   DataPath_RF_BLOCKi_16_Q_reg_9_inst : DFF_X1 port map( D => n3789, CK => CLK,
                           Q => n_3727, QN => 
                           DataPath_RF_bus_reg_dataout_265_port);
   DataPath_RF_BLOCKi_16_Q_reg_8_inst : DFF_X1 port map( D => n3790, CK => CLK,
                           Q => n_3728, QN => 
                           DataPath_RF_bus_reg_dataout_264_port);
   DataPath_RF_BLOCKi_16_Q_reg_7_inst : DFF_X1 port map( D => n3791, CK => CLK,
                           Q => n_3729, QN => 
                           DataPath_RF_bus_reg_dataout_263_port);
   DataPath_RF_BLOCKi_16_Q_reg_6_inst : DFF_X1 port map( D => n3792, CK => CLK,
                           Q => n_3730, QN => 
                           DataPath_RF_bus_reg_dataout_262_port);
   DataPath_RF_BLOCKi_16_Q_reg_5_inst : DFF_X1 port map( D => n3793, CK => CLK,
                           Q => n_3731, QN => 
                           DataPath_RF_bus_reg_dataout_261_port);
   DataPath_RF_BLOCKi_16_Q_reg_4_inst : DFF_X1 port map( D => n3794, CK => CLK,
                           Q => n_3732, QN => 
                           DataPath_RF_bus_reg_dataout_260_port);
   DataPath_RF_BLOCKi_16_Q_reg_3_inst : DFF_X1 port map( D => n3795, CK => CLK,
                           Q => n_3733, QN => 
                           DataPath_RF_bus_reg_dataout_259_port);
   DataPath_RF_BLOCKi_16_Q_reg_2_inst : DFF_X1 port map( D => n3796, CK => CLK,
                           Q => n_3734, QN => 
                           DataPath_RF_bus_reg_dataout_258_port);
   DataPath_RF_BLOCKi_16_Q_reg_1_inst : DFF_X1 port map( D => n3797, CK => CLK,
                           Q => n_3735, QN => 
                           DataPath_RF_bus_reg_dataout_257_port);
   DataPath_RF_BLOCKi_16_Q_reg_0_inst : DFF_X1 port map( D => n3798, CK => CLK,
                           Q => n_3736, QN => 
                           DataPath_RF_bus_reg_dataout_256_port);
   DataPath_RF_BLOCKi_32_Q_reg_31_inst : DFF_X1 port map( D => n4390, CK => CLK
                           , Q => n_3737, QN => 
                           DataPath_RF_bus_reg_dataout_799_port);
   DataPath_RF_BLOCKi_32_Q_reg_30_inst : DFF_X1 port map( D => n4393, CK => CLK
                           , Q => n_3738, QN => 
                           DataPath_RF_bus_reg_dataout_798_port);
   DataPath_RF_BLOCKi_32_Q_reg_29_inst : DFF_X1 port map( D => n4394, CK => CLK
                           , Q => n_3739, QN => 
                           DataPath_RF_bus_reg_dataout_797_port);
   DataPath_RF_BLOCKi_32_Q_reg_28_inst : DFF_X1 port map( D => n4395, CK => CLK
                           , Q => n_3740, QN => 
                           DataPath_RF_bus_reg_dataout_796_port);
   DataPath_RF_BLOCKi_32_Q_reg_27_inst : DFF_X1 port map( D => n4396, CK => CLK
                           , Q => n_3741, QN => 
                           DataPath_RF_bus_reg_dataout_795_port);
   DataPath_RF_BLOCKi_32_Q_reg_26_inst : DFF_X1 port map( D => n4397, CK => CLK
                           , Q => n_3742, QN => 
                           DataPath_RF_bus_reg_dataout_794_port);
   DataPath_RF_BLOCKi_32_Q_reg_25_inst : DFF_X1 port map( D => n4398, CK => CLK
                           , Q => n_3743, QN => 
                           DataPath_RF_bus_reg_dataout_793_port);
   DataPath_RF_BLOCKi_32_Q_reg_24_inst : DFF_X1 port map( D => n4399, CK => CLK
                           , Q => n_3744, QN => 
                           DataPath_RF_bus_reg_dataout_792_port);
   DataPath_RF_BLOCKi_32_Q_reg_23_inst : DFF_X1 port map( D => n4400, CK => CLK
                           , Q => n_3745, QN => 
                           DataPath_RF_bus_reg_dataout_791_port);
   DataPath_RF_BLOCKi_32_Q_reg_22_inst : DFF_X1 port map( D => n4401, CK => CLK
                           , Q => n_3746, QN => 
                           DataPath_RF_bus_reg_dataout_790_port);
   DataPath_RF_BLOCKi_32_Q_reg_21_inst : DFF_X1 port map( D => n4402, CK => CLK
                           , Q => n_3747, QN => 
                           DataPath_RF_bus_reg_dataout_789_port);
   DataPath_RF_BLOCKi_32_Q_reg_20_inst : DFF_X1 port map( D => n4403, CK => CLK
                           , Q => n_3748, QN => 
                           DataPath_RF_bus_reg_dataout_788_port);
   DataPath_RF_BLOCKi_32_Q_reg_19_inst : DFF_X1 port map( D => n4404, CK => CLK
                           , Q => n_3749, QN => 
                           DataPath_RF_bus_reg_dataout_787_port);
   DataPath_RF_BLOCKi_32_Q_reg_18_inst : DFF_X1 port map( D => n4405, CK => CLK
                           , Q => n_3750, QN => 
                           DataPath_RF_bus_reg_dataout_786_port);
   DataPath_RF_BLOCKi_32_Q_reg_17_inst : DFF_X1 port map( D => n4406, CK => CLK
                           , Q => n_3751, QN => 
                           DataPath_RF_bus_reg_dataout_785_port);
   DataPath_RF_BLOCKi_32_Q_reg_16_inst : DFF_X1 port map( D => n4407, CK => CLK
                           , Q => n_3752, QN => 
                           DataPath_RF_bus_reg_dataout_784_port);
   DataPath_RF_BLOCKi_32_Q_reg_15_inst : DFF_X1 port map( D => n4408, CK => CLK
                           , Q => n_3753, QN => 
                           DataPath_RF_bus_reg_dataout_783_port);
   DataPath_RF_BLOCKi_32_Q_reg_14_inst : DFF_X1 port map( D => n4409, CK => CLK
                           , Q => n_3754, QN => 
                           DataPath_RF_bus_reg_dataout_782_port);
   DataPath_RF_BLOCKi_32_Q_reg_13_inst : DFF_X1 port map( D => n4410, CK => CLK
                           , Q => n_3755, QN => 
                           DataPath_RF_bus_reg_dataout_781_port);
   DataPath_RF_BLOCKi_32_Q_reg_12_inst : DFF_X1 port map( D => n4411, CK => CLK
                           , Q => n_3756, QN => 
                           DataPath_RF_bus_reg_dataout_780_port);
   DataPath_RF_BLOCKi_32_Q_reg_11_inst : DFF_X1 port map( D => n4412, CK => CLK
                           , Q => n_3757, QN => 
                           DataPath_RF_bus_reg_dataout_779_port);
   DataPath_RF_BLOCKi_32_Q_reg_9_inst : DFF_X1 port map( D => n4414, CK => CLK,
                           Q => n_3758, QN => 
                           DataPath_RF_bus_reg_dataout_777_port);
   DataPath_RF_BLOCKi_32_Q_reg_8_inst : DFF_X1 port map( D => n4415, CK => CLK,
                           Q => n_3759, QN => 
                           DataPath_RF_bus_reg_dataout_776_port);
   DataPath_RF_BLOCKi_32_Q_reg_7_inst : DFF_X1 port map( D => n4416, CK => CLK,
                           Q => n_3760, QN => 
                           DataPath_RF_bus_reg_dataout_775_port);
   DataPath_RF_BLOCKi_32_Q_reg_6_inst : DFF_X1 port map( D => n4417, CK => CLK,
                           Q => n_3761, QN => 
                           DataPath_RF_bus_reg_dataout_774_port);
   DataPath_RF_BLOCKi_32_Q_reg_5_inst : DFF_X1 port map( D => n4418, CK => CLK,
                           Q => n_3762, QN => 
                           DataPath_RF_bus_reg_dataout_773_port);
   DataPath_RF_BLOCKi_32_Q_reg_4_inst : DFF_X1 port map( D => n4419, CK => CLK,
                           Q => n_3763, QN => 
                           DataPath_RF_bus_reg_dataout_772_port);
   DataPath_RF_BLOCKi_32_Q_reg_3_inst : DFF_X1 port map( D => n4420, CK => CLK,
                           Q => n_3764, QN => 
                           DataPath_RF_bus_reg_dataout_771_port);
   DataPath_RF_BLOCKi_32_Q_reg_2_inst : DFF_X1 port map( D => n4421, CK => CLK,
                           Q => n_3765, QN => 
                           DataPath_RF_bus_reg_dataout_770_port);
   DataPath_RF_BLOCKi_32_Q_reg_1_inst : DFF_X1 port map( D => n4422, CK => CLK,
                           Q => n_3766, QN => 
                           DataPath_RF_bus_reg_dataout_769_port);
   DataPath_RF_BLOCKi_32_Q_reg_0_inst : DFF_X1 port map( D => n4423, CK => CLK,
                           Q => n_3767, QN => 
                           DataPath_RF_bus_reg_dataout_768_port);
   DataPath_RF_BLOCKi_48_Q_reg_31_inst : DFF_X1 port map( D => n4983, CK => CLK
                           , Q => n_3768, QN => 
                           DataPath_RF_bus_reg_dataout_1311_port);
   DataPath_RF_BLOCKi_48_Q_reg_30_inst : DFF_X1 port map( D => n4986, CK => CLK
                           , Q => n_3769, QN => 
                           DataPath_RF_bus_reg_dataout_1310_port);
   DataPath_RF_BLOCKi_48_Q_reg_29_inst : DFF_X1 port map( D => n4987, CK => CLK
                           , Q => n_3770, QN => 
                           DataPath_RF_bus_reg_dataout_1309_port);
   DataPath_RF_BLOCKi_48_Q_reg_28_inst : DFF_X1 port map( D => n4988, CK => CLK
                           , Q => n_3771, QN => 
                           DataPath_RF_bus_reg_dataout_1308_port);
   DataPath_RF_BLOCKi_48_Q_reg_27_inst : DFF_X1 port map( D => n4989, CK => CLK
                           , Q => n_3772, QN => 
                           DataPath_RF_bus_reg_dataout_1307_port);
   DataPath_RF_BLOCKi_48_Q_reg_26_inst : DFF_X1 port map( D => n4990, CK => CLK
                           , Q => n_3773, QN => 
                           DataPath_RF_bus_reg_dataout_1306_port);
   DataPath_RF_BLOCKi_48_Q_reg_25_inst : DFF_X1 port map( D => n4991, CK => CLK
                           , Q => n_3774, QN => 
                           DataPath_RF_bus_reg_dataout_1305_port);
   DataPath_RF_BLOCKi_48_Q_reg_24_inst : DFF_X1 port map( D => n4992, CK => CLK
                           , Q => n_3775, QN => 
                           DataPath_RF_bus_reg_dataout_1304_port);
   DataPath_RF_BLOCKi_48_Q_reg_23_inst : DFF_X1 port map( D => n4993, CK => CLK
                           , Q => n_3776, QN => 
                           DataPath_RF_bus_reg_dataout_1303_port);
   DataPath_RF_BLOCKi_48_Q_reg_22_inst : DFF_X1 port map( D => n4994, CK => CLK
                           , Q => n_3777, QN => 
                           DataPath_RF_bus_reg_dataout_1302_port);
   DataPath_RF_BLOCKi_48_Q_reg_21_inst : DFF_X1 port map( D => n4995, CK => CLK
                           , Q => n_3778, QN => 
                           DataPath_RF_bus_reg_dataout_1301_port);
   DataPath_RF_BLOCKi_48_Q_reg_20_inst : DFF_X1 port map( D => n4996, CK => CLK
                           , Q => n_3779, QN => 
                           DataPath_RF_bus_reg_dataout_1300_port);
   DataPath_RF_BLOCKi_48_Q_reg_19_inst : DFF_X1 port map( D => n4997, CK => CLK
                           , Q => n_3780, QN => 
                           DataPath_RF_bus_reg_dataout_1299_port);
   DataPath_RF_BLOCKi_48_Q_reg_18_inst : DFF_X1 port map( D => n4998, CK => CLK
                           , Q => n_3781, QN => 
                           DataPath_RF_bus_reg_dataout_1298_port);
   DataPath_RF_BLOCKi_48_Q_reg_17_inst : DFF_X1 port map( D => n4999, CK => CLK
                           , Q => n_3782, QN => 
                           DataPath_RF_bus_reg_dataout_1297_port);
   DataPath_RF_BLOCKi_48_Q_reg_16_inst : DFF_X1 port map( D => n5000, CK => CLK
                           , Q => n_3783, QN => 
                           DataPath_RF_bus_reg_dataout_1296_port);
   DataPath_RF_BLOCKi_48_Q_reg_15_inst : DFF_X1 port map( D => n5001, CK => CLK
                           , Q => n_3784, QN => 
                           DataPath_RF_bus_reg_dataout_1295_port);
   DataPath_RF_BLOCKi_48_Q_reg_14_inst : DFF_X1 port map( D => n5002, CK => CLK
                           , Q => n_3785, QN => 
                           DataPath_RF_bus_reg_dataout_1294_port);
   DataPath_RF_BLOCKi_48_Q_reg_13_inst : DFF_X1 port map( D => n5003, CK => CLK
                           , Q => n_3786, QN => 
                           DataPath_RF_bus_reg_dataout_1293_port);
   DataPath_RF_BLOCKi_48_Q_reg_12_inst : DFF_X1 port map( D => n5004, CK => CLK
                           , Q => n_3787, QN => 
                           DataPath_RF_bus_reg_dataout_1292_port);
   DataPath_RF_BLOCKi_48_Q_reg_11_inst : DFF_X1 port map( D => n5005, CK => CLK
                           , Q => n_3788, QN => 
                           DataPath_RF_bus_reg_dataout_1291_port);
   DataPath_RF_BLOCKi_48_Q_reg_9_inst : DFF_X1 port map( D => n5007, CK => CLK,
                           Q => n_3789, QN => 
                           DataPath_RF_bus_reg_dataout_1289_port);
   DataPath_RF_BLOCKi_48_Q_reg_8_inst : DFF_X1 port map( D => n5008, CK => CLK,
                           Q => n_3790, QN => 
                           DataPath_RF_bus_reg_dataout_1288_port);
   DataPath_RF_BLOCKi_48_Q_reg_7_inst : DFF_X1 port map( D => n5009, CK => CLK,
                           Q => n_3791, QN => 
                           DataPath_RF_bus_reg_dataout_1287_port);
   DataPath_RF_BLOCKi_48_Q_reg_6_inst : DFF_X1 port map( D => n5010, CK => CLK,
                           Q => n_3792, QN => 
                           DataPath_RF_bus_reg_dataout_1286_port);
   DataPath_RF_BLOCKi_48_Q_reg_5_inst : DFF_X1 port map( D => n5011, CK => CLK,
                           Q => n_3793, QN => 
                           DataPath_RF_bus_reg_dataout_1285_port);
   DataPath_RF_BLOCKi_48_Q_reg_4_inst : DFF_X1 port map( D => n5012, CK => CLK,
                           Q => n_3794, QN => 
                           DataPath_RF_bus_reg_dataout_1284_port);
   DataPath_RF_BLOCKi_48_Q_reg_3_inst : DFF_X1 port map( D => n5013, CK => CLK,
                           Q => n_3795, QN => 
                           DataPath_RF_bus_reg_dataout_1283_port);
   DataPath_RF_BLOCKi_48_Q_reg_2_inst : DFF_X1 port map( D => n5014, CK => CLK,
                           Q => n_3796, QN => 
                           DataPath_RF_bus_reg_dataout_1282_port);
   DataPath_RF_BLOCKi_48_Q_reg_1_inst : DFF_X1 port map( D => n5015, CK => CLK,
                           Q => n_3797, QN => 
                           DataPath_RF_bus_reg_dataout_1281_port);
   DataPath_RF_BLOCKi_48_Q_reg_0_inst : DFF_X1 port map( D => n5016, CK => CLK,
                           Q => n_3798, QN => 
                           DataPath_RF_bus_reg_dataout_1280_port);
   DataPath_RF_BLOCKi_64_Q_reg_31_inst : DFF_X1 port map( D => n5576, CK => CLK
                           , Q => n_3799, QN => 
                           DataPath_RF_bus_reg_dataout_1823_port);
   DataPath_RF_BLOCKi_64_Q_reg_30_inst : DFF_X1 port map( D => n5579, CK => CLK
                           , Q => n_3800, QN => 
                           DataPath_RF_bus_reg_dataout_1822_port);
   DataPath_RF_BLOCKi_64_Q_reg_29_inst : DFF_X1 port map( D => n5580, CK => CLK
                           , Q => n_3801, QN => 
                           DataPath_RF_bus_reg_dataout_1821_port);
   DataPath_RF_BLOCKi_64_Q_reg_28_inst : DFF_X1 port map( D => n5581, CK => CLK
                           , Q => n_3802, QN => 
                           DataPath_RF_bus_reg_dataout_1820_port);
   DataPath_RF_BLOCKi_64_Q_reg_27_inst : DFF_X1 port map( D => n5582, CK => CLK
                           , Q => n_3803, QN => 
                           DataPath_RF_bus_reg_dataout_1819_port);
   DataPath_RF_BLOCKi_64_Q_reg_26_inst : DFF_X1 port map( D => n5583, CK => CLK
                           , Q => n_3804, QN => 
                           DataPath_RF_bus_reg_dataout_1818_port);
   DataPath_RF_BLOCKi_64_Q_reg_25_inst : DFF_X1 port map( D => n5584, CK => CLK
                           , Q => n_3805, QN => 
                           DataPath_RF_bus_reg_dataout_1817_port);
   DataPath_RF_BLOCKi_64_Q_reg_24_inst : DFF_X1 port map( D => n5585, CK => CLK
                           , Q => n_3806, QN => 
                           DataPath_RF_bus_reg_dataout_1816_port);
   DataPath_RF_BLOCKi_64_Q_reg_23_inst : DFF_X1 port map( D => n5586, CK => CLK
                           , Q => n_3807, QN => 
                           DataPath_RF_bus_reg_dataout_1815_port);
   DataPath_RF_BLOCKi_64_Q_reg_22_inst : DFF_X1 port map( D => n5587, CK => CLK
                           , Q => n_3808, QN => 
                           DataPath_RF_bus_reg_dataout_1814_port);
   DataPath_RF_BLOCKi_64_Q_reg_21_inst : DFF_X1 port map( D => n5588, CK => CLK
                           , Q => n_3809, QN => 
                           DataPath_RF_bus_reg_dataout_1813_port);
   DataPath_RF_BLOCKi_64_Q_reg_20_inst : DFF_X1 port map( D => n5589, CK => CLK
                           , Q => n_3810, QN => 
                           DataPath_RF_bus_reg_dataout_1812_port);
   DataPath_RF_BLOCKi_64_Q_reg_19_inst : DFF_X1 port map( D => n5590, CK => CLK
                           , Q => n_3811, QN => 
                           DataPath_RF_bus_reg_dataout_1811_port);
   DataPath_RF_BLOCKi_64_Q_reg_18_inst : DFF_X1 port map( D => n5591, CK => CLK
                           , Q => n_3812, QN => 
                           DataPath_RF_bus_reg_dataout_1810_port);
   DataPath_RF_BLOCKi_64_Q_reg_17_inst : DFF_X1 port map( D => n5592, CK => CLK
                           , Q => n_3813, QN => 
                           DataPath_RF_bus_reg_dataout_1809_port);
   DataPath_RF_BLOCKi_64_Q_reg_16_inst : DFF_X1 port map( D => n5593, CK => CLK
                           , Q => n_3814, QN => 
                           DataPath_RF_bus_reg_dataout_1808_port);
   DataPath_RF_BLOCKi_64_Q_reg_15_inst : DFF_X1 port map( D => n5594, CK => CLK
                           , Q => n_3815, QN => 
                           DataPath_RF_bus_reg_dataout_1807_port);
   DataPath_RF_BLOCKi_64_Q_reg_14_inst : DFF_X1 port map( D => n5595, CK => CLK
                           , Q => n_3816, QN => 
                           DataPath_RF_bus_reg_dataout_1806_port);
   DataPath_RF_BLOCKi_64_Q_reg_13_inst : DFF_X1 port map( D => n5596, CK => CLK
                           , Q => n_3817, QN => 
                           DataPath_RF_bus_reg_dataout_1805_port);
   DataPath_RF_BLOCKi_64_Q_reg_12_inst : DFF_X1 port map( D => n5597, CK => CLK
                           , Q => n_3818, QN => 
                           DataPath_RF_bus_reg_dataout_1804_port);
   DataPath_RF_BLOCKi_64_Q_reg_11_inst : DFF_X1 port map( D => n5598, CK => CLK
                           , Q => n_3819, QN => 
                           DataPath_RF_bus_reg_dataout_1803_port);
   DataPath_RF_BLOCKi_64_Q_reg_9_inst : DFF_X1 port map( D => n5600, CK => CLK,
                           Q => n_3820, QN => 
                           DataPath_RF_bus_reg_dataout_1801_port);
   DataPath_RF_BLOCKi_64_Q_reg_8_inst : DFF_X1 port map( D => n5601, CK => CLK,
                           Q => n_3821, QN => 
                           DataPath_RF_bus_reg_dataout_1800_port);
   DataPath_RF_BLOCKi_64_Q_reg_7_inst : DFF_X1 port map( D => n5602, CK => CLK,
                           Q => n_3822, QN => 
                           DataPath_RF_bus_reg_dataout_1799_port);
   DataPath_RF_BLOCKi_64_Q_reg_6_inst : DFF_X1 port map( D => n5603, CK => CLK,
                           Q => n_3823, QN => 
                           DataPath_RF_bus_reg_dataout_1798_port);
   DataPath_RF_BLOCKi_64_Q_reg_5_inst : DFF_X1 port map( D => n5604, CK => CLK,
                           Q => n_3824, QN => 
                           DataPath_RF_bus_reg_dataout_1797_port);
   DataPath_RF_BLOCKi_64_Q_reg_4_inst : DFF_X1 port map( D => n5605, CK => CLK,
                           Q => n_3825, QN => 
                           DataPath_RF_bus_reg_dataout_1796_port);
   DataPath_RF_BLOCKi_64_Q_reg_3_inst : DFF_X1 port map( D => n5606, CK => CLK,
                           Q => n_3826, QN => 
                           DataPath_RF_bus_reg_dataout_1795_port);
   DataPath_RF_BLOCKi_64_Q_reg_2_inst : DFF_X1 port map( D => n5607, CK => CLK,
                           Q => n_3827, QN => 
                           DataPath_RF_bus_reg_dataout_1794_port);
   DataPath_RF_BLOCKi_64_Q_reg_1_inst : DFF_X1 port map( D => n5608, CK => CLK,
                           Q => n_3828, QN => 
                           DataPath_RF_bus_reg_dataout_1793_port);
   DataPath_RF_BLOCKi_64_Q_reg_0_inst : DFF_X1 port map( D => n5609, CK => CLK,
                           Q => n_3829, QN => 
                           DataPath_RF_bus_reg_dataout_1792_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_31_inst : DFF_X1 port map( D => n6768, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_63_port,
                           QN => n627);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_30_inst : DFF_X1 port map( D => n6769, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_62_port,
                           QN => n626);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_29_inst : DFF_X1 port map( D => n6770, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_61_port,
                           QN => n625);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_28_inst : DFF_X1 port map( D => n6771, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_60_port,
                           QN => n624);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_27_inst : DFF_X1 port map( D => n6772, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_59_port,
                           QN => n623);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_26_inst : DFF_X1 port map( D => n6773, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_58_port,
                           QN => n622);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_25_inst : DFF_X1 port map( D => n6774, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_57_port,
                           QN => n621);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_24_inst : DFF_X1 port map( D => n6775, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_56_port,
                           QN => n620);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_23_inst : DFF_X1 port map( D => n6776, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_55_port,
                           QN => n619);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_22_inst : DFF_X1 port map( D => n6777, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_54_port,
                           QN => n618);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_21_inst : DFF_X1 port map( D => n6778, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_53_port,
                           QN => n617);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_20_inst : DFF_X1 port map( D => n6779, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_52_port,
                           QN => n616);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_19_inst : DFF_X1 port map( D => n6780, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_51_port,
                           QN => n615);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_18_inst : DFF_X1 port map( D => n6781, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_50_port,
                           QN => n614);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_17_inst : DFF_X1 port map( D => n6782, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_49_port,
                           QN => n613);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_16_inst : DFF_X1 port map( D => n6783, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_48_port,
                           QN => n612);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_15_inst : DFF_X1 port map( D => n6784, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_47_port,
                           QN => n611);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_14_inst : DFF_X1 port map( D => n6785, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_46_port,
                           QN => n610);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_13_inst : DFF_X1 port map( D => n6786, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_45_port,
                           QN => n609);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_12_inst : DFF_X1 port map( D => n6787, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_44_port,
                           QN => n608);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_11_inst : DFF_X1 port map( D => n6788, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_43_port,
                           QN => n607);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_10_inst : DFF_X1 port map( D => n6789, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_42_port,
                           QN => n606);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_9_inst : DFF_X1 port map( D => n6790, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_41_port,
                           QN => n605);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_8_inst : DFF_X1 port map( D => n6791, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_40_port,
                           QN => n604);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_7_inst : DFF_X1 port map( D => n6792, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_39_port,
                           QN => n603);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_6_inst : DFF_X1 port map( D => n6793, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_38_port,
                           QN => n602);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_5_inst : DFF_X1 port map( D => n6794, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_37_port,
                           QN => n601);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_4_inst : DFF_X1 port map( D => n6795, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_36_port,
                           QN => n600);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_3_inst : DFF_X1 port map( D => n6796, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_35_port,
                           QN => n599);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_2_inst : DFF_X1 port map( D => n6797, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_34_port,
                           QN => n598);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_1_inst : DFF_X1 port map( D => n6798, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_33_port,
                           QN => n597);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_0_inst : DFF_X1 port map( D => n6799, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_32_port,
                           QN => n596);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_31_inst : DFF_X1 port map( D => n6800, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_95_port,
                           QN => n659);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_30_inst : DFF_X1 port map( D => n6801, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_94_port,
                           QN => n658);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_29_inst : DFF_X1 port map( D => n6802, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_93_port,
                           QN => n657);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_28_inst : DFF_X1 port map( D => n6803, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_92_port,
                           QN => n656);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_27_inst : DFF_X1 port map( D => n6804, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_91_port,
                           QN => n655);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_26_inst : DFF_X1 port map( D => n6805, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_90_port,
                           QN => n654);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_25_inst : DFF_X1 port map( D => n6806, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_89_port,
                           QN => n653);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_24_inst : DFF_X1 port map( D => n6807, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_88_port,
                           QN => n652);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_23_inst : DFF_X1 port map( D => n6808, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_87_port,
                           QN => n651);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_22_inst : DFF_X1 port map( D => n6809, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_86_port,
                           QN => n650);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_21_inst : DFF_X1 port map( D => n6810, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_85_port,
                           QN => n649);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_20_inst : DFF_X1 port map( D => n6811, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_84_port,
                           QN => n648);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_19_inst : DFF_X1 port map( D => n6812, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_83_port,
                           QN => n647);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_18_inst : DFF_X1 port map( D => n6813, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_82_port,
                           QN => n646);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_17_inst : DFF_X1 port map( D => n6814, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_81_port,
                           QN => n645);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_16_inst : DFF_X1 port map( D => n6815, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_80_port,
                           QN => n644);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_15_inst : DFF_X1 port map( D => n6816, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_79_port,
                           QN => n643);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_14_inst : DFF_X1 port map( D => n6817, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_78_port,
                           QN => n642);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_13_inst : DFF_X1 port map( D => n6818, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_77_port,
                           QN => n641);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_12_inst : DFF_X1 port map( D => n6819, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_76_port,
                           QN => n640);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_11_inst : DFF_X1 port map( D => n6820, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_75_port,
                           QN => n639);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_10_inst : DFF_X1 port map( D => n6821, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_74_port,
                           QN => n638);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_9_inst : DFF_X1 port map( D => n6822, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_73_port,
                           QN => n637);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_8_inst : DFF_X1 port map( D => n6823, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_72_port,
                           QN => n636);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_7_inst : DFF_X1 port map( D => n6824, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_71_port,
                           QN => n635);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_6_inst : DFF_X1 port map( D => n6825, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_70_port,
                           QN => n634);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_5_inst : DFF_X1 port map( D => n6826, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_69_port,
                           QN => n633);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_4_inst : DFF_X1 port map( D => n6827, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_68_port,
                           QN => n632);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_3_inst : DFF_X1 port map( D => n6828, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_67_port,
                           QN => n631);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_2_inst : DFF_X1 port map( D => n6829, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_66_port,
                           QN => n630);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_1_inst : DFF_X1 port map( D => n6830, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_65_port,
                           QN => n629);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_0_inst : DFF_X1 port map( D => n6831, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_64_port,
                           QN => n628);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_31_inst : DFF_X1 port map( D => n6832, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_127_port
                           , QN => n691);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_30_inst : DFF_X1 port map( D => n6833, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_126_port
                           , QN => n690);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_29_inst : DFF_X1 port map( D => n6834, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_125_port
                           , QN => n689);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_28_inst : DFF_X1 port map( D => n6835, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_124_port
                           , QN => n688);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_27_inst : DFF_X1 port map( D => n6836, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_123_port
                           , QN => n687);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_26_inst : DFF_X1 port map( D => n6837, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_122_port
                           , QN => n686);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_25_inst : DFF_X1 port map( D => n6838, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_121_port
                           , QN => n685);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_24_inst : DFF_X1 port map( D => n6839, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_120_port
                           , QN => n684);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_23_inst : DFF_X1 port map( D => n6840, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_119_port
                           , QN => n683);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_22_inst : DFF_X1 port map( D => n6841, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_118_port
                           , QN => n682);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_21_inst : DFF_X1 port map( D => n6842, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_117_port
                           , QN => n681);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_20_inst : DFF_X1 port map( D => n6843, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_116_port
                           , QN => n680);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_19_inst : DFF_X1 port map( D => n6844, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_115_port
                           , QN => n679);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_18_inst : DFF_X1 port map( D => n6845, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_114_port
                           , QN => n678);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_17_inst : DFF_X1 port map( D => n6846, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_113_port
                           , QN => n677);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_16_inst : DFF_X1 port map( D => n6847, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_112_port
                           , QN => n676);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_15_inst : DFF_X1 port map( D => n6848, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_111_port
                           , QN => n675);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_14_inst : DFF_X1 port map( D => n6849, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_110_port
                           , QN => n674);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_13_inst : DFF_X1 port map( D => n6850, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_109_port
                           , QN => n673);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_12_inst : DFF_X1 port map( D => n6851, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_108_port
                           , QN => n672);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_11_inst : DFF_X1 port map( D => n6852, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_107_port
                           , QN => n671);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_10_inst : DFF_X1 port map( D => n6853, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_106_port
                           , QN => n670);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_9_inst : DFF_X1 port map( D => n6854, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_105_port
                           , QN => n669);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_8_inst : DFF_X1 port map( D => n6855, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_104_port
                           , QN => n668);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_7_inst : DFF_X1 port map( D => n6856, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_103_port
                           , QN => n667);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_6_inst : DFF_X1 port map( D => n6857, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_102_port
                           , QN => n666);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_5_inst : DFF_X1 port map( D => n6858, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_101_port
                           , QN => n665);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_4_inst : DFF_X1 port map( D => n6859, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_100_port
                           , QN => n664);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_3_inst : DFF_X1 port map( D => n6860, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_99_port,
                           QN => n663);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_2_inst : DFF_X1 port map( D => n6861, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_98_port,
                           QN => n662);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_1_inst : DFF_X1 port map( D => n6862, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_97_port,
                           QN => n661);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_0_inst : DFF_X1 port map( D => n6863, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_96_port,
                           QN => n660);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_31_inst : DFF_X1 port map( D => n6864, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_159_port
                           , QN => n723);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_30_inst : DFF_X1 port map( D => n6865, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_158_port
                           , QN => n722);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_29_inst : DFF_X1 port map( D => n6866, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_157_port
                           , QN => n721);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_28_inst : DFF_X1 port map( D => n6867, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_156_port
                           , QN => n720);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_27_inst : DFF_X1 port map( D => n6868, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_155_port
                           , QN => n719);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_26_inst : DFF_X1 port map( D => n6869, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_154_port
                           , QN => n718);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_25_inst : DFF_X1 port map( D => n6870, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_153_port
                           , QN => n717);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_24_inst : DFF_X1 port map( D => n6871, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_152_port
                           , QN => n716);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_23_inst : DFF_X1 port map( D => n6872, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_151_port
                           , QN => n715);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_22_inst : DFF_X1 port map( D => n6873, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_150_port
                           , QN => n714);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_21_inst : DFF_X1 port map( D => n6874, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_149_port
                           , QN => n713);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_20_inst : DFF_X1 port map( D => n6875, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_148_port
                           , QN => n712);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_19_inst : DFF_X1 port map( D => n6876, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_147_port
                           , QN => n711);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_18_inst : DFF_X1 port map( D => n6877, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_146_port
                           , QN => n710);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_17_inst : DFF_X1 port map( D => n6878, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_145_port
                           , QN => n709);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_16_inst : DFF_X1 port map( D => n6879, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_144_port
                           , QN => n708);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_15_inst : DFF_X1 port map( D => n6880, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_143_port
                           , QN => n707);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_14_inst : DFF_X1 port map( D => n6881, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_142_port
                           , QN => n706);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_13_inst : DFF_X1 port map( D => n6882, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_141_port
                           , QN => n705);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_12_inst : DFF_X1 port map( D => n6883, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_140_port
                           , QN => n704);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_11_inst : DFF_X1 port map( D => n6884, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_139_port
                           , QN => n703);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_10_inst : DFF_X1 port map( D => n6885, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_138_port
                           , QN => n702);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_9_inst : DFF_X1 port map( D => n6886, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_137_port
                           , QN => n701);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_8_inst : DFF_X1 port map( D => n6887, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_136_port
                           , QN => n700);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_7_inst : DFF_X1 port map( D => n6888, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_135_port
                           , QN => n699);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_6_inst : DFF_X1 port map( D => n6889, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_134_port
                           , QN => n698);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_5_inst : DFF_X1 port map( D => n6890, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_133_port
                           , QN => n697);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_4_inst : DFF_X1 port map( D => n6891, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_132_port
                           , QN => n696);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_3_inst : DFF_X1 port map( D => n6892, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_131_port
                           , QN => n695);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_2_inst : DFF_X1 port map( D => n6893, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_130_port
                           , QN => n694);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_1_inst : DFF_X1 port map( D => n6894, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_129_port
                           , QN => n693);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_0_inst : DFF_X1 port map( D => n6895, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_128_port
                           , QN => n692);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_31_inst : DFF_X1 port map( D => n6896, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_191_port
                           , QN => n755);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_30_inst : DFF_X1 port map( D => n6897, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_190_port
                           , QN => n754);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_29_inst : DFF_X1 port map( D => n6898, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_189_port
                           , QN => n753);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_28_inst : DFF_X1 port map( D => n6899, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_188_port
                           , QN => n752);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_27_inst : DFF_X1 port map( D => n6900, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_187_port
                           , QN => n751);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_26_inst : DFF_X1 port map( D => n6901, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_186_port
                           , QN => n750);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_25_inst : DFF_X1 port map( D => n6902, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_185_port
                           , QN => n749);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_24_inst : DFF_X1 port map( D => n6903, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_184_port
                           , QN => n748);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_23_inst : DFF_X1 port map( D => n6904, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_183_port
                           , QN => n747);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_22_inst : DFF_X1 port map( D => n6905, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_182_port
                           , QN => n746);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_21_inst : DFF_X1 port map( D => n6906, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_181_port
                           , QN => n745);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_20_inst : DFF_X1 port map( D => n6907, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_180_port
                           , QN => n744);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_19_inst : DFF_X1 port map( D => n6908, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_179_port
                           , QN => n743);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_18_inst : DFF_X1 port map( D => n6909, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_178_port
                           , QN => n742);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_17_inst : DFF_X1 port map( D => n6910, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_177_port
                           , QN => n741);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_16_inst : DFF_X1 port map( D => n6911, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_176_port
                           , QN => n740);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_15_inst : DFF_X1 port map( D => n6912, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_175_port
                           , QN => n739);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_14_inst : DFF_X1 port map( D => n6913, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_174_port
                           , QN => n738);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_13_inst : DFF_X1 port map( D => n6914, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_173_port
                           , QN => n737);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_12_inst : DFF_X1 port map( D => n6915, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_172_port
                           , QN => n736);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_11_inst : DFF_X1 port map( D => n6916, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_171_port
                           , QN => n735);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_10_inst : DFF_X1 port map( D => n6917, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_170_port
                           , QN => n734);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_9_inst : DFF_X1 port map( D => n6918, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_169_port
                           , QN => n733);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_8_inst : DFF_X1 port map( D => n6919, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_168_port
                           , QN => n732);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_7_inst : DFF_X1 port map( D => n6920, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_167_port
                           , QN => n731);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_6_inst : DFF_X1 port map( D => n6921, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_166_port
                           , QN => n730);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_5_inst : DFF_X1 port map( D => n6922, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_165_port
                           , QN => n729);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_4_inst : DFF_X1 port map( D => n6923, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_164_port
                           , QN => n728);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_3_inst : DFF_X1 port map( D => n6924, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_163_port
                           , QN => n727);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_2_inst : DFF_X1 port map( D => n6925, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_162_port
                           , QN => n726);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_1_inst : DFF_X1 port map( D => n6926, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_161_port
                           , QN => n725);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_0_inst : DFF_X1 port map( D => n6927, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_160_port
                           , QN => n724);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_31_inst : DFF_X1 port map( D => n6928, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_223_port
                           , QN => n787);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_30_inst : DFF_X1 port map( D => n6929, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_222_port
                           , QN => n786);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_29_inst : DFF_X1 port map( D => n6930, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_221_port
                           , QN => n785);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_28_inst : DFF_X1 port map( D => n6931, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_220_port
                           , QN => n784);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_27_inst : DFF_X1 port map( D => n6932, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_219_port
                           , QN => n783);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_26_inst : DFF_X1 port map( D => n6933, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_218_port
                           , QN => n782);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_25_inst : DFF_X1 port map( D => n6934, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_217_port
                           , QN => n781);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_24_inst : DFF_X1 port map( D => n6935, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_216_port
                           , QN => n780);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_23_inst : DFF_X1 port map( D => n6936, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_215_port
                           , QN => n779);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_22_inst : DFF_X1 port map( D => n6937, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_214_port
                           , QN => n778);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_21_inst : DFF_X1 port map( D => n6938, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_213_port
                           , QN => n777);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_20_inst : DFF_X1 port map( D => n6939, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_212_port
                           , QN => n776);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_19_inst : DFF_X1 port map( D => n6940, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_211_port
                           , QN => n775);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_18_inst : DFF_X1 port map( D => n6941, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_210_port
                           , QN => n774);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_17_inst : DFF_X1 port map( D => n6942, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_209_port
                           , QN => n773);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_16_inst : DFF_X1 port map( D => n6943, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_208_port
                           , QN => n772);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_15_inst : DFF_X1 port map( D => n6944, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_207_port
                           , QN => n771);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_14_inst : DFF_X1 port map( D => n6945, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_206_port
                           , QN => n770);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_13_inst : DFF_X1 port map( D => n6946, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_205_port
                           , QN => n769);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_12_inst : DFF_X1 port map( D => n6947, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_204_port
                           , QN => n768);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_11_inst : DFF_X1 port map( D => n6948, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_203_port
                           , QN => n767);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_10_inst : DFF_X1 port map( D => n6949, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_202_port
                           , QN => n766);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_9_inst : DFF_X1 port map( D => n6950, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_201_port
                           , QN => n765);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_8_inst : DFF_X1 port map( D => n6951, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_200_port
                           , QN => n764);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_7_inst : DFF_X1 port map( D => n6952, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_199_port
                           , QN => n763);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_6_inst : DFF_X1 port map( D => n6953, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_198_port
                           , QN => n762);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_5_inst : DFF_X1 port map( D => n6954, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_197_port
                           , QN => n761);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_4_inst : DFF_X1 port map( D => n6955, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_196_port
                           , QN => n760);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_3_inst : DFF_X1 port map( D => n6956, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_195_port
                           , QN => n759);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_2_inst : DFF_X1 port map( D => n6957, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_194_port
                           , QN => n758);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_1_inst : DFF_X1 port map( D => n6958, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_193_port
                           , QN => n757);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_0_inst : DFF_X1 port map( D => n6959, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_192_port
                           , QN => n756);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_31_inst : DFF_X1 port map( D => n6960, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_255_port
                           , QN => n819);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_30_inst : DFF_X1 port map( D => n6961, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_254_port
                           , QN => n818);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_29_inst : DFF_X1 port map( D => n6962, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_253_port
                           , QN => n817);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_28_inst : DFF_X1 port map( D => n6963, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_252_port
                           , QN => n816);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_27_inst : DFF_X1 port map( D => n6964, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_251_port
                           , QN => n815);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_26_inst : DFF_X1 port map( D => n6965, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_250_port
                           , QN => n814);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_25_inst : DFF_X1 port map( D => n6966, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_249_port
                           , QN => n813);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_24_inst : DFF_X1 port map( D => n6967, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_248_port
                           , QN => n812);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_23_inst : DFF_X1 port map( D => n6968, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_247_port
                           , QN => n811);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_22_inst : DFF_X1 port map( D => n6969, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_246_port
                           , QN => n810);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_21_inst : DFF_X1 port map( D => n6970, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_245_port
                           , QN => n809);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_20_inst : DFF_X1 port map( D => n6971, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_244_port
                           , QN => n808);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_19_inst : DFF_X1 port map( D => n6972, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_243_port
                           , QN => n807);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_18_inst : DFF_X1 port map( D => n6973, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_242_port
                           , QN => n806);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_17_inst : DFF_X1 port map( D => n6974, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_241_port
                           , QN => n805);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_16_inst : DFF_X1 port map( D => n6975, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_240_port
                           , QN => n804);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_15_inst : DFF_X1 port map( D => n6976, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_239_port
                           , QN => n803);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_14_inst : DFF_X1 port map( D => n6977, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_238_port
                           , QN => n802);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_13_inst : DFF_X1 port map( D => n6978, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_237_port
                           , QN => n801);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_12_inst : DFF_X1 port map( D => n6979, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_236_port
                           , QN => n800);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_11_inst : DFF_X1 port map( D => n6980, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_235_port
                           , QN => n799);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_9_inst : DFF_X1 port map( D => n6982, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_233_port
                           , QN => n797);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_8_inst : DFF_X1 port map( D => n6983, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_232_port
                           , QN => n796);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_7_inst : DFF_X1 port map( D => n6984, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_231_port
                           , QN => n795);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_6_inst : DFF_X1 port map( D => n6985, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_230_port
                           , QN => n794);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_5_inst : DFF_X1 port map( D => n6986, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_229_port
                           , QN => n793);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_4_inst : DFF_X1 port map( D => n6987, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_228_port
                           , QN => n792);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_3_inst : DFF_X1 port map( D => n6988, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_227_port
                           , QN => n791);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_2_inst : DFF_X1 port map( D => n6989, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_226_port
                           , QN => n790);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_1_inst : DFF_X1 port map( D => n6990, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_225_port
                           , QN => n789);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_0_inst : DFF_X1 port map( D => n6991, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_224_port
                           , QN => n788);
   DataPath_RF_BLOCKi_8_Q_reg_10_inst : DFF_X1 port map( D => n3472, CK => CLK,
                           Q => n_3830, QN => 
                           DataPath_RF_bus_reg_dataout_10_port);
   DataPath_RF_BLOCKi_9_Q_reg_10_inst : DFF_X1 port map( D => n3522, CK => CLK,
                           Q => n_3831, QN => 
                           DataPath_RF_bus_reg_dataout_42_port);
   DataPath_RF_BLOCKi_10_Q_reg_10_inst : DFF_X1 port map( D => n3560, CK => CLK
                           , Q => n_3832, QN => 
                           DataPath_RF_bus_reg_dataout_74_port);
   DataPath_RF_BLOCKi_11_Q_reg_10_inst : DFF_X1 port map( D => n3598, CK => CLK
                           , Q => n_3833, QN => 
                           DataPath_RF_bus_reg_dataout_106_port);
   DataPath_RF_BLOCKi_12_Q_reg_10_inst : DFF_X1 port map( D => n3636, CK => CLK
                           , Q => n_3834, QN => 
                           DataPath_RF_bus_reg_dataout_138_port);
   DataPath_RF_BLOCKi_13_Q_reg_10_inst : DFF_X1 port map( D => n3674, CK => CLK
                           , Q => n_3835, QN => 
                           DataPath_RF_bus_reg_dataout_170_port);
   DataPath_RF_BLOCKi_14_Q_reg_10_inst : DFF_X1 port map( D => n3712, CK => CLK
                           , Q => n_3836, QN => 
                           DataPath_RF_bus_reg_dataout_202_port);
   DataPath_RF_BLOCKi_15_Q_reg_10_inst : DFF_X1 port map( D => n3750, CK => CLK
                           , Q => n_3837, QN => 
                           DataPath_RF_bus_reg_dataout_234_port);
   DataPath_RF_BLOCKi_16_Q_reg_10_inst : DFF_X1 port map( D => n3788, CK => CLK
                           , Q => n_3838, QN => 
                           DataPath_RF_bus_reg_dataout_266_port);
   DataPath_RF_BLOCKi_17_Q_reg_10_inst : DFF_X1 port map( D => n3823, CK => CLK
                           , Q => n_3839, QN => 
                           DataPath_RF_bus_reg_dataout_298_port);
   DataPath_RF_BLOCKi_18_Q_reg_10_inst : DFF_X1 port map( D => n3858, CK => CLK
                           , Q => n_3840, QN => 
                           DataPath_RF_bus_reg_dataout_330_port);
   DataPath_RF_BLOCKi_19_Q_reg_10_inst : DFF_X1 port map( D => n3893, CK => CLK
                           , Q => n_3841, QN => 
                           DataPath_RF_bus_reg_dataout_362_port);
   DataPath_RF_BLOCKi_20_Q_reg_10_inst : DFF_X1 port map( D => n3928, CK => CLK
                           , Q => n_3842, QN => 
                           DataPath_RF_bus_reg_dataout_394_port);
   DataPath_RF_BLOCKi_21_Q_reg_10_inst : DFF_X1 port map( D => n3963, CK => CLK
                           , Q => n_3843, QN => 
                           DataPath_RF_bus_reg_dataout_426_port);
   DataPath_RF_BLOCKi_22_Q_reg_10_inst : DFF_X1 port map( D => n3998, CK => CLK
                           , Q => n_3844, QN => 
                           DataPath_RF_bus_reg_dataout_458_port);
   DataPath_RF_BLOCKi_23_Q_reg_10_inst : DFF_X1 port map( D => n4054, CK => CLK
                           , Q => n_3845, QN => 
                           DataPath_RF_bus_reg_dataout_490_port);
   DataPath_RF_BLOCKi_24_Q_reg_10_inst : DFF_X1 port map( D => n4121, CK => CLK
                           , Q => n_3846, QN => 
                           DataPath_RF_bus_reg_dataout_522_port);
   DataPath_RF_BLOCKi_25_Q_reg_10_inst : DFF_X1 port map( D => n4168, CK => CLK
                           , Q => n_3847, QN => 
                           DataPath_RF_bus_reg_dataout_554_port);
   DataPath_RF_BLOCKi_26_Q_reg_10_inst : DFF_X1 port map( D => n4203, CK => CLK
                           , Q => n_3848, QN => 
                           DataPath_RF_bus_reg_dataout_586_port);
   DataPath_RF_BLOCKi_27_Q_reg_10_inst : DFF_X1 port map( D => n4238, CK => CLK
                           , Q => n_3849, QN => 
                           DataPath_RF_bus_reg_dataout_618_port);
   DataPath_RF_BLOCKi_28_Q_reg_10_inst : DFF_X1 port map( D => n4273, CK => CLK
                           , Q => n_3850, QN => 
                           DataPath_RF_bus_reg_dataout_650_port);
   DataPath_RF_BLOCKi_29_Q_reg_10_inst : DFF_X1 port map( D => n4308, CK => CLK
                           , Q => n_3851, QN => 
                           DataPath_RF_bus_reg_dataout_682_port);
   DataPath_RF_BLOCKi_30_Q_reg_10_inst : DFF_X1 port map( D => n4343, CK => CLK
                           , Q => n_3852, QN => 
                           DataPath_RF_bus_reg_dataout_714_port);
   DataPath_RF_BLOCKi_31_Q_reg_10_inst : DFF_X1 port map( D => n4378, CK => CLK
                           , Q => n_3853, QN => 
                           DataPath_RF_bus_reg_dataout_746_port);
   DataPath_RF_BLOCKi_32_Q_reg_10_inst : DFF_X1 port map( D => n4413, CK => CLK
                           , Q => n_3854, QN => 
                           DataPath_RF_bus_reg_dataout_778_port);
   DataPath_RF_BLOCKi_33_Q_reg_10_inst : DFF_X1 port map( D => n4448, CK => CLK
                           , Q => n_3855, QN => 
                           DataPath_RF_bus_reg_dataout_810_port);
   DataPath_RF_BLOCKi_34_Q_reg_10_inst : DFF_X1 port map( D => n4483, CK => CLK
                           , Q => n_3856, QN => 
                           DataPath_RF_bus_reg_dataout_842_port);
   DataPath_RF_BLOCKi_35_Q_reg_10_inst : DFF_X1 port map( D => n4518, CK => CLK
                           , Q => n_3857, QN => 
                           DataPath_RF_bus_reg_dataout_874_port);
   DataPath_RF_BLOCKi_36_Q_reg_10_inst : DFF_X1 port map( D => n4553, CK => CLK
                           , Q => n_3858, QN => 
                           DataPath_RF_bus_reg_dataout_906_port);
   DataPath_RF_BLOCKi_37_Q_reg_10_inst : DFF_X1 port map( D => n4588, CK => CLK
                           , Q => n_3859, QN => 
                           DataPath_RF_bus_reg_dataout_938_port);
   DataPath_RF_BLOCKi_38_Q_reg_10_inst : DFF_X1 port map( D => n4623, CK => CLK
                           , Q => n_3860, QN => 
                           DataPath_RF_bus_reg_dataout_970_port);
   DataPath_RF_BLOCKi_39_Q_reg_10_inst : DFF_X1 port map( D => n4658, CK => CLK
                           , Q => n_3861, QN => 
                           DataPath_RF_bus_reg_dataout_1002_port);
   DataPath_RF_BLOCKi_40_Q_reg_10_inst : DFF_X1 port map( D => n4714, CK => CLK
                           , Q => n_3862, QN => 
                           DataPath_RF_bus_reg_dataout_1034_port);
   DataPath_RF_BLOCKi_41_Q_reg_10_inst : DFF_X1 port map( D => n4761, CK => CLK
                           , Q => n_3863, QN => 
                           DataPath_RF_bus_reg_dataout_1066_port);
   DataPath_RF_BLOCKi_42_Q_reg_10_inst : DFF_X1 port map( D => n4796, CK => CLK
                           , Q => n_3864, QN => 
                           DataPath_RF_bus_reg_dataout_1098_port);
   DataPath_RF_BLOCKi_43_Q_reg_10_inst : DFF_X1 port map( D => n4831, CK => CLK
                           , Q => n_3865, QN => 
                           DataPath_RF_bus_reg_dataout_1130_port);
   DataPath_RF_BLOCKi_44_Q_reg_10_inst : DFF_X1 port map( D => n4866, CK => CLK
                           , Q => n_3866, QN => 
                           DataPath_RF_bus_reg_dataout_1162_port);
   DataPath_RF_BLOCKi_45_Q_reg_10_inst : DFF_X1 port map( D => n4901, CK => CLK
                           , Q => n_3867, QN => 
                           DataPath_RF_bus_reg_dataout_1194_port);
   DataPath_RF_BLOCKi_46_Q_reg_10_inst : DFF_X1 port map( D => n4936, CK => CLK
                           , Q => n_3868, QN => 
                           DataPath_RF_bus_reg_dataout_1226_port);
   DataPath_RF_BLOCKi_47_Q_reg_10_inst : DFF_X1 port map( D => n4971, CK => CLK
                           , Q => n_3869, QN => 
                           DataPath_RF_bus_reg_dataout_1258_port);
   DataPath_RF_BLOCKi_48_Q_reg_10_inst : DFF_X1 port map( D => n5006, CK => CLK
                           , Q => n_3870, QN => 
                           DataPath_RF_bus_reg_dataout_1290_port);
   DataPath_RF_BLOCKi_49_Q_reg_10_inst : DFF_X1 port map( D => n5041, CK => CLK
                           , Q => n_3871, QN => 
                           DataPath_RF_bus_reg_dataout_1322_port);
   DataPath_RF_BLOCKi_50_Q_reg_10_inst : DFF_X1 port map( D => n5076, CK => CLK
                           , Q => n_3872, QN => 
                           DataPath_RF_bus_reg_dataout_1354_port);
   DataPath_RF_BLOCKi_51_Q_reg_10_inst : DFF_X1 port map( D => n5111, CK => CLK
                           , Q => n_3873, QN => 
                           DataPath_RF_bus_reg_dataout_1386_port);
   DataPath_RF_BLOCKi_52_Q_reg_10_inst : DFF_X1 port map( D => n5146, CK => CLK
                           , Q => n_3874, QN => 
                           DataPath_RF_bus_reg_dataout_1418_port);
   DataPath_RF_BLOCKi_53_Q_reg_10_inst : DFF_X1 port map( D => n5181, CK => CLK
                           , Q => n_3875, QN => 
                           DataPath_RF_bus_reg_dataout_1450_port);
   DataPath_RF_BLOCKi_54_Q_reg_10_inst : DFF_X1 port map( D => n5216, CK => CLK
                           , Q => n_3876, QN => 
                           DataPath_RF_bus_reg_dataout_1482_port);
   DataPath_RF_BLOCKi_55_Q_reg_10_inst : DFF_X1 port map( D => n5251, CK => CLK
                           , Q => n_3877, QN => 
                           DataPath_RF_bus_reg_dataout_1514_port);
   DataPath_RF_BLOCKi_56_Q_reg_10_inst : DFF_X1 port map( D => n5307, CK => CLK
                           , Q => n_3878, QN => 
                           DataPath_RF_bus_reg_dataout_1546_port);
   DataPath_RF_BLOCKi_57_Q_reg_10_inst : DFF_X1 port map( D => n5354, CK => CLK
                           , Q => n_3879, QN => 
                           DataPath_RF_bus_reg_dataout_1578_port);
   DataPath_RF_BLOCKi_58_Q_reg_10_inst : DFF_X1 port map( D => n5389, CK => CLK
                           , Q => n_3880, QN => 
                           DataPath_RF_bus_reg_dataout_1610_port);
   DataPath_RF_BLOCKi_59_Q_reg_10_inst : DFF_X1 port map( D => n5424, CK => CLK
                           , Q => n_3881, QN => 
                           DataPath_RF_bus_reg_dataout_1642_port);
   DataPath_RF_BLOCKi_60_Q_reg_10_inst : DFF_X1 port map( D => n5459, CK => CLK
                           , Q => n_3882, QN => 
                           DataPath_RF_bus_reg_dataout_1674_port);
   DataPath_RF_BLOCKi_61_Q_reg_10_inst : DFF_X1 port map( D => n5494, CK => CLK
                           , Q => n_3883, QN => 
                           DataPath_RF_bus_reg_dataout_1706_port);
   DataPath_RF_BLOCKi_62_Q_reg_10_inst : DFF_X1 port map( D => n5529, CK => CLK
                           , Q => n_3884, QN => 
                           DataPath_RF_bus_reg_dataout_1738_port);
   DataPath_RF_BLOCKi_63_Q_reg_10_inst : DFF_X1 port map( D => n5564, CK => CLK
                           , Q => n_3885, QN => 
                           DataPath_RF_bus_reg_dataout_1770_port);
   DataPath_RF_BLOCKi_64_Q_reg_10_inst : DFF_X1 port map( D => n5599, CK => CLK
                           , Q => n_3886, QN => 
                           DataPath_RF_bus_reg_dataout_1802_port);
   DataPath_RF_BLOCKi_65_Q_reg_10_inst : DFF_X1 port map( D => n5638, CK => CLK
                           , Q => n_3887, QN => 
                           DataPath_RF_bus_reg_dataout_1834_port);
   DataPath_RF_BLOCKi_66_Q_reg_10_inst : DFF_X1 port map( D => n5674, CK => CLK
                           , Q => n_3888, QN => 
                           DataPath_RF_bus_reg_dataout_1866_port);
   DataPath_RF_BLOCKi_67_Q_reg_10_inst : DFF_X1 port map( D => n5710, CK => CLK
                           , Q => n_3889, QN => 
                           DataPath_RF_bus_reg_dataout_1898_port);
   DataPath_RF_BLOCKi_68_Q_reg_10_inst : DFF_X1 port map( D => n5746, CK => CLK
                           , Q => n_3890, QN => 
                           DataPath_RF_bus_reg_dataout_1930_port);
   DataPath_RF_BLOCKi_69_Q_reg_10_inst : DFF_X1 port map( D => n5782, CK => CLK
                           , Q => n_3891, QN => 
                           DataPath_RF_bus_reg_dataout_1962_port);
   DataPath_RF_BLOCKi_70_Q_reg_10_inst : DFF_X1 port map( D => n5818, CK => CLK
                           , Q => n_3892, QN => 
                           DataPath_RF_bus_reg_dataout_1994_port);
   DataPath_RF_BLOCKi_71_Q_reg_10_inst : DFF_X1 port map( D => n5854, CK => CLK
                           , Q => n_3893, QN => 
                           DataPath_RF_bus_reg_dataout_2026_port);
   DataPath_RF_BLOCKi_79_Q_reg_10_inst : DFF_X1 port map( D => n891, CK => CLK,
                           Q => n_3894, QN => 
                           DataPath_RF_bus_reg_dataout_2282_port);
   DataPath_RF_BLOCKi_80_Q_reg_10_inst : DFF_X1 port map( D => n952, CK => CLK,
                           Q => n_3895, QN => 
                           DataPath_RF_bus_reg_dataout_2314_port);
   DataPath_RF_BLOCKi_81_Q_reg_10_inst : DFF_X1 port map( D => n989, CK => CLK,
                           Q => n_3896, QN => 
                           DataPath_RF_bus_reg_dataout_2346_port);
   DataPath_RF_BLOCKi_82_Q_reg_10_inst : DFF_X1 port map( D => n1026, CK => CLK
                           , Q => n_3897, QN => 
                           DataPath_RF_bus_reg_dataout_2378_port);
   DataPath_RF_BLOCKi_83_Q_reg_10_inst : DFF_X1 port map( D => n1063, CK => CLK
                           , Q => n_3898, QN => 
                           DataPath_RF_bus_reg_dataout_2410_port);
   DataPath_RF_BLOCKi_84_Q_reg_10_inst : DFF_X1 port map( D => n1100, CK => CLK
                           , Q => n_3899, QN => 
                           DataPath_RF_bus_reg_dataout_2442_port);
   DataPath_RF_BLOCKi_85_Q_reg_10_inst : DFF_X1 port map( D => n1137, CK => CLK
                           , Q => n_3900, QN => 
                           DataPath_RF_bus_reg_dataout_2474_port);
   DataPath_RF_BLOCKi_86_Q_reg_10_inst : DFF_X1 port map( D => n1174, CK => CLK
                           , Q => n_3901, QN => 
                           DataPath_RF_bus_reg_dataout_2506_port);
   DataPath_RF_BLOCKi_87_Q_reg_10_inst : DFF_X1 port map( D => n1211, CK => CLK
                           , Q => n_3902, QN => 
                           DataPath_RF_bus_reg_dataout_2538_port);
   DataPath_RF_BLOCKi_72_Q_reg_10_inst : DFF_X1 port map( D => n5890, CK => CLK
                           , Q => n_3903, QN => 
                           DataPath_RF_bus_reg_dataout_2058_port);
   DataPath_RF_BLOCKi_73_Q_reg_10_inst : DFF_X1 port map( D => n5928, CK => CLK
                           , Q => n_3904, QN => 
                           DataPath_RF_bus_reg_dataout_2090_port);
   DataPath_RF_BLOCKi_74_Q_reg_10_inst : DFF_X1 port map( D => n5965, CK => CLK
                           , Q => n_3905, QN => 
                           DataPath_RF_bus_reg_dataout_2122_port);
   DataPath_RF_BLOCKi_75_Q_reg_10_inst : DFF_X1 port map( D => n6002, CK => CLK
                           , Q => n_3906, QN => 
                           DataPath_RF_bus_reg_dataout_2154_port);
   DataPath_RF_BLOCKi_76_Q_reg_10_inst : DFF_X1 port map( D => n6039, CK => CLK
                           , Q => n_3907, QN => 
                           DataPath_RF_bus_reg_dataout_2186_port);
   DataPath_RF_BLOCKi_77_Q_reg_10_inst : DFF_X1 port map( D => n6076, CK => CLK
                           , Q => n_3908, QN => 
                           DataPath_RF_bus_reg_dataout_2218_port);
   DataPath_RF_BLOCKi_78_Q_reg_10_inst : DFF_X1 port map( D => n6113, CK => CLK
                           , Q => n_3909, QN => 
                           DataPath_RF_bus_reg_dataout_2250_port);
   IR_reg_28_inst : DFFS_X1 port map( D => n7107, CK => CLK, SN => n8693, Q => 
                           n8503, QN => n181);
   PC_reg_30_inst : DFFS_X1 port map( D => n8477, CK => CLK, SN => n8696, Q => 
                           n8393, QN => IRAM_ADDRESS_30_port);
   PC_reg_31_inst : DFFS_X1 port map( D => n8476, CK => CLK, SN => n8696, Q => 
                           n8430, QN => IRAM_ADDRESS_31_port);
   CU_I_aluOpcode1_reg_4_inst : DFF_X1 port map( D => n7083, CK => CLK, Q => 
                           n8385, QN => n368);
   DataPath_RF_CWP_Q_reg_0_inst : DFF_X2 port map( D => n7073, CK => CLK, Q => 
                           DataPath_RF_c_win_0_port, QN => n8299);
   DataPath_REG_ALU_OUT_Q_reg_31_inst : DFF_X1 port map( D => n6992, CK => CLK,
                           Q => DRAM_ADDRESS_31_port, QN => n516);
   DataPath_WRF_CUhw_curr_addr_reg_29_inst : DFF_X1 port map( D => n8482, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_29_port, QN =>
                           n_3910);
   DataPath_WRF_CUhw_curr_addr_reg_30_inst : DFF_X1 port map( D => n8481, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_30_port, QN =>
                           n_3911);
   DP_OP_1090J1_126_7243_U28 : FA_X1 port map( A => DP_OP_1090J1_126_7243_n72, 
                           B => DataPath_WRF_CUhw_curr_addr_5_port, CI => 
                           DP_OP_1090J1_126_7243_n28, CO => 
                           DP_OP_1090J1_126_7243_n27, S => C620_DATA2_5);
   DP_OP_1090J1_126_7243_U27 : FA_X1 port map( A => DP_OP_1090J1_126_7243_n72, 
                           B => DataPath_WRF_CUhw_curr_addr_6_port, CI => 
                           DP_OP_1090J1_126_7243_n27, CO => 
                           DP_OP_1090J1_126_7243_n26, S => C620_DATA2_6);
   DP_OP_1090J1_126_7243_U26 : FA_X1 port map( A => DP_OP_1090J1_126_7243_n72, 
                           B => DataPath_WRF_CUhw_curr_addr_7_port, CI => 
                           DP_OP_1090J1_126_7243_n26, CO => 
                           DP_OP_1090J1_126_7243_n25, S => C620_DATA2_7);
   DP_OP_1090J1_126_7243_U25 : FA_X1 port map( A => DP_OP_1090J1_126_7243_n72, 
                           B => DataPath_WRF_CUhw_curr_addr_8_port, CI => 
                           DP_OP_1090J1_126_7243_n25, CO => 
                           DP_OP_1090J1_126_7243_n24, S => C620_DATA2_8);
   DP_OP_1090J1_126_7243_U24 : FA_X1 port map( A => DP_OP_1090J1_126_7243_n72, 
                           B => DataPath_WRF_CUhw_curr_addr_9_port, CI => 
                           DP_OP_1090J1_126_7243_n24, CO => 
                           DP_OP_1090J1_126_7243_n23, S => C620_DATA2_9);
   DP_OP_1090J1_126_7243_U23 : FA_X1 port map( A => DP_OP_1090J1_126_7243_n72, 
                           B => DataPath_WRF_CUhw_curr_addr_10_port, CI => 
                           DP_OP_1090J1_126_7243_n23, CO => 
                           DP_OP_1090J1_126_7243_n22, S => C620_DATA2_10);
   DP_OP_1090J1_126_7243_U13 : FA_X1 port map( A => DP_OP_1090J1_126_7243_n72, 
                           B => DataPath_WRF_CUhw_curr_addr_20_port, CI => 
                           DP_OP_1090J1_126_7243_n13, CO => 
                           DP_OP_1090J1_126_7243_n12, S => C620_DATA2_20);
   DP_OP_1090J1_126_7243_U12 : FA_X1 port map( A => DP_OP_1090J1_126_7243_n72, 
                           B => DataPath_WRF_CUhw_curr_addr_21_port, CI => 
                           DP_OP_1090J1_126_7243_n12, CO => 
                           DP_OP_1090J1_126_7243_n11, S => C620_DATA2_21);
   DP_OP_1090J1_126_7243_U2 : XOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72,
                           B => DataPath_WRF_CUhw_curr_addr_31_port, Z => 
                           DP_OP_1090J1_126_7243_n1);
   DP_OP_751_130_5637_U244 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n31, B 
                           => n8283, ZN => DataPath_ALUhw_i_Q_EXTENDED_34_port)
                           ;
   DP_OP_751_130_5637_U248 : NAND2_X1 port map( A1 => n8281, A2 => 
                           DP_OP_751_130_5637_n191, ZN => 
                           DP_OP_751_130_5637_n31);
   DP_OP_751_130_5637_U192 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n24, B 
                           => DP_OP_751_130_5637_n162, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_41_port);
   DP_OP_751_130_5637_U197 : NAND2_X1 port map( A1 => n8270, A2 => 
                           DP_OP_751_130_5637_n161, ZN => 
                           DP_OP_751_130_5637_n24);
   DP_OP_751_130_5637_U184 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n23, B 
                           => DP_OP_751_130_5637_n156, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_42_port);
   DP_OP_751_130_5637_U188 : NAND2_X1 port map( A1 => n8279, A2 => 
                           DP_OP_751_130_5637_n155, ZN => 
                           DP_OP_751_130_5637_n23);
   DP_OP_751_130_5637_U170 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n21, B 
                           => DP_OP_751_130_5637_n148, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_44_port);
   DP_OP_751_130_5637_U174 : NAND2_X1 port map( A1 => n8278, A2 => 
                           DP_OP_751_130_5637_n147, ZN => 
                           DP_OP_751_130_5637_n21);
   DP_OP_751_130_5637_U166 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n218, 
                           A2 => DP_OP_751_130_5637_n142, ZN => 
                           DP_OP_751_130_5637_n20);
   DP_OP_751_130_5637_U149 : XOR2_X1 port map( A => DP_OP_751_130_5637_n18, B 
                           => DP_OP_751_130_5637_n135, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_47_port);
   DP_OP_751_130_5637_U152 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n216, 
                           A2 => DP_OP_751_130_5637_n134, ZN => 
                           DP_OP_751_130_5637_n18);
   DP_OP_751_130_5637_U143 : XOR2_X1 port map( A => DP_OP_751_130_5637_n17, B 
                           => DP_OP_751_130_5637_n131, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_48_port);
   DP_OP_751_130_5637_U145 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n215, 
                           A2 => DP_OP_751_130_5637_n130, ZN => 
                           DP_OP_751_130_5637_n17);
   DP_OP_751_130_5637_U135 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n16, B 
                           => DP_OP_751_130_5637_n128, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_49_port);
   DP_OP_751_130_5637_U139 : NAND2_X1 port map( A1 => n8276, A2 => 
                           DP_OP_751_130_5637_n127, ZN => 
                           DP_OP_751_130_5637_n16);
   DP_OP_751_130_5637_U129 : XOR2_X1 port map( A => DP_OP_751_130_5637_n15, B 
                           => DP_OP_751_130_5637_n123, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_50_port);
   DP_OP_751_130_5637_U131 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n213, 
                           A2 => DP_OP_751_130_5637_n122, ZN => 
                           DP_OP_751_130_5637_n15);
   DP_OP_751_130_5637_U121 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n14, B 
                           => n7682, ZN => DataPath_ALUhw_i_Q_EXTENDED_51_port)
                           ;
   DP_OP_751_130_5637_U125 : NAND2_X1 port map( A1 => n8275, A2 => 
                           DP_OP_751_130_5637_n119, ZN => 
                           DP_OP_751_130_5637_n14);
   DP_OP_751_130_5637_U115 : XOR2_X1 port map( A => DP_OP_751_130_5637_n13, B 
                           => DP_OP_751_130_5637_n115, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_52_port);
   DP_OP_751_130_5637_U117 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n211, 
                           A2 => DP_OP_751_130_5637_n114, ZN => 
                           DP_OP_751_130_5637_n13);
   DP_OP_751_130_5637_U107 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n12, B 
                           => n7853, ZN => DataPath_ALUhw_i_Q_EXTENDED_53_port)
                           ;
   DP_OP_751_130_5637_U111 : NAND2_X1 port map( A1 => n8274, A2 => 
                           DP_OP_751_130_5637_n111, ZN => 
                           DP_OP_751_130_5637_n12);
   DP_OP_751_130_5637_U101 : XOR2_X1 port map( A => DP_OP_751_130_5637_n11, B 
                           => n8053, Z => DataPath_ALUhw_i_Q_EXTENDED_54_port);
   DP_OP_751_130_5637_U103 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n209, 
                           A2 => DP_OP_751_130_5637_n106, ZN => 
                           DP_OP_751_130_5637_n11);
   DP_OP_751_130_5637_U92 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n10, B 
                           => DP_OP_751_130_5637_n104, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_55_port);
   DP_OP_751_130_5637_U84 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n9, B =>
                           n7743, ZN => DataPath_ALUhw_i_Q_EXTENDED_56_port);
   DP_OP_751_130_5637_U88 : NAND2_X1 port map( A1 => n8272, A2 => 
                           DP_OP_751_130_5637_n97, ZN => DP_OP_751_130_5637_n9)
                           ;
   DP_OP_751_130_5637_U80 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n206, 
                           A2 => DP_OP_751_130_5637_n92, ZN => 
                           DP_OP_751_130_5637_n8);
   DP_OP_751_130_5637_U74 : NAND2_X1 port map( A1 => n8271, A2 => 
                           DP_OP_751_130_5637_n89, ZN => DP_OP_751_130_5637_n7)
                           ;
   DP_OP_751_130_5637_U64 : XOR2_X1 port map( A => DP_OP_751_130_5637_n6, B => 
                           n7683, Z => DataPath_ALUhw_i_Q_EXTENDED_59_port);
   DP_OP_751_130_5637_U56 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n5, B =>
                           DP_OP_751_130_5637_n82, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_60_port);
   DP_OP_751_130_5637_U48 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n298, 
                           A2 => DP_OP_751_130_5637_n396, ZN => 
                           DP_OP_751_130_5637_n72);
   DP_OP_751_130_5637_U55 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n398, 
                           A2 => DP_OP_751_130_5637_n399, ZN => 
                           DP_OP_751_130_5637_n76);
   DP_OP_751_130_5637_U65 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n83, B2
                           => DP_OP_751_130_5637_n85, A => 
                           DP_OP_751_130_5637_n84, ZN => DP_OP_751_130_5637_n82
                           );
   DP_OP_751_130_5637_U69 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n500, 
                           A2 => DP_OP_751_130_5637_n501, ZN => 
                           DP_OP_751_130_5637_n84);
   DP_OP_751_130_5637_U83 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n602, 
                           A2 => DP_OP_751_130_5637_n603, ZN => 
                           DP_OP_751_130_5637_n92);
   DP_OP_751_130_5637_U106 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n706, 
                           A2 => DP_OP_751_130_5637_n804, ZN => 
                           DP_OP_751_130_5637_n106);
   DP_OP_751_130_5637_U114 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n806, 
                           A2 => DP_OP_751_130_5637_n807, ZN => 
                           DP_OP_751_130_5637_n111);
   DP_OP_751_130_5637_U120 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n808, 
                           A2 => DP_OP_751_130_5637_n906, ZN => 
                           DP_OP_751_130_5637_n114);
   DP_OP_751_130_5637_U122 : AOI21_X1 port map( B1 => n8275, B2 => 
                           DP_OP_751_130_5637_n120, A => 
                           DP_OP_751_130_5637_n117, ZN => 
                           DP_OP_751_130_5637_n115);
   DP_OP_751_130_5637_U128 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n908, 
                           A2 => DP_OP_751_130_5637_n909, ZN => 
                           DP_OP_751_130_5637_n119);
   DP_OP_751_130_5637_U130 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n121, 
                           B2 => DP_OP_751_130_5637_n123, A => 
                           DP_OP_751_130_5637_n122, ZN => 
                           DP_OP_751_130_5637_n120);
   DP_OP_751_130_5637_U134 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n910, 
                           A2 => DP_OP_751_130_5637_n1008, ZN => 
                           DP_OP_751_130_5637_n122);
   DP_OP_751_130_5637_U136 : AOI21_X1 port map( B1 => n8276, B2 => 
                           DP_OP_751_130_5637_n128, A => 
                           DP_OP_751_130_5637_n125, ZN => 
                           DP_OP_751_130_5637_n123);
   DP_OP_751_130_5637_U142 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1010,
                           A2 => DP_OP_751_130_5637_n1011, ZN => 
                           DP_OP_751_130_5637_n127);
   DP_OP_751_130_5637_U148 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1012,
                           A2 => DP_OP_751_130_5637_n1110, ZN => 
                           DP_OP_751_130_5637_n130);
   DP_OP_751_130_5637_U155 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1112,
                           A2 => DP_OP_751_130_5637_n1113, ZN => 
                           DP_OP_751_130_5637_n134);
   DP_OP_751_130_5637_U163 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1114,
                           A2 => DP_OP_751_130_5637_n1212, ZN => 
                           DP_OP_751_130_5637_n139);
   DP_OP_751_130_5637_U169 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1214,
                           A2 => DP_OP_751_130_5637_n1215, ZN => 
                           DP_OP_751_130_5637_n142);
   DP_OP_751_130_5637_U171 : AOI21_X1 port map( B1 => n8278, B2 => 
                           DP_OP_751_130_5637_n148, A => 
                           DP_OP_751_130_5637_n145, ZN => 
                           DP_OP_751_130_5637_n143);
   DP_OP_751_130_5637_U177 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1216,
                           A2 => DP_OP_751_130_5637_n1314, ZN => 
                           DP_OP_751_130_5637_n147);
   DP_OP_751_130_5637_U179 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n149, 
                           B2 => DP_OP_751_130_5637_n151, A => 
                           DP_OP_751_130_5637_n150, ZN => 
                           DP_OP_751_130_5637_n148);
   DP_OP_751_130_5637_U183 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1316,
                           A2 => DP_OP_751_130_5637_n1317, ZN => 
                           DP_OP_751_130_5637_n150);
   DP_OP_751_130_5637_U185 : AOI21_X1 port map( B1 => n8279, B2 => 
                           DP_OP_751_130_5637_n156, A => 
                           DP_OP_751_130_5637_n153, ZN => 
                           DP_OP_751_130_5637_n151);
   DP_OP_751_130_5637_U191 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1318,
                           A2 => DP_OP_751_130_5637_n1416, ZN => 
                           DP_OP_751_130_5637_n155);
   DP_OP_751_130_5637_U200 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1418,
                           A2 => DP_OP_751_130_5637_n1419, ZN => 
                           DP_OP_751_130_5637_n161);
   DP_OP_751_130_5637_U206 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1420,
                           A2 => DP_OP_751_130_5637_n1518, ZN => 
                           DP_OP_751_130_5637_n164);
   DP_OP_751_130_5637_U208 : AOI21_X1 port map( B1 => n8280, B2 => 
                           DP_OP_751_130_5637_n170, A => 
                           DP_OP_751_130_5637_n167, ZN => 
                           DP_OP_751_130_5637_n165);
   DP_OP_751_130_5637_U214 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1520,
                           A2 => DP_OP_751_130_5637_n1521, ZN => 
                           DP_OP_751_130_5637_n169);
   DP_OP_751_130_5637_U220 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1522,
                           A2 => DP_OP_751_130_5637_n1620, ZN => 
                           DP_OP_751_130_5637_n172);
   DP_OP_751_130_5637_U222 : AOI21_X1 port map( B1 => n8282, B2 => 
                           DP_OP_751_130_5637_n178, A => 
                           DP_OP_751_130_5637_n175, ZN => 
                           DP_OP_751_130_5637_n173);
   DP_OP_751_130_5637_U228 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1622,
                           A2 => DP_OP_751_130_5637_n1623, ZN => 
                           DP_OP_751_130_5637_n177);
   DP_OP_751_130_5637_U237 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1624,
                           A2 => DP_OP_751_130_5637_n1722, ZN => 
                           DP_OP_751_130_5637_n183);
   DP_OP_751_130_5637_U239 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n185, 
                           B2 => DP_OP_751_130_5637_n187, A => 
                           DP_OP_751_130_5637_n186, ZN => 
                           DP_OP_751_130_5637_n184);
   DP_OP_751_130_5637_U243 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1724,
                           A2 => DP_OP_751_130_5637_n1725, ZN => 
                           DP_OP_751_130_5637_n186);
   DP_OP_751_130_5637_U245 : AOI21_X1 port map( B1 => n8281, B2 => n8283, A => 
                           DP_OP_751_130_5637_n189, ZN => 
                           DP_OP_751_130_5637_n187);
   DP_OP_751_130_5637_U251 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1726,
                           A2 => DP_OP_751_130_5637_n1792, ZN => 
                           DP_OP_751_130_5637_n191);
   DP_OP_751_130_5637_U264 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1795,
                           A2 => n8076, ZN => DP_OP_751_130_5637_n198);
   DP_OP_751_130_5637_U1348 : MUX2_X1 port map( A => DP_OP_751_130_5637_n1828, 
                           B => DataPath_ALUhw_MULT_mux_out_0_1_port, S => 
                           n8264, Z => DP_OP_751_130_5637_n194);
   DP_OP_751_130_5637_U242 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n1724, 
                           A2 => DP_OP_751_130_5637_n1725, ZN => 
                           DP_OP_751_130_5637_n185);
   DP_OP_751_130_5637_U1314 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_1_3_port, B => n8263, Z 
                           => DP_OP_751_130_5637_n1725);
   DP_OP_751_130_5637_U219 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n1522, 
                           A2 => DP_OP_751_130_5637_n1620, ZN => 
                           DP_OP_751_130_5637_n171);
   DP_OP_751_130_5637_U1242 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_5_port, B => n8262, Z 
                           => DP_OP_751_130_5637_n1657);
   DP_OP_751_130_5637_U205 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n1420, 
                           A2 => DP_OP_751_130_5637_n1518, ZN => 
                           DP_OP_751_130_5637_n163);
   DP_OP_751_130_5637_U1172 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_7_port, B => n8260, Z 
                           => DP_OP_751_130_5637_n1555);
   DP_OP_751_130_5637_U1241 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_6_port, B => n8262, Z 
                           => DP_OP_751_130_5637_n1656);
   DP_OP_751_130_5637_U182 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n1316, 
                           A2 => DP_OP_751_130_5637_n1317, ZN => 
                           DP_OP_751_130_5637_n149);
   DP_OP_751_130_5637_U1102 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_9_port, B => n7798, Z 
                           => DP_OP_751_130_5637_n1453);
   DP_OP_751_130_5637_U1171 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_8_port, B => n8261, Z 
                           => DP_OP_751_130_5637_n1554);
   DP_OP_751_130_5637_U1240 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_7_port, B => n8262, Z 
                           => DP_OP_751_130_5637_n1655);
   DP_OP_751_130_5637_U1033 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_10_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1352);
   DP_OP_751_130_5637_U168 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n1214, 
                           A2 => DP_OP_751_130_5637_n1215, ZN => 
                           DP_OP_751_130_5637_n141);
   DP_OP_751_130_5637_U1032 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_11_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1351);
   DP_OP_751_130_5637_U1101 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_10_port, B => n7798, Z
                           => DP_OP_751_130_5637_n1452);
   DP_OP_751_130_5637_U1170 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_9_port, B => n8261, Z 
                           => DP_OP_751_130_5637_n1553);
   DP_OP_751_130_5637_U1239 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_8_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1654);
   DP_OP_751_130_5637_U154 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n1112, 
                           A2 => DP_OP_751_130_5637_n1113, ZN => 
                           DP_OP_751_130_5637_n133);
   DP_OP_751_130_5637_U962 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_13_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1249);
   DP_OP_751_130_5637_U1031 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_12_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1350);
   DP_OP_751_130_5637_U1100 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_11_port, B => n7798, Z
                           => DP_OP_751_130_5637_n1451);
   DP_OP_751_130_5637_U1169 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_10_port, B => n8261, Z
                           => DP_OP_751_130_5637_n1552);
   DP_OP_751_130_5637_U1238 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_9_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1653);
   DP_OP_751_130_5637_U892 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_15_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1147);
   DP_OP_751_130_5637_U961 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_14_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1248);
   DP_OP_751_130_5637_U1030 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_13_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1349);
   DP_OP_751_130_5637_U1099 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_12_port, B => n7798, Z
                           => DP_OP_751_130_5637_n1450);
   DP_OP_751_130_5637_U1168 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_11_port, B => n8261, Z
                           => DP_OP_751_130_5637_n1551);
   DP_OP_751_130_5637_U1237 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_10_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1652);
   DP_OP_751_130_5637_U823 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_16_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1046);
   DP_OP_751_130_5637_U133 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n910, 
                           A2 => DP_OP_751_130_5637_n1008, ZN => 
                           DP_OP_751_130_5637_n121);
   DP_OP_751_130_5637_U822 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_17_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1045);
   DP_OP_751_130_5637_U891 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_16_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1146);
   DP_OP_751_130_5637_U960 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_15_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1247);
   DP_OP_751_130_5637_U1029 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_14_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1348);
   DP_OP_751_130_5637_U1098 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_13_port, B => n7798, Z
                           => DP_OP_751_130_5637_n1449);
   DP_OP_751_130_5637_U1167 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_12_port, B => n8261, Z
                           => DP_OP_751_130_5637_n1550);
   DP_OP_751_130_5637_U1236 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_11_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1651);
   DP_OP_751_130_5637_U119 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n808, 
                           A2 => DP_OP_751_130_5637_n906, ZN => 
                           DP_OP_751_130_5637_n113);
   DP_OP_751_130_5637_U752 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_19_port, B => n8267, Z
                           => DP_OP_751_130_5637_n943);
   DP_OP_751_130_5637_U821 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_18_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1044);
   DP_OP_751_130_5637_U890 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_17_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1145);
   DP_OP_751_130_5637_U959 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_16_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1246);
   DP_OP_751_130_5637_U1028 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_15_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1347);
   DP_OP_751_130_5637_U1097 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_14_port, B => n7798, Z
                           => DP_OP_751_130_5637_n1448);
   DP_OP_751_130_5637_U1166 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_13_port, B => n8261, Z
                           => DP_OP_751_130_5637_n1549);
   DP_OP_751_130_5637_U1235 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_12_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1650);
   DP_OP_751_130_5637_U683 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_20_port, B => n8268, 
                           Z => DP_OP_751_130_5637_n842);
   DP_OP_751_130_5637_U682 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_21_port, B => n8268, 
                           Z => DP_OP_751_130_5637_n841);
   DP_OP_751_130_5637_U751 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_20_port, B => n8267, Z
                           => DP_OP_751_130_5637_n942);
   DP_OP_751_130_5637_U820 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_19_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1043);
   DP_OP_751_130_5637_U889 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_18_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1144);
   DP_OP_751_130_5637_U958 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_17_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1245);
   DP_OP_751_130_5637_U1027 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_16_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1346);
   DP_OP_751_130_5637_U1096 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_15_port, B => n7798, Z
                           => DP_OP_751_130_5637_n1447);
   DP_OP_751_130_5637_U1165 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_14_port, B => n8261, Z
                           => DP_OP_751_130_5637_n1548);
   DP_OP_751_130_5637_U1234 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_13_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1649);
   DP_OP_751_130_5637_U613 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_22_port, B => 
                           DP_OP_751_130_5637_n741, Z => 
                           DP_OP_751_130_5637_n740);
   DP_OP_751_130_5637_U612 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_23_port, B => 
                           DP_OP_751_130_5637_n741, Z => 
                           DP_OP_751_130_5637_n739);
   DP_OP_751_130_5637_U681 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_22_port, B => n8268, 
                           Z => DP_OP_751_130_5637_n840);
   DP_OP_751_130_5637_U750 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_21_port, B => n8267, Z
                           => DP_OP_751_130_5637_n941);
   DP_OP_751_130_5637_U819 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_20_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1042);
   DP_OP_751_130_5637_U888 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_19_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1143);
   DP_OP_751_130_5637_U957 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_18_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1244);
   DP_OP_751_130_5637_U1026 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_17_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1345);
   DP_OP_751_130_5637_U1095 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_16_port, B => n8259, Z
                           => DP_OP_751_130_5637_n1446);
   DP_OP_751_130_5637_U1164 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_15_port, B => n8261, Z
                           => DP_OP_751_130_5637_n1547);
   DP_OP_751_130_5637_U1233 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_14_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1648);
   DP_OP_751_130_5637_U1336 : MUX2_X1 port map( A => DP_OP_751_130_5637_n1816, 
                           B => DataPath_ALUhw_MULT_mux_out_0_13_port, S => 
                           n8265, Z => DP_OP_751_130_5637_n1781);
   DP_OP_751_130_5637_U1304 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_1_13_port, B => n8263, Z
                           => DP_OP_751_130_5637_n1750);
   DP_OP_751_130_5637_U543 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_24_port, B => 
                           DP_OP_751_130_5637_n639, Z => 
                           DP_OP_751_130_5637_n638);
   DP_OP_751_130_5637_U68 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n500, A2
                           => DP_OP_751_130_5637_n501, ZN => 
                           DP_OP_751_130_5637_n83);
   DP_OP_751_130_5637_U542 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_25_port, B => 
                           DP_OP_751_130_5637_n639, Z => 
                           DP_OP_751_130_5637_n637);
   DP_OP_751_130_5637_U611 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_24_port, B => 
                           DP_OP_751_130_5637_n741, Z => 
                           DP_OP_751_130_5637_n738);
   DP_OP_751_130_5637_U680 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_23_port, B => n8268, 
                           Z => DP_OP_751_130_5637_n839);
   DP_OP_751_130_5637_U749 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_22_port, B => n8267, Z
                           => DP_OP_751_130_5637_n940);
   DP_OP_751_130_5637_U818 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_21_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1041);
   DP_OP_751_130_5637_U887 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_20_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1142);
   DP_OP_751_130_5637_U956 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_19_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1243);
   DP_OP_751_130_5637_U1025 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_18_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1344);
   DP_OP_751_130_5637_U1094 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_17_port, B => n8259, Z
                           => DP_OP_751_130_5637_n1445);
   DP_OP_751_130_5637_U1163 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_16_port, B => n8261, Z
                           => DP_OP_751_130_5637_n1546);
   DP_OP_751_130_5637_U1232 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_15_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1647);
   DP_OP_751_130_5637_U1335 : MUX2_X1 port map( A => DP_OP_751_130_5637_n1815, 
                           B => DataPath_ALUhw_MULT_mux_out_0_14_port, S => 
                           n8265, Z => DP_OP_751_130_5637_n1780);
   DP_OP_751_130_5637_U1303 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_1_14_port, B => n8263, Z
                           => DP_OP_751_130_5637_n1749);
   DP_OP_751_130_5637_U473 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_13_26_port, B => 
                           DP_OP_751_130_5637_n537, Z => 
                           DP_OP_751_130_5637_n536);
   DP_OP_751_130_5637_U472 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_13_27_port, B => 
                           DP_OP_751_130_5637_n537, Z => 
                           DP_OP_751_130_5637_n535);
   DP_OP_751_130_5637_U541 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_26_port, B => 
                           DP_OP_751_130_5637_n639, Z => 
                           DP_OP_751_130_5637_n636);
   DP_OP_751_130_5637_U610 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_25_port, B => 
                           DP_OP_751_130_5637_n741, Z => 
                           DP_OP_751_130_5637_n737);
   DP_OP_751_130_5637_U679 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_24_port, B => n8268, 
                           Z => DP_OP_751_130_5637_n838);
   DP_OP_751_130_5637_U748 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_23_port, B => n8267, Z
                           => DP_OP_751_130_5637_n939);
   DP_OP_751_130_5637_U817 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_22_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1040);
   DP_OP_751_130_5637_U886 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_21_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1141);
   DP_OP_751_130_5637_U955 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_20_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1242);
   DP_OP_751_130_5637_U1024 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_19_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1343);
   DP_OP_751_130_5637_U1093 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_18_port, B => n8259, Z
                           => DP_OP_751_130_5637_n1444);
   DP_OP_751_130_5637_U1162 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_17_port, B => n8261, Z
                           => DP_OP_751_130_5637_n1545);
   DP_OP_751_130_5637_U1231 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_16_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1646);
   DP_OP_751_130_5637_U1334 : MUX2_X1 port map( A => DP_OP_751_130_5637_n1814, 
                           B => DataPath_ALUhw_MULT_mux_out_0_15_port, S => 
                           n8265, Z => DP_OP_751_130_5637_n1779);
   DP_OP_751_130_5637_U1302 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_1_15_port, B => n8263, Z
                           => DP_OP_751_130_5637_n1748);
   DP_OP_751_130_5637_U403 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_14_28_port, B => 
                           DP_OP_751_130_5637_n435, Z => 
                           DP_OP_751_130_5637_n434);
   DP_OP_751_130_5637_U47 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n396, A2
                           => DP_OP_751_130_5637_n298, ZN => 
                           DP_OP_751_130_5637_n71);
   DP_OP_751_130_5637_U402 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_14_29_port, B => 
                           DP_OP_751_130_5637_n435, Z => 
                           DP_OP_751_130_5637_n433);
   DP_OP_751_130_5637_U471 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_13_28_port, B => 
                           DP_OP_751_130_5637_n537, Z => 
                           DP_OP_751_130_5637_n534);
   DP_OP_751_130_5637_U540 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_27_port, B => 
                           DP_OP_751_130_5637_n639, Z => 
                           DP_OP_751_130_5637_n635);
   DP_OP_751_130_5637_U609 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_26_port, B => 
                           DP_OP_751_130_5637_n741, Z => 
                           DP_OP_751_130_5637_n736);
   DP_OP_751_130_5637_U678 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_25_port, B => n8268, 
                           Z => DP_OP_751_130_5637_n837);
   DP_OP_751_130_5637_U747 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_24_port, B => n8267, Z
                           => DP_OP_751_130_5637_n938);
   DP_OP_751_130_5637_U816 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_23_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1039);
   DP_OP_751_130_5637_U885 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_22_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1140);
   DP_OP_751_130_5637_U954 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_21_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1241);
   DP_OP_751_130_5637_U1023 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_20_port, B => 
                           DP_OP_751_130_5637_n1353, Z => 
                           DP_OP_751_130_5637_n1342);
   DP_OP_751_130_5637_U1092 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_19_port, B => n8259, Z
                           => DP_OP_751_130_5637_n1443);
   DP_OP_751_130_5637_U1161 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_18_port, B => n8261, Z
                           => DP_OP_751_130_5637_n1544);
   DP_OP_751_130_5637_U1230 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_17_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1645);
   DP_OP_751_130_5637_U1333 : MUX2_X1 port map( A => DP_OP_751_130_5637_n1813, 
                           B => DataPath_ALUhw_MULT_mux_out_0_16_port, S => 
                           n8265, Z => DP_OP_751_130_5637_n1778);
   DP_OP_751_130_5637_U1301 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_1_16_port, B => n8263, Z
                           => DP_OP_751_130_5637_n1747);
   DP_OP_751_130_5637_U333 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_15_30_port, B => 
                           DP_OP_751_130_5637_n333, Z => 
                           DP_OP_751_130_5637_n332);
   DP_OP_751_130_5637_U1318 : MUX2_X1 port map( A => DP_OP_751_130_5637_n1798, 
                           B => DataPath_ALUhw_MULT_mux_out_0_31_port, S => 
                           n7979, Z => DP_OP_751_130_5637_n1763);
   DP_OP_751_130_5637_U1286 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_1_31_port, B => n8263, Z
                           => DP_OP_751_130_5637_n1732);
   DP_OP_751_130_5637_U1216 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_31_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1631);
   DP_OP_751_130_5637_U1148 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_31_port, B => n8261, Z
                           => DP_OP_751_130_5637_n1531);
   DP_OP_751_130_5637_U1080 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_31_port, B => n7798, Z
                           => DP_OP_751_130_5637_n1431);
   DP_OP_751_130_5637_U1012 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_31_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1331);
   DP_OP_751_130_5637_U944 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_31_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1231);
   DP_OP_751_130_5637_U876 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_31_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1131);
   DP_OP_751_130_5637_U808 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_31_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1031);
   DP_OP_751_130_5637_U740 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_31_port, B => n8267, Z
                           => DP_OP_751_130_5637_n931);
   DP_OP_751_130_5637_U672 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_31_port, B => n8268, 
                           Z => DP_OP_751_130_5637_n831);
   DP_OP_751_130_5637_U604 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_31_port, B => 
                           DP_OP_751_130_5637_n741, Z => 
                           DP_OP_751_130_5637_n731);
   DP_OP_751_130_5637_U536 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_31_port, B => 
                           DP_OP_751_130_5637_n639, Z => 
                           DP_OP_751_130_5637_n631);
   DP_OP_751_130_5637_U468 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_13_31_port, B => 
                           DP_OP_751_130_5637_n537, Z => 
                           DP_OP_751_130_5637_n531);
   DP_OP_751_130_5637_U400 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_14_31_port, B => 
                           DP_OP_751_130_5637_n435, Z => 
                           DP_OP_751_130_5637_n431);
   DP_OP_751_130_5637_U1217 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_30_port, B => n8262, Z
                           => DP_OP_751_130_5637_n1632);
   DP_OP_751_130_5637_U1149 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_30_port, B => n8261, Z
                           => DP_OP_751_130_5637_n1532);
   DP_OP_751_130_5637_U1081 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_30_port, B => n8259, Z
                           => DP_OP_751_130_5637_n1432);
   DP_OP_751_130_5637_U1013 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_30_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1332);
   DP_OP_751_130_5637_U945 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_30_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1232);
   DP_OP_751_130_5637_U877 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_30_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1132);
   DP_OP_751_130_5637_U809 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_30_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1032);
   DP_OP_751_130_5637_U741 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_30_port, B => n8267, Z
                           => DP_OP_751_130_5637_n932);
   DP_OP_751_130_5637_U673 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_30_port, B => n8268, 
                           Z => DP_OP_751_130_5637_n832);
   DP_OP_751_130_5637_U605 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_30_port, B => 
                           DP_OP_751_130_5637_n741, Z => 
                           DP_OP_751_130_5637_n732);
   DP_OP_751_130_5637_U537 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_30_port, B => 
                           DP_OP_751_130_5637_n639, Z => 
                           DP_OP_751_130_5637_n632);
   DP_OP_751_130_5637_U469 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_13_30_port, B => 
                           DP_OP_751_130_5637_n537, Z => 
                           DP_OP_751_130_5637_n532);
   DP_OP_751_130_5637_U401 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_14_30_port, B => 
                           DP_OP_751_130_5637_n435, Z => 
                           DP_OP_751_130_5637_n432);
   DP_OP_751_130_5637_U1218 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_29_port, B => n8262, Z
                           => DP_OP_751_130_5637_n1633);
   DP_OP_751_130_5637_U1150 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_29_port, B => 
                           DP_OP_751_130_5637_n1557, Z => 
                           DP_OP_751_130_5637_n1533);
   DP_OP_751_130_5637_U1082 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_29_port, B => n8259, Z
                           => DP_OP_751_130_5637_n1433);
   DP_OP_751_130_5637_U1014 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_29_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1333);
   DP_OP_751_130_5637_U946 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_29_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1233);
   DP_OP_751_130_5637_U878 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_29_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1133);
   DP_OP_751_130_5637_U810 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_29_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1033);
   DP_OP_751_130_5637_U742 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_29_port, B => n8267, Z
                           => DP_OP_751_130_5637_n933);
   DP_OP_751_130_5637_U674 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_29_port, B => n8268, 
                           Z => DP_OP_751_130_5637_n833);
   DP_OP_751_130_5637_U606 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_29_port, B => 
                           DP_OP_751_130_5637_n741, Z => 
                           DP_OP_751_130_5637_n733);
   DP_OP_751_130_5637_U538 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_29_port, B => 
                           DP_OP_751_130_5637_n639, Z => 
                           DP_OP_751_130_5637_n633);
   DP_OP_751_130_5637_U470 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_13_29_port, B => 
                           DP_OP_751_130_5637_n537, Z => 
                           DP_OP_751_130_5637_n533);
   DP_OP_751_130_5637_U1219 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_28_port, B => n8262, Z
                           => DP_OP_751_130_5637_n1634);
   DP_OP_751_130_5637_U1151 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_28_port, B => n8260, Z
                           => DP_OP_751_130_5637_n1534);
   DP_OP_751_130_5637_U1083 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_28_port, B => n8259, Z
                           => DP_OP_751_130_5637_n1434);
   DP_OP_751_130_5637_U1015 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_28_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1334);
   DP_OP_751_130_5637_U947 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_28_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1234);
   DP_OP_751_130_5637_U879 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_28_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1134);
   DP_OP_751_130_5637_U811 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_28_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1034);
   DP_OP_751_130_5637_U743 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_28_port, B => n8267, Z
                           => DP_OP_751_130_5637_n934);
   DP_OP_751_130_5637_U675 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_28_port, B => n8268, 
                           Z => DP_OP_751_130_5637_n834);
   DP_OP_751_130_5637_U607 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_28_port, B => 
                           DP_OP_751_130_5637_n741, Z => 
                           DP_OP_751_130_5637_n734);
   DP_OP_751_130_5637_U539 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_28_port, B => 
                           DP_OP_751_130_5637_n639, Z => 
                           DP_OP_751_130_5637_n634);
   DP_OP_751_130_5637_U1220 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_27_port, B => n8262, Z
                           => DP_OP_751_130_5637_n1635);
   DP_OP_751_130_5637_U1152 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_27_port, B => n8260, Z
                           => DP_OP_751_130_5637_n1535);
   DP_OP_751_130_5637_U1084 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_27_port, B => n7798, Z
                           => DP_OP_751_130_5637_n1435);
   DP_OP_751_130_5637_U1016 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_27_port, B => 
                           DP_OP_751_130_5637_n1353, Z => 
                           DP_OP_751_130_5637_n1335);
   DP_OP_751_130_5637_U948 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_27_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1235);
   DP_OP_751_130_5637_U880 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_27_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1135);
   DP_OP_751_130_5637_U812 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_27_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1035);
   DP_OP_751_130_5637_U744 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_27_port, B => n8267, Z
                           => DP_OP_751_130_5637_n935);
   DP_OP_751_130_5637_U676 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_27_port, B => n8268, 
                           Z => DP_OP_751_130_5637_n835);
   DP_OP_751_130_5637_U608 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_27_port, B => 
                           DP_OP_751_130_5637_n741, Z => 
                           DP_OP_751_130_5637_n735);
   DP_OP_751_130_5637_U1221 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_26_port, B => n8262, Z
                           => DP_OP_751_130_5637_n1636);
   DP_OP_751_130_5637_U1153 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_26_port, B => 
                           DP_OP_751_130_5637_n1557, Z => 
                           DP_OP_751_130_5637_n1536);
   DP_OP_751_130_5637_U1085 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_26_port, B => n7798, Z
                           => DP_OP_751_130_5637_n1436);
   DP_OP_751_130_5637_U1017 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_26_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1336);
   DP_OP_751_130_5637_U949 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_26_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1236);
   DP_OP_751_130_5637_U881 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_26_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1136);
   DP_OP_751_130_5637_U813 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_26_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1036);
   DP_OP_751_130_5637_U745 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_26_port, B => n8267, Z
                           => DP_OP_751_130_5637_n936);
   DP_OP_751_130_5637_U677 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_26_port, B => n8268, 
                           Z => DP_OP_751_130_5637_n836);
   DP_OP_751_130_5637_U1222 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_25_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1637);
   DP_OP_751_130_5637_U1086 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_25_port, B => n7798, Z
                           => DP_OP_751_130_5637_n1437);
   DP_OP_751_130_5637_U1018 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_25_port, B => 
                           DP_OP_751_130_5637_n1353, Z => 
                           DP_OP_751_130_5637_n1337);
   DP_OP_751_130_5637_U950 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_25_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1237);
   DP_OP_751_130_5637_U882 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_25_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1137);
   DP_OP_751_130_5637_U814 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_25_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1037);
   DP_OP_751_130_5637_U746 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_25_port, B => n8267, Z
                           => DP_OP_751_130_5637_n937);
   DP_OP_751_130_5637_U1223 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_24_port, B => n8262, Z
                           => DP_OP_751_130_5637_n1638);
   DP_OP_751_130_5637_U1155 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_24_port, B => 
                           DP_OP_751_130_5637_n1557, Z => 
                           DP_OP_751_130_5637_n1538);
   DP_OP_751_130_5637_U1087 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_24_port, B => n7798, Z
                           => DP_OP_751_130_5637_n1438);
   DP_OP_751_130_5637_U1019 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_24_port, B => 
                           DP_OP_751_130_5637_n1353, Z => 
                           DP_OP_751_130_5637_n1338);
   DP_OP_751_130_5637_U951 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_24_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1238);
   DP_OP_751_130_5637_U883 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_24_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1138);
   DP_OP_751_130_5637_U815 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_24_port, B => n8266, Z
                           => DP_OP_751_130_5637_n1038);
   DP_OP_751_130_5637_U1224 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_23_port, B => n8262, Z
                           => DP_OP_751_130_5637_n1639);
   DP_OP_751_130_5637_U1156 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_23_port, B => n8260, Z
                           => DP_OP_751_130_5637_n1539);
   DP_OP_751_130_5637_U1088 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_23_port, B => n8259, Z
                           => DP_OP_751_130_5637_n1439);
   DP_OP_751_130_5637_U1020 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_23_port, B => 
                           DP_OP_751_130_5637_n1353, Z => 
                           DP_OP_751_130_5637_n1339);
   DP_OP_751_130_5637_U952 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_23_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1239);
   DP_OP_751_130_5637_U884 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_23_port, B => n7770, Z
                           => DP_OP_751_130_5637_n1139);
   DP_OP_751_130_5637_U1327 : MUX2_X1 port map( A => DP_OP_751_130_5637_n1807, 
                           B => DataPath_ALUhw_MULT_mux_out_0_22_port, S => 
                           n7979, Z => DP_OP_751_130_5637_n1772);
   DP_OP_751_130_5637_U1225 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_22_port, B => n8262, Z
                           => DP_OP_751_130_5637_n1640);
   DP_OP_751_130_5637_U1157 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_22_port, B => 
                           DP_OP_751_130_5637_n1557, Z => 
                           DP_OP_751_130_5637_n1540);
   DP_OP_751_130_5637_U1089 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_22_port, B => n8259, Z
                           => DP_OP_751_130_5637_n1440);
   DP_OP_751_130_5637_U1021 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_22_port, B => 
                           DP_OP_751_130_5637_n1353, Z => 
                           DP_OP_751_130_5637_n1340);
   DP_OP_751_130_5637_U953 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_22_port, B => 
                           DP_OP_751_130_5637_n1251, Z => 
                           DP_OP_751_130_5637_n1240);
   DP_OP_751_130_5637_U1158 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_21_port, B => n8260, Z
                           => DP_OP_751_130_5637_n1541);
   DP_OP_751_130_5637_U1090 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_21_port, B => n8259, Z
                           => DP_OP_751_130_5637_n1441);
   DP_OP_751_130_5637_U1022 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_21_port, B => n8258, Z
                           => DP_OP_751_130_5637_n1341);
   DP_OP_751_130_5637_U1329 : MUX2_X1 port map( A => DP_OP_751_130_5637_n1809, 
                           B => DataPath_ALUhw_MULT_mux_out_0_20_port, S => 
                           n7979, Z => DP_OP_751_130_5637_n1774);
   DP_OP_751_130_5637_U1227 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_20_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1642);
   DP_OP_751_130_5637_U1159 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_20_port, B => n8260, Z
                           => DP_OP_751_130_5637_n1542);
   DP_OP_751_130_5637_U1091 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_20_port, B => n8259, Z
                           => DP_OP_751_130_5637_n1442);
   DP_OP_751_130_5637_U1330 : MUX2_X1 port map( A => DP_OP_751_130_5637_n1810, 
                           B => DataPath_ALUhw_MULT_mux_out_0_19_port, S => 
                           n8265, Z => DP_OP_751_130_5637_n1775);
   DP_OP_751_130_5637_U1228 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_19_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1643);
   DP_OP_751_130_5637_U1160 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_19_port, B => n8261, Z
                           => DP_OP_751_130_5637_n1543);
   DP_OP_751_130_5637_U1331 : MUX2_X1 port map( A => DP_OP_751_130_5637_n1811, 
                           B => DataPath_ALUhw_MULT_mux_out_0_18_port, S => 
                           n8265, Z => DP_OP_751_130_5637_n1776);
   DP_OP_751_130_5637_U1229 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_18_port, B => 
                           DP_OP_751_130_5637_n1659, Z => 
                           DP_OP_751_130_5637_n1644);
   DP_OP_751_130_5637_U1332 : MUX2_X1 port map( A => DP_OP_751_130_5637_n1812, 
                           B => DataPath_ALUhw_MULT_mux_out_0_17_port, S => 
                           n8265, Z => DP_OP_751_130_5637_n1777);
   DP_OP_751_130_5637_U1281 : HA_X1 port map( A => DP_OP_751_130_5637_n1760, B 
                           => n8263, CO => DP_OP_751_130_5637_n1727, S => 
                           DP_OP_751_130_5637_n1726);
   DP_OP_751_130_5637_U1270 : HA_X1 port map( A => DP_OP_751_130_5637_n1750, B 
                           => DP_OP_751_130_5637_n1781, CO => 
                           DP_OP_751_130_5637_n1703, S => 
                           DP_OP_751_130_5637_n1704);
   DP_OP_751_130_5637_U1269 : HA_X1 port map( A => DP_OP_751_130_5637_n1749, B 
                           => DP_OP_751_130_5637_n1780, CO => 
                           DP_OP_751_130_5637_n1701, S => 
                           DP_OP_751_130_5637_n1702);
   DP_OP_751_130_5637_U1268 : HA_X1 port map( A => DP_OP_751_130_5637_n1748, B 
                           => DP_OP_751_130_5637_n1779, CO => 
                           DP_OP_751_130_5637_n1699, S => 
                           DP_OP_751_130_5637_n1700);
   DP_OP_751_130_5637_U1267 : HA_X1 port map( A => DP_OP_751_130_5637_n1747, B 
                           => DP_OP_751_130_5637_n1778, CO => 
                           DP_OP_751_130_5637_n1697, S => 
                           DP_OP_751_130_5637_n1698);
   DP_OP_751_130_5637_U1266 : HA_X1 port map( A => DP_OP_751_130_5637_n1746, B 
                           => DP_OP_751_130_5637_n1777, CO => 
                           DP_OP_751_130_5637_n1695, S => 
                           DP_OP_751_130_5637_n1696);
   DP_OP_751_130_5637_U1265 : HA_X1 port map( A => DP_OP_751_130_5637_n1745, B 
                           => DP_OP_751_130_5637_n1776, CO => 
                           DP_OP_751_130_5637_n1693, S => 
                           DP_OP_751_130_5637_n1694);
   DP_OP_751_130_5637_U1263 : HA_X1 port map( A => DP_OP_751_130_5637_n1743, B 
                           => DP_OP_751_130_5637_n1774, CO => 
                           DP_OP_751_130_5637_n1689, S => 
                           DP_OP_751_130_5637_n1690);
   DP_OP_751_130_5637_U1258 : HA_X1 port map( A => DP_OP_751_130_5637_n1738, B 
                           => DP_OP_751_130_5637_n1769, CO => 
                           DP_OP_751_130_5637_n1679, S => 
                           DP_OP_751_130_5637_n1680);
   DP_OP_751_130_5637_U1254 : HA_X1 port map( A => DP_OP_751_130_5637_n1734, B 
                           => DP_OP_751_130_5637_n1765, CO => 
                           DP_OP_751_130_5637_n1671, S => 
                           DP_OP_751_130_5637_n1672);
   DP_OP_751_130_5637_U1252 : HA_X1 port map( A => DP_OP_751_130_5637_n1732, B 
                           => DP_OP_751_130_5637_n1763, CO => n_3912, S => 
                           DP_OP_751_130_5637_n1668);
   DP_OP_751_130_5637_U1208 : FA_X1 port map( A => DP_OP_751_130_5637_n1721, B 
                           => DP_OP_751_130_5637_n1657, CI => 
                           DP_OP_751_130_5637_n1720, CO => 
                           DP_OP_751_130_5637_n1621, S => 
                           DP_OP_751_130_5637_n1622);
   DP_OP_751_130_5637_U1207 : FA_X1 port map( A => DP_OP_751_130_5637_n1719, B 
                           => DP_OP_751_130_5637_n1656, CI => 
                           DP_OP_751_130_5637_n1718, CO => 
                           DP_OP_751_130_5637_n1619, S => 
                           DP_OP_751_130_5637_n1620);
   DP_OP_751_130_5637_U1206 : FA_X1 port map( A => DP_OP_751_130_5637_n1717, B 
                           => DP_OP_751_130_5637_n1655, CI => 
                           DP_OP_751_130_5637_n1716, CO => 
                           DP_OP_751_130_5637_n1617, S => 
                           DP_OP_751_130_5637_n1618);
   DP_OP_751_130_5637_U1205 : FA_X1 port map( A => DP_OP_751_130_5637_n1715, B 
                           => DP_OP_751_130_5637_n1654, CI => 
                           DP_OP_751_130_5637_n1714, CO => 
                           DP_OP_751_130_5637_n1615, S => 
                           DP_OP_751_130_5637_n1616);
   DP_OP_751_130_5637_U1204 : FA_X1 port map( A => DP_OP_751_130_5637_n1713, B 
                           => DP_OP_751_130_5637_n1653, CI => 
                           DP_OP_751_130_5637_n1712, CO => 
                           DP_OP_751_130_5637_n1613, S => 
                           DP_OP_751_130_5637_n1614);
   DP_OP_751_130_5637_U1203 : FA_X1 port map( A => DP_OP_751_130_5637_n1711, B 
                           => DP_OP_751_130_5637_n1652, CI => 
                           DP_OP_751_130_5637_n1710, CO => 
                           DP_OP_751_130_5637_n1611, S => 
                           DP_OP_751_130_5637_n1612);
   DP_OP_751_130_5637_U1202 : FA_X1 port map( A => DP_OP_751_130_5637_n1709, B 
                           => DP_OP_751_130_5637_n1651, CI => 
                           DP_OP_751_130_5637_n1708, CO => 
                           DP_OP_751_130_5637_n1609, S => 
                           DP_OP_751_130_5637_n1610);
   DP_OP_751_130_5637_U1201 : FA_X1 port map( A => DP_OP_751_130_5637_n1707, B 
                           => DP_OP_751_130_5637_n1650, CI => 
                           DP_OP_751_130_5637_n1706, CO => 
                           DP_OP_751_130_5637_n1607, S => 
                           DP_OP_751_130_5637_n1608);
   DP_OP_751_130_5637_U1200 : FA_X1 port map( A => DP_OP_751_130_5637_n1705, B 
                           => DP_OP_751_130_5637_n1649, CI => 
                           DP_OP_751_130_5637_n1704, CO => 
                           DP_OP_751_130_5637_n1605, S => 
                           DP_OP_751_130_5637_n1606);
   DP_OP_751_130_5637_U1199 : FA_X1 port map( A => DP_OP_751_130_5637_n1703, B 
                           => DP_OP_751_130_5637_n1648, CI => 
                           DP_OP_751_130_5637_n1702, CO => 
                           DP_OP_751_130_5637_n1603, S => 
                           DP_OP_751_130_5637_n1604);
   DP_OP_751_130_5637_U1198 : FA_X1 port map( A => DP_OP_751_130_5637_n1701, B 
                           => DP_OP_751_130_5637_n1647, CI => 
                           DP_OP_751_130_5637_n1700, CO => 
                           DP_OP_751_130_5637_n1601, S => 
                           DP_OP_751_130_5637_n1602);
   DP_OP_751_130_5637_U1197 : FA_X1 port map( A => DP_OP_751_130_5637_n1699, B 
                           => DP_OP_751_130_5637_n1646, CI => 
                           DP_OP_751_130_5637_n1698, CO => 
                           DP_OP_751_130_5637_n1599, S => 
                           DP_OP_751_130_5637_n1600);
   DP_OP_751_130_5637_U1196 : FA_X1 port map( A => DP_OP_751_130_5637_n1697, B 
                           => DP_OP_751_130_5637_n1645, CI => 
                           DP_OP_751_130_5637_n1696, CO => 
                           DP_OP_751_130_5637_n1597, S => 
                           DP_OP_751_130_5637_n1598);
   DP_OP_751_130_5637_U1195 : FA_X1 port map( A => DP_OP_751_130_5637_n1695, B 
                           => DP_OP_751_130_5637_n1644, CI => 
                           DP_OP_751_130_5637_n1694, CO => 
                           DP_OP_751_130_5637_n1595, S => 
                           DP_OP_751_130_5637_n1596);
   DP_OP_751_130_5637_U1194 : FA_X1 port map( A => DP_OP_751_130_5637_n1693, B 
                           => DP_OP_751_130_5637_n1643, CI => 
                           DP_OP_751_130_5637_n1692, CO => 
                           DP_OP_751_130_5637_n1593, S => 
                           DP_OP_751_130_5637_n1594);
   DP_OP_751_130_5637_U1193 : FA_X1 port map( A => DP_OP_751_130_5637_n1691, B 
                           => DP_OP_751_130_5637_n1642, CI => 
                           DP_OP_751_130_5637_n1690, CO => 
                           DP_OP_751_130_5637_n1591, S => 
                           DP_OP_751_130_5637_n1592);
   DP_OP_751_130_5637_U1191 : FA_X1 port map( A => DP_OP_751_130_5637_n1687, B 
                           => DP_OP_751_130_5637_n1640, CI => 
                           DP_OP_751_130_5637_n1686, CO => 
                           DP_OP_751_130_5637_n1587, S => 
                           DP_OP_751_130_5637_n1588);
   DP_OP_751_130_5637_U1189 : FA_X1 port map( A => DP_OP_751_130_5637_n1638, B 
                           => DP_OP_751_130_5637_n1683, CI => 
                           DP_OP_751_130_5637_n1682, CO => 
                           DP_OP_751_130_5637_n1583, S => 
                           DP_OP_751_130_5637_n1584);
   DP_OP_751_130_5637_U1187 : FA_X1 port map( A => DP_OP_751_130_5637_n1679, B 
                           => DP_OP_751_130_5637_n1636, CI => 
                           DP_OP_751_130_5637_n1678, CO => 
                           DP_OP_751_130_5637_n1579, S => 
                           DP_OP_751_130_5637_n1580);
   DP_OP_751_130_5637_U1185 : FA_X1 port map( A => DP_OP_751_130_5637_n1675, B 
                           => DP_OP_751_130_5637_n1634, CI => 
                           DP_OP_751_130_5637_n1674, CO => 
                           DP_OP_751_130_5637_n1575, S => 
                           DP_OP_751_130_5637_n1576);
   DP_OP_751_130_5637_U1184 : FA_X1 port map( A => DP_OP_751_130_5637_n1673, B 
                           => DP_OP_751_130_5637_n1633, CI => 
                           DP_OP_751_130_5637_n1672, CO => 
                           DP_OP_751_130_5637_n1573, S => 
                           DP_OP_751_130_5637_n1574);
   DP_OP_751_130_5637_U1183 : FA_X1 port map( A => DP_OP_751_130_5637_n1671, B 
                           => DP_OP_751_130_5637_n1632, CI => 
                           DP_OP_751_130_5637_n1670, CO => 
                           DP_OP_751_130_5637_n1571, S => 
                           DP_OP_751_130_5637_n1572);
   DP_OP_751_130_5637_U1138 : FA_X1 port map( A => DP_OP_751_130_5637_n1619, B 
                           => DP_OP_751_130_5637_n1555, CI => 
                           DP_OP_751_130_5637_n1618, CO => 
                           DP_OP_751_130_5637_n1519, S => 
                           DP_OP_751_130_5637_n1520);
   DP_OP_751_130_5637_U1137 : FA_X1 port map( A => DP_OP_751_130_5637_n1617, B 
                           => DP_OP_751_130_5637_n1554, CI => 
                           DP_OP_751_130_5637_n1616, CO => 
                           DP_OP_751_130_5637_n1517, S => 
                           DP_OP_751_130_5637_n1518);
   DP_OP_751_130_5637_U1136 : FA_X1 port map( A => DP_OP_751_130_5637_n1615, B 
                           => DP_OP_751_130_5637_n1553, CI => 
                           DP_OP_751_130_5637_n1614, CO => 
                           DP_OP_751_130_5637_n1515, S => 
                           DP_OP_751_130_5637_n1516);
   DP_OP_751_130_5637_U1135 : FA_X1 port map( A => DP_OP_751_130_5637_n1613, B 
                           => DP_OP_751_130_5637_n1552, CI => 
                           DP_OP_751_130_5637_n1612, CO => 
                           DP_OP_751_130_5637_n1513, S => 
                           DP_OP_751_130_5637_n1514);
   DP_OP_751_130_5637_U1134 : FA_X1 port map( A => DP_OP_751_130_5637_n1611, B 
                           => DP_OP_751_130_5637_n1551, CI => 
                           DP_OP_751_130_5637_n1610, CO => 
                           DP_OP_751_130_5637_n1511, S => 
                           DP_OP_751_130_5637_n1512);
   DP_OP_751_130_5637_U1133 : FA_X1 port map( A => DP_OP_751_130_5637_n1609, B 
                           => DP_OP_751_130_5637_n1550, CI => 
                           DP_OP_751_130_5637_n1608, CO => 
                           DP_OP_751_130_5637_n1509, S => 
                           DP_OP_751_130_5637_n1510);
   DP_OP_751_130_5637_U1132 : FA_X1 port map( A => DP_OP_751_130_5637_n1607, B 
                           => DP_OP_751_130_5637_n1549, CI => 
                           DP_OP_751_130_5637_n1606, CO => 
                           DP_OP_751_130_5637_n1507, S => 
                           DP_OP_751_130_5637_n1508);
   DP_OP_751_130_5637_U1131 : FA_X1 port map( A => DP_OP_751_130_5637_n1605, B 
                           => DP_OP_751_130_5637_n1548, CI => 
                           DP_OP_751_130_5637_n1604, CO => 
                           DP_OP_751_130_5637_n1505, S => 
                           DP_OP_751_130_5637_n1506);
   DP_OP_751_130_5637_U1130 : FA_X1 port map( A => DP_OP_751_130_5637_n1603, B 
                           => DP_OP_751_130_5637_n1547, CI => 
                           DP_OP_751_130_5637_n1602, CO => 
                           DP_OP_751_130_5637_n1503, S => 
                           DP_OP_751_130_5637_n1504);
   DP_OP_751_130_5637_U1129 : FA_X1 port map( A => DP_OP_751_130_5637_n1601, B 
                           => DP_OP_751_130_5637_n1546, CI => 
                           DP_OP_751_130_5637_n1600, CO => 
                           DP_OP_751_130_5637_n1501, S => 
                           DP_OP_751_130_5637_n1502);
   DP_OP_751_130_5637_U1128 : FA_X1 port map( A => DP_OP_751_130_5637_n1599, B 
                           => DP_OP_751_130_5637_n1545, CI => 
                           DP_OP_751_130_5637_n1598, CO => 
                           DP_OP_751_130_5637_n1499, S => 
                           DP_OP_751_130_5637_n1500);
   DP_OP_751_130_5637_U1127 : FA_X1 port map( A => DP_OP_751_130_5637_n1597, B 
                           => DP_OP_751_130_5637_n1544, CI => 
                           DP_OP_751_130_5637_n1596, CO => 
                           DP_OP_751_130_5637_n1497, S => 
                           DP_OP_751_130_5637_n1498);
   DP_OP_751_130_5637_U1126 : FA_X1 port map( A => DP_OP_751_130_5637_n1595, B 
                           => DP_OP_751_130_5637_n1543, CI => 
                           DP_OP_751_130_5637_n1594, CO => 
                           DP_OP_751_130_5637_n1495, S => 
                           DP_OP_751_130_5637_n1496);
   DP_OP_751_130_5637_U1114 : FA_X1 port map( A => DP_OP_751_130_5637_n1571, B 
                           => DP_OP_751_130_5637_n1531, CI => 
                           DP_OP_751_130_5637_n1570, CO => n_3913, S => 
                           DP_OP_751_130_5637_n1472);
   DP_OP_751_130_5637_U1068 : FA_X1 port map( A => DP_OP_751_130_5637_n1517, B 
                           => DP_OP_751_130_5637_n1453, CI => 
                           DP_OP_751_130_5637_n1516, CO => 
                           DP_OP_751_130_5637_n1417, S => 
                           DP_OP_751_130_5637_n1418);
   DP_OP_751_130_5637_U1067 : FA_X1 port map( A => DP_OP_751_130_5637_n1515, B 
                           => DP_OP_751_130_5637_n1452, CI => 
                           DP_OP_751_130_5637_n1514, CO => 
                           DP_OP_751_130_5637_n1415, S => 
                           DP_OP_751_130_5637_n1416);
   DP_OP_751_130_5637_U1066 : FA_X1 port map( A => DP_OP_751_130_5637_n1513, B 
                           => DP_OP_751_130_5637_n1451, CI => 
                           DP_OP_751_130_5637_n1512, CO => 
                           DP_OP_751_130_5637_n1413, S => 
                           DP_OP_751_130_5637_n1414);
   DP_OP_751_130_5637_U1065 : FA_X1 port map( A => DP_OP_751_130_5637_n1511, B 
                           => DP_OP_751_130_5637_n1450, CI => 
                           DP_OP_751_130_5637_n1510, CO => 
                           DP_OP_751_130_5637_n1411, S => 
                           DP_OP_751_130_5637_n1412);
   DP_OP_751_130_5637_U1064 : FA_X1 port map( A => DP_OP_751_130_5637_n1509, B 
                           => DP_OP_751_130_5637_n1449, CI => 
                           DP_OP_751_130_5637_n1508, CO => 
                           DP_OP_751_130_5637_n1409, S => 
                           DP_OP_751_130_5637_n1410);
   DP_OP_751_130_5637_U1063 : FA_X1 port map( A => DP_OP_751_130_5637_n1507, B 
                           => DP_OP_751_130_5637_n1448, CI => 
                           DP_OP_751_130_5637_n1506, CO => 
                           DP_OP_751_130_5637_n1407, S => 
                           DP_OP_751_130_5637_n1408);
   DP_OP_751_130_5637_U1062 : FA_X1 port map( A => DP_OP_751_130_5637_n1505, B 
                           => DP_OP_751_130_5637_n1447, CI => 
                           DP_OP_751_130_5637_n1504, CO => 
                           DP_OP_751_130_5637_n1405, S => 
                           DP_OP_751_130_5637_n1406);
   DP_OP_751_130_5637_U1061 : FA_X1 port map( A => DP_OP_751_130_5637_n1503, B 
                           => DP_OP_751_130_5637_n1446, CI => 
                           DP_OP_751_130_5637_n1502, CO => 
                           DP_OP_751_130_5637_n1403, S => 
                           DP_OP_751_130_5637_n1404);
   DP_OP_751_130_5637_U1060 : FA_X1 port map( A => DP_OP_751_130_5637_n1501, B 
                           => DP_OP_751_130_5637_n1445, CI => 
                           DP_OP_751_130_5637_n1500, CO => 
                           DP_OP_751_130_5637_n1401, S => 
                           DP_OP_751_130_5637_n1402);
   DP_OP_751_130_5637_U1059 : FA_X1 port map( A => DP_OP_751_130_5637_n1499, B 
                           => DP_OP_751_130_5637_n1444, CI => 
                           DP_OP_751_130_5637_n1498, CO => 
                           DP_OP_751_130_5637_n1399, S => 
                           DP_OP_751_130_5637_n1400);
   DP_OP_751_130_5637_U1058 : FA_X1 port map( A => DP_OP_751_130_5637_n1497, B 
                           => DP_OP_751_130_5637_n1443, CI => 
                           DP_OP_751_130_5637_n1496, CO => 
                           DP_OP_751_130_5637_n1397, S => 
                           DP_OP_751_130_5637_n1398);
   DP_OP_751_130_5637_U1057 : FA_X1 port map( A => DP_OP_751_130_5637_n1495, B 
                           => DP_OP_751_130_5637_n1442, CI => 
                           DP_OP_751_130_5637_n1494, CO => 
                           DP_OP_751_130_5637_n1395, S => 
                           DP_OP_751_130_5637_n1396);
   DP_OP_751_130_5637_U1056 : FA_X1 port map( A => DP_OP_751_130_5637_n1493, B 
                           => DP_OP_751_130_5637_n1441, CI => 
                           DP_OP_751_130_5637_n1492, CO => 
                           DP_OP_751_130_5637_n1393, S => 
                           DP_OP_751_130_5637_n1394);
   DP_OP_751_130_5637_U1053 : FA_X1 port map( A => DP_OP_751_130_5637_n1487, B 
                           => DP_OP_751_130_5637_n1438, CI => 
                           DP_OP_751_130_5637_n1486, CO => 
                           DP_OP_751_130_5637_n1387, S => 
                           DP_OP_751_130_5637_n1388);
   DP_OP_751_130_5637_U1052 : FA_X1 port map( A => DP_OP_751_130_5637_n1485, B 
                           => DP_OP_751_130_5637_n1437, CI => 
                           DP_OP_751_130_5637_n1484, CO => 
                           DP_OP_751_130_5637_n1385, S => 
                           DP_OP_751_130_5637_n1386);
   DP_OP_751_130_5637_U998 : FA_X1 port map( A => DP_OP_751_130_5637_n1415, B 
                           => DP_OP_751_130_5637_n1351, CI => 
                           DP_OP_751_130_5637_n1414, CO => 
                           DP_OP_751_130_5637_n1315, S => 
                           DP_OP_751_130_5637_n1316);
   DP_OP_751_130_5637_U997 : FA_X1 port map( A => DP_OP_751_130_5637_n1413, B 
                           => DP_OP_751_130_5637_n1350, CI => 
                           DP_OP_751_130_5637_n1412, CO => 
                           DP_OP_751_130_5637_n1313, S => 
                           DP_OP_751_130_5637_n1314);
   DP_OP_751_130_5637_U996 : FA_X1 port map( A => DP_OP_751_130_5637_n1411, B 
                           => DP_OP_751_130_5637_n1349, CI => 
                           DP_OP_751_130_5637_n1410, CO => 
                           DP_OP_751_130_5637_n1311, S => 
                           DP_OP_751_130_5637_n1312);
   DP_OP_751_130_5637_U995 : FA_X1 port map( A => DP_OP_751_130_5637_n1409, B 
                           => DP_OP_751_130_5637_n1348, CI => 
                           DP_OP_751_130_5637_n1408, CO => 
                           DP_OP_751_130_5637_n1309, S => 
                           DP_OP_751_130_5637_n1310);
   DP_OP_751_130_5637_U994 : FA_X1 port map( A => DP_OP_751_130_5637_n1407, B 
                           => DP_OP_751_130_5637_n1347, CI => 
                           DP_OP_751_130_5637_n1406, CO => 
                           DP_OP_751_130_5637_n1307, S => 
                           DP_OP_751_130_5637_n1308);
   DP_OP_751_130_5637_U993 : FA_X1 port map( A => DP_OP_751_130_5637_n1405, B 
                           => DP_OP_751_130_5637_n1346, CI => 
                           DP_OP_751_130_5637_n1404, CO => 
                           DP_OP_751_130_5637_n1305, S => 
                           DP_OP_751_130_5637_n1306);
   DP_OP_751_130_5637_U992 : FA_X1 port map( A => DP_OP_751_130_5637_n1403, B 
                           => DP_OP_751_130_5637_n1345, CI => 
                           DP_OP_751_130_5637_n1402, CO => 
                           DP_OP_751_130_5637_n1303, S => 
                           DP_OP_751_130_5637_n1304);
   DP_OP_751_130_5637_U991 : FA_X1 port map( A => DP_OP_751_130_5637_n1401, B 
                           => DP_OP_751_130_5637_n1344, CI => 
                           DP_OP_751_130_5637_n1400, CO => 
                           DP_OP_751_130_5637_n1301, S => 
                           DP_OP_751_130_5637_n1302);
   DP_OP_751_130_5637_U990 : FA_X1 port map( A => DP_OP_751_130_5637_n1399, B 
                           => DP_OP_751_130_5637_n1343, CI => 
                           DP_OP_751_130_5637_n1398, CO => 
                           DP_OP_751_130_5637_n1299, S => 
                           DP_OP_751_130_5637_n1300);
   DP_OP_751_130_5637_U989 : FA_X1 port map( A => DP_OP_751_130_5637_n1397, B 
                           => DP_OP_751_130_5637_n1342, CI => 
                           DP_OP_751_130_5637_n1396, CO => 
                           DP_OP_751_130_5637_n1297, S => 
                           DP_OP_751_130_5637_n1298);
   DP_OP_751_130_5637_U988 : FA_X1 port map( A => DP_OP_751_130_5637_n1395, B 
                           => DP_OP_751_130_5637_n1341, CI => 
                           DP_OP_751_130_5637_n1394, CO => 
                           DP_OP_751_130_5637_n1295, S => 
                           DP_OP_751_130_5637_n1296);
   DP_OP_751_130_5637_U985 : FA_X1 port map( A => DP_OP_751_130_5637_n1389, B 
                           => DP_OP_751_130_5637_n1338, CI => 
                           DP_OP_751_130_5637_n1388, CO => 
                           DP_OP_751_130_5637_n1289, S => 
                           DP_OP_751_130_5637_n1290);
   DP_OP_751_130_5637_U984 : FA_X1 port map( A => DP_OP_751_130_5637_n1387, B 
                           => DP_OP_751_130_5637_n1337, CI => 
                           DP_OP_751_130_5637_n1386, CO => 
                           DP_OP_751_130_5637_n1287, S => 
                           DP_OP_751_130_5637_n1288);
   DP_OP_751_130_5637_U983 : FA_X1 port map( A => DP_OP_751_130_5637_n1385, B 
                           => DP_OP_751_130_5637_n1336, CI => 
                           DP_OP_751_130_5637_n1384, CO => 
                           DP_OP_751_130_5637_n1285, S => 
                           DP_OP_751_130_5637_n1286);
   DP_OP_751_130_5637_U981 : FA_X1 port map( A => DP_OP_751_130_5637_n1381, B 
                           => DP_OP_751_130_5637_n1334, CI => 
                           DP_OP_751_130_5637_n1380, CO => 
                           DP_OP_751_130_5637_n1281, S => 
                           DP_OP_751_130_5637_n1282);
   DP_OP_751_130_5637_U978 : FA_X1 port map( A => DP_OP_751_130_5637_n1375, B 
                           => DP_OP_751_130_5637_n1331, CI => 
                           DP_OP_751_130_5637_n1374, CO => n_3914, S => 
                           DP_OP_751_130_5637_n1276);
   DP_OP_751_130_5637_U928 : FA_X1 port map( A => DP_OP_751_130_5637_n1313, B 
                           => DP_OP_751_130_5637_n1249, CI => 
                           DP_OP_751_130_5637_n1312, CO => 
                           DP_OP_751_130_5637_n1213, S => 
                           DP_OP_751_130_5637_n1214);
   DP_OP_751_130_5637_U927 : FA_X1 port map( A => DP_OP_751_130_5637_n1311, B 
                           => DP_OP_751_130_5637_n1248, CI => 
                           DP_OP_751_130_5637_n1310, CO => 
                           DP_OP_751_130_5637_n1211, S => 
                           DP_OP_751_130_5637_n1212);
   DP_OP_751_130_5637_U926 : FA_X1 port map( A => DP_OP_751_130_5637_n1309, B 
                           => DP_OP_751_130_5637_n1247, CI => 
                           DP_OP_751_130_5637_n1308, CO => 
                           DP_OP_751_130_5637_n1209, S => 
                           DP_OP_751_130_5637_n1210);
   DP_OP_751_130_5637_U925 : FA_X1 port map( A => DP_OP_751_130_5637_n1307, B 
                           => DP_OP_751_130_5637_n1246, CI => 
                           DP_OP_751_130_5637_n1306, CO => 
                           DP_OP_751_130_5637_n1207, S => 
                           DP_OP_751_130_5637_n1208);
   DP_OP_751_130_5637_U924 : FA_X1 port map( A => DP_OP_751_130_5637_n1305, B 
                           => DP_OP_751_130_5637_n1245, CI => 
                           DP_OP_751_130_5637_n1304, CO => 
                           DP_OP_751_130_5637_n1205, S => 
                           DP_OP_751_130_5637_n1206);
   DP_OP_751_130_5637_U923 : FA_X1 port map( A => DP_OP_751_130_5637_n1303, B 
                           => DP_OP_751_130_5637_n1244, CI => 
                           DP_OP_751_130_5637_n1302, CO => 
                           DP_OP_751_130_5637_n1203, S => 
                           DP_OP_751_130_5637_n1204);
   DP_OP_751_130_5637_U922 : FA_X1 port map( A => DP_OP_751_130_5637_n1301, B 
                           => DP_OP_751_130_5637_n1243, CI => 
                           DP_OP_751_130_5637_n1300, CO => 
                           DP_OP_751_130_5637_n1201, S => 
                           DP_OP_751_130_5637_n1202);
   DP_OP_751_130_5637_U921 : FA_X1 port map( A => DP_OP_751_130_5637_n1299, B 
                           => DP_OP_751_130_5637_n1242, CI => 
                           DP_OP_751_130_5637_n1298, CO => 
                           DP_OP_751_130_5637_n1199, S => 
                           DP_OP_751_130_5637_n1200);
   DP_OP_751_130_5637_U920 : FA_X1 port map( A => DP_OP_751_130_5637_n1297, B 
                           => DP_OP_751_130_5637_n1241, CI => 
                           DP_OP_751_130_5637_n1296, CO => 
                           DP_OP_751_130_5637_n1197, S => 
                           DP_OP_751_130_5637_n1198);
   DP_OP_751_130_5637_U919 : FA_X1 port map( A => DP_OP_751_130_5637_n1295, B 
                           => DP_OP_751_130_5637_n1240, CI => 
                           DP_OP_751_130_5637_n1294, CO => 
                           DP_OP_751_130_5637_n1195, S => 
                           DP_OP_751_130_5637_n1196);
   DP_OP_751_130_5637_U918 : FA_X1 port map( A => DP_OP_751_130_5637_n1293, B 
                           => DP_OP_751_130_5637_n1239, CI => 
                           DP_OP_751_130_5637_n1292, CO => 
                           DP_OP_751_130_5637_n1193, S => 
                           DP_OP_751_130_5637_n1194);
   DP_OP_751_130_5637_U917 : FA_X1 port map( A => DP_OP_751_130_5637_n1291, B 
                           => DP_OP_751_130_5637_n1238, CI => 
                           DP_OP_751_130_5637_n1290, CO => 
                           DP_OP_751_130_5637_n1191, S => 
                           DP_OP_751_130_5637_n1192);
   DP_OP_751_130_5637_U916 : FA_X1 port map( A => DP_OP_751_130_5637_n1289, B 
                           => DP_OP_751_130_5637_n1237, CI => 
                           DP_OP_751_130_5637_n1288, CO => 
                           DP_OP_751_130_5637_n1189, S => 
                           DP_OP_751_130_5637_n1190);
   DP_OP_751_130_5637_U915 : FA_X1 port map( A => DP_OP_751_130_5637_n1287, B 
                           => DP_OP_751_130_5637_n1236, CI => 
                           DP_OP_751_130_5637_n1286, CO => 
                           DP_OP_751_130_5637_n1187, S => 
                           DP_OP_751_130_5637_n1188);
   DP_OP_751_130_5637_U914 : FA_X1 port map( A => DP_OP_751_130_5637_n1285, B 
                           => DP_OP_751_130_5637_n1235, CI => 
                           DP_OP_751_130_5637_n1284, CO => 
                           DP_OP_751_130_5637_n1185, S => 
                           DP_OP_751_130_5637_n1186);
   DP_OP_751_130_5637_U912 : FA_X1 port map( A => DP_OP_751_130_5637_n1281, B 
                           => DP_OP_751_130_5637_n1233, CI => 
                           DP_OP_751_130_5637_n1280, CO => 
                           DP_OP_751_130_5637_n1181, S => 
                           DP_OP_751_130_5637_n1182);
   DP_OP_751_130_5637_U910 : FA_X1 port map( A => DP_OP_751_130_5637_n1277, B 
                           => DP_OP_751_130_5637_n1231, CI => 
                           DP_OP_751_130_5637_n1276, CO => n_3915, S => 
                           DP_OP_751_130_5637_n1178);
   DP_OP_751_130_5637_U858 : FA_X1 port map( A => DP_OP_751_130_5637_n1211, B 
                           => DP_OP_751_130_5637_n1147, CI => 
                           DP_OP_751_130_5637_n1210, CO => 
                           DP_OP_751_130_5637_n1111, S => 
                           DP_OP_751_130_5637_n1112);
   DP_OP_751_130_5637_U857 : FA_X1 port map( A => DP_OP_751_130_5637_n1209, B 
                           => DP_OP_751_130_5637_n1146, CI => 
                           DP_OP_751_130_5637_n1208, CO => 
                           DP_OP_751_130_5637_n1109, S => 
                           DP_OP_751_130_5637_n1110);
   DP_OP_751_130_5637_U856 : FA_X1 port map( A => DP_OP_751_130_5637_n1207, B 
                           => DP_OP_751_130_5637_n1145, CI => 
                           DP_OP_751_130_5637_n1206, CO => 
                           DP_OP_751_130_5637_n1107, S => 
                           DP_OP_751_130_5637_n1108);
   DP_OP_751_130_5637_U855 : FA_X1 port map( A => DP_OP_751_130_5637_n1205, B 
                           => DP_OP_751_130_5637_n1144, CI => 
                           DP_OP_751_130_5637_n1204, CO => 
                           DP_OP_751_130_5637_n1105, S => 
                           DP_OP_751_130_5637_n1106);
   DP_OP_751_130_5637_U854 : FA_X1 port map( A => DP_OP_751_130_5637_n1203, B 
                           => DP_OP_751_130_5637_n1143, CI => 
                           DP_OP_751_130_5637_n1202, CO => 
                           DP_OP_751_130_5637_n1103, S => 
                           DP_OP_751_130_5637_n1104);
   DP_OP_751_130_5637_U853 : FA_X1 port map( A => DP_OP_751_130_5637_n1201, B 
                           => DP_OP_751_130_5637_n1142, CI => 
                           DP_OP_751_130_5637_n1200, CO => 
                           DP_OP_751_130_5637_n1101, S => 
                           DP_OP_751_130_5637_n1102);
   DP_OP_751_130_5637_U852 : FA_X1 port map( A => DP_OP_751_130_5637_n1199, B 
                           => DP_OP_751_130_5637_n1141, CI => 
                           DP_OP_751_130_5637_n1198, CO => 
                           DP_OP_751_130_5637_n1099, S => 
                           DP_OP_751_130_5637_n1100);
   DP_OP_751_130_5637_U851 : FA_X1 port map( A => DP_OP_751_130_5637_n1197, B 
                           => DP_OP_751_130_5637_n1140, CI => 
                           DP_OP_751_130_5637_n1196, CO => 
                           DP_OP_751_130_5637_n1097, S => 
                           DP_OP_751_130_5637_n1098);
   DP_OP_751_130_5637_U850 : FA_X1 port map( A => DP_OP_751_130_5637_n1195, B 
                           => DP_OP_751_130_5637_n1139, CI => 
                           DP_OP_751_130_5637_n1194, CO => 
                           DP_OP_751_130_5637_n1095, S => 
                           DP_OP_751_130_5637_n1096);
   DP_OP_751_130_5637_U848 : FA_X1 port map( A => DP_OP_751_130_5637_n1191, B 
                           => DP_OP_751_130_5637_n1137, CI => 
                           DP_OP_751_130_5637_n1190, CO => 
                           DP_OP_751_130_5637_n1091, S => 
                           DP_OP_751_130_5637_n1092);
   DP_OP_751_130_5637_U847 : FA_X1 port map( A => DP_OP_751_130_5637_n1189, B 
                           => DP_OP_751_130_5637_n1136, CI => 
                           DP_OP_751_130_5637_n1188, CO => 
                           DP_OP_751_130_5637_n1089, S => 
                           DP_OP_751_130_5637_n1090);
   DP_OP_751_130_5637_U846 : FA_X1 port map( A => DP_OP_751_130_5637_n1187, B 
                           => DP_OP_751_130_5637_n1135, CI => 
                           DP_OP_751_130_5637_n1186, CO => 
                           DP_OP_751_130_5637_n1087, S => 
                           DP_OP_751_130_5637_n1088);
   DP_OP_751_130_5637_U845 : FA_X1 port map( A => DP_OP_751_130_5637_n1185, B 
                           => DP_OP_751_130_5637_n1134, CI => 
                           DP_OP_751_130_5637_n1184, CO => 
                           DP_OP_751_130_5637_n1085, S => 
                           DP_OP_751_130_5637_n1086);
   DP_OP_751_130_5637_U844 : FA_X1 port map( A => DP_OP_751_130_5637_n1183, B 
                           => DP_OP_751_130_5637_n1133, CI => 
                           DP_OP_751_130_5637_n1182, CO => 
                           DP_OP_751_130_5637_n1083, S => 
                           DP_OP_751_130_5637_n1084);
   DP_OP_751_130_5637_U843 : FA_X1 port map( A => DP_OP_751_130_5637_n1181, B 
                           => DP_OP_751_130_5637_n1132, CI => 
                           DP_OP_751_130_5637_n1180, CO => 
                           DP_OP_751_130_5637_n1081, S => 
                           DP_OP_751_130_5637_n1082);
   DP_OP_751_130_5637_U789 : FA_X1 port map( A => DP_OP_751_130_5637_n1046, B 
                           => n8266, CI => DP_OP_751_130_5637_n1111, CO => 
                           DP_OP_751_130_5637_n1011, S => 
                           DP_OP_751_130_5637_n1012);
   DP_OP_751_130_5637_U788 : FA_X1 port map( A => DP_OP_751_130_5637_n1109, B 
                           => DP_OP_751_130_5637_n1045, CI => 
                           DP_OP_751_130_5637_n1108, CO => 
                           DP_OP_751_130_5637_n1009, S => 
                           DP_OP_751_130_5637_n1010);
   DP_OP_751_130_5637_U787 : FA_X1 port map( A => DP_OP_751_130_5637_n1107, B 
                           => DP_OP_751_130_5637_n1044, CI => 
                           DP_OP_751_130_5637_n1106, CO => 
                           DP_OP_751_130_5637_n1007, S => 
                           DP_OP_751_130_5637_n1008);
   DP_OP_751_130_5637_U786 : FA_X1 port map( A => DP_OP_751_130_5637_n1105, B 
                           => DP_OP_751_130_5637_n1043, CI => 
                           DP_OP_751_130_5637_n1104, CO => 
                           DP_OP_751_130_5637_n1005, S => 
                           DP_OP_751_130_5637_n1006);
   DP_OP_751_130_5637_U785 : FA_X1 port map( A => DP_OP_751_130_5637_n1103, B 
                           => DP_OP_751_130_5637_n1042, CI => 
                           DP_OP_751_130_5637_n1102, CO => 
                           DP_OP_751_130_5637_n1003, S => 
                           DP_OP_751_130_5637_n1004);
   DP_OP_751_130_5637_U784 : FA_X1 port map( A => DP_OP_751_130_5637_n1101, B 
                           => DP_OP_751_130_5637_n1041, CI => 
                           DP_OP_751_130_5637_n1100, CO => 
                           DP_OP_751_130_5637_n1001, S => 
                           DP_OP_751_130_5637_n1002);
   DP_OP_751_130_5637_U783 : FA_X1 port map( A => DP_OP_751_130_5637_n1099, B 
                           => DP_OP_751_130_5637_n1040, CI => 
                           DP_OP_751_130_5637_n1098, CO => 
                           DP_OP_751_130_5637_n999, S => 
                           DP_OP_751_130_5637_n1000);
   DP_OP_751_130_5637_U782 : FA_X1 port map( A => DP_OP_751_130_5637_n1097, B 
                           => DP_OP_751_130_5637_n1039, CI => 
                           DP_OP_751_130_5637_n1096, CO => 
                           DP_OP_751_130_5637_n997, S => 
                           DP_OP_751_130_5637_n998);
   DP_OP_751_130_5637_U781 : FA_X1 port map( A => DP_OP_751_130_5637_n1095, B 
                           => DP_OP_751_130_5637_n1038, CI => 
                           DP_OP_751_130_5637_n1094, CO => 
                           DP_OP_751_130_5637_n995, S => 
                           DP_OP_751_130_5637_n996);
   DP_OP_751_130_5637_U780 : FA_X1 port map( A => DP_OP_751_130_5637_n1093, B 
                           => DP_OP_751_130_5637_n1037, CI => 
                           DP_OP_751_130_5637_n1092, CO => 
                           DP_OP_751_130_5637_n993, S => 
                           DP_OP_751_130_5637_n994);
   DP_OP_751_130_5637_U779 : FA_X1 port map( A => DP_OP_751_130_5637_n1091, B 
                           => DP_OP_751_130_5637_n1036, CI => 
                           DP_OP_751_130_5637_n1090, CO => 
                           DP_OP_751_130_5637_n991, S => 
                           DP_OP_751_130_5637_n992);
   DP_OP_751_130_5637_U778 : FA_X1 port map( A => DP_OP_751_130_5637_n1089, B 
                           => DP_OP_751_130_5637_n1035, CI => 
                           DP_OP_751_130_5637_n1088, CO => 
                           DP_OP_751_130_5637_n989, S => 
                           DP_OP_751_130_5637_n990);
   DP_OP_751_130_5637_U776 : FA_X1 port map( A => DP_OP_751_130_5637_n1085, B 
                           => DP_OP_751_130_5637_n1033, CI => 
                           DP_OP_751_130_5637_n1084, CO => 
                           DP_OP_751_130_5637_n985, S => 
                           DP_OP_751_130_5637_n986);
   DP_OP_751_130_5637_U775 : FA_X1 port map( A => DP_OP_751_130_5637_n1083, B 
                           => DP_OP_751_130_5637_n1032, CI => 
                           DP_OP_751_130_5637_n1082, CO => 
                           DP_OP_751_130_5637_n983, S => 
                           DP_OP_751_130_5637_n984);
   DP_OP_751_130_5637_U774 : FA_X1 port map( A => DP_OP_751_130_5637_n1081, B 
                           => DP_OP_751_130_5637_n1031, CI => 
                           DP_OP_751_130_5637_n1080, CO => n_3916, S => 
                           DP_OP_751_130_5637_n982);
   DP_OP_751_130_5637_U718 : FA_X1 port map( A => DP_OP_751_130_5637_n1007, B 
                           => DP_OP_751_130_5637_n943, CI => 
                           DP_OP_751_130_5637_n1006, CO => 
                           DP_OP_751_130_5637_n907, S => 
                           DP_OP_751_130_5637_n908);
   DP_OP_751_130_5637_U717 : FA_X1 port map( A => DP_OP_751_130_5637_n1005, B 
                           => DP_OP_751_130_5637_n942, CI => 
                           DP_OP_751_130_5637_n1004, CO => 
                           DP_OP_751_130_5637_n905, S => 
                           DP_OP_751_130_5637_n906);
   DP_OP_751_130_5637_U716 : FA_X1 port map( A => DP_OP_751_130_5637_n1003, B 
                           => DP_OP_751_130_5637_n941, CI => 
                           DP_OP_751_130_5637_n1002, CO => 
                           DP_OP_751_130_5637_n903, S => 
                           DP_OP_751_130_5637_n904);
   DP_OP_751_130_5637_U715 : FA_X1 port map( A => DP_OP_751_130_5637_n1001, B 
                           => DP_OP_751_130_5637_n940, CI => 
                           DP_OP_751_130_5637_n1000, CO => 
                           DP_OP_751_130_5637_n901, S => 
                           DP_OP_751_130_5637_n902);
   DP_OP_751_130_5637_U714 : FA_X1 port map( A => DP_OP_751_130_5637_n999, B =>
                           DP_OP_751_130_5637_n939, CI => 
                           DP_OP_751_130_5637_n998, CO => 
                           DP_OP_751_130_5637_n899, S => 
                           DP_OP_751_130_5637_n900);
   DP_OP_751_130_5637_U713 : FA_X1 port map( A => DP_OP_751_130_5637_n997, B =>
                           DP_OP_751_130_5637_n938, CI => 
                           DP_OP_751_130_5637_n996, CO => 
                           DP_OP_751_130_5637_n897, S => 
                           DP_OP_751_130_5637_n898);
   DP_OP_751_130_5637_U712 : FA_X1 port map( A => DP_OP_751_130_5637_n995, B =>
                           DP_OP_751_130_5637_n937, CI => 
                           DP_OP_751_130_5637_n994, CO => 
                           DP_OP_751_130_5637_n895, S => 
                           DP_OP_751_130_5637_n896);
   DP_OP_751_130_5637_U711 : FA_X1 port map( A => DP_OP_751_130_5637_n993, B =>
                           DP_OP_751_130_5637_n936, CI => 
                           DP_OP_751_130_5637_n992, CO => 
                           DP_OP_751_130_5637_n893, S => 
                           DP_OP_751_130_5637_n894);
   DP_OP_751_130_5637_U710 : FA_X1 port map( A => DP_OP_751_130_5637_n991, B =>
                           DP_OP_751_130_5637_n935, CI => 
                           DP_OP_751_130_5637_n990, CO => 
                           DP_OP_751_130_5637_n891, S => 
                           DP_OP_751_130_5637_n892);
   DP_OP_751_130_5637_U709 : FA_X1 port map( A => DP_OP_751_130_5637_n989, B =>
                           DP_OP_751_130_5637_n934, CI => 
                           DP_OP_751_130_5637_n988, CO => 
                           DP_OP_751_130_5637_n889, S => 
                           DP_OP_751_130_5637_n890);
   DP_OP_751_130_5637_U707 : FA_X1 port map( A => DP_OP_751_130_5637_n985, B =>
                           DP_OP_751_130_5637_n932, CI => 
                           DP_OP_751_130_5637_n984, CO => 
                           DP_OP_751_130_5637_n885, S => 
                           DP_OP_751_130_5637_n886);
   DP_OP_751_130_5637_U706 : FA_X1 port map( A => DP_OP_751_130_5637_n983, B =>
                           DP_OP_751_130_5637_n931, CI => 
                           DP_OP_751_130_5637_n982, CO => n_3917, S => 
                           DP_OP_751_130_5637_n884);
   DP_OP_751_130_5637_U648 : FA_X1 port map( A => DP_OP_751_130_5637_n905, B =>
                           DP_OP_751_130_5637_n841, CI => 
                           DP_OP_751_130_5637_n904, CO => 
                           DP_OP_751_130_5637_n805, S => 
                           DP_OP_751_130_5637_n806);
   DP_OP_751_130_5637_U647 : FA_X1 port map( A => DP_OP_751_130_5637_n903, B =>
                           DP_OP_751_130_5637_n840, CI => 
                           DP_OP_751_130_5637_n902, CO => 
                           DP_OP_751_130_5637_n803, S => 
                           DP_OP_751_130_5637_n804);
   DP_OP_751_130_5637_U646 : FA_X1 port map( A => DP_OP_751_130_5637_n901, B =>
                           DP_OP_751_130_5637_n839, CI => 
                           DP_OP_751_130_5637_n900, CO => 
                           DP_OP_751_130_5637_n801, S => 
                           DP_OP_751_130_5637_n802);
   DP_OP_751_130_5637_U645 : FA_X1 port map( A => DP_OP_751_130_5637_n899, B =>
                           DP_OP_751_130_5637_n838, CI => 
                           DP_OP_751_130_5637_n898, CO => 
                           DP_OP_751_130_5637_n799, S => 
                           DP_OP_751_130_5637_n800);
   DP_OP_751_130_5637_U643 : FA_X1 port map( A => DP_OP_751_130_5637_n895, B =>
                           DP_OP_751_130_5637_n836, CI => 
                           DP_OP_751_130_5637_n894, CO => 
                           DP_OP_751_130_5637_n795, S => 
                           DP_OP_751_130_5637_n796);
   DP_OP_751_130_5637_U642 : FA_X1 port map( A => DP_OP_751_130_5637_n893, B =>
                           DP_OP_751_130_5637_n835, CI => 
                           DP_OP_751_130_5637_n892, CO => 
                           DP_OP_751_130_5637_n793, S => 
                           DP_OP_751_130_5637_n794);
   DP_OP_751_130_5637_U640 : FA_X1 port map( A => DP_OP_751_130_5637_n889, B =>
                           DP_OP_751_130_5637_n833, CI => 
                           DP_OP_751_130_5637_n888, CO => 
                           DP_OP_751_130_5637_n789, S => 
                           DP_OP_751_130_5637_n790);
   DP_OP_751_130_5637_U639 : FA_X1 port map( A => DP_OP_751_130_5637_n887, B =>
                           DP_OP_751_130_5637_n832, CI => 
                           DP_OP_751_130_5637_n886, CO => 
                           DP_OP_751_130_5637_n787, S => 
                           DP_OP_751_130_5637_n788);
   DP_OP_751_130_5637_U638 : FA_X1 port map( A => DP_OP_751_130_5637_n885, B =>
                           DP_OP_751_130_5637_n831, CI => 
                           DP_OP_751_130_5637_n884, CO => n_3918, S => 
                           DP_OP_751_130_5637_n786);
   DP_OP_751_130_5637_U578 : FA_X1 port map( A => DP_OP_751_130_5637_n803, B =>
                           DP_OP_751_130_5637_n739, CI => 
                           DP_OP_751_130_5637_n802, CO => 
                           DP_OP_751_130_5637_n703, S => 
                           DP_OP_751_130_5637_n704);
   DP_OP_751_130_5637_U577 : FA_X1 port map( A => DP_OP_751_130_5637_n801, B =>
                           DP_OP_751_130_5637_n738, CI => 
                           DP_OP_751_130_5637_n800, CO => 
                           DP_OP_751_130_5637_n701, S => 
                           DP_OP_751_130_5637_n702);
   DP_OP_751_130_5637_U576 : FA_X1 port map( A => DP_OP_751_130_5637_n799, B =>
                           DP_OP_751_130_5637_n737, CI => 
                           DP_OP_751_130_5637_n798, CO => 
                           DP_OP_751_130_5637_n699, S => 
                           DP_OP_751_130_5637_n700);
   DP_OP_751_130_5637_U575 : FA_X1 port map( A => DP_OP_751_130_5637_n797, B =>
                           DP_OP_751_130_5637_n736, CI => 
                           DP_OP_751_130_5637_n796, CO => 
                           DP_OP_751_130_5637_n697, S => 
                           DP_OP_751_130_5637_n698);
   DP_OP_751_130_5637_U574 : FA_X1 port map( A => DP_OP_751_130_5637_n795, B =>
                           DP_OP_751_130_5637_n735, CI => 
                           DP_OP_751_130_5637_n794, CO => 
                           DP_OP_751_130_5637_n695, S => 
                           DP_OP_751_130_5637_n696);
   DP_OP_751_130_5637_U573 : FA_X1 port map( A => DP_OP_751_130_5637_n793, B =>
                           DP_OP_751_130_5637_n734, CI => 
                           DP_OP_751_130_5637_n792, CO => 
                           DP_OP_751_130_5637_n693, S => 
                           DP_OP_751_130_5637_n694);
   DP_OP_751_130_5637_U570 : FA_X1 port map( A => DP_OP_751_130_5637_n787, B =>
                           DP_OP_751_130_5637_n731, CI => 
                           DP_OP_751_130_5637_n786, CO => n_3919, S => 
                           DP_OP_751_130_5637_n688);
   DP_OP_751_130_5637_U508 : FA_X1 port map( A => DP_OP_751_130_5637_n701, B =>
                           DP_OP_751_130_5637_n637, CI => 
                           DP_OP_751_130_5637_n700, CO => 
                           DP_OP_751_130_5637_n601, S => 
                           DP_OP_751_130_5637_n602);
   DP_OP_751_130_5637_U507 : FA_X1 port map( A => DP_OP_751_130_5637_n699, B =>
                           DP_OP_751_130_5637_n636, CI => 
                           DP_OP_751_130_5637_n698, CO => 
                           DP_OP_751_130_5637_n599, S => 
                           DP_OP_751_130_5637_n600);
   DP_OP_751_130_5637_U506 : FA_X1 port map( A => DP_OP_751_130_5637_n697, B =>
                           DP_OP_751_130_5637_n635, CI => 
                           DP_OP_751_130_5637_n696, CO => 
                           DP_OP_751_130_5637_n597, S => 
                           DP_OP_751_130_5637_n598);
   DP_OP_751_130_5637_U505 : FA_X1 port map( A => DP_OP_751_130_5637_n695, B =>
                           DP_OP_751_130_5637_n634, CI => 
                           DP_OP_751_130_5637_n694, CO => 
                           DP_OP_751_130_5637_n595, S => 
                           DP_OP_751_130_5637_n596);
   DP_OP_751_130_5637_U504 : FA_X1 port map( A => DP_OP_751_130_5637_n693, B =>
                           DP_OP_751_130_5637_n633, CI => 
                           DP_OP_751_130_5637_n692, CO => 
                           DP_OP_751_130_5637_n593, S => 
                           DP_OP_751_130_5637_n594);
   DP_OP_751_130_5637_U502 : FA_X1 port map( A => DP_OP_751_130_5637_n689, B =>
                           DP_OP_751_130_5637_n631, CI => 
                           DP_OP_751_130_5637_n688, CO => n_3920, S => 
                           DP_OP_751_130_5637_n590);
   DP_OP_751_130_5637_U438 : FA_X1 port map( A => DP_OP_751_130_5637_n599, B =>
                           DP_OP_751_130_5637_n535, CI => 
                           DP_OP_751_130_5637_n598, CO => 
                           DP_OP_751_130_5637_n499, S => 
                           DP_OP_751_130_5637_n500);
   DP_OP_751_130_5637_U437 : FA_X1 port map( A => DP_OP_751_130_5637_n597, B =>
                           DP_OP_751_130_5637_n534, CI => 
                           DP_OP_751_130_5637_n596, CO => 
                           DP_OP_751_130_5637_n497, S => 
                           DP_OP_751_130_5637_n498);
   DP_OP_751_130_5637_U435 : FA_X1 port map( A => DP_OP_751_130_5637_n593, B =>
                           DP_OP_751_130_5637_n532, CI => 
                           DP_OP_751_130_5637_n592, CO => 
                           DP_OP_751_130_5637_n493, S => 
                           DP_OP_751_130_5637_n494);
   DP_OP_751_130_5637_U366 : FA_X1 port map( A => DP_OP_751_130_5637_n493, B =>
                           DP_OP_751_130_5637_n431, CI => 
                           DP_OP_751_130_5637_n492, CO => n_3921, S => 
                           DP_OP_751_130_5637_n394);
   DataPath_RF_CWP_Q_reg_1_inst : DFF_X1 port map( D => n7072, CK => CLK, Q => 
                           DataPath_RF_c_win_1_port, QN => n8442);
   PC_reg_29_inst : DFFS_X2 port map( D => n8475, CK => CLK, SN => n8696, Q => 
                           n8389, QN => IRAM_ADDRESS_29_port);
   IR_reg_26_inst : DFFS_X1 port map( D => n7109, CK => CLK, SN => n8693, Q => 
                           IR_26_port, QN => n8501);
   IR_reg_30_inst : DFFS_X1 port map( D => n7105, CK => CLK, SN => n8693, Q => 
                           IR_30_port, QN => n8308);
   IR_reg_31_inst : DFFS_X1 port map( D => n8479, CK => CLK, SN => n8696, Q => 
                           n171, QN => n10771);
   IR_reg_29_inst : DFFS_X1 port map( D => n8478, CK => CLK, SN => n8696, Q => 
                           n176, QN => n10744);
   CU_I_CW_EX_reg_16_inst : DFF_X1 port map( D => n7854, CK => CLK, Q => n8684,
                           QN => i_S2);
   DataPath_RF_CWP_Q_reg_2_inst : DFF_X1 port map( D => n7071, CK => CLK, Q => 
                           DataPath_RF_c_win_2_port, QN => n_3922);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_14_inst : DFF_X1 port map( D => n7742,
                           CK => CLK, Q => n8401, QN => n866);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_13_inst : DFF_X1 port map( D => n7741,
                           CK => CLK, Q => n8426, QN => n865);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_12_inst : DFF_X1 port map( D => n7740,
                           CK => CLK, Q => n8415, QN => n864);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_11_inst : DFF_X1 port map( D => n7739,
                           CK => CLK, Q => n8425, QN => n863);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_10_inst : DFF_X1 port map( D => n7738,
                           CK => CLK, Q => n8414, QN => n862);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_9_inst : DFF_X1 port map( D => n7737, 
                           CK => CLK, Q => n8424, QN => n861);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_8_inst : DFF_X1 port map( D => n7736, 
                           CK => CLK, Q => n8423, QN => n860);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_7_inst : DFF_X1 port map( D => n7735, 
                           CK => CLK, Q => n8422, QN => n859);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_6_inst : DFF_X1 port map( D => n7734, 
                           CK => CLK, Q => n8421, QN => n858);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_5_inst : DFF_X1 port map( D => n7733, 
                           CK => CLK, Q => n8420, QN => n857);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_4_inst : DFF_X1 port map( D => n7732, 
                           CK => CLK, Q => n8419, QN => n856);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_3_inst : DFF_X1 port map( D => n7731, 
                           CK => CLK, Q => n8418, QN => n855);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_2_inst : DFF_X1 port map( D => n7730, 
                           CK => CLK, Q => n8417, QN => n854);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_1_inst : DFF_X1 port map( D => n7729, 
                           CK => CLK, Q => n8416, QN => n853);
   DataPath_WRF_CUhw_curr_addr_reg_2_inst : DFF_X1 port map( D => n7728, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_2_port, QN => 
                           n_3923);
   DataPath_WRF_CUhw_curr_addr_reg_3_inst : DFF_X1 port map( D => n7727, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_3_port, QN => 
                           n_3924);
   DataPath_WRF_CUhw_curr_addr_reg_4_inst : DFF_X1 port map( D => n7726, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_4_port, QN => 
                           n_3925);
   DataPath_WRF_CUhw_curr_addr_reg_5_inst : DFF_X1 port map( D => n7725, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_5_port, QN => 
                           n_3926);
   DataPath_WRF_CUhw_curr_addr_reg_6_inst : DFF_X1 port map( D => n7724, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_6_port, QN => 
                           n_3927);
   DataPath_WRF_CUhw_curr_addr_reg_7_inst : DFF_X1 port map( D => n7723, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_7_port, QN => 
                           n_3928);
   DataPath_WRF_CUhw_curr_addr_reg_8_inst : DFF_X1 port map( D => n7722, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_8_port, QN => 
                           n_3929);
   DataPath_WRF_CUhw_curr_addr_reg_9_inst : DFF_X1 port map( D => n7721, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_9_port, QN => 
                           n_3930);
   DataPath_WRF_CUhw_curr_addr_reg_10_inst : DFF_X1 port map( D => n7720, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_10_port, QN =>
                           n_3931);
   DataPath_WRF_CUhw_curr_addr_reg_11_inst : DFF_X1 port map( D => n7719, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_11_port, QN =>
                           n_3932);
   DataPath_WRF_CUhw_curr_addr_reg_12_inst : DFF_X1 port map( D => n7718, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_12_port, QN =>
                           n_3933);
   DataPath_WRF_CUhw_curr_addr_reg_13_inst : DFF_X1 port map( D => n7717, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_13_port, QN =>
                           n_3934);
   DataPath_WRF_CUhw_curr_addr_reg_14_inst : DFF_X1 port map( D => n7716, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_14_port, QN =>
                           n_3935);
   DataPath_WRF_CUhw_curr_addr_reg_15_inst : DFF_X1 port map( D => n7715, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_15_port, QN =>
                           n_3936);
   DataPath_WRF_CUhw_curr_addr_reg_16_inst : DFF_X1 port map( D => n7714, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_16_port, QN =>
                           n_3937);
   DataPath_WRF_CUhw_curr_addr_reg_19_inst : DFF_X1 port map( D => n7713, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_19_port, QN =>
                           n8187);
   DataPath_WRF_CUhw_curr_addr_reg_17_inst : DFF_X1 port map( D => n7712, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_17_port, QN =>
                           n_3938);
   DataPath_WRF_CUhw_curr_addr_reg_18_inst : DFF_X1 port map( D => n7711, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_18_port, QN =>
                           n_3939);
   DataPath_WRF_CUhw_curr_addr_reg_20_inst : DFF_X1 port map( D => n7710, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_20_port, QN =>
                           n_3940);
   DataPath_WRF_CUhw_curr_addr_reg_21_inst : DFF_X1 port map( D => n7709, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_21_port, QN =>
                           n_3941);
   DataPath_WRF_CUhw_curr_addr_reg_22_inst : DFF_X1 port map( D => n7708, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_22_port, QN =>
                           n_3942);
   DataPath_WRF_CUhw_curr_addr_reg_26_inst : DFF_X1 port map( D => n7707, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_26_port, QN =>
                           n_3943);
   DataPath_WRF_CUhw_curr_addr_reg_23_inst : DFF_X1 port map( D => n7706, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_23_port, QN =>
                           n_3944);
   DataPath_WRF_CUhw_curr_addr_reg_24_inst : DFF_X1 port map( D => n7705, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_24_port, QN =>
                           n_3945);
   DataPath_WRF_CUhw_curr_addr_reg_27_inst : DFF_X1 port map( D => n7704, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_27_port, QN =>
                           n_3946);
   DataPath_WRF_CUhw_curr_addr_reg_28_inst : DFF_X1 port map( D => n7703, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_28_port, QN =>
                           n8203);
   DataPath_WRF_CUhw_curr_addr_reg_25_inst : DFF_X1 port map( D => n7702, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_25_port, QN =>
                           n8229);
   IR_reg_0_inst : DFFR_X1 port map( D => n48, CK => CLK, RN => n8691, Q => 
                           n8427, QN => n210);
   IR_reg_2_inst : DFFR_X1 port map( D => n50, CK => CLK, RN => n8689, Q => 
                           IR_2_port, QN => n8428);
   IR_reg_14_inst : DFFR_X1 port map( D => n7121, CK => CLK, RN => n8688, Q => 
                           n8391, QN => n195);
   IR_reg_12_inst : DFFR_X1 port map( D => n57, CK => CLK, RN => n8694, Q => 
                           n8306, QN => n196);
   IR_reg_24_inst : DFFR_X1 port map( D => n7111, CK => CLK, RN => n8690, Q => 
                           n8305, QN => n185);
   IR_reg_4_inst : DFFR_X1 port map( D => n52, CK => CLK, RN => n8691, Q => 
                           IR_4_port, QN => n8317);
   IR_reg_1_inst : DFFR_X1 port map( D => n49, CK => CLK, RN => n8689, Q => 
                           IR_1_port, QN => n8315);
   IR_reg_9_inst : DFFR_X1 port map( D => n7122, CK => CLK, RN => n8688, Q => 
                           IR_9_port, QN => n8407);
   IR_reg_7_inst : DFFR_X1 port map( D => n55, CK => CLK, RN => n8690, Q => 
                           IR_7_port, QN => n8332);
   IR_reg_6_inst : DFFR_X1 port map( D => n54, CK => CLK, RN => n8691, Q => 
                           IR_6_port, QN => n8307);
   IR_reg_5_inst : DFFR_X1 port map( D => n53, CK => CLK, RN => n8689, Q => 
                           IR_5_port, QN => n8320);
   IR_reg_3_inst : DFFR_X1 port map( D => n51, CK => CLK, RN => n8688, Q => 
                           IR_3_port, QN => n8318);
   IR_reg_27_inst : DFFR_X1 port map( D => n7108, CK => CLK, RN => n8690, Q => 
                           n8312, QN => n8502);
   IR_reg_15_inst : DFFR_X1 port map( D => n7120, CK => CLK, RN => n8690, Q => 
                           n8304, QN => n194);
   IR_reg_11_inst : DFFR_X1 port map( D => n56, CK => CLK, RN => n8691, Q => 
                           n8302, QN => n197);
   IR_reg_25_inst : DFFR_X1 port map( D => n7110, CK => CLK, RN => n8689, Q => 
                           n8399, QN => n184);
   IR_reg_23_inst : DFFR_X1 port map( D => n7112, CK => CLK, RN => n8688, Q => 
                           n8397, QN => n186);
   IR_reg_22_inst : DFFR_X1 port map( D => n7113, CK => CLK, RN => n8690, Q => 
                           n8396, QN => n187);
   IR_reg_21_inst : DFFR_X1 port map( D => n7114, CK => CLK, RN => n8691, Q => 
                           n8395, QN => n188);
   PC_reg_6_inst : DFFR_X1 port map( D => n7053, CK => CLK, RN => n8689, Q => 
                           IRAM_ADDRESS_6_port, QN => n8366);
   PC_reg_3_inst : DFFR_X1 port map( D => n7056, CK => CLK, RN => n8690, Q => 
                           IRAM_ADDRESS_3_port, QN => n8326);
   PC_reg_4_inst : DFFR_X1 port map( D => n7055, CK => CLK, RN => n8691, Q => 
                           IRAM_ADDRESS_4_port, QN => n8325);
   PC_reg_2_inst : DFFR_X1 port map( D => n7057, CK => CLK, RN => n8689, Q => 
                           IRAM_ADDRESS_2_port, QN => intadd_1_A_1_port);
   PC_reg_1_inst : DFFR_X1 port map( D => n7058, CK => CLK, RN => n8690, Q => 
                           IRAM_ADDRESS_1_port, QN => intadd_1_A_0_port);
   PC_reg_5_inst : DFFR_X1 port map( D => n7054, CK => CLK, RN => n8691, Q => 
                           IRAM_ADDRESS_5_port, QN => n226);
   PC_reg_0_inst : DFFR_X1 port map( D => n7059, CK => CLK, RN => n8689, Q => 
                           IRAM_ADDRESS_0_port, QN => n230);
   PC_reg_9_inst : DFFR_X1 port map( D => n7050, CK => CLK, RN => n8691, Q => 
                           IRAM_ADDRESS_9_port, QN => n224);
   PC_reg_10_inst : DFFR_X1 port map( D => n7049, CK => CLK, RN => n8690, Q => 
                           IRAM_ADDRESS_10_port, QN => n8429);
   PC_reg_11_inst : DFFR_X1 port map( D => n7048, CK => CLK, RN => n8689, Q => 
                           IRAM_ADDRESS_11_port, QN => n8383);
   PC_reg_12_inst : DFFR_X1 port map( D => n7047, CK => CLK, RN => n8690, Q => 
                           IRAM_ADDRESS_12_port, QN => n222);
   PC_reg_13_inst : DFFR_X1 port map( D => n7046, CK => CLK, RN => n8691, Q => 
                           IRAM_ADDRESS_13_port, QN => n8398);
   PC_reg_14_inst : DFFR_X1 port map( D => n7045, CK => CLK, RN => n8689, Q => 
                           IRAM_ADDRESS_14_port, QN => n8384);
   PC_reg_15_inst : DFFR_X1 port map( D => n7044, CK => CLK, RN => n8691, Q => 
                           IRAM_ADDRESS_15_port, QN => n8381);
   PC_reg_16_inst : DFFR_X1 port map( D => n7043, CK => CLK, RN => n8690, Q => 
                           IRAM_ADDRESS_16_port, QN => n220);
   PC_reg_28_inst : DFFR_X1 port map( D => n7031, CK => CLK, RN => n8689, Q => 
                           IRAM_ADDRESS_28_port, QN => n8156);
   PC_reg_20_inst : DFFR_X1 port map( D => n7039, CK => CLK, RN => n8690, Q => 
                           IRAM_ADDRESS_20_port, QN => intadd_0_A_0_port);
   PC_reg_22_inst : DFFR_X1 port map( D => n7037, CK => CLK, RN => n8691, Q => 
                           IRAM_ADDRESS_22_port, QN => n8390);
   PC_reg_21_inst : DFFR_X1 port map( D => n7038, CK => CLK, RN => n8691, Q => 
                           IRAM_ADDRESS_21_port, QN => n8387);
   PC_reg_19_inst : DFFR_X1 port map( D => n7040, CK => CLK, RN => n8690, Q => 
                           IRAM_ADDRESS_19_port, QN => n8392);
   PC_reg_24_inst : DFFR_X1 port map( D => n7035, CK => CLK, RN => n8690, Q => 
                           IRAM_ADDRESS_24_port, QN => n8377);
   PC_reg_23_inst : DFFR_X1 port map( D => n7036, CK => CLK, RN => n8691, Q => 
                           IRAM_ADDRESS_23_port, QN => n8394);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_2_inst : DFF_X1 port map( D => 
                           n11974, CK => CLK, Q => n_3947, QN => 
                           DECODEhw_i_tickcounter_2_port);
   DataPath_RF_SWP_Q_reg_4_inst : DFF_X2 port map( D => n7062, CK => CLK, Q => 
                           DataPath_RF_c_swin_4_port, QN => n824);
   CU_I_CW_MEM_reg_5_inst : DFF_X2 port map( D => n385, CK => CLK, Q => 
                           i_DATAMEM_RM, QN => n_3948);
   CU_I_aluOpcode1_reg_2_inst : DFF_X2 port map( D => n7085, CK => CLK, Q => 
                           i_ALU_OP_2_port, QN => n8300);
   DataPath_RF_CWP_Q_reg_3_inst : DFF_X2 port map( D => n7070, CK => CLK, Q => 
                           DataPath_RF_c_win_3_port, QN => n577);
   DataPath_WRF_CUhw_curr_addr_reg_31_inst : DFF_X1 port map( D => n8480, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_31_port, QN =>
                           n_3949);
   U7526 : OAI33_X1 port map( A1 => n7652, A2 => DataPath_i_LGET_0_port, A3 => 
                           n7650, B1 => n7651, B2 => n494, B3 => n235, ZN => 
                           n7653);
   U7527 : AND2_X1 port map( A1 => n8457, A2 => n8122, ZN => n7688);
   U7528 : NAND2_X1 port map( A1 => n476, A2 => n477, ZN => n10730);
   U7529 : OR2_X1 port map( A1 => n10580, A2 => n8155, ZN => n10576);
   U7530 : INV_X1 port map( A => n10044, ZN => n7769);
   U7531 : INV_X1 port map( A => n10223, ZN => n7767);
   U7532 : BUF_X1 port map( A => n10492, Z => n8578);
   U7533 : AND2_X1 port map( A1 => n10702, A2 => n10577, ZN => n8303);
   U7534 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n22, B => n8019, ZN =>
                           C620_DATA2_11);
   U7535 : INV_X1 port map( A => n7745, ZN => DP_OP_1090J1_126_7243_n18);
   U7536 : CLKBUF_X3 port map( A => n8505, Z => n7757);
   U7537 : OAI21_X1 port map( B1 => n10144, B2 => n10124, A => n9499, ZN => 
                           n9500);
   U7538 : AND4_X1 port map( A1 => n9189, A2 => n9190, A3 => n9198, A4 => n9195
                           , ZN => n7744);
   U7539 : BUF_X2 port map( A => n9207, Z => n7698);
   U7540 : INV_X1 port map( A => n7744, ZN => n9191);
   U7541 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_7_port, B => 
                           n8263, ZN => n7174);
   U7542 : OAI22_X1 port map( A1 => n7754, A2 => n7787, B1 => n9659, B2 => 
                           n7796, ZN => n7175);
   U7543 : XOR2_X1 port map( A => n8264, B => n7175, Z => n7176);
   U7544 : XOR2_X1 port map( A => n7174, B => n7176, Z => 
                           DP_OP_751_130_5637_n1716);
   U7545 : NOR2_X1 port map( A1 => n7174, A2 => n7176, ZN => 
                           DP_OP_751_130_5637_n1715);
   U7546 : OAI22_X1 port map( A1 => n8299, A2 => n11838, B1 => n8441, B2 => 
                           n11839, ZN => n7177);
   U7547 : AOI211_X1 port map( C1 => n8964, C2 => n8971, A => RST, B => n7177, 
                           ZN => n11841);
   U7548 : AOI22_X1 port map( A1 => n10231, A2 => n10091, B1 => n10089, B2 => 
                           n9767, ZN => n7178);
   U7549 : AOI22_X1 port map( A1 => n10086, A2 => n10232, B1 => n7781, B2 => 
                           n9820, ZN => n7179);
   U7550 : INV_X1 port map( A => n9771, ZN => n7180);
   U7551 : AOI22_X1 port map( A1 => n9816, A2 => n9748, B1 => n10090, B2 => 
                           n7180, ZN => n7181);
   U7552 : NAND3_X1 port map( A1 => n7178, A2 => n7179, A3 => n7181, ZN => 
                           n9829);
   U7553 : INV_X1 port map( A => n8552, ZN => n7182);
   U7554 : OAI21_X1 port map( B1 => n9411, B2 => n7182, A => n9889, ZN => n9575
                           );
   U7555 : NAND2_X1 port map( A1 => n8277, A2 => DP_OP_751_130_5637_n139, ZN =>
                           n7183);
   U7556 : XNOR2_X1 port map( A => n7183, B => DP_OP_751_130_5637_n140, ZN => 
                           n7184);
   U7557 : INV_X1 port map( A => n10368, ZN => n7185);
   U7558 : INV_X1 port map( A => n10370, ZN => n7186);
   U7559 : AOI221_X1 port map( B1 => n10368, B2 => n10370, C1 => n7185, C2 => 
                           n7186, A => n10381, ZN => n7187);
   U7560 : INV_X1 port map( A => n10377, ZN => n7188);
   U7561 : AOI22_X1 port map( A1 => n10377, A2 => n10468, B1 => n10469, B2 => 
                           n7188, ZN => n7189);
   U7562 : XOR2_X1 port map( A => n10370, B => n10369, Z => n7190);
   U7563 : OAI22_X1 port map( A1 => n10432, A2 => n10376, B1 => n10374, B2 => 
                           n10505, ZN => n7191);
   U7564 : AOI21_X1 port map( B1 => n10440, B2 => n10493, A => n7191, ZN => 
                           n7192);
   U7565 : OAI22_X1 port map( A1 => n10371, A2 => n10460, B1 => n10443, B2 => 
                           n10442, ZN => n7193);
   U7566 : OAI22_X1 port map( A1 => n10372, A2 => n10507, B1 => n10373, B2 => 
                           n10388, ZN => n7194);
   U7567 : AOI211_X1 port map( C1 => n10495, C2 => n10402, A => n7193, B => 
                           n7194, ZN => n7195);
   U7568 : OAI211_X1 port map( C1 => n10375, C2 => n10479, A => n7192, B => 
                           n7195, ZN => n7196);
   U7569 : INV_X1 port map( A => n10452, ZN => n7197);
   U7570 : AOI22_X1 port map( A1 => n7190, A2 => n10380, B1 => n7196, B2 => 
                           n7197, ZN => n7198);
   U7571 : INV_X1 port map( A => n7789, ZN => n7199);
   U7572 : OAI221_X1 port map( B1 => n7789, B2 => n10458, C1 => n7199, C2 => 
                           n10468, A => n10379, ZN => n7200);
   U7573 : OAI211_X1 port map( C1 => n7189, C2 => n10379, A => n7198, B => 
                           n7200, ZN => n7201);
   U7574 : AOI211_X1 port map( C1 => n8578, C2 => n7184, A => n7187, B => n7201
                           , ZN => n7202);
   U7575 : OAI22_X1 port map( A1 => n503, A2 => n12092, B1 => n12093, B2 => 
                           n7202, ZN => n7009);
   U7576 : AND2_X1 port map( A1 => n8695, A2 => 
                           DataPath_RF_internal_out1_22_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N26);
   U7577 : AND2_X1 port map( A1 => n8694, A2 => 
                           DataPath_RF_internal_out2_21_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N25);
   U7578 : OAI22_X1 port map( A1 => n8441, A2 => n11847, B1 => n577, B2 => 
                           n11848, ZN => n7203);
   U7579 : AOI211_X1 port map( C1 => n8967, C2 => n8771, A => RST, B => n7203, 
                           ZN => n11410);
   U7580 : OAI22_X1 port map( A1 => n9452, A2 => n9560, B1 => n10511, B2 => 
                           n8562, ZN => n7204);
   U7581 : XNOR2_X1 port map( A => n8263, B => n7204, ZN => n7205);
   U7582 : OAI22_X1 port map( A1 => n7755, A2 => n9721, B1 => n7796, B2 => 
                           n8496, ZN => n7206);
   U7583 : XOR2_X1 port map( A => n8264, B => n7206, Z => n7207);
   U7584 : NOR2_X1 port map( A1 => n7205, A2 => n7207, ZN => 
                           DP_OP_751_130_5637_n1721);
   U7585 : XOR2_X1 port map( A => n7205, B => n7207, Z => 
                           DP_OP_751_130_5637_n1722);
   U7586 : AOI22_X1 port map( A1 => n8681, A2 => n7772, B1 => n7800, B2 => 
                           n10445, ZN => n7208);
   U7587 : INV_X1 port map( A => n7208, ZN => n9987);
   U7588 : INV_X1 port map( A => n9918, ZN => n7209);
   U7589 : OAI21_X1 port map( B1 => n10197, B2 => n9411, A => n7209, ZN => 
                           n9542);
   U7590 : NAND3_X1 port map( A1 => n9816, A2 => DP_OP_751_130_5637_n435, A3 =>
                           n10458, ZN => n7210);
   U7591 : NAND3_X1 port map( A1 => n9817, A2 => n10469, A3 => n9815, ZN => 
                           n7211);
   U7592 : INV_X1 port map( A => n9854, ZN => n7212);
   U7593 : OAI221_X1 port map( B1 => n9813, B2 => n9856, C1 => n9813, C2 => 
                           n9814, A => n7212, ZN => n7213);
   U7594 : AOI21_X1 port map( B1 => n9814, B2 => n9855, A => n9842, ZN => n7214
                           );
   U7595 : OAI21_X1 port map( B1 => n9814, B2 => n9855, A => n7214, ZN => n7215
                           );
   U7596 : NAND4_X1 port map( A1 => n7210, A2 => n7211, A3 => n7213, A4 => 
                           n7215, ZN => n7949);
   U7597 : AOI22_X1 port map( A1 => n10439, A2 => n10495, B1 => n10461, B2 => 
                           n10389, ZN => n7216);
   U7598 : AOI22_X1 port map( A1 => n10440, A2 => n10502, B1 => n10476, B2 => 
                           n10387, ZN => n7217);
   U7599 : AOI22_X1 port map( A1 => n10475, A2 => n10503, B1 => n10498, B2 => 
                           n10428, ZN => n7218);
   U7600 : OAI211_X1 port map( C1 => n10441, C2 => n10388, A => n7217, B => 
                           n7218, ZN => n7219);
   U7601 : AOI21_X1 port map( B1 => n10499, B2 => n10427, A => n7219, ZN => 
                           n7220);
   U7602 : OAI211_X1 port map( C1 => n10481, C2 => n10444, A => n7216, B => 
                           n7220, ZN => n7221);
   U7603 : INV_X1 port map( A => DP_OP_751_130_5637_n149, ZN => n7222);
   U7604 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n150, A2 => n7222, ZN =>
                           n7223);
   U7605 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n151, B2 => n7223, A => 
                           n8578, ZN => n7224);
   U7606 : AOI21_X1 port map( B1 => DP_OP_751_130_5637_n151, B2 => n7223, A => 
                           n7224, ZN => n7225);
   U7607 : XNOR2_X1 port map( A => n8090, B => n10384, ZN => n7226);
   U7608 : XNOR2_X1 port map( A => n7226, B => n10383, ZN => n7227);
   U7609 : NOR2_X1 port map( A1 => n8090, A2 => DP_OP_751_130_5637_n1353, ZN =>
                           n7228);
   U7610 : AOI22_X1 port map( A1 => n8090, A2 => DP_OP_751_130_5637_n1353, B1 
                           => n7228, B2 => n10488, ZN => n7229);
   U7611 : OAI21_X1 port map( B1 => n7228, B2 => n10468, A => n7229, ZN => 
                           n7230);
   U7612 : OR3_X1 port map( A1 => n8677, A2 => n10489, A3 => n10386, ZN => 
                           n7231);
   U7613 : OAI211_X1 port map( C1 => n10421, C2 => n7227, A => n7230, B => 
                           n7231, ZN => n7232);
   U7614 : AOI211_X1 port map( C1 => n10390, C2 => n7221, A => n7225, B => 
                           n7232, ZN => n7233);
   U7615 : OAI22_X1 port map( A1 => n501, A2 => n12092, B1 => n12093, B2 => 
                           n7233, ZN => n7012);
   U7616 : AND2_X1 port map( A1 => n8692, A2 => 
                           DataPath_RF_internal_out1_13_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N17);
   U7617 : AND2_X1 port map( A1 => n8694, A2 => 
                           DataPath_RF_internal_out2_20_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N24);
   U7618 : OAI22_X1 port map( A1 => n7754, A2 => n9874, B1 => n7796, B2 => 
                           n10114, ZN => n7234);
   U7619 : XNOR2_X1 port map( A => n7979, B => n7234, ZN => n8175);
   U7620 : OAI22_X1 port map( A1 => n11848, A2 => n11596, B1 => n577, B2 => 
                           n11847, ZN => n7235);
   U7621 : AOI211_X1 port map( C1 => n8967, C2 => n8803, A => RST, B => n7235, 
                           ZN => n11475);
   U7622 : AOI211_X1 port map( C1 => n9603, C2 => n12089, A => n9375, B => 
                           n12072, ZN => n9798);
   U7623 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_B_3_port, A2 => n8684, B1
                           => DataPath_i_PIPLIN_IN2_3_port, B2 => i_S2, ZN => 
                           n7236);
   U7624 : INV_X1 port map( A => n7236, ZN => DP_OP_751_130_5637_n1761);
   U7625 : NAND2_X1 port map( A1 => n8011, A2 => DP_OP_751_130_5637_n1557, ZN 
                           => n7237);
   U7626 : NAND2_X1 port map( A1 => n10465, A2 => n7237, ZN => n7238);
   U7627 : OAI221_X1 port map( B1 => n7237, B2 => n10458, C1 => n8011, C2 => 
                           DP_OP_751_130_5637_n1557, A => n7238, ZN => n7239);
   U7628 : INV_X1 port map( A => n10839, ZN => n7240);
   U7629 : XNOR2_X1 port map( A => n9658, B => n8011, ZN => n7241);
   U7630 : OAI21_X1 port map( B1 => n7240, B2 => n12083, A => n9653, ZN => 
                           n7242);
   U7631 : XOR2_X1 port map( A => n7242, B => n7241, Z => n7243);
   U7632 : NAND2_X1 port map( A1 => n8280, A2 => DP_OP_751_130_5637_n169, ZN =>
                           n7244);
   U7633 : XNOR2_X1 port map( A => n7244, B => DP_OP_751_130_5637_n170, ZN => 
                           n7245);
   U7634 : AOI22_X1 port map( A1 => n10837, A2 => n7243, B1 => n8578, B2 => 
                           n7245, ZN => n7246);
   U7635 : NAND3_X1 port map( A1 => n415, A2 => n10469, A3 => n9659, ZN => 
                           n7247);
   U7636 : AOI21_X1 port map( B1 => n9657, B2 => n7241, A => n12084, ZN => 
                           n7248);
   U7637 : OAI21_X1 port map( B1 => n9657, B2 => n7241, A => n7248, ZN => n7249
                           );
   U7638 : NAND4_X1 port map( A1 => n7239, A2 => n7246, A3 => n7247, A4 => 
                           n7249, ZN => n7250);
   U7639 : OAI22_X1 port map( A1 => n10506, A2 => n10442, B1 => n10508, B2 => 
                           n10462, ZN => n7251);
   U7640 : OAI22_X1 port map( A1 => n10431, A2 => n10388, B1 => n10443, B2 => 
                           n10507, ZN => n7252);
   U7641 : AOI211_X1 port map( C1 => n10493, C2 => n10500, A => n7251, B => 
                           n7252, ZN => n7253);
   U7642 : AOI22_X1 port map( A1 => n10474, A2 => n10502, B1 => n10461, B2 => 
                           n10440, ZN => n7254);
   U7643 : AOI22_X1 port map( A1 => n10439, A2 => n10499, B1 => n10498, B2 => 
                           n10403, ZN => n7255);
   U7644 : NAND3_X1 port map( A1 => n7253, A2 => n7254, A3 => n7255, ZN => 
                           n7256);
   U7645 : AOI222_X1 port map( A1 => n7250, A2 => n10841, B1 => n7782, B2 => 
                           DRAM_ADDRESS_7_port, C1 => n7256, C2 => n10840, ZN 
                           => n2106);
   U7646 : AND2_X1 port map( A1 => n8695, A2 => 
                           DataPath_RF_internal_out1_20_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N24);
   U7647 : AND2_X1 port map( A1 => n8694, A2 => 
                           DataPath_RF_internal_out2_13_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N17);
   U7648 : OAI22_X1 port map( A1 => n8485, A2 => n8491, B1 => n8563, B2 => 
                           n9560, ZN => n7257);
   U7649 : XNOR2_X1 port map( A => n8263, B => n7257, ZN => n7258);
   U7650 : OAI22_X1 port map( A1 => n7755, A2 => n10466, B1 => n7796, B2 => 
                           n10457, ZN => n7259);
   U7651 : XOR2_X1 port map( A => n8264, B => n7259, Z => n7260);
   U7652 : XOR2_X1 port map( A => n7258, B => n7260, Z => 
                           DP_OP_751_130_5637_n1720);
   U7653 : NOR2_X1 port map( A1 => n7258, A2 => n7260, ZN => 
                           DP_OP_751_130_5637_n1719);
   U7654 : OAI22_X1 port map( A1 => n11596, A2 => n11847, B1 => n8442, B2 => 
                           n11848, ZN => n7261);
   U7655 : AOI211_X1 port map( C1 => n8967, C2 => n8852, A => RST, B => n7261, 
                           ZN => n11593);
   U7656 : OAI21_X1 port map( B1 => n10021, B2 => n9780, A => n9714, ZN => 
                           n9748);
   U7657 : NOR2_X1 port map( A1 => n7786, A2 => n8489, ZN => n7262);
   U7658 : XOR2_X1 port map( A => DP_OP_751_130_5637_n1723, B => n7262, Z => 
                           DP_OP_751_130_5637_n1624);
   U7659 : NOR2_X1 port map( A1 => n7786, A2 => n8489, ZN => n7263);
   U7660 : MUX2_X1 port map( A => n8262, B => DP_OP_751_130_5637_n1723, S => 
                           n7263, Z => DP_OP_751_130_5637_n1623);
   U7661 : AOI21_X1 port map( B1 => n368, B2 => i_ALU_OP_2_port, A => n10182, 
                           ZN => n9433);
   U7662 : INV_X1 port map( A => n10445, ZN => n7264);
   U7663 : AOI22_X1 port map( A1 => n10445, A2 => n10489, B1 => n10465, B2 => 
                           n7264, ZN => n7265);
   U7664 : INV_X1 port map( A => n8559, ZN => n7266);
   U7665 : AOI221_X1 port map( B1 => n10488, B2 => n8559, C1 => n10465, C2 => 
                           n7266, A => n10446, ZN => n7267);
   U7666 : AOI22_X1 port map( A1 => n10440, A2 => n10499, B1 => n10510, B2 => 
                           n10439, ZN => n7268);
   U7667 : AOI22_X1 port map( A1 => n10498, A2 => n10475, B1 => n10474, B2 => 
                           n10495, ZN => n7269);
   U7668 : OAI211_X1 port map( C1 => n10441, C2 => n10507, A => n7268, B => 
                           n7269, ZN => n7270);
   U7669 : OAI22_X1 port map( A1 => n10443, A2 => n10505, B1 => n10508, B2 => 
                           n10442, ZN => n7271);
   U7670 : OAI22_X1 port map( A1 => n10481, A2 => n10479, B1 => n10506, B2 => 
                           n10444, ZN => n7272);
   U7671 : NOR3_X1 port map( A1 => n7270, A2 => n7271, A3 => n7272, ZN => n7273
                           );
   U7672 : INV_X1 port map( A => DP_OP_751_130_5637_n163, ZN => n7274);
   U7673 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n164, A2 => n7274, ZN =>
                           n7275);
   U7674 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n165, A2 => n7275, ZN =>
                           n7276);
   U7675 : OAI211_X1 port map( C1 => DP_OP_751_130_5637_n165, C2 => n7275, A =>
                           n8578, B => n7276, ZN => n7277);
   U7676 : XNOR2_X1 port map( A => n10447, B => n8559, ZN => n7278);
   U7677 : INV_X1 port map( A => n10448, ZN => n7279);
   U7678 : OAI21_X1 port map( B1 => n10449, B2 => n7279, A => n10451, ZN => 
                           n7280);
   U7679 : OAI211_X1 port map( C1 => n10451, C2 => n7278, A => n10450, B => 
                           n7280, ZN => n7281);
   U7680 : OAI211_X1 port map( C1 => n7273, C2 => n10452, A => n7277, B => 
                           n7281, ZN => n7282);
   U7681 : AOI211_X1 port map( C1 => n7265, C2 => n10446, A => n7267, B => 
                           n7282, ZN => n7283);
   U7682 : OAI22_X1 port map( A1 => n12093, A2 => n7283, B1 => n499, B2 => 
                           n12092, ZN => n7015);
   U7683 : AND2_X1 port map( A1 => n8695, A2 => 
                           DataPath_RF_internal_out1_9_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N13);
   U7684 : AND2_X1 port map( A1 => n8694, A2 => 
                           DataPath_RF_internal_out2_11_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N15);
   U7685 : OAI22_X1 port map( A1 => n8299, A2 => n11848, B1 => n8442, B2 => 
                           n11847, ZN => n7284);
   U7686 : AOI211_X1 port map( C1 => n8967, C2 => n8901, A => RST, B => n7284, 
                           ZN => n11713);
   U7687 : OAI22_X1 port map( A1 => n7754, A2 => n9560, B1 => n7796, B2 => 
                           n9721, ZN => n7285);
   U7688 : XNOR2_X1 port map( A => n8264, B => n7285, ZN => n7286);
   U7689 : AND2_X1 port map( A1 => n7286, A2 => DP_OP_751_130_5637_n1727, ZN =>
                           DP_OP_751_130_5637_n1723);
   U7690 : XOR2_X1 port map( A => n7286, B => DP_OP_751_130_5637_n1727, Z => 
                           DP_OP_751_130_5637_n1724);
   U7691 : NOR2_X1 port map( A1 => n9798, A2 => n9714, ZN => n7287);
   U7692 : OAI22_X1 port map( A1 => n10059, A2 => n9379, B1 => n9434, B2 => 
                           n10057, ZN => n7288);
   U7693 : AOI211_X1 port map( C1 => n10288, C2 => n9605, A => n7287, B => 
                           n7288, ZN => n7289);
   U7694 : AOI22_X1 port map( A1 => n9603, A2 => n9374, B1 => n7785, B2 => 
                           n9602, ZN => n7290);
   U7695 : OAI211_X1 port map( C1 => n9761, C2 => n9419, A => n7289, B => n7290
                           , ZN => n10509);
   U7696 : AND2_X1 port map( A1 => n8697, A2 => 
                           DataPath_RF_internal_out1_11_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N15);
   U7697 : AND2_X1 port map( A1 => n8694, A2 => 
                           DataPath_RF_internal_out2_9_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N13);
   U7698 : OAI22_X1 port map( A1 => n7755, A2 => n10457, B1 => n7796, B2 => 
                           n8490, ZN => n7291);
   U7699 : XOR2_X1 port map( A => n8264, B => n7291, Z => n7292);
   U7700 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_6_port, B => 
                           n8263, ZN => n7293);
   U7701 : NOR2_X1 port map( A1 => n7292, A2 => n7293, ZN => 
                           DP_OP_751_130_5637_n1717);
   U7702 : XOR2_X1 port map( A => n7292, B => n7293, Z => 
                           DP_OP_751_130_5637_n1718);
   U7703 : OAI22_X1 port map( A1 => n8299, A2 => n11847, B1 => n8441, B2 => 
                           n11848, ZN => n7294);
   U7704 : AOI211_X1 port map( C1 => n8967, C2 => n8544, A => RST, B => n7294, 
                           ZN => n11850);
   U7705 : OAI21_X1 port map( B1 => n9603, B2 => n8681, A => n9604, ZN => n9797
                           );
   U7706 : NOR2_X1 port map( A1 => n12087, A2 => n9917, ZN => n7295);
   U7707 : AOI211_X1 port map( C1 => n10286, C2 => n10185, A => n10182, B => 
                           n7295, ZN => n7296);
   U7708 : AOI21_X1 port map( B1 => n9918, B2 => n10231, A => n7296, ZN => 
                           n7297);
   U7709 : AOI22_X1 port map( A1 => n9919, A2 => n9920, B1 => n7885, B2 => 
                           n9983, ZN => n7298);
   U7710 : NAND2_X1 port map( A1 => n9922, A2 => n7785, ZN => n7299);
   U7711 : OAI211_X1 port map( C1 => n10286, C2 => n10190, A => n10113, B => 
                           n10188, ZN => n7300);
   U7712 : NAND4_X1 port map( A1 => n7297, A2 => n7298, A3 => n7299, A4 => 
                           n7300, ZN => n10158);
   U7713 : INV_X1 port map( A => n8493, ZN => n7301);
   U7714 : NOR2_X1 port map( A1 => n9670, A2 => n7301, ZN => n10343);
   U7715 : NAND2_X1 port map( A1 => n8282, A2 => DP_OP_751_130_5637_n177, ZN =>
                           n7302);
   U7716 : XNOR2_X1 port map( A => n7302, B => DP_OP_751_130_5637_n178, ZN => 
                           n7303);
   U7717 : NAND3_X1 port map( A1 => n8676, A2 => n10469, A3 => n10457, ZN => 
                           n7304);
   U7718 : NAND3_X1 port map( A1 => n10458, A2 => DP_OP_751_130_5637_n1659, A3 
                           => n7818, ZN => n7305);
   U7719 : INV_X1 port map( A => n10456, ZN => n7306);
   U7720 : INV_X1 port map( A => n10454, ZN => n7307);
   U7721 : OAI211_X1 port map( C1 => n7306, C2 => n7307, A => n10471, B => 
                           n10455, ZN => n7308);
   U7722 : INV_X1 port map( A => n10472, ZN => n7309);
   U7723 : OAI221_X1 port map( B1 => n10456, B2 => n7309, C1 => n7306, C2 => 
                           n10472, A => n10837, ZN => n7310);
   U7724 : NAND4_X1 port map( A1 => n7304, A2 => n7305, A3 => n7308, A4 => 
                           n7310, ZN => n7311);
   U7725 : AOI21_X1 port map( B1 => n7303, B2 => n8578, A => n7311, ZN => n7312
                           );
   U7726 : OAI22_X1 port map( A1 => n10459, A2 => n10507, B1 => n10481, B2 => 
                           n10460, ZN => n7313);
   U7727 : AOI22_X1 port map( A1 => n10510, A2 => n10474, B1 => n10475, B2 => 
                           n10461, ZN => n7314);
   U7728 : OAI21_X1 port map( B1 => n10480, B2 => n10462, A => n7314, ZN => 
                           n7315);
   U7729 : AOI211_X1 port map( C1 => n10509, C2 => n10503, A => n7313, B => 
                           n7315, ZN => n7316);
   U7730 : AOI22_X1 port map( A1 => n10502, A2 => n10477, B1 => n10498, B2 => 
                           n10478, ZN => n7317);
   U7731 : NAND2_X1 port map( A1 => n10493, A2 => n10497, ZN => n7318);
   U7732 : NAND3_X1 port map( A1 => n7318, A2 => n7316, A3 => n7317, ZN => 
                           n7319);
   U7733 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1659, B => n7818, ZN => 
                           n7320);
   U7734 : OAI22_X1 port map( A1 => n10512, A2 => n7320, B1 => n8434, B2 => 
                           n12092, ZN => n7321);
   U7735 : AOI21_X1 port map( B1 => n10840, B2 => n7319, A => n7321, ZN => 
                           n7322);
   U7736 : OAI21_X1 port map( B1 => n10513, B2 => n7312, A => n7322, ZN => 
                           n7017);
   U7737 : AND2_X1 port map( A1 => n8695, A2 => 
                           DataPath_RF_internal_out1_7_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N11);
   U7738 : AND2_X1 port map( A1 => n8694, A2 => 
                           DataPath_RF_internal_out2_8_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N12);
   U7739 : OAI22_X1 port map( A1 => n8441, A2 => n11851, B1 => n577, B2 => 
                           n11852, ZN => n7323);
   U7740 : AOI211_X1 port map( C1 => n8969, C2 => n7762, A => RST, B => n7323, 
                           ZN => n11412);
   U7741 : OAI22_X1 port map( A1 => n7796, A2 => n9560, B1 => n7755, B2 => 
                           n10511, ZN => n7324);
   U7742 : XNOR2_X1 port map( A => n8264, B => n7324, ZN => 
                           DP_OP_751_130_5637_n1792);
   U7743 : INV_X1 port map( A => n9951, ZN => n7325);
   U7744 : AOI22_X1 port map( A1 => n7767, A2 => n9983, B1 => n10229, B2 => 
                           n7325, ZN => n7326);
   U7745 : NOR2_X1 port map( A1 => n9953, A2 => n10286, ZN => n7327);
   U7746 : AOI211_X1 port map( C1 => n9952, C2 => n12087, A => n10182, B => 
                           n7327, ZN => n7328);
   U7747 : AOI21_X1 port map( B1 => n9954, B2 => n10231, A => n7328, ZN => 
                           n7329);
   U7748 : AOI22_X1 port map( A1 => n9955, A2 => n7785, B1 => n9950, B2 => 
                           n10113, ZN => n7330);
   U7749 : NAND3_X1 port map( A1 => n7326, A2 => n7329, A3 => n7330, ZN => 
                           n10227);
   U7750 : INV_X1 port map( A => n10416, ZN => n7331);
   U7751 : NOR2_X1 port map( A1 => n10416, A2 => n10423, ZN => n7332);
   U7752 : OAI22_X1 port map( A1 => n10415, A2 => n7332, B1 => n9664, B2 => 
                           n7331, ZN => n10384);
   U7753 : INV_X1 port map( A => n7787, ZN => n7333);
   U7754 : AOI221_X1 port map( B1 => n10488, B2 => n7787, C1 => n10465, C2 => 
                           n7333, A => n9626, ZN => n7334);
   U7755 : OAI21_X1 port map( B1 => n10839, B2 => n12083, A => n10837, ZN => 
                           n7335);
   U7756 : AOI21_X1 port map( B1 => n10839, B2 => n12083, A => n7335, ZN => 
                           n7336);
   U7757 : INV_X1 port map( A => n12083, ZN => n7337);
   U7758 : INV_X1 port map( A => n10838, ZN => n7338);
   U7759 : AOI221_X1 port map( B1 => n12083, B2 => n10838, C1 => n7337, C2 => 
                           n7338, A => n12084, ZN => n7339);
   U7760 : OAI22_X1 port map( A1 => n10459, A2 => n10505, B1 => n10481, B2 => 
                           n10388, ZN => n7340);
   U7761 : INV_X1 port map( A => n10507, ZN => n7341);
   U7762 : OAI22_X1 port map( A1 => n10506, A2 => n10462, B1 => n10508, B2 => 
                           n10479, ZN => n7342);
   U7763 : OAI22_X1 port map( A1 => n10431, A2 => n10460, B1 => n10480, B2 => 
                           n10442, ZN => n7343);
   U7764 : AOI211_X1 port map( C1 => n10440, C2 => n7341, A => n7342, B => 
                           n7343, ZN => n7344);
   U7765 : OAI21_X1 port map( B1 => n10400, B2 => n10376, A => n7344, ZN => 
                           n7345);
   U7766 : AOI211_X1 port map( C1 => n10509, C2 => n10493, A => n7340, B => 
                           n7345, ZN => n7346);
   U7767 : OAI221_X1 port map( B1 => n7787, B2 => n10458, C1 => n7333, C2 => 
                           n10468, A => n9626, ZN => n7347);
   U7768 : INV_X1 port map( A => DP_OP_751_130_5637_n171, ZN => n7348);
   U7769 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n172, A2 => n7348, ZN =>
                           n7349);
   U7770 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n173, A2 => n7349, ZN =>
                           n7350);
   U7771 : OAI211_X1 port map( C1 => DP_OP_751_130_5637_n173, C2 => n7349, A =>
                           n10492, B => n7350, ZN => n7351);
   U7772 : OAI211_X1 port map( C1 => n10452, C2 => n7346, A => n7347, B => 
                           n7351, ZN => n7352);
   U7773 : NOR4_X1 port map( A1 => n7334, A2 => n7336, A3 => n7339, A4 => n7352
                           , ZN => n7353);
   U7774 : OAI22_X1 port map( A1 => n12093, A2 => n7353, B1 => n498, B2 => 
                           n12092, ZN => n7016);
   U7775 : AND2_X1 port map( A1 => n8695, A2 => 
                           DataPath_RF_internal_out1_8_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N12);
   U7776 : AND2_X1 port map( A1 => n8693, A2 => 
                           DataPath_RF_internal_out2_7_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N11);
   U7777 : XOR2_X1 port map( A => n7828, B => 
                           DataPath_ALUhw_MULT_mux_out_1_12_port, Z => n7354);
   U7778 : OAI22_X1 port map( A1 => n7754, A2 => n10386, B1 => n8487, B2 => 
                           n8492, ZN => n7355);
   U7779 : XOR2_X1 port map( A => n8265, B => n7355, Z => n7356);
   U7780 : NOR2_X1 port map( A1 => n7354, A2 => n7356, ZN => 
                           DP_OP_751_130_5637_n1705);
   U7781 : XOR2_X1 port map( A => n7354, B => n7356, Z => 
                           DP_OP_751_130_5637_n1706);
   U7782 : OAI22_X1 port map( A1 => n11852, A2 => n11596, B1 => n577, B2 => 
                           n11851, ZN => n7357);
   U7783 : AOI211_X1 port map( C1 => n8969, C2 => n8803, A => RST, B => n7357, 
                           ZN => n11477);
   U7784 : AOI211_X1 port map( C1 => n10487, C2 => n12089, A => n9340, B => 
                           n12072, ZN => n7358);
   U7785 : INV_X1 port map( A => n7358, ZN => n9953);
   U7786 : INV_X1 port map( A => n9434, ZN => n7359);
   U7787 : AOI222_X1 port map( A1 => n7359, A2 => n10089, B1 => n9620, B2 => 
                           n10288, C1 => n10090, C2 => n9983, ZN => n7360);
   U7788 : INV_X1 port map( A => n9433, ZN => n7361);
   U7789 : NOR2_X1 port map( A1 => n9747, A2 => n7361, ZN => n7362);
   U7790 : AOI21_X1 port map( B1 => n9423, B2 => n9980, A => n10457, ZN => 
                           n7363);
   U7791 : AOI211_X1 port map( C1 => n7785, C2 => n9820, A => n7362, B => n7363
                           , ZN => n7364);
   U7792 : OAI211_X1 port map( C1 => n9817, C2 => n9419, A => n7360, B => n7364
                           , ZN => n10497);
   U7793 : AND2_X1 port map( A1 => n8695, A2 => 
                           DataPath_RF_internal_out1_5_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N9);
   U7794 : AND2_X1 port map( A1 => n8694, A2 => 
                           DataPath_RF_internal_out2_6_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N10);
   U7795 : XOR2_X1 port map( A => DP_OP_751_130_5637_n1736, B => 
                           DP_OP_751_130_5637_n1767, Z => 
                           DP_OP_751_130_5637_n1676);
   U7796 : OAI22_X1 port map( A1 => n9452, A2 => n10395, B1 => n8560, B2 => 
                           n8559, ZN => n7365);
   U7797 : XNOR2_X1 port map( A => n8263, B => n7365, ZN => n7366);
   U7798 : XOR2_X1 port map( A => n8265, B => 
                           DataPath_ALUhw_MULT_mux_out_0_11_port, Z => n7367);
   U7799 : XOR2_X1 port map( A => n7366, B => n7367, Z => 
                           DP_OP_751_130_5637_n1708);
   U7800 : NOR2_X1 port map( A1 => n7366, A2 => n7367, ZN => 
                           DP_OP_751_130_5637_n1707);
   U7801 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, B2 => 
                           n8716, ZN => n7368);
   U7802 : INV_X1 port map( A => n7368, ZN => n8719);
   U7803 : NOR2_X1 port map( A1 => n10590, A2 => IRAM_ADDRESS_27_port, ZN => 
                           n7369);
   U7804 : NOR3_X1 port map( A1 => n7369, A2 => n10587, A3 => n10572, ZN => 
                           n8122);
   U7805 : OAI22_X1 port map( A1 => n11596, A2 => n11851, B1 => n8442, B2 => 
                           n11852, ZN => n7370);
   U7806 : AOI211_X1 port map( C1 => n8969, C2 => n7761, A => RST, B => n7370, 
                           ZN => n11595);
   U7807 : NOR2_X1 port map( A1 => n9494, A2 => n8489, ZN => n7371);
   U7808 : XOR2_X1 port map( A => DP_OP_751_130_5637_n1009, B => n7371, Z => 
                           DP_OP_751_130_5637_n910);
   U7809 : NOR2_X1 port map( A1 => n9494, A2 => n8489, ZN => n7372);
   U7810 : MUX2_X1 port map( A => n8267, B => DP_OP_751_130_5637_n1009, S => 
                           n7372, Z => DP_OP_751_130_5637_n909);
   U7811 : NOR2_X1 port map( A1 => n9482, A2 => n8488, ZN => n7373);
   U7812 : XOR2_X1 port map( A => DP_OP_751_130_5637_n1213, B => n7373, Z => 
                           DP_OP_751_130_5637_n1114);
   U7813 : NOR2_X1 port map( A1 => n9482, A2 => n8488, ZN => n7374);
   U7814 : MUX2_X1 port map( A => n7770, B => DP_OP_751_130_5637_n1213, S => 
                           n7374, Z => DP_OP_751_130_5637_n1113);
   U7815 : AOI211_X1 port map( C1 => n8016, C2 => n12089, A => n9365, B => 
                           n12072, ZN => n7375);
   U7816 : INV_X1 port map( A => n7375, ZN => n9885);
   U7817 : NOR2_X1 port map( A1 => n8455, A2 => n8501, ZN => n7376);
   U7818 : NAND3_X1 port map( A1 => n8255, A2 => IR_30_port, A3 => n7376, ZN =>
                           n10709);
   U7819 : AND2_X1 port map( A1 => n8693, A2 => 
                           DataPath_RF_internal_out1_6_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N10);
   U7820 : AND2_X1 port map( A1 => n8693, A2 => 
                           DataPath_RF_internal_out2_5_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N9);
   U7821 : NAND2_X1 port map( A1 => n7879, A2 => n7927, ZN => n7377);
   U7822 : INV_X1 port map( A => n8072, ZN => n7378);
   U7823 : OAI21_X1 port map( B1 => n8072, B2 => DP_OP_751_130_5637_n1335, A =>
                           n7377, ZN => n7379);
   U7824 : OAI21_X1 port map( B1 => n7826, B2 => n7378, A => n7379, ZN => 
                           DP_OP_751_130_5637_n1283);
   U7825 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_14_port, B2 => 
                           n8716, ZN => n10891);
   U7826 : OAI22_X1 port map( A1 => n8487, A2 => n10181, B1 => n7755, B2 => 
                           n9944, ZN => n7380);
   U7827 : XNOR2_X1 port map( A => n7979, B => n7380, ZN => 
                           DP_OP_751_130_5637_n1768);
   U7828 : INV_X1 port map( A => DataPath_RF_c_win_0_port, ZN => n7381);
   U7829 : INV_X1 port map( A => DataPath_RF_c_win_4_port, ZN => n7382);
   U7830 : OAI22_X1 port map( A1 => n7381, A2 => DataPath_RF_c_swin_2_port, B1 
                           => n7382, B2 => DataPath_RF_c_swin_1_port, ZN => 
                           n7383);
   U7831 : AOI221_X1 port map( B1 => n7381, B2 => DataPath_RF_c_swin_2_port, C1
                           => DataPath_RF_c_swin_1_port, C2 => n7382, A => 
                           n7383, ZN => n7384);
   U7832 : OAI22_X1 port map( A1 => DataPath_RF_c_win_1_port, A2 => n823, B1 =>
                           DataPath_RF_c_win_2_port, B2 => n824, ZN => n7385);
   U7833 : AOI221_X1 port map( B1 => DataPath_RF_c_win_1_port, B2 => n823, C1 
                           => n824, C2 => DataPath_RF_c_win_2_port, A => n7385,
                           ZN => n7386);
   U7834 : XNOR2_X1 port map( A => DataPath_RF_c_swin_0_port, B => 
                           DataPath_RF_c_win_3_port, ZN => n7387);
   U7835 : NAND3_X1 port map( A1 => n7386, A2 => n7384, A3 => n7387, ZN => 
                           n8978);
   U7836 : OR3_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_23_port, A3 => n8121, ZN
                           => n7942);
   U7837 : NAND2_X1 port map( A1 => n8229, A2 => n7799, ZN => n7388);
   U7838 : OAI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n72, B2 => 
                           DataPath_WRF_CUhw_curr_addr_24_port, A => n7388, ZN 
                           => n8228);
   U7839 : OAI22_X1 port map( A1 => n11856, A2 => n11596, B1 => n577, B2 => 
                           n11855, ZN => n7389);
   U7840 : AOI211_X1 port map( C1 => n8972, C2 => n8803, A => RST, B => n7389, 
                           ZN => n11511);
   U7841 : INV_X1 port map( A => n10006, ZN => n7390);
   U7842 : NAND2_X1 port map( A1 => n7390, A2 => n9694, ZN => n7391);
   U7843 : OAI21_X1 port map( B1 => n10004, B2 => n7391, A => n10007, ZN => 
                           n7392);
   U7844 : AOI21_X1 port map( B1 => n10001, B2 => n7392, A => n10002, ZN => 
                           n9868);
   U7845 : NOR2_X1 port map( A1 => n7694, A2 => n8489, ZN => n7393);
   U7846 : XOR2_X1 port map( A => DP_OP_751_130_5637_n1519, B => n7393, Z => 
                           DP_OP_751_130_5637_n1420);
   U7847 : NOR2_X1 port map( A1 => n7694, A2 => n8489, ZN => n7394);
   U7848 : MUX2_X1 port map( A => n7798, B => DP_OP_751_130_5637_n1519, S => 
                           n7394, Z => DP_OP_751_130_5637_n1419);
   U7849 : INV_X1 port map( A => n10576, ZN => n7395);
   U7850 : NAND3_X1 port map( A1 => n8393, A2 => n8389, A3 => n7395, ZN => 
                           n8474);
   U7851 : AOI22_X1 port map( A1 => n10026, A2 => n10229, B1 => n10027, B2 => 
                           n10113, ZN => n7396);
   U7852 : OAI21_X1 port map( B1 => n10182, B2 => n10024, A => n10180, ZN => 
                           n7397);
   U7853 : AOI22_X1 port map( A1 => n10028, A2 => n10288, B1 => n10025, B2 => 
                           n7397, ZN => n7398);
   U7854 : NAND3_X1 port map( A1 => n10023, A2 => n10022, A3 => n10084, ZN => 
                           n7399);
   U7855 : NAND3_X1 port map( A1 => n7396, A2 => n7398, A3 => n7399, ZN => 
                           n10294);
   U7856 : AOI22_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_16_port,
                           B1 => DataPath_i_PIPLIN_B_16_port, B2 => n8165, ZN 
                           => n7400);
   U7857 : INV_X1 port map( A => n7400, ZN => n10313);
   U7858 : AOI21_X1 port map( B1 => n7691, B2 => n10648, A => n7759, ZN => 
                           n7401);
   U7859 : AOI222_X1 port map( A1 => n10650, A2 => n7401, B1 => n10835, B2 => 
                           IRAM_ADDRESS_13_port, C1 => i_RD1_13_port, C2 => 
                           n12070, ZN => n7402);
   U7860 : INV_X1 port map( A => n7402, ZN => n7046);
   U7861 : NAND2_X1 port map( A1 => n7751, A2 => DP_OP_751_130_5637_n183, ZN =>
                           n7403);
   U7862 : XNOR2_X1 port map( A => n7403, B => DP_OP_751_130_5637_n184, ZN => 
                           n7404);
   U7863 : INV_X1 port map( A => n8015, ZN => n7405);
   U7864 : AOI22_X1 port map( A1 => n8015, A2 => n10468, B1 => n10469, B2 => 
                           n7405, ZN => n7406);
   U7865 : NAND2_X1 port map( A1 => n10471, A2 => n10470, ZN => n7407);
   U7866 : AOI21_X1 port map( B1 => n7407, B2 => n7406, A => n10473, ZN => 
                           n7408);
   U7867 : INV_X1 port map( A => n12084, ZN => n7409);
   U7868 : INV_X1 port map( A => n10470, ZN => n7410);
   U7869 : AOI22_X1 port map( A1 => n8015, A2 => n10489, B1 => n10465, B2 => 
                           n7405, ZN => n7411);
   U7870 : AOI221_X1 port map( B1 => n10837, B2 => n10470, C1 => n7409, C2 => 
                           n7410, A => n7411, ZN => n7412);
   U7871 : INV_X1 port map( A => n10837, ZN => n7413);
   U7872 : OAI22_X1 port map( A1 => n8495, A2 => n7412, B1 => n10472, B2 => 
                           n7413, ZN => n7414);
   U7873 : AOI211_X1 port map( C1 => n7404, C2 => n8578, A => n7408, B => n7414
                           , ZN => n7415);
   U7874 : AOI22_X1 port map( A1 => n10498, A2 => n10477, B1 => n10510, B2 => 
                           n10478, ZN => n7416);
   U7875 : AOI22_X1 port map( A1 => n10499, A2 => n10474, B1 => n10475, B2 => 
                           n10476, ZN => n7417);
   U7876 : AOI22_X1 port map( A1 => n10493, A2 => n10501, B1 => n10503, B2 => 
                           n10497, ZN => n7418);
   U7877 : NAND3_X1 port map( A1 => n7416, A2 => n7417, A3 => n7418, ZN => 
                           n7419);
   U7878 : OAI22_X1 port map( A1 => n10480, A2 => n10479, B1 => n10481, B2 => 
                           n10505, ZN => n7420);
   U7879 : AOI211_X1 port map( C1 => n10495, C2 => n10509, A => n7419, B => 
                           n7420, ZN => n7421);
   U7880 : OAI222_X1 port map( A1 => n12093, A2 => n7415, B1 => n12092, B2 => 
                           n497, C1 => n10482, C2 => n7421, ZN => n7018);
   U7881 : AND2_X1 port map( A1 => n8695, A2 => 
                           DataPath_RF_internal_out1_3_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N7);
   U7882 : AND2_X1 port map( A1 => n8693, A2 => 
                           DataPath_RF_internal_out2_4_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N8);
   U7883 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n987, B2 => 
                           DP_OP_751_130_5637_n933, A => 
                           DP_OP_751_130_5637_n986, ZN => n7821);
   U7884 : NAND2_X1 port map( A1 => n7825, A2 => n7879, ZN => n7422);
   U7885 : OAI221_X1 port map( B1 => n7826, B2 => n7927, C1 => n7826, C2 => 
                           n7879, A => n7422, ZN => n8073);
   U7886 : INV_X1 port map( A => n8179, ZN => n7423);
   U7887 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n432, A2 => n7423, ZN => 
                           n7895);
   U7888 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, B2 => 
                           n8716, ZN => n10889);
   U7889 : OR2_X1 port map( A1 => n8290, A2 => n8295, ZN => n8232);
   U7890 : OAI22_X1 port map( A1 => n11596, A2 => n11855, B1 => n8442, B2 => 
                           n11856, ZN => n7424);
   U7891 : AOI211_X1 port map( C1 => n8972, C2 => n8852, A => RST, B => n7424, 
                           ZN => n11630);
   U7892 : INV_X1 port map( A => DP_OP_751_130_5637_n536, ZN => n7425);
   U7893 : INV_X1 port map( A => DP_OP_751_130_5637_n537, ZN => n7426);
   U7894 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n537, B2 => 
                           DP_OP_751_130_5637_n536, A => 
                           DP_OP_751_130_5637_n601, ZN => n7427);
   U7895 : OAI21_X1 port map( B1 => n7425, B2 => n7426, A => n7427, ZN => 
                           DP_OP_751_130_5637_n501);
   U7896 : AOI21_X1 port map( B1 => n12082, B2 => n10487, A => n9340, ZN => 
                           n7428);
   U7897 : INV_X1 port map( A => n7428, ZN => n9954);
   U7898 : NOR2_X1 port map( A1 => n9458, A2 => n8489, ZN => n7429);
   U7899 : XOR2_X1 port map( A => DP_OP_751_130_5637_n1621, B => n7429, Z => 
                           DP_OP_751_130_5637_n1522);
   U7900 : NOR2_X1 port map( A1 => n9458, A2 => n8489, ZN => n7430);
   U7901 : MUX2_X1 port map( A => n8260, B => DP_OP_751_130_5637_n1621, S => 
                           n7430, Z => DP_OP_751_130_5637_n1521);
   U7902 : AOI22_X1 port map( A1 => n7767, A2 => n7800, B1 => n8681, B2 => 
                           n8093, ZN => n7431);
   U7903 : INV_X1 port map( A => n7431, ZN => n9730);
   U7904 : INV_X1 port map( A => n8446, ZN => n7432);
   U7905 : AOI21_X1 port map( B1 => n7760, B2 => n8218, A => n7432, ZN => n8216
                           );
   U7906 : INV_X1 port map( A => n7942, ZN => n7433);
   U7907 : AOI21_X1 port map( B1 => n7943, B2 => n8088, A => n7433, ZN => 
                           DP_OP_1090J1_126_7243_n9);
   U7908 : INV_X1 port map( A => n9563, ZN => n7434);
   U7909 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_I2, A2 => n8081, ZN => 
                           n7435);
   U7910 : OAI21_X1 port map( B1 => n7434, B2 => DP_OP_751_130_5637_n1761, A =>
                           n7435, ZN => n9451);
   U7911 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n333, A2 => n9742, ZN =>
                           n7436);
   U7912 : NAND2_X1 port map( A1 => n10465, A2 => n7436, ZN => n7437);
   U7913 : OAI221_X1 port map( B1 => n7436, B2 => n10458, C1 => 
                           DP_OP_751_130_5637_n333, C2 => n9742, A => n7437, ZN
                           => n7438);
   U7914 : OAI21_X1 port map( B1 => n9742, B2 => n8681, A => n12091, ZN => 
                           n7439);
   U7915 : XNOR2_X1 port map( A => n7439, B => DP_OP_751_130_5637_n333, ZN => 
                           n7440);
   U7916 : NOR2_X1 port map( A1 => n9650, A2 => n9761, ZN => n7441);
   U7917 : AOI21_X1 port map( B1 => n9791, B2 => n9792, A => n7441, ZN => n7442
                           );
   U7918 : AOI21_X1 port map( B1 => n7440, B2 => n7442, A => n9854, ZN => n7443
                           );
   U7919 : OAI21_X1 port map( B1 => n7440, B2 => n7442, A => n7443, ZN => n7444
                           );
   U7920 : AOI21_X1 port map( B1 => n9792, B2 => n9793, A => n7441, ZN => n7445
                           );
   U7921 : NAND2_X1 port map( A1 => n7440, A2 => n7445, ZN => n7446);
   U7922 : OAI211_X1 port map( C1 => n7440, C2 => n7445, A => n9838, B => n7446
                           , ZN => n7447);
   U7923 : INV_X1 port map( A => DP_OP_751_130_5637_n333, ZN => n7448);
   U7924 : NAND3_X1 port map( A1 => n10024, A2 => n10469, A3 => n7448, ZN => 
                           n7449);
   U7925 : NAND4_X1 port map( A1 => n7438, A2 => n7444, A3 => n7447, A4 => 
                           n7449, ZN => n9712);
   U7926 : INV_X1 port map( A => n10181, ZN => n7450);
   U7927 : OAI21_X1 port map( B1 => n9702, B2 => n7450, A => n9871, ZN => n9905
                           );
   U7928 : AOI222_X1 port map( A1 => n10110, A2 => n10288, B1 => n10111, B2 => 
                           n10229, C1 => n10112, C2 => n10113, ZN => n7451);
   U7929 : INV_X1 port map( A => n10115, ZN => n7452);
   U7930 : INV_X1 port map( A => n10114, ZN => n7453);
   U7931 : OAI221_X1 port map( B1 => n10115, B2 => n10116, C1 => n7452, C2 => 
                           n7453, A => n10232, ZN => n7454);
   U7932 : OAI211_X1 port map( C1 => n10109, C2 => n10292, A => n7451, B => 
                           n7454, ZN => n7455);
   U7933 : AOI21_X1 port map( B1 => n7785, B2 => n10108, A => n7455, ZN => 
                           n10371);
   U7934 : XNOR2_X1 port map( A => n8264, B => 
                           DataPath_ALUhw_MULT_mux_out_0_0_port, ZN => 
                           DP_OP_751_130_5637_n1795);
   U7935 : NOR2_X1 port map( A1 => n10716, A2 => n10771, ZN => n7456);
   U7936 : OAI21_X1 port map( B1 => n8255, B2 => n7456, A => n8185, ZN => 
                           n10715);
   U7937 : AOI211_X1 port map( C1 => n7687, C2 => n7686, A => n8156, B => 
                           n10590, ZN => n7457);
   U7938 : INV_X1 port map( A => n7457, ZN => n7458);
   U7939 : AOI21_X1 port map( B1 => n10576, B2 => n7458, A => n10835, ZN => 
                           n7459);
   U7940 : NOR3_X1 port map( A1 => n12070, A2 => n7459, A3 => n8389, ZN => 
                           n7460);
   U7941 : NAND3_X1 port map( A1 => n7459, A2 => n8389, A3 => n10577, ZN => 
                           n7461);
   U7942 : OAI21_X1 port map( B1 => n8549, B2 => n10578, A => n7461, ZN => 
                           n7462);
   U7943 : NOR2_X1 port map( A1 => n7460, A2 => n7462, ZN => n8475);
   U7944 : NAND2_X1 port map( A1 => n8016, A2 => n8263, ZN => n7463);
   U7945 : NAND2_X1 port map( A1 => n10465, A2 => n7463, ZN => n7464);
   U7946 : OAI221_X1 port map( B1 => n7463, B2 => n10458, C1 => n8016, C2 => 
                           n8263, A => n7464, ZN => n7465);
   U7947 : XNOR2_X1 port map( A => n8016, B => n9597, ZN => n7466);
   U7948 : NAND2_X1 port map( A1 => n9573, A2 => n9591, ZN => n7467);
   U7949 : OAI21_X1 port map( B1 => n7467, B2 => n10491, A => n9595, ZN => 
                           n7468);
   U7950 : NAND2_X1 port map( A1 => n12080, A2 => n7468, ZN => n7469);
   U7951 : OAI21_X1 port map( B1 => n7466, B2 => n7469, A => n10842, ZN => 
                           n7470);
   U7952 : AOI21_X1 port map( B1 => n7466, B2 => n7469, A => n7470, ZN => n7471
                           );
   U7953 : XNOR2_X1 port map( A => n7466, B => n7468, ZN => n7472);
   U7954 : AOI21_X1 port map( B1 => n7472, B2 => n10490, A => n7471, ZN => 
                           n7473);
   U7955 : INV_X1 port map( A => DP_OP_751_130_5637_n185, ZN => n7474);
   U7956 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n186, A2 => n7474, ZN =>
                           n7475);
   U7957 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n187, A2 => n7475, ZN =>
                           n7476);
   U7958 : OAI211_X1 port map( C1 => DP_OP_751_130_5637_n187, C2 => n7475, A =>
                           n10492, B => n7476, ZN => n7477);
   U7959 : NAND3_X1 port map( A1 => n9721, A2 => n10469, A3 => n7828, ZN => 
                           n7478);
   U7960 : NAND4_X1 port map( A1 => n7465, A2 => n7473, A3 => n7477, A4 => 
                           n7478, ZN => n7479);
   U7961 : AOI22_X1 port map( A1 => n10510, A2 => n10477, B1 => n10499, B2 => 
                           n10478, ZN => n7480);
   U7962 : NAND2_X1 port map( A1 => n10503, A2 => n10501, ZN => n7481);
   U7963 : OAI21_X1 port map( B1 => n10376, B2 => n10480, A => n7481, ZN => 
                           n7482);
   U7964 : AOI21_X1 port map( B1 => n10502, B2 => n10509, A => n7482, ZN => 
                           n7483);
   U7965 : AOI22_X1 port map( A1 => n10497, A2 => n10495, B1 => n10493, B2 => 
                           n10496, ZN => n7484);
   U7966 : AOI22_X1 port map( A1 => n10474, A2 => n10461, B1 => n10476, B2 => 
                           n10403, ZN => n7485);
   U7967 : NAND4_X1 port map( A1 => n7480, A2 => n7483, A3 => n7484, A4 => 
                           n7485, ZN => n7486);
   U7968 : AOI222_X1 port map( A1 => n7479, A2 => n10841, B1 => n7764, B2 => 
                           DRAM_ADDRESS_3_port, C1 => n7486, C2 => n10840, ZN 
                           => n2228);
   U7969 : AND2_X1 port map( A1 => n8695, A2 => 
                           DataPath_RF_internal_out1_4_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N8);
   U7970 : AND2_X1 port map( A1 => n8694, A2 => 
                           DataPath_RF_internal_out2_3_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N7);
   U7971 : NAND2_X1 port map( A1 => n8077, A2 => n7917, ZN => n7487);
   U7972 : OAI21_X1 port map( B1 => n7487, B2 => DP_OP_751_130_5637_n1435, A =>
                           DP_OP_751_130_5637_n1480, ZN => n8071);
   U7973 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n595, B2 => 
                           DP_OP_751_130_5637_n533, A => 
                           DP_OP_751_130_5637_n594, ZN => n7930);
   U7974 : OAI22_X1 port map( A1 => n9452, A2 => n9659, B1 => n8562, B2 => 
                           n7787, ZN => n7488);
   U7975 : XNOR2_X1 port map( A => n8263, B => n7488, ZN => n7489);
   U7976 : OAI22_X1 port map( A1 => n7755, A2 => n8559, B1 => n7796, B2 => 
                           n10395, ZN => n7490);
   U7977 : XOR2_X1 port map( A => n8265, B => n7490, Z => n7491);
   U7978 : XOR2_X1 port map( A => n7489, B => n7491, Z => 
                           DP_OP_751_130_5637_n1712);
   U7979 : NOR2_X1 port map( A1 => n7489, A2 => n7491, ZN => 
                           DP_OP_751_130_5637_n1711);
   U7980 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, B2 => 
                           n8716, ZN => n10890);
   U7981 : INV_X1 port map( A => DP_OP_751_130_5637_n333, ZN => n7492);
   U7982 : AOI22_X1 port map( A1 => DP_OP_751_130_5637_n333, A2 => n9794, B1 =>
                           n9815, B2 => n7492, ZN => n7493);
   U7983 : OAI21_X1 port map( B1 => n9794, B2 => n9815, A => n7493, ZN => n7494
                           );
   U7984 : OAI22_X1 port map( A1 => n10511, A2 => n9526, B1 => n8488, B2 => 
                           n7494, ZN => n7495);
   U7985 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n333, B => n7495, ZN => 
                           n7753);
   U7986 : INV_X1 port map( A => n7791, ZN => n7496);
   U7987 : NAND2_X1 port map( A1 => n8286, A2 => n7496, ZN => n8242);
   U7988 : NOR4_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_17_port, A3 => n8290, A4
                           => n8295, ZN => n8231);
   U7989 : OAI22_X1 port map( A1 => n8299, A2 => n11856, B1 => n8442, B2 => 
                           n11855, ZN => n7497);
   U7990 : AOI211_X1 port map( C1 => n8972, C2 => n8532, A => RST, B => n7497, 
                           ZN => n11749);
   U7991 : AOI211_X1 port map( C1 => n8011, C2 => n12089, A => n9387, B => 
                           n12072, ZN => n9774);
   U7992 : NOR2_X1 port map( A1 => n9475, A2 => n8488, ZN => n7498);
   U7993 : XOR2_X1 port map( A => DP_OP_751_130_5637_n1315, B => n7498, Z => 
                           DP_OP_751_130_5637_n1216);
   U7994 : NOR2_X1 port map( A1 => n9475, A2 => n8488, ZN => n7499);
   U7995 : MUX2_X1 port map( A => DP_OP_751_130_5637_n1251, B => 
                           DP_OP_751_130_5637_n1315, S => n7499, Z => 
                           DP_OP_751_130_5637_n1215);
   U7996 : AOI22_X1 port map( A1 => n8681, A2 => n7769, B1 => n7800, B2 => 
                           n10377, ZN => n7500);
   U7997 : INV_X1 port map( A => n7500, ZN => n9799);
   U7998 : AOI21_X1 port map( B1 => n10642, B2 => n10643, A => n7775, ZN => 
                           n8218);
   U7999 : AOI221_X1 port map( B1 => n8723, B2 => n8256, C1 => n10876, C2 => 
                           n8256, A => n10846, ZN => n8981);
   U8000 : INV_X1 port map( A => n8298, ZN => n7501);
   U8001 : OAI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n72, B2 => n7501, A 
                           => DataPath_WRF_CUhw_curr_addr_25_port, ZN => n7502)
                           ;
   U8002 : OAI21_X1 port map( B1 => n8298, B2 => n7799, A => n7502, ZN => n7503
                           );
   U8003 : NOR3_X1 port map( A1 => n7943, A2 => n8228, A3 => n7941, ZN => n7504
                           );
   U8004 : NOR2_X1 port map( A1 => n7504, A2 => n7503, ZN => n7939);
   U8005 : OAI21_X1 port map( B1 => n10569, B2 => n192, A => n10571, ZN => 
                           n12065);
   U8006 : INV_X1 port map( A => n10573, ZN => n7505);
   U8007 : NAND2_X1 port map( A1 => n8122, A2 => n7505, ZN => n7687);
   U8008 : AOI222_X1 port map( A1 => n10112, A2 => n10231, B1 => n9983, B2 => 
                           n10122, C1 => n10111, C2 => n9844, ZN => n7506);
   U8009 : AOI22_X1 port map( A1 => n9845, A2 => n9920, B1 => n10116, B2 => 
                           n9985, ZN => n7507);
   U8010 : INV_X1 port map( A => n9846, ZN => n7508);
   U8011 : AOI22_X1 port map( A1 => n10110, A2 => n10282, B1 => n7785, B2 => 
                           n7508, ZN => n7509);
   U8012 : NAND3_X1 port map( A1 => n7506, A2 => n7507, A3 => n7509, ZN => 
                           n7510);
   U8013 : AOI21_X1 port map( B1 => n10108, B2 => n10288, A => n7510, ZN => 
                           n10064);
   U8014 : INV_X1 port map( A => n8550, ZN => n7511);
   U8015 : OAI21_X1 port map( B1 => n9681, B2 => n7511, A => n10213, ZN => 
                           n10174);
   U8016 : INV_X1 port map( A => n7772, ZN => n7512);
   U8017 : NOR2_X1 port map( A1 => n9680, A2 => n7512, ZN => n10304);
   U8018 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n184, A2 => n7751, ZN =>
                           n7513);
   U8019 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n183, A2 => n7513, ZN =>
                           DP_OP_751_130_5637_n178);
   U8020 : NAND3_X1 port map( A1 => n8084, A2 => n10857, A3 => n10744, ZN => 
                           n10751);
   U8021 : XOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_23_port, Z => n7514);
   U8022 : NAND2_X1 port map( A1 => n8088, A2 => n8087, ZN => n7515);
   U8023 : OAI21_X1 port map( B1 => n7514, B2 => n7515, A => n10730, ZN => 
                           n7516);
   U8024 : AOI21_X1 port map( B1 => n7514, B2 => n7515, A => n7516, ZN => 
                           DRAMRF_ADDRESS_23_port);
   U8025 : INV_X1 port map( A => n10740, ZN => n7517);
   U8026 : AOI22_X1 port map( A1 => n10740, A2 => n8420, B1 => n5686, B2 => 
                           n7517, ZN => n9641);
   U8027 : AOI22_X2 port map( A1 => n8314, A2 => DataPath_i_PIPLIN_IN1_15_port,
                           B1 => n8674, B2 => DataPath_i_PIPLIN_A_15_port, ZN 
                           => n8554);
   U8028 : NOR2_X1 port map( A1 => n8080, A2 => n10832, ZN => n7518);
   U8029 : AOI21_X1 port map( B1 => IRAM_DATA(31), B2 => n8580, A => n7518, ZN 
                           => n8479);
   U8030 : NAND2_X1 port map( A1 => n8474, A2 => n8473, ZN => n7519);
   U8031 : XNOR2_X1 port map( A => n7519, B => n8430, ZN => n7520);
   U8032 : AOI222_X1 port map( A1 => n7520, A2 => n8303, B1 => n10835, B2 => 
                           IRAM_ADDRESS_31_port, C1 => i_RD1_31_port, C2 => 
                           n12070, ZN => n8476);
   U8033 : AOI22_X1 port map( A1 => n10490, A2 => n10483, B1 => n10842, B2 => 
                           n10485, ZN => n7521);
   U8034 : INV_X1 port map( A => n10486, ZN => n7522);
   U8035 : NOR3_X1 port map( A1 => n10511, A2 => n7979, A3 => n10489, ZN => 
                           n7523);
   U8036 : OAI33_X1 port map( A1 => n10485, A2 => n10486, A3 => n10484, B1 => 
                           n8076, B2 => n10487, B3 => n10488, ZN => n7524);
   U8037 : AOI211_X1 port map( C1 => n10490, C2 => n10491, A => n7523, B => 
                           n7524, ZN => n7525);
   U8038 : OAI21_X1 port map( B1 => n7521, B2 => n7522, A => n7525, ZN => n7526
                           );
   U8039 : XOR2_X1 port map( A => DP_OP_751_130_5637_n196, B => 
                           DP_OP_751_130_5637_n194, Z => n7527);
   U8040 : AOI21_X1 port map( B1 => n7527, B2 => n8578, A => n7526, ZN => n7528
                           );
   U8041 : AOI22_X1 port map( A1 => n10496, A2 => n10495, B1 => n10494, B2 => 
                           n10493, ZN => n7529);
   U8042 : AOI22_X1 port map( A1 => n10500, A2 => n10499, B1 => n10498, B2 => 
                           n10497, ZN => n7530);
   U8043 : AOI22_X1 port map( A1 => n10504, A2 => n10503, B1 => n10502, B2 => 
                           n10501, ZN => n7531);
   U8044 : OAI22_X1 port map( A1 => n10508, A2 => n10507, B1 => n10506, B2 => 
                           n10505, ZN => n7532);
   U8045 : AOI21_X1 port map( B1 => n10510, B2 => n10509, A => n7532, ZN => 
                           n7533);
   U8046 : NAND4_X1 port map( A1 => n7529, A2 => n7530, A3 => n7531, A4 => 
                           n7533, ZN => n7534);
   U8047 : XNOR2_X1 port map( A => n10511, B => n7979, ZN => n7535);
   U8048 : OAI22_X1 port map( A1 => n10512, A2 => n7535, B1 => n496, B2 => 
                           n12092, ZN => n7536);
   U8049 : AOI21_X1 port map( B1 => n10840, B2 => n7534, A => n7536, ZN => 
                           n7537);
   U8050 : OAI21_X1 port map( B1 => n10513, B2 => n7528, A => n7537, ZN => 
                           n7019);
   U8051 : AND2_X1 port map( A1 => n8695, A2 => 
                           DataPath_RF_internal_out1_2_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N6);
   U8052 : AND2_X1 port map( A1 => n8694, A2 => 
                           DataPath_RF_internal_out2_1_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N5);
   U8053 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1283, B2 => 
                           DP_OP_751_130_5637_n1234, A => 
                           DP_OP_751_130_5637_n1282, ZN => n7888);
   U8054 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, B2 => 
                           n8716, ZN => n10888);
   U8055 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1087, B2 => 
                           DP_OP_751_130_5637_n1034, A => 
                           DP_OP_751_130_5637_n1086, ZN => n7538);
   U8056 : OAI21_X1 port map( B1 => n7539, B2 => n7540, A => n7538, ZN => 
                           DP_OP_751_130_5637_n987);
   U8057 : INV_X1 port map( A => DP_OP_751_130_5637_n1034, ZN => n7539);
   U8058 : INV_X1 port map( A => DP_OP_751_130_5637_n1087, ZN => n7540);
   U8059 : OAI22_X1 port map( A1 => n7754, A2 => n9659, B1 => n7796, B2 => 
                           n8559, ZN => n7541);
   U8060 : XOR2_X1 port map( A => n8265, B => n7541, Z => n7542);
   U8061 : XNOR2_X1 port map( A => n8263, B => 
                           DataPath_ALUhw_MULT_mux_out_1_8_port, ZN => n7543);
   U8062 : NOR2_X1 port map( A1 => n7542, A2 => n7543, ZN => 
                           DP_OP_751_130_5637_n1713);
   U8063 : XOR2_X1 port map( A => n7542, B => n7543, Z => 
                           DP_OP_751_130_5637_n1714);
   U8064 : INV_X1 port map( A => n10884, ZN => n7544);
   U8065 : NAND2_X1 port map( A1 => n7544, A2 => n10879, ZN => n7545);
   U8066 : OAI21_X1 port map( B1 => n10881, B2 => n7545, A => n10910, ZN => 
                           n10911);
   U8067 : NAND3_X1 port map( A1 => n8313, A2 => n10734, A3 => n477, ZN => 
                           n8452);
   U8068 : NOR3_X1 port map( A1 => n8290, A2 => 
                           DataPath_WRF_CUhw_curr_addr_18_port, A3 => 
                           DP_OP_1090J1_126_7243_n72, ZN => n8233);
   U8069 : INV_X1 port map( A => DP_OP_751_130_5637_n435, ZN => n7546);
   U8070 : NAND2_X1 port map( A1 => n9839, A2 => n9875, ZN => n7547);
   U8071 : OAI221_X1 port map( B1 => n9839, B2 => DP_OP_751_130_5637_n435, C1 
                           => n9875, C2 => n7546, A => n7547, ZN => n9522);
   U8072 : INV_X1 port map( A => n8216, ZN => n7548);
   U8073 : NOR2_X1 port map( A1 => n10553, A2 => n7548, ZN => n8215);
   U8074 : NOR2_X1 port map( A1 => n7779, A2 => n11753, ZN => n7549);
   U8075 : AOI21_X1 port map( B1 => n11754, B2 => n7761, A => n7549, ZN => 
                           n11519);
   U8076 : INV_X1 port map( A => n11632, ZN => n7550);
   U8077 : INV_X1 port map( A => n8531, ZN => n7551);
   U8078 : AOI22_X1 port map( A1 => n8531, A2 => n11633, B1 => n7550, B2 => 
                           n7551, ZN => n11643);
   U8079 : INV_X1 port map( A => DP_OP_751_130_5637_n703, ZN => n7552);
   U8080 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n703, B2 => 
                           DP_OP_751_130_5637_n639, A => 
                           DP_OP_751_130_5637_n638, ZN => n7553);
   U8081 : OAI21_X1 port map( B1 => n7790, B2 => n7552, A => n7553, ZN => 
                           DP_OP_751_130_5637_n603);
   U8082 : INV_X1 port map( A => DP_OP_751_130_5637_n740, ZN => n7554);
   U8083 : INV_X1 port map( A => DP_OP_751_130_5637_n741, ZN => n7555);
   U8084 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n741, B2 => 
                           DP_OP_751_130_5637_n740, A => 
                           DP_OP_751_130_5637_n805, ZN => n7556);
   U8085 : OAI21_X1 port map( B1 => n7554, B2 => n7555, A => n7556, ZN => 
                           DP_OP_751_130_5637_n705);
   U8086 : OAI21_X1 port map( B1 => n10185, B2 => n10869, A => n9753, ZN => 
                           n9922);
   U8087 : AOI21_X1 port map( B1 => n10143, B2 => n7800, A => n9720, ZN => 
                           n7557);
   U8088 : INV_X1 port map( A => n7557, ZN => n10160);
   U8089 : AOI21_X1 port map( B1 => n8011, B2 => n12082, A => n9387, ZN => 
                           n7558);
   U8090 : INV_X1 port map( A => n7558, ZN => n10027);
   U8091 : NAND2_X1 port map( A1 => n8978, A2 => n8979, ZN => n7559);
   U8092 : OAI21_X1 port map( B1 => n7559, B2 => n7685, A => n12208, ZN => 
                           n8980);
   U8093 : OAI22_X1 port map( A1 => n8441, A2 => n11855, B1 => n577, B2 => 
                           n11856, ZN => n7560);
   U8094 : AOI211_X1 port map( C1 => n8972, C2 => n7762, A => RST, B => n7560, 
                           ZN => n11416);
   U8095 : OAI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n72, B2 => 
                           DataPath_WRF_CUhw_curr_addr_24_port, A => 
                           DP_OP_1090J1_126_7243_n9, ZN => n7561);
   U8096 : NAND2_X1 port map( A1 => n7561, A2 => n8298, ZN => n8257);
   U8097 : INV_X1 port map( A => n8284, ZN => n7562);
   U8098 : AOI21_X1 port map( B1 => n8241, B2 => n7562, A => n8205, ZN => n7563
                           );
   U8099 : OAI21_X1 port map( B1 => n8241, B2 => n7562, A => n7563, ZN => n7564
                           );
   U8100 : NAND3_X1 port map( A1 => n8202, A2 => n8289, A3 => n8237, ZN => 
                           n7565);
   U8101 : OAI211_X1 port map( C1 => n8238, C2 => n8202, A => n7564, B => n7565
                           , ZN => C620_DATA2_30);
   U8102 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n500, B2 => 
                           DP_OP_751_130_5637_n501, A => DP_OP_751_130_5637_n84
                           , ZN => DP_OP_751_130_5637_n6);
   U8103 : INV_X1 port map( A => n10087, ZN => n7566);
   U8104 : OAI22_X1 port map( A1 => n10182, A2 => n10088, B1 => n10284, B2 => 
                           n7566, ZN => n7567);
   U8105 : AOI21_X1 port map( B1 => n10089, B2 => n10229, A => n7567, ZN => 
                           n7568);
   U8106 : AOI22_X1 port map( A1 => n10090, A2 => n10288, B1 => n10091, B2 => 
                           n7781, ZN => n7569);
   U8107 : OAI21_X1 port map( B1 => n10086, B2 => n10085, A => n10084, ZN => 
                           n7570);
   U8108 : NAND3_X1 port map( A1 => n7568, A2 => n7569, A3 => n7570, ZN => 
                           n10358);
   U8109 : OAI21_X1 port map( B1 => n10451, B2 => n10449, A => n10448, ZN => 
                           n7571);
   U8110 : INV_X1 port map( A => n10395, ZN => n7572);
   U8111 : AOI222_X1 port map( A1 => n10392, A2 => n7571, B1 => n10392, B2 => 
                           n8093, C1 => n7571, C2 => n7572, ZN => n10416);
   U8112 : INV_X1 port map( A => n9586, ZN => n7573);
   U8113 : AOI21_X1 port map( B1 => n9652, B2 => n10472, A => n7573, ZN => 
                           n10839);
   U8114 : INV_X1 port map( A => n8218, ZN => n7574);
   U8115 : OAI221_X1 port map( B1 => n7574, B2 => n10645, C1 => n7574, C2 => 
                           n10642, A => n8448, ZN => n10632);
   U8116 : XOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_17_port, Z => n7575);
   U8117 : OAI21_X1 port map( B1 => n8189, B2 => n7575, A => n10730, ZN => 
                           n7576);
   U8118 : AOI21_X1 port map( B1 => n8189, B2 => n7575, A => n7576, ZN => 
                           DRAMRF_ADDRESS_17_port);
   U8119 : XOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_26_port, Z => n7577);
   U8120 : OAI21_X1 port map( B1 => n8088, B2 => n7940, A => n7939, ZN => n7578
                           );
   U8121 : OAI21_X1 port map( B1 => n7577, B2 => n7578, A => n10730, ZN => 
                           n7579);
   U8122 : AOI21_X1 port map( B1 => n7577, B2 => n7578, A => n7579, ZN => 
                           DRAMRF_ADDRESS_26_port);
   U8123 : INV_X1 port map( A => n10740, ZN => n7580);
   U8124 : AOI22_X1 port map( A1 => n10740, A2 => n8415, B1 => n6015, B2 => 
                           n7580, ZN => n8966);
   U8125 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_A_14_port, A2 => n8674, 
                           B1 => DataPath_i_PIPLIN_IN1_14_port, B2 => n8314, ZN
                           => n7581);
   U8126 : INV_X1 port map( A => n7581, ZN => n10377);
   U8127 : OR4_X1 port map( A1 => IR_9_port, A2 => IR_10_port, A3 => IR_6_port,
                           A4 => IR_8_port, ZN => n7582);
   U8128 : NOR2_X1 port map( A1 => IR_7_port, A2 => n7582, ZN => n10742);
   U8129 : NOR2_X1 port map( A1 => n8455, A2 => n10832, ZN => n7583);
   U8130 : AOI21_X1 port map( B1 => IRAM_DATA(29), B2 => n8580, A => n7583, ZN 
                           => n8478);
   U8131 : NAND2_X1 port map( A1 => n10710, A2 => n8185, ZN => n7584);
   U8132 : NAND3_X1 port map( A1 => n7584, A2 => n10541, A3 => n10542, ZN => 
                           CU_I_CW_16_port);
   U8133 : AND2_X1 port map( A1 => n8694, A2 => 
                           DataPath_RF_internal_out2_0_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N4);
   U8134 : AND2_X1 port map( A1 => n8695, A2 => 
                           DataPath_RF_internal_out1_31_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N35);
   U8135 : OAI22_X1 port map( A1 => n8485, A2 => n8559, B1 => n9659, B2 => 
                           n8562, ZN => n7585);
   U8136 : XNOR2_X1 port map( A => n8263, B => n7585, ZN => n7586);
   U8137 : XOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_10_port, B => 
                           n8265, Z => n7587);
   U8138 : XOR2_X1 port map( A => n7586, B => n7587, Z => 
                           DP_OP_751_130_5637_n1710);
   U8139 : NOR2_X1 port map( A1 => n7586, A2 => n7587, ZN => 
                           DP_OP_751_130_5637_n1709);
   U8140 : INV_X1 port map( A => n10884, ZN => n7588);
   U8141 : AOI21_X1 port map( B1 => n10881, B2 => n7588, A => n10882, ZN => 
                           n7589);
   U8142 : NOR2_X1 port map( A1 => n10883, A2 => n7589, ZN => n7590);
   U8143 : AOI221_X1 port map( B1 => n7590, B2 => n10885, C1 => n10886, C2 => 
                           n10885, A => n10880, ZN => n7591);
   U8144 : NOR2_X1 port map( A1 => n7591, A2 => n10887, ZN => n10920);
   U8145 : OAI21_X1 port map( B1 => n8011, B2 => n8681, A => n9629, ZN => n9781
                           );
   U8146 : INV_X1 port map( A => n8247, ZN => n7592);
   U8147 : OAI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n72, B2 => 
                           DataPath_WRF_CUhw_curr_addr_30_port, A => n8241, ZN 
                           => n7593);
   U8148 : NAND2_X1 port map( A1 => n7593, A2 => n7592, ZN => n8243);
   U8149 : OAI22_X1 port map( A1 => n8299, A2 => n11852, B1 => n8442, B2 => 
                           n11851, ZN => n7594);
   U8150 : AOI211_X1 port map( C1 => n8969, C2 => n8531, A => RST, B => n7594, 
                           ZN => n11715);
   U8151 : NOR2_X1 port map( A1 => n8901, A2 => n11753, ZN => n7595);
   U8152 : AOI21_X1 port map( B1 => n11754, B2 => n8531, A => n7595, ZN => 
                           n11642);
   U8153 : INV_X1 port map( A => DP_OP_751_130_5637_n842, ZN => n7596);
   U8154 : INV_X1 port map( A => n8268, ZN => n7597);
   U8155 : OAI21_X1 port map( B1 => n8268, B2 => DP_OP_751_130_5637_n842, A => 
                           DP_OP_751_130_5637_n907, ZN => n7598);
   U8156 : OAI21_X1 port map( B1 => n7596, B2 => n7597, A => n7598, ZN => 
                           DP_OP_751_130_5637_n807);
   U8157 : INV_X1 port map( A => n10197, ZN => n7599);
   U8158 : OAI21_X1 port map( B1 => n9679, B2 => n7599, A => n9683, ZN => n9682
                           );
   U8159 : NOR2_X1 port map( A1 => n7762, A2 => n11632, ZN => n7600);
   U8160 : AOI21_X1 port map( B1 => n11633, B2 => n8771, A => n7600, ZN => 
                           n12098);
   U8161 : NOR2_X1 port map( A1 => n7762, A2 => n11931, ZN => n7601);
   U8162 : AOI21_X1 port map( B1 => n11631, B2 => n8771, A => n7601, ZN => 
                           n12097);
   U8163 : OAI21_X1 port map( B1 => n8681, B2 => n7818, A => n9619, ZN => n7602
                           );
   U8164 : INV_X1 port map( A => n7602, ZN => n10091);
   U8165 : OAI21_X1 port map( B1 => n9562, B2 => n8681, A => n9540, ZN => n9921
                           );
   U8166 : OAI22_X1 port map( A1 => n7796, A2 => n10010, B1 => n7755, B2 => 
                           n10044, ZN => n7603);
   U8167 : XNOR2_X1 port map( A => n7979, B => n7603, ZN => 
                           DP_OP_751_130_5637_n1771);
   U8168 : INV_X1 port map( A => n8326, ZN => n7604);
   U8169 : NOR2_X1 port map( A1 => n9282, A2 => n7604, ZN => n10687);
   U8170 : NAND3_X1 port map( A1 => IRAM_ADDRESS_28_port, A2 => 
                           IRAM_ADDRESS_29_port, A3 => n10580, ZN => n7605);
   U8171 : NOR2_X1 port map( A1 => n10590, A2 => n7605, ZN => n10833);
   U8172 : NOR2_X1 port map( A1 => n7792, A2 => n9794, ZN => n7606);
   U8173 : NAND2_X1 port map( A1 => n7792, A2 => n9794, ZN => n7607);
   U8174 : AOI22_X1 port map( A1 => n7606, A2 => n10469, B1 => n7608, B2 => 
                           n10458, ZN => n7609);
   U8175 : INV_X1 port map( A => n7607, ZN => n7608);
   U8176 : OAI211_X1 port map( C1 => n7792, C2 => n9794, A => n10468, B => 
                           n7607, ZN => n7610);
   U8177 : AOI21_X1 port map( B1 => n9793, B2 => n9792, A => n9842, ZN => n7611
                           );
   U8178 : OAI21_X1 port map( B1 => n9793, B2 => n9792, A => n7611, ZN => n7612
                           );
   U8179 : AOI21_X1 port map( B1 => n9792, B2 => n9791, A => n9854, ZN => n7613
                           );
   U8180 : OAI21_X1 port map( B1 => n9792, B2 => n9791, A => n7613, ZN => n7614
                           );
   U8181 : NAND4_X1 port map( A1 => n7609, A2 => n7610, A3 => n7612, A4 => 
                           n7614, ZN => n8164);
   U8182 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n604, A2 => 
                           DP_OP_751_130_5637_n702, ZN => n8272);
   U8183 : NOR2_X1 port map( A1 => n8683, A2 => n8344, ZN => n7615);
   U8184 : AOI21_X1 port map( B1 => n8683, B2 => DataPath_i_PIPLIN_IN2_13_port,
                           A => n7615, ZN => n7793);
   U8185 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n162, A2 => n8270, ZN =>
                           n7616);
   U8186 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n161, A2 => n7616, ZN =>
                           DP_OP_751_130_5637_n156);
   U8187 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_A_1_port, A2 => n8671, B1
                           => DataPath_i_PIPLIN_IN1_1_port, B2 => n8314, ZN => 
                           n7617);
   U8188 : INV_X1 port map( A => n7617, ZN => n10487);
   U8189 : NAND3_X1 port map( A1 => DRAMRF_READY, A2 => n8979, A3 => n8712, ZN 
                           => n7618);
   U8190 : OAI21_X1 port map( B1 => n10868, B2 => n8713, A => n7618, ZN => 
                           n10734);
   U8191 : NAND3_X1 port map( A1 => DataPath_RF_POP_ADDRGEN_curr_addr_15_port, 
                           A2 => n10852, A3 => DRAMRF_READY, ZN => n12058);
   U8192 : INV_X1 port map( A => n210, ZN => n7619);
   U8193 : OR3_X1 port map( A1 => n10780, A2 => n12029, A3 => n7619, ZN => 
                           n12027);
   U8194 : XOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_16_port, Z => n7620);
   U8195 : OAI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n17, B2 => n7620, A 
                           => n10730, ZN => n7621);
   U8196 : AOI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n17, B2 => n7620, A 
                           => n7621, ZN => DRAMRF_ADDRESS_16_port);
   U8197 : AOI221_X1 port map( B1 => DP_OP_1090J1_126_7243_n72, B2 => n8189, C1
                           => DataPath_WRF_CUhw_curr_addr_17_port, C2 => n8189,
                           A => n8295, ZN => n7622);
   U8198 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_18_port, ZN => n7623);
   U8199 : OAI21_X1 port map( B1 => n7622, B2 => n7623, A => n10730, ZN => 
                           n7624);
   U8200 : AOI21_X1 port map( B1 => n7622, B2 => n7623, A => n7624, ZN => 
                           DRAMRF_ADDRESS_18_port);
   U8201 : XOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_19_port, Z => n7625);
   U8202 : OAI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n14, B2 => n7625, A 
                           => n10730, ZN => n7626);
   U8203 : AOI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n14, B2 => n7625, A 
                           => n7626, ZN => DRAMRF_ADDRESS_19_port);
   U8204 : XOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_22_port, Z => n7627);
   U8205 : OAI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n11, B2 => n7627, A 
                           => n10730, ZN => n7628);
   U8206 : AOI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n11, B2 => n7627, A 
                           => n7628, ZN => DRAMRF_ADDRESS_22_port);
   U8207 : XOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_24_port, Z => n7629);
   U8208 : OAI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n9, B2 => n7629, A =>
                           n10730, ZN => n7630);
   U8209 : AOI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n9, B2 => n7629, A =>
                           n7630, ZN => DRAMRF_ADDRESS_24_port);
   U8210 : XOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_25_port, Z => n7631);
   U8211 : OAI21_X1 port map( B1 => n8257, B2 => n7631, A => n10730, ZN => 
                           n7632);
   U8212 : AOI21_X1 port map( B1 => n8257, B2 => n7631, A => n7632, ZN => 
                           DRAMRF_ADDRESS_25_port);
   U8213 : AOI21_X1 port map( B1 => n8204, B2 => n7935, A => n7766, ZN => n7633
                           );
   U8214 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_28_port, ZN => n7634);
   U8215 : NOR2_X1 port map( A1 => n7633, A2 => n7634, ZN => n7635);
   U8216 : AOI211_X1 port map( C1 => n7633, C2 => n7634, A => n7773, B => n7635
                           , ZN => DRAMRF_ADDRESS_28_port);
   U8217 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n435, B2 => 
                           DP_OP_751_130_5637_n434, A => n7680, ZN => n7636);
   U8218 : OAI21_X1 port map( B1 => n7637, B2 => n7638, A => n7636, ZN => 
                           DP_OP_751_130_5637_n399);
   U8219 : INV_X1 port map( A => DP_OP_751_130_5637_n434, ZN => n7637);
   U8220 : INV_X1 port map( A => DP_OP_751_130_5637_n435, ZN => n7638);
   U8221 : INV_X1 port map( A => n10740, ZN => n7639);
   U8222 : AOI22_X1 port map( A1 => n10740, A2 => n8414, B1 => n6089, B2 => 
                           n7639, ZN => n8963);
   U8223 : NAND2_X1 port map( A1 => n10011, A2 => n9969, ZN => n7640);
   U8224 : OAI221_X1 port map( B1 => n7790, B2 => n10011, C1 => n9969, C2 => 
                           DP_OP_751_130_5637_n639, A => n7640, ZN => n9511);
   U8225 : AOI22_X1 port map( A1 => n8682, A2 => DataPath_i_PIPLIN_IN2_6_port, 
                           B1 => DataPath_i_PIPLIN_B_6_port, B2 => n8165, ZN =>
                           n7641);
   U8226 : INV_X1 port map( A => n7641, ZN => n9626);
   U8227 : AOI211_X1 port map( C1 => n10421, C2 => n10465, A => n8488, B => 
                           n8167, ZN => n7642);
   U8228 : NAND2_X1 port map( A1 => n10465, A2 => n10484, ZN => n7643);
   U8229 : INV_X1 port map( A => n7796, ZN => n7644);
   U8230 : INV_X1 port map( A => n9533, ZN => n7645);
   U8231 : OAI221_X1 port map( B1 => n7796, B2 => n7643, C1 => n7644, C2 => 
                           n10469, A => n7645, ZN => n7646);
   U8232 : OAI211_X1 port map( C1 => DP_OP_751_130_5637_n1795, C2 => n8076, A 
                           => n8578, B => DP_OP_751_130_5637_n198, ZN => n7647)
                           ;
   U8233 : OAI211_X1 port map( C1 => n10483, C2 => n9572, A => n7646, B => 
                           n7647, ZN => n7648);
   U8234 : AOI211_X1 port map( C1 => DataPath_ALUhw_MULT_mux_out_0_0_port, C2 
                           => n10458, A => n7642, B => n7648, ZN => n7649);
   U8235 : INV_X1 port map( A => n8438, ZN => n7650);
   U8236 : INV_X1 port map( A => DataPath_i_LGET_0_port, ZN => n7651);
   n7652 <= '0';
   U8238 : AOI22_X1 port map( A1 => i_SEL_LGET_0_port, A2 => n8378, B1 => 
                           i_SEL_LGET_1_port, B2 => n494, ZN => n7654);
   U8239 : AOI22_X1 port map( A1 => i_SEL_LGET_0_port, A2 => n8386, B1 => n7654
                           , B2 => DataPath_i_LGET_0_port, ZN => n7655);
   U8240 : AOI22_X1 port map( A1 => n8378, A2 => n7653, B1 => n7655, B2 => n235
                           , ZN => n7656);
   U8241 : INV_X1 port map( A => n8380, ZN => n7657);
   U8242 : AOI22_X1 port map( A1 => n8380, A2 => n7649, B1 => n7656, B2 => 
                           n7657, ZN => n7658);
   U8243 : AOI22_X1 port map( A1 => n10281, A2 => n9628, B1 => n7785, B2 => 
                           n9440, ZN => n7659);
   U8244 : INV_X1 port map( A => n10291, ZN => n7660);
   U8245 : INV_X1 port map( A => n10288, ZN => n7661);
   U8246 : AOI21_X1 port map( B1 => n8558, B2 => n10283, A => n7661, ZN => 
                           n7662);
   U8247 : OAI22_X1 port map( A1 => n9980, A2 => n8489, B1 => n9434, B2 => 
                           n10274, ZN => n7663);
   U8248 : AOI211_X1 port map( C1 => n9433, C2 => n7660, A => n7662, B => n7663
                           , ZN => n7664);
   U8249 : INV_X1 port map( A => n10493, ZN => n7665);
   U8250 : AOI21_X1 port map( B1 => n7659, B2 => n7664, A => n7665, ZN => n7666
                           );
   U8251 : AOI22_X1 port map( A1 => n10510, A2 => n10497, B1 => n10498, B2 => 
                           n10501, ZN => n7667);
   U8252 : OAI21_X1 port map( B1 => n10480, B2 => n10505, A => n7667, ZN => 
                           n7668);
   U8253 : AOI211_X1 port map( C1 => n10477, C2 => n10476, A => n7666, B => 
                           n7668, ZN => n7669);
   U8254 : AOI22_X1 port map( A1 => n10504, A2 => n10495, B1 => n10503, B2 => 
                           n10494, ZN => n7670);
   U8255 : AOI22_X1 port map( A1 => n10509, A2 => n10499, B1 => n10502, B2 => 
                           n10496, ZN => n7671);
   U8256 : NAND3_X1 port map( A1 => n7669, A2 => n7670, A3 => n7671, ZN => 
                           n7672);
   U8257 : AOI22_X1 port map( A1 => n10848, A2 => n7658, B1 => n10840, B2 => 
                           n7672, ZN => n7673);
   U8258 : OAI21_X1 port map( B1 => n495, B2 => n12092, A => n7673, ZN => n7020
                           );
   U8259 : OAI211_X1 port map( C1 => CU_I_CW_6_port, C2 => n10541, A => n10715,
                           B => n10542, ZN => n7674);
   U8260 : AND3_X1 port map( A1 => n8080, A2 => n10543, A3 => n8308, ZN => 
                           n7675);
   U8261 : NOR2_X1 port map( A1 => n7675, A2 => n7674, ZN => n8440);
   U8262 : NAND3_X1 port map( A1 => n9324, A2 => n9321, A3 => n10632, ZN => 
                           n7676);
   U8263 : OAI211_X1 port map( C1 => n9321, C2 => n9324, A => n7676, B => 
                           n10554, ZN => n7677);
   U8264 : AOI22_X1 port map( A1 => n10835, A2 => IRAM_ADDRESS_17_port, B1 => 
                           i_RD1_17_port, B2 => n12070, ZN => n7678);
   U8265 : OAI21_X1 port map( B1 => n7759, B2 => n7677, A => n7678, ZN => n7042
                           );
   U8266 : AND2_X1 port map( A1 => n8695, A2 => 
                           DataPath_RF_internal_out1_0_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N4);
   U8267 : AND2_X1 port map( A1 => n8694, A2 => 
                           DataPath_RF_internal_out2_31_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N35);
   U8268 : INV_X1 port map( A => n8564, ZN => n8567);
   U8269 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n398, A2 => 
                           DP_OP_751_130_5637_n399, ZN => n7679);
   U8270 : BUF_X1 port map( A => DP_OP_751_130_5637_n499, Z => n7680);
   U8271 : BUF_X1 port map( A => DP_OP_751_130_5637_n75, Z => n7681);
   U8272 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n398, A2 => 
                           DP_OP_751_130_5637_n399, ZN => 
                           DP_OP_751_130_5637_n75);
   U8273 : BUF_X1 port map( A => DP_OP_751_130_5637_n120, Z => n7682);
   U8274 : BUF_X1 port map( A => DP_OP_751_130_5637_n85, Z => n7683);
   U8275 : INV_X2 port map( A => n9450, ZN => n8485);
   U8276 : AND2_X1 port map( A1 => n10574, A2 => n7687, ZN => n7684);
   U8277 : NAND2_X1 port map( A1 => n9271, A2 => n8699, ZN => n7685);
   U8278 : NAND2_X1 port map( A1 => n8456, A2 => n7688, ZN => n7686);
   U8279 : BUF_X1 port map( A => n9232, Z => n7689);
   U8280 : BUF_X1 port map( A => n7696, Z => n7690);
   U8281 : BUF_X1 port map( A => n10649, Z => n7691);
   U8282 : INV_X1 port map( A => n9108, ZN => n7692);
   U8283 : NOR2_X1 port map( A1 => n8985, A2 => n9008, ZN => n7693);
   U8284 : INV_X2 port map( A => n9092, ZN => n9108);
   U8285 : INV_X2 port map( A => n9450, ZN => n9452);
   U8286 : OR2_X2 port map( A1 => DP_OP_751_130_5637_I2, A2 => n9587, ZN => 
                           n9447);
   U8287 : INV_X2 port map( A => n10409, ZN => n10395);
   U8288 : OAI21_X2 port map( B1 => n8088, B2 => n7938, A => n7936, ZN => n7935
                           );
   U8289 : INV_X2 port map( A => n10082, ZN => n8556);
   U8290 : NAND2_X2 port map( A1 => DataPath_i_PIPLIN_A_19_port, A2 => n8672, 
                           ZN => n10143);
   U8291 : INV_X2 port map( A => n10385, ZN => n10386);
   U8292 : NOR2_X2 port map( A1 => n8702, A2 => n185, ZN => n10859);
   U8293 : INV_X2 port map( A => n9919, ZN => n10181);
   U8294 : INV_X2 port map( A => n8561, ZN => n8563);
   U8295 : BUF_X2 port map( A => n9207, Z => n7697);
   U8296 : INV_X4 port map( A => n10463, ZN => n10457);
   U8297 : INV_X2 port map( A => n9596, ZN => n9721);
   U8298 : INV_X2 port map( A => i_ALU_OP_2_port, ZN => n8681);
   U8299 : INV_X4 port map( A => n10487, ZN => n10511);
   U8300 : INV_X2 port map( A => n9664, ZN => n10423);
   U8301 : NOR2_X2 port map( A1 => n8502, A2 => n181, ZN => n8255);
   U8302 : AND2_X4 port map( A1 => n8982, A2 => DataPath_RF_c_swin_4_port, ZN 
                           => n8803);
   U8303 : AND2_X1 port map( A1 => n8982, A2 => DataPath_RF_c_swin_0_port, ZN 
                           => n8771);
   U8304 : BUF_X1 port map( A => n10847, Z => n7764);
   U8305 : AND2_X1 port map( A1 => n8982, A2 => DataPath_RF_c_swin_3_port, ZN 
                           => n8852);
   U8306 : BUF_X1 port map( A => n8852, Z => n7779);
   U8307 : BUF_X1 port map( A => n8852, Z => n7761);
   U8308 : NAND2_X2 port map( A1 => n8673, A2 => DataPath_i_PIPLIN_A_18_port, 
                           ZN => n10197);
   U8309 : INV_X1 port map( A => n10841, ZN => n12093);
   U8310 : XOR2_X1 port map( A => DP_OP_751_130_5637_n1557, B => n10446, Z => 
                           n8575);
   U8311 : INV_X2 port map( A => n8575, ZN => n7694);
   U8312 : CLKBUF_X1 port map( A => n10522, Z => n7695);
   U8313 : NAND2_X1 port map( A1 => n10520, A2 => n9004, ZN => n7696);
   U8314 : NAND2_X1 port map( A1 => n7693, A2 => n8986, ZN => n9207);
   U8315 : NOR2_X1 port map( A1 => n12207, A2 => n10519, ZN => n10522);
   U8316 : AOI21_X2 port map( B1 => n10658, B2 => n9309, A => n9308, ZN => 
                           n10653);
   U8317 : NOR2_X2 port map( A1 => n10716, A2 => n8102, ZN => n10770);
   U8318 : AND2_X4 port map( A1 => n9431, A2 => n9430, ZN => n8559);
   U8319 : AND2_X4 port map( A1 => n9398, A2 => n9397, ZN => n8555);
   U8320 : NAND2_X1 port map( A1 => n10520, A2 => n9004, ZN => n7699);
   U8321 : BUF_X2 port map( A => n8571, Z => n7700);
   U8322 : BUF_X2 port map( A => n8571, Z => n7701);
   DRAMRF_ADDRESS_0_port <= '0';
   DRAMRF_ADDRESS_1_port <= '0';
   U8325 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_25_port, A2 => n8691, ZN => 
                           n7702);
   U8326 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_28_port, A2 => n8690, ZN => 
                           n7703);
   U8327 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_27_port, A2 => n8696, ZN => 
                           n7704);
   U8328 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_24_port, A2 => n8696, ZN => 
                           n7705);
   U8329 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_23_port, A2 => n8698, ZN => 
                           n7706);
   U8330 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_26_port, A2 => n8697, ZN => 
                           n7707);
   U8331 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_22_port, A2 => n8692, ZN => 
                           n7708);
   U8332 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_21_port, A2 => n8689, ZN => 
                           n7709);
   U8333 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_20_port, A2 => n8695, ZN => 
                           n7710);
   U8334 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_18_port, A2 => n8691, ZN => 
                           n7711);
   U8335 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_17_port, A2 => n8690, ZN => 
                           n7712);
   U8336 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_19_port, A2 => n8696, ZN => 
                           n7713);
   U8337 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_16_port, A2 => n8698, ZN => 
                           n7714);
   U8338 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_15_port, A2 => n8697, ZN => 
                           n7715);
   U8339 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_14_port, A2 => n8696, ZN => 
                           n7716);
   U8340 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_13_port, A2 => n8696, ZN => 
                           n7717);
   U8341 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_12_port, A2 => n8692, ZN => 
                           n7718);
   U8342 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_11_port, A2 => n8689, ZN => 
                           n7719);
   U8343 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_10_port, A2 => n8696, ZN => 
                           n7720);
   U8344 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_9_port, A2 => n8688, ZN => 
                           n7721);
   U8345 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_8_port, A2 => n8694, ZN => 
                           n7722);
   U8346 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_7_port, A2 => n8695, ZN => 
                           n7723);
   U8347 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_6_port, A2 => n8693, ZN => 
                           n7724);
   U8348 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_5_port, A2 => n8696, ZN => 
                           n7725);
   U8349 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_4_port, A2 => n8691, ZN => 
                           n7726);
   U8350 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_3_port, A2 => n8690, ZN => 
                           n7727);
   U8351 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_2_port, A2 => n8698, ZN => 
                           n7728);
   U8352 : AND2_X1 port map( A1 => n8688, A2 => n5830, ZN => n7729);
   U8353 : AND2_X1 port map( A1 => n8688, A2 => n5794, ZN => n7730);
   U8354 : AND2_X1 port map( A1 => n8688, A2 => n5758, ZN => n7731);
   U8355 : AND2_X1 port map( A1 => n8688, A2 => n5722, ZN => n7732);
   U8356 : AND2_X1 port map( A1 => n8688, A2 => n5686, ZN => n7733);
   U8357 : AND2_X1 port map( A1 => n8688, A2 => n5650, ZN => n7734);
   U8358 : AND2_X1 port map( A1 => n8688, A2 => n5614, ZN => n7735);
   U8359 : AND2_X1 port map( A1 => n8689, A2 => n6146, ZN => n7736);
   U8360 : AND2_X1 port map( A1 => n8688, A2 => n6126, ZN => n7737);
   U8361 : AND2_X1 port map( A1 => n8689, A2 => n6089, ZN => n7738);
   U8362 : AND2_X1 port map( A1 => n8689, A2 => n6052, ZN => n7739);
   U8363 : AND2_X1 port map( A1 => n8689, A2 => n6015, ZN => n7740);
   U8364 : AND2_X1 port map( A1 => n8688, A2 => n5978, ZN => n7741);
   U8365 : AND2_X1 port map( A1 => n8688, A2 => n5941, ZN => n7742);
   U8366 : OR2_X2 port map( A1 => DP_OP_751_130_5637_n400, A2 => 
                           DP_OP_751_130_5637_n498, ZN => n8273);
   U8367 : NOR2_X2 port map( A1 => n10752, A2 => n8503, ZN => n10543);
   U8368 : BUF_X1 port map( A => DP_OP_751_130_5637_n98, Z => n7743);
   U8369 : AOI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n19, B2 => n7746, A 
                           => n7747, ZN => n7745);
   U8370 : OR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_14_port, ZN => n7746);
   U8371 : AND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_14_port, ZN => n7747);
   U8372 : AOI21_X1 port map( B1 => n7743, B2 => n8272, A => n7871, ZN => n7748
                           );
   U8373 : OAI21_X1 port map( B1 => n7935, B2 => n7766, A => n8209, ZN => n8289
                           );
   U8374 : INV_X1 port map( A => DP_OP_751_130_5637_n1794, ZN => n7749);
   U8375 : OAI21_X1 port map( B1 => i_S2, B2 => DataPath_i_PIPLIN_B_1_port, A 
                           => n7831, ZN => DP_OP_751_130_5637_I2);
   U8376 : NOR2_X2 port map( A1 => n9281, A2 => IRAM_ADDRESS_2_port, ZN => 
                           n10692);
   U8377 : NOR2_X2 port map( A1 => i_HAZARD_SIG_CU, A2 => n9274, ZN => n10823);
   U8378 : NOR2_X2 port map( A1 => n8700, A2 => n189, ZN => n10863);
   U8379 : OR2_X1 port map( A1 => n7796, A2 => n9761, ZN => n7750);
   U8380 : INV_X2 port map( A => n8684, ZN => n8683);
   U8381 : INV_X2 port map( A => n8263, ZN => n7828);
   U8382 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1624, A2 => 
                           DP_OP_751_130_5637_n1722, ZN => n7751);
   U8383 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1761, A2 => 
                           DP_OP_751_130_5637_n1794, ZN => n7752);
   U8384 : BUF_X4 port map( A => DP_OP_751_130_5637_n1761, Z => n8263);
   U8385 : OAI21_X2 port map( B1 => DP_OP_751_130_5637_n1047, B2 => n10313, A 
                           => n9485, ZN => n9486);
   U8386 : OAI21_X4 port map( B1 => n415, B2 => n10446, A => n9463, ZN => n8574
                           );
   U8387 : OAI21_X2 port map( B1 => n10217, B2 => n10198, A => n9492, ZN => 
                           n9493);
   U8388 : BUF_X2 port map( A => n9447, Z => n7754);
   U8389 : BUF_X2 port map( A => n9447, Z => n7755);
   U8390 : INV_X2 port map( A => n9651, ZN => n9659);
   U8391 : AND2_X4 port map( A1 => n9351, A2 => n9350, ZN => n9560);
   U8392 : BUF_X2 port map( A => n8505, Z => n7756);
   U8393 : AOI21_X2 port map( B1 => DP_OP_751_130_5637_n82, B2 => n8273, A => 
                           DP_OP_751_130_5637_n79, ZN => DP_OP_751_130_5637_n77
                           );
   U8394 : BUF_X1 port map( A => DP_OP_1090J1_126_7243_n16, Z => n8189);
   U8395 : CLKBUF_X1 port map( A => n10653, Z => n8040);
   U8396 : INV_X1 port map( A => n10552, ZN => n7758);
   U8397 : AND2_X1 port map( A1 => n10702, A2 => i_NPC_SEL, ZN => n12070);
   U8398 : INV_X2 port map( A => n8303, ZN => n7759);
   U8399 : INV_X1 port map( A => n10642, ZN => n7760);
   U8400 : NAND2_X1 port map( A1 => n8192, A2 => n10794, ZN => n10702);
   U8401 : BUF_X2 port map( A => n8579, Z => n8580);
   U8402 : AND2_X1 port map( A1 => n9147, A2 => n7778, ZN => n7964);
   U8403 : NAND2_X1 port map( A1 => n9239, A2 => n9234, ZN => n8105);
   U8404 : NOR2_X1 port map( A1 => n10926, A2 => n10922, ZN => n8595);
   U8405 : NOR2_X1 port map( A1 => n10927, A2 => n10913, ZN => n8581);
   U8406 : NOR2_X1 port map( A1 => n10924, A2 => n10922, ZN => n8597);
   U8407 : NOR2_X1 port map( A1 => n10924, A2 => n10922, ZN => n8598);
   U8408 : INV_X2 port map( A => n11402, ZN => n11401);
   U8409 : INV_X2 port map( A => n11467, ZN => n11466);
   U8410 : INV_X2 port map( A => n11846, ZN => n11845);
   U8411 : INV_X2 port map( A => n11837, ZN => n11836);
   U8412 : INV_X2 port map( A => n11705, ZN => n11704);
   U8413 : INV_X2 port map( A => n11408, ZN => n11407);
   U8414 : INV_X2 port map( A => n11711, ZN => n11710);
   U8415 : NOR2_X1 port map( A1 => RST, A2 => n8657, ZN => n12114);
   U8416 : NOR2_X1 port map( A1 => RST, A2 => n8664, ZN => n12157);
   U8417 : INV_X2 port map( A => n11473, ZN => n11472);
   U8418 : BUF_X2 port map( A => n11820, Z => n7804);
   U8419 : BUF_X2 port map( A => n11814, Z => n7805);
   U8420 : BUF_X2 port map( A => n11781, Z => n7803);
   U8421 : BUF_X2 port map( A => n11426, Z => n7801);
   U8422 : BUF_X2 port map( A => n11765, Z => n7802);
   U8423 : BUF_X2 port map( A => n11821, Z => n7806);
   U8424 : AND2_X2 port map( A1 => n8982, A2 => DataPath_RF_c_swin_1_port, ZN 
                           => n8971);
   U8425 : BUF_X2 port map( A => n8771, Z => n7762);
   U8426 : AND2_X2 port map( A1 => n8982, A2 => DataPath_RF_c_swin_2_port, ZN 
                           => n8901);
   U8427 : NOR2_X1 port map( A1 => n7780, A2 => n10197, ZN => n7887);
   U8428 : INV_X1 port map( A => i_SEL_CMPB, ZN => n8687);
   U8429 : BUF_X2 port map( A => n9474, Z => n7763);
   U8430 : NAND2_X1 port map( A1 => n10520, A2 => n9004, ZN => n8505);
   U8431 : INV_X1 port map( A => n10847, ZN => n12092);
   U8432 : BUF_X1 port map( A => n10847, Z => n7782);
   U8433 : BUF_X1 port map( A => n8572, Z => n7783);
   U8434 : BUF_X1 port map( A => n9625, Z => n8490);
   U8435 : BUF_X2 port map( A => n8572, Z => n7784);
   U8436 : INV_X1 port map( A => n8677, ZN => DP_OP_751_130_5637_n1353);
   U8437 : NOR2_X2 port map( A1 => n8094, A2 => n8681, ZN => n9983);
   U8438 : BUF_X1 port map( A => n10378, Z => n7789);
   U8439 : BUF_X4 port map( A => n12204, Z => n7765);
   U8440 : BUF_X1 port map( A => n9455, Z => n7786);
   U8441 : BUF_X1 port map( A => n10240, Z => n7785);
   U8442 : AOI21_X1 port map( B1 => n8210, B2 => n8291, A => n7799, ZN => n8209
                           );
   U8443 : INV_X2 port map( A => n7793, ZN => DP_OP_751_130_5637_n1251);
   U8444 : BUF_X1 port map( A => n9208, Z => n8106);
   U8445 : OR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_19_port, ZN => n8188);
   U8446 : INV_X1 port map( A => n8291, ZN => n7766);
   U8447 : BUF_X1 port map( A => DP_OP_751_130_5637_n1455, Z => n7798);
   U8448 : INV_X2 port map( A => n9938, ZN => n9944);
   U8449 : BUF_X2 port map( A => n10123, Z => n7795);
   U8450 : OAI21_X1 port map( B1 => n8363, B2 => n8673, A => n9407, ZN => n9669
                           );
   U8451 : INV_X1 port map( A => n9816, ZN => n9817);
   U8452 : OAI21_X2 port map( B1 => n8352, B2 => n8682, A => n9502, ZN => 
                           DP_OP_751_130_5637_n741);
   U8453 : INV_X1 port map( A => n10877, ZN => n7768);
   U8454 : AND2_X2 port map( A1 => n9456, A2 => n7980, ZN => n415);
   U8455 : NAND2_X2 port map( A1 => DataPath_i_PIPLIN_A_23_port, A2 => n8672, 
                           ZN => n10010);
   U8456 : BUF_X2 port map( A => DP_OP_751_130_5637_n1149, Z => n7770);
   U8457 : INV_X1 port map( A => DP_OP_751_130_5637_n1455, ZN => n7771);
   U8458 : INV_X2 port map( A => n10312, ZN => n7772);
   U8459 : NOR2_X1 port map( A1 => n10711, A2 => n8084, ZN => n9275);
   U8460 : INV_X1 port map( A => n10730, ZN => n7773);
   U8461 : INV_X4 port map( A => n8316, ZN => DP_OP_1090J1_126_7243_n72);
   U8462 : INV_X1 port map( A => n8681, ZN => n7800);
   U8463 : INV_X1 port map( A => n8578, ZN => n7774);
   U8464 : BUF_X2 port map( A => n10825, Z => n8185);
   U8465 : INV_X2 port map( A => n8684, ZN => n8682);
   U8466 : NAND2_X1 port map( A1 => n171, A2 => n176, ZN => n10711);
   U8467 : BUF_X2 port map( A => IR_30_port, Z => n8084);
   U8468 : BUF_X1 port map( A => n10592, Z => n8096);
   U8469 : OAI21_X1 port map( B1 => n10645, B2 => n8217, A => n8216, ZN => 
                           n10554);
   U8470 : NAND2_X1 port map( A1 => n10650, A2 => n9314, ZN => n10645);
   U8471 : AND2_X1 port map( A1 => n8444, A2 => n8220, ZN => n8219);
   U8472 : AOI21_X1 port map( B1 => n8216, B2 => n8214, A => n7758, ZN => n8213
                           );
   U8473 : INV_X1 port map( A => n8223, ZN => n8222);
   U8474 : NAND2_X1 port map( A1 => n8223, A2 => n8221, ZN => n8220);
   U8475 : AND2_X1 port map( A1 => n8227, A2 => n8224, ZN => n8223);
   U8476 : NOR2_X1 port map( A1 => n10553, A2 => n8218, ZN => n8214);
   U8477 : AOI21_X1 port map( B1 => n10551, B2 => n10550, A => n8030, ZN => 
                           n10552);
   U8478 : NAND2_X1 port map( A1 => n10590, A2 => n8156, ZN => n8155);
   U8479 : INV_X1 port map( A => n8218, ZN => n8217);
   U8480 : INV_X1 port map( A => n8225, ZN => n8221);
   U8481 : NAND2_X1 port map( A1 => n8225, A2 => n10648, ZN => n8224);
   U8482 : INV_X1 port map( A => n12070, ZN => n8549);
   U8483 : AND2_X1 port map( A1 => n9314, A2 => n8226, ZN => n8225);
   U8484 : INV_X1 port map( A => n10643, ZN => n8226);
   U8485 : NAND2_X1 port map( A1 => n10571, A2 => n10570, ZN => n10590);
   U8486 : AND2_X1 port map( A1 => n10549, A2 => IRAM_ADDRESS_19_port, ZN => 
                           n8030);
   U8487 : INV_X1 port map( A => n8451, ZN => n7775);
   U8488 : INV_X1 port map( A => n10702, ZN => n10835);
   U8489 : NAND2_X1 port map( A1 => n9287, A2 => n226, ZN => n10674);
   U8490 : INV_X1 port map( A => n9303, ZN => n7776);
   U8491 : AND2_X1 port map( A1 => C620_DATA2_27, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_27_port);
   U8492 : OR2_X1 port map( A1 => n8208, A2 => n8203, ZN => n8202);
   U8493 : INV_X1 port map( A => n10668, ZN => n7777);
   U8494 : BUF_X1 port map( A => n8484, Z => n8192);
   U8495 : OR2_X1 port map( A1 => n9315, A2 => n194, ZN => n10638);
   U8496 : NOR2_X1 port map( A1 => n8177, A2 => n10794, ZN => n8579);
   U8497 : BUF_X1 port map( A => n10796, Z => n8177);
   U8498 : BUF_X2 port map( A => n9315, Z => n8484);
   U8499 : BUF_X1 port map( A => DP_OP_751_130_5637_n90, Z => n8056);
   U8500 : NAND2_X1 port map( A1 => n8250, A2 => n9260, ZN => n10523);
   U8501 : XNOR2_X1 port map( A => n7929, B => DP_OP_751_130_5637_n494, ZN => 
                           DP_OP_751_130_5637_n396);
   U8502 : AND2_X1 port map( A1 => n8147, A2 => n8146, ZN => 
                           DP_OP_751_130_5637_n297);
   U8503 : XNOR2_X1 port map( A => n7847, B => DP_OP_751_130_5637_n590, ZN => 
                           DP_OP_751_130_5637_n492);
   U8504 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n591, B => 
                           DP_OP_751_130_5637_n531, ZN => n7847);
   U8505 : NAND2_X1 port map( A1 => n7823, A2 => n8148, ZN => n8147);
   U8506 : NAND2_X1 port map( A1 => n7958, A2 => n7962, ZN => n9193);
   U8507 : NAND2_X1 port map( A1 => n7934, A2 => DP_OP_751_130_5637_n432, ZN =>
                           n7931);
   U8508 : INV_X1 port map( A => DP_OP_751_130_5637_n79, ZN => n7824);
   U8509 : NAND2_X1 port map( A1 => n7969, A2 => n7968, ZN => 
                           DP_OP_751_130_5637_n591);
   U8510 : AND2_X1 port map( A1 => DP_OP_751_130_5637_n400, A2 => 
                           DP_OP_751_130_5637_n498, ZN => 
                           DP_OP_751_130_5637_n79);
   U8511 : OAI21_X1 port map( B1 => n7973, B2 => DP_OP_751_130_5637_n632, A => 
                           n7970, ZN => n7969);
   U8512 : NAND2_X1 port map( A1 => n7930, A2 => n7895, ZN => n7933);
   U8513 : NAND2_X1 port map( A1 => n7973, A2 => DP_OP_751_130_5637_n632, ZN =>
                           n7968);
   U8514 : BUF_X1 port map( A => DP_OP_751_130_5637_n112, Z => n7853);
   U8515 : NAND2_X1 port map( A1 => n7966, A2 => n7965, ZN => 
                           DP_OP_751_130_5637_n689);
   U8516 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n732, B2 => 
                           DP_OP_751_130_5637_n789, A => 
                           DP_OP_751_130_5637_n788, ZN => n7966);
   U8517 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n18, B => n8168, ZN =>
                           C620_DATA2_15);
   U8518 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n790, B => n7967, ZN => 
                           DP_OP_751_130_5637_n692);
   U8519 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n789, A2 => 
                           DP_OP_751_130_5637_n732, ZN => n7965);
   U8520 : NAND2_X1 port map( A1 => n7821, A2 => n7820, ZN => 
                           DP_OP_751_130_5637_n887);
   U8521 : AND2_X1 port map( A1 => n7840, A2 => n7839, ZN => n7842);
   U8522 : AOI21_X1 port map( B1 => n7959, B2 => n9213, A => n9255, ZN => n7957
                           );
   U8523 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n791, B => 
                           DP_OP_751_130_5637_n733, ZN => n7967);
   U8524 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n20, B => n8160, ZN =>
                           C620_DATA2_13);
   U8525 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n19, B => n8166, ZN =>
                           C620_DATA2_14);
   U8526 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n791, A2 => 
                           DP_OP_751_130_5637_n733, ZN => n7974);
   U8527 : AND2_X1 port map( A1 => n7964, A2 => n9192, ZN => n7961);
   U8528 : AOI21_X1 port map( B1 => n8105, B2 => n9114, A => n7841, ZN => n7840
                           );
   U8529 : AOI21_X1 port map( B1 => n9226, B2 => n9225, A => n9224, ZN => n9227
                           );
   U8530 : AND2_X1 port map( A1 => n9201, A2 => n9200, ZN => n9213);
   U8531 : AND2_X1 port map( A1 => n9163, A2 => n7963, ZN => n7962);
   U8532 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n987, A2 => 
                           DP_OP_751_130_5637_n933, ZN => n7820);
   U8533 : NOR2_X1 port map( A1 => n7894, A2 => DP_OP_751_130_5637_n137, ZN => 
                           DP_OP_751_130_5637_n135);
   U8534 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n21, B => n8135, ZN =>
                           C620_DATA2_12);
   U8535 : OAI21_X1 port map( B1 => n7893, B2 => n7894, A => n7892, ZN => 
                           DP_OP_751_130_5637_n131);
   U8536 : INV_X1 port map( A => n9114, ZN => n7843);
   U8537 : INV_X1 port map( A => n9192, ZN => n7960);
   U8538 : INV_X1 port map( A => n9212, ZN => n9215);
   U8539 : NOR3_X1 port map( A1 => n9130, A2 => n9131, A3 => n9139, ZN => n8191
                           );
   U8540 : AND2_X1 port map( A1 => n9223, A2 => n8992, ZN => n9212);
   U8541 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n704, A2 => 
                           DP_OP_751_130_5637_n705, ZN => 
                           DP_OP_751_130_5637_n101);
   U8542 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n897, A2 => 
                           DP_OP_751_130_5637_n837, ZN => n8005);
   U8543 : AND2_X1 port map( A1 => n9051, A2 => n9050, ZN => n8163);
   U8544 : OR3_X1 port map( A1 => n9140, A2 => n9133, A3 => n9141, ZN => n9130)
                           ;
   U8545 : INV_X1 port map( A => n9103, ZN => n7846);
   U8546 : OR2_X1 port map( A1 => n9237, A2 => n9146, ZN => n7963);
   U8547 : OAI22_X1 port map( A1 => i_RD1_13_port, A2 => n9102, B1 => n9097, B2
                           => i_RD1_12_port, ZN => n9103);
   U8548 : INV_X1 port map( A => n9237, ZN => n7778);
   U8549 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n806, A2 => 
                           DP_OP_751_130_5637_n807, ZN => n8274);
   U8550 : NAND2_X1 port map( A1 => n9113, A2 => i_RD1_15_port, ZN => n9238);
   U8551 : OR2_X1 port map( A1 => n9150, A2 => i_RD1_20_port, ZN => n9146);
   U8552 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1283, A2 => 
                           DP_OP_751_130_5637_n1234, ZN => n7889);
   U8553 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1283, B => 
                           DP_OP_751_130_5637_n1234, ZN => n7890);
   U8554 : OR2_X1 port map( A1 => i_RD1_6_port, A2 => n9019, ZN => n9020);
   U8555 : INV_X1 port map( A => n10808, ZN => n10832);
   U8556 : OR2_X1 port map( A1 => n10808, A2 => n12020, ZN => n10794);
   U8557 : NOR2_X2 port map( A1 => n10922, A2 => n10913, ZN => n11239);
   U8558 : NOR2_X2 port map( A1 => n10924, A2 => n10927, ZN => n11247);
   U8559 : NOR2_X2 port map( A1 => n10922, A2 => n10913, ZN => n8583);
   U8560 : NOR2_X2 port map( A1 => n10924, A2 => n10927, ZN => n8594);
   U8561 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_2_port, ZN => n9027
                           );
   U8562 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1279, A2 => 
                           DP_OP_751_130_5637_n1232, ZN => n8043);
   U8563 : NOR2_X2 port map( A1 => n10925, A2 => n10912, ZN => n11236);
   U8564 : NAND2_X1 port map( A1 => n10823, A2 => n9277, ZN => n10808);
   U8565 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1193, A2 => 
                           DP_OP_751_130_5637_n1138, ZN => n8024);
   U8566 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n907, B => n7819, ZN => 
                           DP_OP_751_130_5637_n808);
   U8567 : NOR2_X2 port map( A1 => n10925, A2 => n10912, ZN => n8591);
   U8568 : NAND2_X1 port map( A1 => n8042, A2 => n8041, ZN => 
                           DP_OP_751_130_5637_n1277);
   U8569 : NAND2_X1 port map( A1 => n8071, A2 => n8070, ZN => 
                           DP_OP_751_130_5637_n1381);
   U8570 : NOR2_X2 port map( A1 => n10923, A2 => n10912, ZN => n11241);
   U8571 : NAND2_X1 port map( A1 => n7864, A2 => n7863, ZN => 
                           DP_OP_751_130_5637_n1291);
   U8572 : NOR2_X2 port map( A1 => n10923, A2 => n10912, ZN => n8584);
   U8573 : BUF_X1 port map( A => n11766, Z => n8635);
   U8574 : NAND2_X1 port map( A1 => n7984, A2 => n7983, ZN => 
                           DP_OP_751_130_5637_n1293);
   U8575 : BUF_X1 port map( A => n11425, Z => n8611);
   U8576 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1391, B2 => 
                           DP_OP_751_130_5637_n1339, A => n7865, ZN => n7864);
   U8577 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1481, A2 => 
                           DP_OP_751_130_5637_n1435, ZN => n8070);
   U8578 : NAND2_X1 port map( A1 => n7924, A2 => DP_OP_751_130_5637_n1333, ZN 
                           => n7920);
   U8579 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1332, B2 => 
                           DP_OP_751_130_5637_n1377, A => 
                           DP_OP_751_130_5637_n1376, ZN => n8042);
   U8580 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1377, A2 => 
                           DP_OP_751_130_5637_n1332, ZN => n8041);
   U8581 : OAI21_X1 port map( B1 => n9811, B2 => n10482, A => n8104, ZN => 
                           n8103);
   U8582 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n29, B => n8126, ZN =>
                           C620_DATA2_4);
   U8583 : OAI21_X1 port map( B1 => n9789, B2 => n10482, A => n8128, ZN => 
                           n8127);
   U8584 : NAND2_X1 port map( A1 => n7990, A2 => n7989, ZN => 
                           DP_OP_751_130_5637_n1377);
   U8585 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1393, A2 => 
                           DP_OP_751_130_5637_n1340, ZN => n7983);
   U8586 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1391, A2 => 
                           DP_OP_751_130_5637_n1339, ZN => n7863);
   U8587 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1393, B2 => 
                           DP_OP_751_130_5637_n1340, A => n7985, ZN => n7984);
   U8588 : INV_X1 port map( A => n11817, ZN => n8640);
   U8589 : BUF_X1 port map( A => n11817, Z => n8497);
   U8590 : BUF_X1 port map( A => n11454, Z => n8615);
   U8591 : BUF_X1 port map( A => n12114, Z => n8658);
   U8592 : BUF_X1 port map( A => n11457, Z => n8616);
   U8593 : BUF_X1 port map( A => n12111, Z => n8656);
   U8594 : BUF_X1 port map( A => n11423, Z => n8610);
   U8595 : BUF_X1 port map( A => n12176, Z => n8667);
   U8596 : BUF_X1 port map( A => n11635, Z => n8627);
   U8597 : BUF_X1 port map( A => n12157, Z => n8665);
   U8598 : BUF_X1 port map( A => n11513, Z => n8617);
   U8599 : AND2_X1 port map( A1 => n7927, A2 => n7826, ZN => n7825);
   U8600 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1489, A2 => 
                           DP_OP_751_130_5637_n1439, ZN => n8150);
   U8601 : NAND2_X1 port map( A1 => n7982, A2 => n7981, ZN => 
                           DP_OP_751_130_5637_n1391);
   U8602 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1433, B2 => 
                           DP_OP_751_130_5637_n1477, A => 
                           DP_OP_751_130_5637_n1476, ZN => n7990);
   U8603 : BUF_X1 port map( A => n11431, Z => n8613);
   U8604 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1477, A2 => 
                           DP_OP_751_130_5637_n1433, ZN => n7989);
   U8605 : INV_X1 port map( A => n7811, ZN => DP_OP_751_130_5637_n1317);
   U8606 : BUF_X1 port map( A => n11419, Z => n8609);
   U8607 : BUF_X1 port map( A => n11452, Z => n8614);
   U8608 : BUF_X1 port map( A => n11813, Z => n8638);
   U8609 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1417, B => n7813, ZN => 
                           DP_OP_751_130_5637_n1318);
   U8610 : INV_X2 port map( A => n11429, ZN => n11428);
   U8611 : BUF_X1 port map( A => n11493, Z => n7807);
   U8612 : AOI22_X1 port map( A1 => DP_OP_751_130_5637_n1417, A2 => n7812, B1 
                           => DP_OP_751_130_5637_n1352, B2 => n8258, ZN => 
                           n7811);
   U8613 : BUF_X1 port map( A => n11533, Z => n8620);
   U8614 : BUF_X1 port map( A => n12108, Z => n8654);
   U8615 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1483, A2 => 
                           DP_OP_751_130_5637_n1436, ZN => n7927);
   U8616 : BUF_X1 port map( A => n11873, Z => n7808);
   U8617 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1479, A2 => 
                           DP_OP_751_130_5637_n1434, ZN => n8049);
   U8618 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1475, A2 => 
                           DP_OP_751_130_5637_n1432, ZN => n8065);
   U8619 : BUF_X1 port map( A => n11780, Z => n8636);
   U8620 : NAND2_X1 port map( A1 => n8064, A2 => n8063, ZN => 
                           DP_OP_751_130_5637_n1473);
   U8621 : AND2_X1 port map( A1 => n8697, A2 => n11796, ZN => n11812);
   U8622 : NAND2_X1 port map( A1 => n8060, A2 => n8059, ZN => 
                           DP_OP_751_130_5637_n1475);
   U8623 : BUF_X1 port map( A => n12116, Z => n8659);
   U8624 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1577, A2 => 
                           DP_OP_751_130_5637_n1534, ZN => n8047);
   U8625 : BUF_X1 port map( A => n11430, Z => n8512);
   U8626 : AND2_X2 port map( A1 => n8698, A2 => n11537, ZN => n11535);
   U8627 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1491, A2 => 
                           DP_OP_751_130_5637_n1440, ZN => n7981);
   U8628 : AND2_X2 port map( A1 => n8697, A2 => n11656, ZN => n11659);
   U8629 : NAND2_X1 port map( A1 => n8117, A2 => n8116, ZN => 
                           DP_OP_751_130_5637_n1479);
   U8630 : BUF_X1 port map( A => n12119, Z => n8661);
   U8631 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1581, A2 => 
                           DP_OP_751_130_5637_n1536, ZN => n8077);
   U8632 : BUF_X1 port map( A => n11514, Z => n8522);
   U8633 : AND2_X2 port map( A1 => n8698, A2 => n11584, ZN => n11583);
   U8634 : BUF_X1 port map( A => n11545, Z => n8524);
   U8635 : BUF_X1 port map( A => n11539, Z => n8523);
   U8636 : BUF_X1 port map( A => n12110, Z => n8655);
   U8637 : BUF_X1 port map( A => n11664, Z => n8537);
   U8638 : BUF_X1 port map( A => n12174, Z => n8666);
   U8639 : AND2_X2 port map( A1 => n8697, A2 => n11692, ZN => n11695);
   U8640 : BUF_X1 port map( A => n11662, Z => n8536);
   U8641 : BUF_X1 port map( A => n11422, Z => n8511);
   U8642 : BUF_X1 port map( A => n11634, Z => n8533);
   U8643 : AND2_X2 port map( A1 => n8698, A2 => n11542, ZN => n11541);
   U8644 : AND2_X1 port map( A1 => n8697, A2 => n11774, ZN => n11779);
   U8645 : AND2_X2 port map( A1 => n8698, A2 => n11530, ZN => n11529);
   U8646 : AND2_X2 port map( A1 => n8697, A2 => n11638, ZN => n11652);
   U8647 : BUF_X1 port map( A => n11512, Z => n8521);
   U8648 : AND2_X2 port map( A1 => n8696, A2 => n12153, ZN => n12152);
   U8649 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n37, B => n8145, ZN =>
                           C620_DATA2_2);
   U8650 : NAND2_X1 port map( A1 => n8115, A2 => n8114, ZN => 
                           DP_OP_751_130_5637_n1577);
   U8651 : NAND2_X1 port map( A1 => n8130, A2 => n8129, ZN => 
                           DP_OP_751_130_5637_n1581);
   U8652 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1538, A2 => n7869, ZN 
                           => n7867);
   U8653 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1589, A2 => 
                           DP_OP_751_130_5637_n1540, ZN => n7849);
   U8654 : XNOR2_X1 port map( A => n7817, B => n7816, ZN => 
                           DP_OP_751_130_5637_n1488);
   U8655 : NAND2_X1 port map( A1 => n8000, A2 => n7999, ZN => 
                           DP_OP_751_130_5637_n1491);
   U8656 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1532, A2 => 
                           DP_OP_751_130_5637_n1573, ZN => n8063);
   U8657 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1575, A2 => 
                           DP_OP_751_130_5637_n1533, ZN => n8059);
   U8658 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1668, B => n8058, ZN => 
                           DP_OP_751_130_5637_n1570);
   U8659 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1532, B2 => 
                           DP_OP_751_130_5637_n1573, A => 
                           DP_OP_751_130_5637_n1572, ZN => n8064);
   U8660 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1587, B => 
                           DP_OP_751_130_5637_n1539, ZN => n7817);
   U8661 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1591, A2 => 
                           DP_OP_751_130_5637_n1541, ZN => n7999);
   U8662 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1593, A2 => 
                           DP_OP_751_130_5637_n1542, ZN => n7836);
   U8663 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1587, A2 => 
                           DP_OP_751_130_5637_n1539, ZN => n7814);
   U8664 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1593, B => 
                           DP_OP_751_130_5637_n1542, ZN => n7835);
   U8665 : BUF_X1 port map( A => n8971, Z => n8544);
   U8666 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1579, A2 => 
                           DP_OP_751_130_5637_n1535, ZN => n8116);
   U8667 : BUF_X1 port map( A => n8901, Z => n8532);
   U8668 : NOR2_X1 port map( A1 => n7937, A2 => n8183, ZN => n7936);
   U8669 : BUF_X1 port map( A => n8901, Z => n8531);
   U8670 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1669, B => 
                           DP_OP_751_130_5637_n1631, ZN => n8058);
   U8671 : AOI21_X1 port map( B1 => n9922, B2 => n10113, A => n7887, ZN => 
                           n9754);
   U8672 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1689, B2 => 
                           DP_OP_751_130_5637_n1641, A => 
                           DP_OP_751_130_5637_n1688, ZN => n7998);
   U8673 : OR2_X1 port map( A1 => n7940, A2 => n8184, ZN => n7938);
   U8674 : INV_X1 port map( A => DP_OP_751_130_5637_n1335, ZN => n7826);
   U8675 : NOR2_X1 port map( A1 => n7939, A2 => n8184, ZN => n7937);
   U8676 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1681, A2 => 
                           DP_OP_751_130_5637_n1637, ZN => n8129);
   U8677 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1677, A2 => 
                           DP_OP_751_130_5637_n1635, ZN => n8114);
   U8678 : AND2_X1 port map( A1 => DP_OP_751_130_5637_n1736, A2 => 
                           DP_OP_751_130_5637_n1767, ZN => 
                           DP_OP_751_130_5637_n1675);
   U8679 : AND2_X1 port map( A1 => DP_OP_751_130_5637_n1764, A2 => 
                           DP_OP_751_130_5637_n1733, ZN => 
                           DP_OP_751_130_5637_n1669);
   U8680 : AND2_X1 port map( A1 => DP_OP_751_130_5637_n1737, A2 => 
                           DP_OP_751_130_5637_n1768, ZN => 
                           DP_OP_751_130_5637_n1677);
   U8681 : NOR2_X1 port map( A1 => n7877, A2 => n7878, ZN => 
                           DP_OP_751_130_5637_n1691);
   U8682 : NAND2_X1 port map( A1 => n8724, A2 => n11375, ZN => n8982);
   U8683 : AND2_X1 port map( A1 => DP_OP_751_130_5637_n1739, A2 => 
                           DP_OP_751_130_5637_n1770, ZN => 
                           DP_OP_751_130_5637_n1681);
   U8684 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1689, A2 => 
                           DP_OP_751_130_5637_n1641, ZN => n7997);
   U8685 : AND2_X1 port map( A1 => DP_OP_751_130_5637_n1742, A2 => 
                           DP_OP_751_130_5637_n1773, ZN => 
                           DP_OP_751_130_5637_n1687);
   U8686 : INV_X1 port map( A => n8686, ZN => n8685);
   U8687 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_26_port, B => 
                           n7828, ZN => DP_OP_751_130_5637_n1737);
   U8688 : INV_X1 port map( A => DP_OP_751_130_5637_n1439, ZN => n8153);
   U8689 : AND2_X1 port map( A1 => n8443, A2 => n8713, ZN => n10740);
   U8690 : OR2_X1 port map( A1 => n8228, A2 => n7941, ZN => n7940);
   U8691 : OR2_X1 port map( A1 => n12092, A2 => n516, ZN => n8128);
   U8692 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n740, B => 
                           DP_OP_751_130_5637_n741, ZN => n8033);
   U8693 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n536, B => 
                           DP_OP_751_130_5637_n537, ZN => n8157);
   U8694 : NAND2_X1 port map( A1 => n8239, A2 => n8207, ZN => n8206);
   U8695 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1352, B => n8258, ZN => 
                           n7813);
   U8696 : INV_X1 port map( A => n9766, ZN => n7780);
   U8697 : OR2_X1 port map( A1 => n8231, A2 => n8233, ZN => n8038);
   U8698 : NOR2_X1 port map( A1 => n9009, A2 => n7995, ZN => n10514);
   U8699 : OR2_X1 port map( A1 => n12092, A2 => n515, ZN => n8104);
   U8700 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n332, A2 => 
                           DP_OP_751_130_5637_n333, ZN => n8148);
   U8701 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1352, A2 => n8258, ZN => 
                           n7812);
   U8702 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n434, B => 
                           DP_OP_751_130_5637_n435, ZN => n8173);
   U8703 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n842, B => n8268, ZN => 
                           n7819);
   U8704 : AND2_X1 port map( A1 => n7696, A2 => IRAM_ADDRESS_4_port, ZN => 
                           n7995);
   U8705 : INV_X1 port map( A => n8701, ZN => n8702);
   U8706 : OR2_X1 port map( A1 => n12093, A2 => n7774, ZN => n7954);
   U8707 : INV_X1 port map( A => n10180, ZN => n7781);
   U8708 : NAND2_X1 port map( A1 => n7886, A2 => n7884, ZN => n10199);
   U8709 : INV_X1 port map( A => n7757, ZN => n8711);
   U8710 : NOR2_X1 port map( A1 => n8242, A2 => n8240, ZN => n8239);
   U8711 : NOR2_X1 port map( A1 => n8242, A2 => n8284, ZN => n8237);
   U8712 : AND2_X1 port map( A1 => n8235, A2 => n8243, ZN => n8234);
   U8713 : BUF_X1 port map( A => n8572, Z => n8573);
   U8714 : NOR2_X1 port map( A1 => n8101, A2 => n9105, ZN => n8701);
   U8715 : OR2_X1 port map( A1 => n7883, A2 => n7979, ZN => n8004);
   U8716 : NAND2_X1 port map( A1 => n8244, A2 => n8236, ZN => n8235);
   U8717 : NAND2_X1 port map( A1 => n10468, A2 => n10197, ZN => n7886);
   U8718 : BUF_X2 port map( A => n10378, Z => n8494);
   U8719 : OAI22_X1 port map( A1 => n7755, A2 => n10123, B1 => n8487, B2 => 
                           n8556, ZN => n8017);
   U8720 : BUF_X1 port map( A => n9301, Z => n8101);
   U8721 : INV_X1 port map( A => n7942, ZN => n7941);
   U8722 : NOR2_X1 port map( A1 => n8247, A2 => n8245, ZN => n8244);
   U8723 : OR2_X1 port map( A1 => n8139, A2 => n550, ZN => n8069);
   U8724 : OR2_X1 port map( A1 => n8139, A2 => n546, ZN => n8091);
   U8725 : NAND2_X1 port map( A1 => n8209, A2 => n7766, ZN => n8207);
   U8726 : NAND2_X1 port map( A1 => n8241, A2 => n8284, ZN => n8238);
   U8727 : NAND2_X1 port map( A1 => n9301, A2 => n10720, ZN => n10520);
   U8728 : NAND2_X1 port map( A1 => n9679, A2 => n7885, ZN => n9683);
   U8729 : NOR2_X1 port map( A1 => n8121, A2 => n7944, ZN => n7943);
   U8730 : BUF_X2 port map( A => n10326, Z => n8492);
   U8731 : NAND2_X1 port map( A1 => n10458, A2 => n7885, ZN => n7884);
   U8732 : BUF_X1 port map( A => n9008, Z => n8190);
   U8733 : INV_X2 port map( A => n9208, ZN => n9105);
   U8734 : NAND2_X1 port map( A1 => n8286, A2 => n8288, ZN => n8245);
   U8735 : INV_X1 port map( A => n8284, ZN => n8240);
   U8736 : NAND2_X1 port map( A1 => n8286, A2 => n8246, ZN => n8241);
   U8737 : AND2_X2 port map( A1 => CU_I_CW_MEM_2_port, A2 => n10857, ZN => 
                           n12203);
   U8738 : INV_X1 port map( A => n8087, ZN => n7944);
   U8739 : OR2_X1 port map( A1 => n8186, A2 => n8187, ZN => n8036);
   U8740 : NAND2_X1 port map( A1 => n8288, A2 => n8236, ZN => n8211);
   U8741 : BUF_X2 port map( A => n9625, Z => n7787);
   U8742 : BUF_X2 port map( A => n9454, Z => n7788);
   U8743 : INV_X1 port map( A => n415, ZN => DP_OP_751_130_5637_n1557);
   U8744 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1659, B => n9626, ZN => 
                           n9458);
   U8745 : BUF_X1 port map( A => n10385, Z => n8090);
   U8746 : BUF_X1 port map( A => n9596, Z => n8016);
   U8747 : BUF_X1 port map( A => n8504, Z => n8139);
   U8748 : OR2_X1 port map( A1 => n8487, A2 => n10044, ZN => n7891);
   U8749 : BUF_X1 port map( A => n10409, Z => n8093);
   U8750 : OR2_X1 port map( A1 => n9208, A2 => n548, ZN => n8108);
   U8751 : INV_X1 port map( A => n10197, ZN => n7885);
   U8752 : BUF_X1 port map( A => n10463, Z => n7818);
   U8753 : INV_X1 port map( A => n8263, ZN => n8068);
   U8754 : BUF_X1 port map( A => n9651, Z => n8011);
   U8755 : OR2_X1 port map( A1 => n9208, A2 => n544, ZN => n8107);
   U8756 : BUF_X1 port map( A => n10273, Z => n8094);
   U8757 : INV_X1 port map( A => n7754, ZN => n9446);
   U8758 : INV_X1 port map( A => DP_OP_751_130_5637_n639, ZN => n7790);
   U8759 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_12_port, ZN => n8135);
   U8760 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_13_port, ZN => n8160);
   U8761 : AND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_26_port, ZN => n8183);
   U8762 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_14_port, ZN => n8166);
   U8763 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_15_port, ZN => n8168);
   U8764 : OR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_3_port, ZN => n8201);
   U8765 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_4_port, ZN => n8126);
   U8766 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_2_port, ZN => n8145);
   U8767 : NOR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_27_port, ZN => n8210);
   U8768 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_11_port, ZN => n8019);
   U8769 : AND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_12_port, ZN => n8136);
   U8770 : OR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_12_port, ZN => n8137);
   U8771 : BUF_X1 port map( A => n11933, Z => n11632);
   U8772 : NOR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_16_port, ZN => n8176);
   U8773 : AND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_17_port, ZN => n8295);
   U8774 : AND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_18_port, ZN => n8290);
   U8775 : BUF_X1 port map( A => n11932, Z => n11753);
   U8776 : AND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_23_port, ZN => n8121);
   U8777 : NOR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_26_port, ZN => n8184);
   U8778 : INV_X1 port map( A => n8288, ZN => n7791);
   U8779 : NOR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_28_port, ZN => n8236);
   U8780 : NOR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_29_port, ZN => n8246);
   U8781 : AND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_30_port, ZN => n8247);
   U8782 : BUF_X1 port map( A => n9530, Z => n8487);
   U8783 : BUF_X1 port map( A => DP_OP_751_130_5637_I2, Z => n7979);
   U8784 : NAND2_X1 port map( A1 => n10770, A2 => n10824, ZN => n9208);
   U8785 : NOR2_X1 port map( A1 => n10757, A2 => n8080, ZN => n10824);
   U8786 : INV_X1 port map( A => n9761, ZN => n7792);
   U8787 : OR2_X1 port map( A1 => n12194, A2 => DRAM_READY, ZN => n10877);
   U8788 : BUF_X1 port map( A => n9275, Z => n8110);
   U8789 : NAND2_X2 port map( A1 => n8693, A2 => n11910, ZN => n11911);
   U8790 : NAND2_X2 port map( A1 => n8693, A2 => n11906, ZN => n11907);
   U8791 : NAND3_X1 port map( A1 => n10710, A2 => n8185, A3 => n181, ZN => 
                           n9004);
   U8792 : NAND2_X2 port map( A1 => n8693, A2 => n11915, ZN => n11947);
   U8793 : NAND2_X2 port map( A1 => n8693, A2 => n11890, ZN => n11891);
   U8794 : NAND2_X2 port map( A1 => n8693, A2 => n11902, ZN => n11903);
   U8795 : INV_X1 port map( A => DP_OP_751_130_5637_n1149, ZN => n7794);
   U8796 : BUF_X1 port map( A => n9563, Z => n8099);
   U8797 : NAND2_X2 port map( A1 => n8693, A2 => n11898, ZN => n11899);
   U8798 : BUF_X2 port map( A => n9530, Z => n7796);
   U8799 : NAND2_X2 port map( A1 => n8693, A2 => n11894, ZN => n11895);
   U8800 : AND2_X2 port map( A1 => DataPath_i_PIPLIN_A_21_port, A2 => n8673, ZN
                           => n10082);
   U8801 : INV_X1 port map( A => n9874, ZN => n7797);
   U8802 : BUF_X1 port map( A => n10467, Z => n8015);
   U8803 : INV_X1 port map( A => DP_OP_1090J1_126_7243_n72, ZN => n7799);
   U8804 : BUF_X1 port map( A => IR_26_port, Z => n8062);
   U8805 : OR2_X1 port map( A1 => n8138, A2 => n8339, ZN => n7980);
   U8806 : CLKBUF_X1 port map( A => DataPath_RF_c_win_4_port, Z => n8678);
   U8807 : OR2_X1 port map( A1 => IR_26_port, A2 => n8312, ZN => n10752);
   U8808 : BUF_X1 port map( A => i_S2, Z => n8138);
   U8809 : BUF_X1 port map( A => n8684, Z => n8165);
   U8810 : BUF_X1 port map( A => n171, Z => n8080);
   U8811 : AND2_X1 port map( A1 => n176, A2 => IR_30_port, ZN => n10825);
   U8812 : OR2_X1 port map( A1 => IR_26_port, A2 => n181, ZN => n10716);
   U8813 : BUF_X1 port map( A => n8312, Z => n8102);
   U8814 : NOR3_X2 port map( A1 => i_ADD_WB_3_port, A2 => n8310, A3 => n8409, 
                           ZN => n11456);
   U8815 : BUF_X1 port map( A => n11819, Z => n8641);
   U8816 : BUF_X1 port map( A => n11663, Z => n8633);
   U8817 : BUF_X1 port map( A => n12113, Z => n8657);
   U8818 : BUF_X1 port map( A => n12156, Z => n8664);
   U8819 : BUF_X1 port map( A => n11655, Z => n8630);
   U8820 : BUF_X1 port map( A => n11782, Z => n8637);
   U8821 : BUF_X1 port map( A => n11661, Z => n8632);
   U8822 : BUF_X1 port map( A => n11637, Z => n8628);
   U8823 : BUF_X1 port map( A => n12117, Z => n8660);
   U8824 : BUF_X1 port map( A => n11538, Z => n8622);
   U8825 : BUF_X1 port map( A => n11544, Z => n8624);
   U8826 : BUF_X1 port map( A => n11815, Z => n8639);
   U8827 : BUF_X1 port map( A => n11822, Z => n8642);
   U8828 : INV_X1 port map( A => n11818, ZN => n11817);
   U8829 : BUF_X1 port map( A => n12120, Z => n8662);
   U8830 : NOR2_X2 port map( A1 => RST, A2 => n11646, ZN => n11737);
   U8831 : NOR2_X2 port map( A1 => RST, A2 => n11640, ZN => n11728);
   U8832 : NOR2_X2 port map( A1 => RST, A2 => n11647, ZN => n11738);
   U8833 : NOR2_X2 port map( A1 => RST, A2 => n11645, ZN => n11736);
   U8834 : NOR2_X2 port map( A1 => RST, A2 => n11641, ZN => n11731);
   U8835 : NOR2_X2 port map( A1 => RST, A2 => n11643, ZN => n11733);
   U8836 : NOR2_X2 port map( A1 => RST, A2 => n11639, ZN => n11726);
   U8837 : NOR2_X2 port map( A1 => RST, A2 => n11642, ZN => n11732);
   U8838 : NOR2_X2 port map( A1 => RST, A2 => n11644, ZN => n11735);
   U8839 : NOR3_X2 port map( A1 => n8376, A2 => n11270, A3 => n11260, ZN => 
                           n11304);
   U8840 : INV_X2 port map( A => DataPath_RF_c_win_2_port, ZN => n11596);
   U8841 : NOR2_X2 port map( A1 => RST, A2 => n11772, ZN => n11877);
   U8842 : NOR2_X2 port map( A1 => RST, A2 => n11768, ZN => n11868);
   U8843 : BUF_X1 port map( A => n11636, Z => n8534);
   U8844 : OAI22_X2 port map( A1 => n9637, A2 => n8900, B1 => n12109, B2 => 
                           n8442, ZN => n11636);
   U8845 : BUF_X1 port map( A => n11458, Z => n8514);
   U8846 : OAI22_X2 port map( A1 => n9644, A2 => n8802, B1 => n577, B2 => 
                           n12158, ZN => n11458);
   U8847 : BUF_X1 port map( A => n11453, Z => n8513);
   U8848 : OAI22_X2 port map( A1 => n9642, A2 => n8802, B1 => n577, B2 => 
                           n12155, ZN => n11453);
   U8849 : OAI22_X2 port map( A1 => n9637, A2 => n8802, B1 => n577, B2 => 
                           n12109, ZN => n11422);
   U8850 : INV_X1 port map( A => n8793, ZN => n9637);
   U8851 : BUF_X1 port map( A => n11654, Z => n8535);
   U8852 : OAI22_X2 port map( A1 => n9639, A2 => n8900, B1 => n12115, B2 => 
                           n8442, ZN => n11654);
   U8853 : OAI22_X2 port map( A1 => n9640, A2 => n8802, B1 => n577, B2 => 
                           n12118, ZN => n11430);
   U8854 : INV_X1 port map( A => n8796, ZN => n9640);
   U8855 : OAI22_X2 port map( A1 => n9642, A2 => n8900, B1 => n12155, B2 => 
                           n8442, ZN => n11664);
   U8856 : INV_X1 port map( A => n8797, ZN => n9642);
   U8857 : AOI22_X2 port map( A1 => n8932, A2 => n3340, B1 => n11933, B2 => 
                           n8965, ZN => n11875);
   U8858 : AOI22_X2 port map( A1 => n8932, A2 => n3350, B1 => n11923, B2 => 
                           n8965, ZN => n11865);
   U8859 : AOI22_X2 port map( A1 => n8791, A2 => n3337, B1 => n11936, B2 => 
                           n8802, ZN => n11498);
   U8860 : AOI22_X2 port map( A1 => n8791, A2 => n3335, B1 => n11938, B2 => 
                           n8802, ZN => n11500);
   U8861 : AOI22_X2 port map( A1 => n8791, A2 => n3341, B1 => n11932, B2 => 
                           n8802, ZN => n11494);
   U8862 : AOI22_X2 port map( A1 => n8791, A2 => n3345, B1 => n11928, B2 => 
                           n8802, ZN => n11490);
   U8863 : AOI22_X2 port map( A1 => n8791, A2 => n3347, B1 => n11926, B2 => 
                           n8802, ZN => n11488);
   U8864 : AOI22_X2 port map( A1 => n8791, A2 => n3332, B1 => n11941, B2 => 
                           n8802, ZN => n11503);
   U8865 : OAI22_X2 port map( A1 => n8791, A2 => n11945, B1 => n3328, B2 => 
                           n8802, ZN => n11507);
   U8866 : OAI22_X2 port map( A1 => n8791, A2 => n11933, B1 => n3340, B2 => 
                           n8802, ZN => n11495);
   U8867 : OAI22_X2 port map( A1 => n8791, A2 => n11937, B1 => n3336, B2 => 
                           n8802, ZN => n11499);
   U8868 : OAI22_X2 port map( A1 => n8791, A2 => n11935, B1 => n3338, B2 => 
                           n8802, ZN => n11497);
   U8869 : OAI22_X2 port map( A1 => n8791, A2 => n11946, B1 => n3327, B2 => 
                           n8802, ZN => n11508);
   U8870 : INV_X8 port map( A => n12207, ZN => n10872);
   U8871 : INV_X8 port map( A => n12206, ZN => n10871);
   U8872 : AOI211_X2 port map( C1 => n10232, C2 => n10276, A => n9719, B => 
                           n9718, ZN => n9946);
   U8873 : BUF_X1 port map( A => n11591, Z => n8626);
   U8874 : BUF_X1 port map( A => n11515, Z => n8618);
   U8875 : NOR2_X2 port map( A1 => RST, A2 => n11651, ZN => n11746);
   U8876 : NOR2_X2 port map( A1 => RST, A2 => n11649, ZN => n11743);
   U8877 : NOR2_X2 port map( A1 => RST, A2 => n11648, ZN => n11741);
   U8878 : NOR2_X2 port map( A1 => RST, A2 => n11528, ZN => n11627);
   U8879 : NOR2_X2 port map( A1 => n12093, A2 => n10452, ZN => n10840);
   U8880 : AOI221_X2 port map( B1 => n495, B2 => n11331, C1 => n11261, C2 => 
                           n11331, A => n11305, ZN => n11307);
   U8881 : NOR2_X2 port map( A1 => RST, A2 => n11776, ZN => n11885);
   U8882 : NOR2_X2 port map( A1 => RST, A2 => n11778, ZN => n11888);
   U8883 : NOR2_X2 port map( A1 => RST, A2 => n11777, ZN => n11887);
   U8884 : NOR2_X2 port map( A1 => RST, A2 => n11775, ZN => n11883);
   U8885 : NOR2_X2 port map( A1 => RST, A2 => n11773, ZN => n11879);
   U8886 : NOR2_X2 port map( A1 => RST, A2 => n11769, ZN => n11870);
   U8887 : NOR2_X2 port map( A1 => RST, A2 => n12105, ZN => n12173);
   U8888 : NOR2_X2 port map( A1 => RST, A2 => n11650, ZN => n11745);
   U8889 : NOR2_X2 port map( A1 => RST, A2 => n12099, ZN => n12162);
   U8890 : NOR2_X2 port map( A1 => RST, A2 => n12095, ZN => n12187);
   U8891 : NOR2_X2 port map( A1 => RST, A2 => n12103, ZN => n12170);
   U8892 : NOR2_X2 port map( A1 => RST, A2 => n12096, ZN => n12189);
   U8893 : NOR2_X2 port map( A1 => RST, A2 => n12097, ZN => n12192);
   U8894 : NOR2_X2 port map( A1 => RST, A2 => n12098, ZN => n12160);
   U8895 : NOR2_X2 port map( A1 => RST, A2 => n12102, ZN => n12165);
   U8896 : NOR2_X2 port map( A1 => RST, A2 => n12104, ZN => n12172);
   U8897 : NOR3_X2 port map( A1 => n7800, A2 => i_ALU_OP_3_port, A3 => n368, ZN
                           => n12089);
   U8898 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n332, A2 => 
                           DP_OP_751_130_5637_n333, ZN => n8146);
   U8899 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n332, B => 
                           DP_OP_751_130_5637_n333, ZN => n8149);
   U8900 : NOR2_X2 port map( A1 => n10855, A2 => n12045, ZN => n11391);
   U8901 : NOR2_X2 port map( A1 => RST, A2 => n11798, ZN => n11878);
   U8902 : NOR2_X2 port map( A1 => RST, A2 => n11770, ZN => n11874);
   U8903 : NOR2_X2 port map( A1 => RST, A2 => n11801, ZN => n11880);
   U8904 : NOR2_X2 port map( A1 => RST, A2 => n12140, ZN => n12164);
   U8905 : NOR2_X2 port map( A1 => RST, A2 => n12100, ZN => n12163);
   U8906 : NOR2_X2 port map( A1 => RST, A2 => n12145, ZN => n12168);
   U8907 : OAI22_X2 port map( A1 => n9644, A2 => n8851, B1 => n11596, B2 => 
                           n12158, ZN => n11545);
   U8908 : INV_X1 port map( A => n8852, ZN => n8851);
   U8909 : INV_X1 port map( A => n8798, ZN => n9644);
   U8910 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n638, B => 
                           DP_OP_751_130_5637_n639, ZN => n8100);
   U8911 : AOI22_X2 port map( A1 => DataPath_RF_POP_ADDRGEN_curr_state_0_port, 
                           A2 => n851, B1 => n10852, B2 => n12047, ZN => n11376
                           );
   U8912 : INV_X1 port map( A => n11377, ZN => n12047);
   U8913 : OAI21_X2 port map( B1 => n9643, B2 => n3324, A => n8749, ZN => 
                           n12175);
   U8914 : NOR2_X2 port map( A1 => n10284, A2 => n12087, ZN => n10288);
   U8915 : OAI22_X2 port map( A1 => n9641, A2 => n8900, B1 => n12121, B2 => 
                           n8442, ZN => n11662);
   U8916 : OAI22_X2 port map( A1 => n9636, A2 => n8900, B1 => n12094, B2 => 
                           n8442, ZN => n11634);
   U8917 : INV_X1 port map( A => n8901, ZN => n8900);
   U8918 : INV_X1 port map( A => n8772, ZN => n9636);
   U8919 : AOI22_X2 port map( A1 => n8932, A2 => n3339, B1 => n11934, B2 => 
                           n8965, ZN => n11876);
   U8920 : INV_X1 port map( A => n8971, ZN => n8965);
   U8921 : OAI22_X2 port map( A1 => n8791, A2 => n11943, B1 => n3330, B2 => 
                           n8802, ZN => n11505);
   U8922 : OAI22_X2 port map( A1 => n8727, A2 => n11932, B1 => n3341, B2 => 
                           n9643, ZN => n12159);
   U8923 : INV_X1 port map( A => n8771, ZN => n9643);
   U8924 : OAI21_X2 port map( B1 => n8402, B2 => n8683, A => n9520, ZN => 
                           DP_OP_751_130_5637_n435);
   U8925 : OAI21_X2 port map( B1 => n8355, B2 => n8683, A => n9513, ZN => 
                           DP_OP_751_130_5637_n537);
   U8926 : XNOR2_X1 port map( A => n7809, B => DP_OP_751_130_5637_n594, ZN => 
                           n8181);
   U8927 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n595, B => 
                           DP_OP_751_130_5637_n533, ZN => n7809);
   U8928 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n497, B2 => 
                           DP_OP_751_130_5637_n433, A => n8181, ZN => n7827);
   U8929 : XNOR2_X1 port map( A => n7810, B => n7830, ZN => 
                           DP_OP_751_130_5637_n1686);
   U8930 : XNOR2_X1 port map( A => n7829, B => n7828, ZN => n7830);
   U8931 : INV_X1 port map( A => DP_OP_751_130_5637_n1772, ZN => n7810);
   U8932 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_2_port, B => 
                           n8068, ZN => DP_OP_751_130_5637_n1760);
   U8933 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1685, A2 => 
                           DP_OP_751_130_5637_n1639, ZN => n8012);
   U8934 : OAI21_X1 port map( B1 => n7962, B2 => n7960, A => n7744, ZN => n7959
                           );
   U8935 : AND2_X1 port map( A1 => DP_OP_751_130_5637_n1740, A2 => 
                           DP_OP_751_130_5637_n1771, ZN => 
                           DP_OP_751_130_5637_n1683);
   U8936 : OAI22_X1 port map( A1 => n9454, A2 => n10143, B1 => n7795, B2 => 
                           n8569, ZN => DataPath_ALUhw_MULT_mux_out_2_24_port);
   U8937 : XNOR2_X1 port map( A => n7852, B => DP_OP_751_130_5637_n1588, ZN => 
                           DP_OP_751_130_5637_n1490);
   U8938 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1440, B2 => 
                           DP_OP_751_130_5637_n1491, A => 
                           DP_OP_751_130_5637_n1490, ZN => n7982);
   U8939 : OAI22_X1 port map( A1 => n8569, A2 => n8556, B1 => n9454, B2 => 
                           n7795, ZN => DataPath_ALUhw_MULT_mux_out_2_25_port);
   U8940 : INV_X1 port map( A => DP_OP_751_130_5637_n1775, ZN => n7877);
   U8941 : NAND2_X1 port map( A1 => n7815, A2 => n7814, ZN => 
                           DP_OP_751_130_5637_n1487);
   U8942 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1539, B2 => 
                           DP_OP_751_130_5637_n1587, A => n7816, ZN => n7815);
   U8943 : XNOR2_X1 port map( A => n8013, B => DP_OP_751_130_5637_n1684, ZN => 
                           n7816);
   U8944 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_18_port, B => 
                           n8068, ZN => DP_OP_751_130_5637_n1745);
   U8945 : NAND2_X1 port map( A1 => n7998, A2 => n7997, ZN => 
                           DP_OP_751_130_5637_n1589);
   U8946 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1589, B => 
                           DP_OP_751_130_5637_n1540, ZN => n7852);
   U8947 : NAND3_X1 port map( A1 => DP_OP_751_130_5637_n77, A2 => 
                           DP_OP_751_130_5637_n72, A3 => DP_OP_751_130_5637_n76
                           , ZN => n7910);
   U8948 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n986, B => n7822, ZN => 
                           DP_OP_751_130_5637_n888);
   U8949 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n987, B => 
                           DP_OP_751_130_5637_n933, ZN => n7822);
   U8950 : XNOR2_X1 port map( A => n7823, B => n8149, ZN => 
                           DP_OP_751_130_5637_n298);
   U8951 : NAND2_X1 port map( A1 => n7827, A2 => n8180, ZN => n7823);
   U8952 : NAND2_X1 port map( A1 => n8273, A2 => n7824, ZN => 
                           DP_OP_751_130_5637_n5);
   U8953 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n499, B => n8173, ZN => 
                           DP_OP_751_130_5637_n400);
   U8954 : OAI22_X1 port map( A1 => n8566, A2 => n10143, B1 => n7795, B2 => 
                           n9452, ZN => n7829);
   U8955 : AND2_X1 port map( A1 => DP_OP_751_130_5637_n1772, A2 => n7830, ZN =>
                           DP_OP_751_130_5637_n1685);
   U8956 : NAND2_X1 port map( A1 => n8333, A2 => i_S2, ZN => n7831);
   U8957 : NAND2_X1 port map( A1 => n7832, A2 => n7836, ZN => 
                           DP_OP_751_130_5637_n1493);
   U8958 : NAND2_X1 port map( A1 => n7833, A2 => DP_OP_751_130_5637_n1592, ZN 
                           => n7832);
   U8959 : NAND2_X1 port map( A1 => n7834, A2 => n7837, ZN => n7833);
   U8960 : INV_X1 port map( A => DP_OP_751_130_5637_n1593, ZN => n7834);
   U8961 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1592, B => n7835, ZN => 
                           DP_OP_751_130_5637_n1494);
   U8962 : INV_X1 port map( A => DP_OP_751_130_5637_n1542, ZN => n7837);
   U8963 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n104, A2 => n8269, ZN =>
                           n8039);
   U8964 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n704, A2 => 
                           DP_OP_751_130_5637_n705, ZN => n8269);
   U8965 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n107, B2 => 
                           DP_OP_751_130_5637_n105, A => 
                           DP_OP_751_130_5637_n106, ZN => 
                           DP_OP_751_130_5637_n104);
   U8966 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n804, A2 => 
                           DP_OP_751_130_5637_n706, ZN => 
                           DP_OP_751_130_5637_n105);
   U8967 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n805, B => n8033, ZN => 
                           DP_OP_751_130_5637_n706);
   U8968 : AOI21_X1 port map( B1 => n8274, B2 => DP_OP_751_130_5637_n112, A => 
                           n7838, ZN => DP_OP_751_130_5637_n107);
   U8969 : INV_X1 port map( A => DP_OP_751_130_5637_n111, ZN => n7838);
   U8970 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n113, B2 => 
                           DP_OP_751_130_5637_n115, A => 
                           DP_OP_751_130_5637_n114, ZN => 
                           DP_OP_751_130_5637_n112);
   U8971 : INV_X1 port map( A => n9238, ZN => n7841);
   U8972 : NAND3_X1 port map( A1 => n9089, A2 => n7846, A3 => n9114, ZN => 
                           n7839);
   U8973 : OAI21_X1 port map( B1 => n7844, B2 => n7843, A => n7842, ZN => n8134
                           );
   U8974 : NAND2_X1 port map( A1 => n9091, A2 => n7845, ZN => n7844);
   U8975 : AND2_X1 port map( A1 => n9090, A2 => n7846, ZN => n7845);
   U8976 : NAND2_X1 port map( A1 => n7848, A2 => n8153, ZN => n8152);
   U8977 : INV_X1 port map( A => DP_OP_751_130_5637_n1489, ZN => n7848);
   U8978 : NAND2_X1 port map( A1 => n7850, A2 => n7849, ZN => 
                           DP_OP_751_130_5637_n1489);
   U8979 : NAND2_X1 port map( A1 => n7851, A2 => DP_OP_751_130_5637_n1588, ZN 
                           => n7850);
   U8980 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1589, A2 => 
                           DP_OP_751_130_5637_n1540, ZN => n7851);
   U8981 : INV_X1 port map( A => n7078, ZN => n7854);
   U8982 : NAND2_X1 port map( A1 => n7867, A2 => n7855, ZN => 
                           DP_OP_751_130_5637_n1485);
   U8983 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1538, B2 => n7869, A =>
                           DP_OP_751_130_5637_n1584, ZN => n7855);
   U8984 : NAND2_X1 port map( A1 => n7856, A2 => n8012, ZN => n7869);
   U8985 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1685, B2 => 
                           DP_OP_751_130_5637_n1639, A => 
                           DP_OP_751_130_5637_n1684, ZN => n7856);
   U8986 : OR2_X1 port map( A1 => n7914, A2 => DP_OP_751_130_5637_n297, ZN => 
                           DP_OP_751_130_5637_n69);
   U8987 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n394, B => n7857, ZN => 
                           n7914);
   U8988 : XNOR2_X1 port map( A => n7874, B => n7753, ZN => n7857);
   U8989 : NAND2_X1 port map( A1 => n7859, A2 => n7858, ZN => 
                           DP_OP_751_130_5637_n1483);
   U8990 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1583, A2 => 
                           DP_OP_751_130_5637_n1537, ZN => n7858);
   U8991 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1537, B2 => 
                           DP_OP_751_130_5637_n1583, A => n8132, ZN => n7859);
   U8992 : XNOR2_X1 port map( A => n7860, B => DP_OP_751_130_5637_n1680, ZN => 
                           n8132);
   U8993 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1681, B => 
                           DP_OP_751_130_5637_n1637, ZN => n7860);
   U8994 : XNOR2_X1 port map( A => n7862, B => n7861, ZN => 
                           DP_OP_751_130_5637_n1537);
   U8995 : INV_X1 port map( A => n8261, ZN => n7861);
   U8996 : OAI22_X1 port map( A1 => n7783, A2 => n10197, B1 => n10143, B2 => 
                           n7701, ZN => n7862);
   U8997 : XNOR2_X1 port map( A => n7866, B => n7865, ZN => 
                           DP_OP_751_130_5637_n1292);
   U8998 : XNOR2_X1 port map( A => n8154, B => DP_OP_751_130_5637_n1488, ZN => 
                           n7865);
   U8999 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1391, B => 
                           DP_OP_751_130_5637_n1339, ZN => n7866);
   U9000 : AND2_X2 port map( A1 => n9451, A2 => n8095, ZN => n8564);
   U9001 : NAND2_X1 port map( A1 => n7930, A2 => n8179, ZN => n7934);
   U9002 : XNOR2_X1 port map( A => n7868, B => DP_OP_751_130_5637_n1584, ZN => 
                           DP_OP_751_130_5637_n1486);
   U9003 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1538, B => n7869, ZN => 
                           n7868);
   U9004 : XNOR2_X1 port map( A => n8079, B => DP_OP_751_130_5637_n1740, ZN => 
                           DP_OP_751_130_5637_n1684);
   U9005 : AOI21_X1 port map( B1 => DP_OP_751_130_5637_n90, B2 => n8271, A => 
                           n7870, ZN => DP_OP_751_130_5637_n85);
   U9006 : INV_X1 port map( A => DP_OP_751_130_5637_n89, ZN => n7870);
   U9007 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n600, A2 => 
                           DP_OP_751_130_5637_n502, ZN => 
                           DP_OP_751_130_5637_n89);
   U9008 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n601, B => n8157, ZN => 
                           DP_OP_751_130_5637_n502);
   U9009 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n93, B2 => 
                           DP_OP_751_130_5637_n91, A => DP_OP_751_130_5637_n92,
                           ZN => DP_OP_751_130_5637_n90);
   U9010 : AOI21_X1 port map( B1 => DP_OP_751_130_5637_n98, B2 => n8272, A => 
                           n7871, ZN => DP_OP_751_130_5637_n93);
   U9011 : INV_X1 port map( A => DP_OP_751_130_5637_n97, ZN => n7871);
   U9012 : NAND2_X1 port map( A1 => n8039, A2 => DP_OP_751_130_5637_n101, ZN =>
                           DP_OP_751_130_5637_n98);
   U9013 : XNOR2_X1 port map( A => n7872, B => DP_OP_751_130_5637_n1480, ZN => 
                           n8072);
   U9014 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1481, B => 
                           DP_OP_751_130_5637_n1435, ZN => n7872);
   U9015 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n101, A2 => n8269, ZN =>
                           DP_OP_751_130_5637_n10);
   U9016 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1192, B => n7873, ZN => 
                           DP_OP_751_130_5637_n1094);
   U9017 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1193, B => 
                           DP_OP_751_130_5637_n1138, ZN => n7873);
   U9018 : NAND2_X1 port map( A1 => n7932, A2 => n7931, ZN => n7874);
   U9019 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1591, B2 => 
                           DP_OP_751_130_5637_n1541, A => n8001, ZN => n8000);
   U9020 : XNOR2_X1 port map( A => n7875, B => DP_OP_751_130_5637_n1688, ZN => 
                           n8001);
   U9021 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1689, B => 
                           DP_OP_751_130_5637_n1641, ZN => n7875);
   U9022 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_2_21_port, B => 
                           n7876, ZN => DP_OP_751_130_5637_n1641);
   U9023 : INV_X1 port map( A => DP_OP_751_130_5637_n1659, ZN => n7876);
   U9024 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n604, A2 => 
                           DP_OP_751_130_5637_n702, ZN => 
                           DP_OP_751_130_5637_n97);
   U9025 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n703, B => n8100, ZN => 
                           DP_OP_751_130_5637_n604);
   U9026 : XNOR2_X1 port map( A => n7878, B => DP_OP_751_130_5637_n1775, ZN => 
                           DP_OP_751_130_5637_n1692);
   U9027 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_19_port, B => 
                           n8263, ZN => n7878);
   U9028 : NAND2_X1 port map( A1 => n7880, A2 => n7928, ZN => n7879);
   U9029 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1483, A2 => 
                           DP_OP_751_130_5637_n1436, ZN => n7880);
   U9030 : XNOR2_X1 port map( A => n8078, B => DP_OP_751_130_5637_n1580, ZN => 
                           n7928);
   U9031 : XNOR2_X1 port map( A => n7881, B => DP_OP_751_130_5637_n1131, ZN => 
                           n7905);
   U9032 : NAND2_X1 port map( A1 => n7882, A2 => n8043, ZN => n7881);
   U9033 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1232, B2 => 
                           DP_OP_751_130_5637_n1279, A => n8044, ZN => n7882);
   U9034 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n602, A2 => 
                           DP_OP_751_130_5637_n603, ZN => 
                           DP_OP_751_130_5637_n91);
   U9035 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1483, B => 
                           DP_OP_751_130_5637_n1436, ZN => n7926);
   U9036 : NAND2_X1 port map( A1 => n7979, A2 => n7883, ZN => n8003);
   U9037 : OAI22_X1 port map( A1 => n7755, A2 => n9979, B1 => n7796, B2 => 
                           n9944, ZN => n7883);
   U9038 : NAND2_X1 port map( A1 => n7889, A2 => n7888, ZN => 
                           DP_OP_751_130_5637_n1183);
   U9039 : XNOR2_X1 port map( A => n7890, B => DP_OP_751_130_5637_n1282, ZN => 
                           DP_OP_751_130_5637_n1184);
   U9040 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_27_port, B => 
                           n7979, ZN => DP_OP_751_130_5637_n1767);
   U9041 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_22_port, ZN => 
                           DP_OP_751_130_5637_n1807);
   U9042 : OAI21_X1 port map( B1 => n8556, B2 => n7755, A => n7891, ZN => 
                           DataPath_ALUhw_MULT_mux_out_0_22_port);
   U9043 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n133, A2 => 
                           DP_OP_751_130_5637_n134, ZN => n7892);
   U9044 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n139, A2 => 
                           DP_OP_751_130_5637_n134, ZN => n7893);
   U9045 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n129, B2 => 
                           DP_OP_751_130_5637_n131, A => 
                           DP_OP_751_130_5637_n130, ZN => 
                           DP_OP_751_130_5637_n128);
   U9046 : AND2_X1 port map( A1 => n8277, A2 => DP_OP_751_130_5637_n140, ZN => 
                           n7894);
   U9047 : NOR2_X1 port map( A1 => DP_OP_751_130_5637_n1012, A2 => 
                           DP_OP_751_130_5637_n1110, ZN => 
                           DP_OP_751_130_5637_n129);
   U9048 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n595, A2 => 
                           DP_OP_751_130_5637_n533, ZN => n8179);
   U9049 : NAND2_X1 port map( A1 => n7897, A2 => n7896, ZN => 
                           DP_OP_751_130_5637_n791);
   U9050 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n891, A2 => 
                           DP_OP_751_130_5637_n834, ZN => n7896);
   U9051 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n834, B2 => 
                           DP_OP_751_130_5637_n891, A => 
                           DP_OP_751_130_5637_n890, ZN => n7897);
   U9052 : XNOR2_X1 port map( A => n7898, B => DP_OP_751_130_5637_n890, ZN => 
                           DP_OP_751_130_5637_n792);
   U9053 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n891, B => 
                           DP_OP_751_130_5637_n834, ZN => n7898);
   U9054 : NAND2_X1 port map( A1 => n7900, A2 => n7899, ZN => n6993);
   U9055 : AOI21_X1 port map( B1 => n8164, B2 => n10841, A => n8103, ZN => 
                           n7899);
   U9056 : NAND2_X1 port map( A1 => n7902, A2 => n7901, ZN => n7900);
   U9057 : NOR2_X1 port map( A1 => n12093, A2 => n7774, ZN => n7901);
   U9058 : XNOR2_X1 port map( A => n7903, B => n7904, ZN => n7902);
   U9059 : OAI21_X1 port map( B1 => n7681, B2 => DP_OP_751_130_5637_n77, A => 
                           DP_OP_751_130_5637_n76, ZN => n7903);
   U9060 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n201, A2 => 
                           DP_OP_751_130_5637_n72, ZN => n7904);
   U9061 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1178, B => n7905, ZN => 
                           DP_OP_751_130_5637_n1080);
   U9062 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1279, B => 
                           DP_OP_751_130_5637_n1232, ZN => n8046);
   U9063 : NAND2_X1 port map( A1 => n7920, A2 => n7906, ZN => 
                           DP_OP_751_130_5637_n1279);
   U9064 : OAI21_X1 port map( B1 => n7924, B2 => DP_OP_751_130_5637_n1333, A =>
                           n7921, ZN => n7906);
   U9065 : XNOR2_X1 port map( A => n7922, B => DP_OP_751_130_5637_n1476, ZN => 
                           n7921);
   U9066 : NAND2_X1 port map( A1 => n8065, A2 => n7907, ZN => 
                           DP_OP_751_130_5637_n1375);
   U9067 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1475, B2 => 
                           DP_OP_751_130_5637_n1432, A => n8066, ZN => n7907);
   U9068 : XNOR2_X1 port map( A => n7908, B => DP_OP_751_130_5637_n1572, ZN => 
                           n8066);
   U9069 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1573, B => 
                           DP_OP_751_130_5637_n1532, ZN => n7908);
   U9070 : OAI211_X1 port map( C1 => n7955, C2 => n7911, A => n7910, B => n7909
                           , ZN => n7915);
   U9071 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n72, A2 => 
                           DP_OP_751_130_5637_n71, ZN => n7909);
   U9072 : INV_X1 port map( A => DP_OP_751_130_5637_n72, ZN => n7911);
   U9073 : XNOR2_X1 port map( A => n7915, B => n7912, ZN => n7945);
   U9074 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n69, A2 => n7913, ZN => 
                           n7912);
   U9075 : NAND2_X1 port map( A1 => n7914, A2 => DP_OP_751_130_5637_n297, ZN =>
                           n7913);
   U9076 : NAND2_X1 port map( A1 => n7917, A2 => n8077, ZN => 
                           DP_OP_751_130_5637_n1481);
   U9077 : NAND2_X1 port map( A1 => n7916, A2 => DP_OP_751_130_5637_n1580, ZN 
                           => n7917);
   U9078 : NAND2_X1 port map( A1 => n7919, A2 => n7918, ZN => n7916);
   U9079 : INV_X1 port map( A => DP_OP_751_130_5637_n1536, ZN => n7918);
   U9080 : INV_X1 port map( A => DP_OP_751_130_5637_n1581, ZN => n7919);
   U9081 : XNOR2_X1 port map( A => n7923, B => n7921, ZN => 
                           DP_OP_751_130_5637_n1280);
   U9082 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1477, B => 
                           DP_OP_751_130_5637_n1433, ZN => n7922);
   U9083 : NAND2_X1 port map( A1 => n8048, A2 => n8047, ZN => 
                           DP_OP_751_130_5637_n1477);
   U9084 : XNOR2_X1 port map( A => n7924, B => DP_OP_751_130_5637_n1333, ZN => 
                           n7923);
   U9085 : NAND2_X1 port map( A1 => n8049, A2 => n7925, ZN => n7924);
   U9086 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1479, B2 => 
                           DP_OP_751_130_5637_n1434, A => n8050, ZN => n7925);
   U9087 : XNOR2_X1 port map( A => n8051, B => DP_OP_751_130_5637_n1576, ZN => 
                           n8050);
   U9088 : XNOR2_X1 port map( A => n7926, B => n7928, ZN => 
                           DP_OP_751_130_5637_n1384);
   U9089 : XNOR2_X1 port map( A => n7934, B => DP_OP_751_130_5637_n432, ZN => 
                           n7929);
   U9090 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n494, A2 => n7933, ZN =>
                           n7932);
   U9091 : OAI21_X1 port map( B1 => n7945, B2 => n7954, A => n7953, ZN => n6992
                           );
   U9092 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1086, B => n7946, ZN => 
                           DP_OP_751_130_5637_n988);
   U9093 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1087, B => 
                           DP_OP_751_130_5637_n1034, ZN => n7946);
   U9094 : OAI21_X1 port map( B1 => n7948, B2 => n10513, A => n7947, ZN => 
                           n6994);
   U9095 : AND2_X1 port map( A1 => n9834, A2 => n9835, ZN => n7947);
   U9096 : AOI21_X1 port map( B1 => n7950, B2 => n8578, A => n7949, ZN => n7948
                           );
   U9097 : XNOR2_X1 port map( A => n7952, B => n7951, ZN => n7950);
   U9098 : INV_X1 port map( A => DP_OP_751_130_5637_n77, ZN => n7951);
   U9099 : NAND2_X1 port map( A1 => n7679, A2 => DP_OP_751_130_5637_n76, ZN => 
                           n7952);
   U9100 : AOI21_X1 port map( B1 => n9712, B2 => n10841, A => n8127, ZN => 
                           n7953);
   U9101 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n76, A2 => 
                           DP_OP_751_130_5637_n75, ZN => n7955);
   U9102 : NAND2_X1 port map( A1 => n9232, A2 => n7964, ZN => n7958);
   U9103 : NAND2_X1 port map( A1 => n7956, A2 => n7957, ZN => n9228);
   U9104 : NAND3_X1 port map( A1 => n9232, A2 => n7961, A3 => n9213, ZN => 
                           n7956);
   U9105 : XNOR2_X1 port map( A => n7972, B => n7970, ZN => 
                           DP_OP_751_130_5637_n592);
   U9106 : XNOR2_X1 port map( A => n7971, B => DP_OP_751_130_5637_n788, ZN => 
                           n7970);
   U9107 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n789, B => 
                           DP_OP_751_130_5637_n732, ZN => n7971);
   U9108 : XNOR2_X1 port map( A => n7973, B => DP_OP_751_130_5637_n632, ZN => 
                           n7972);
   U9109 : NAND2_X1 port map( A1 => n7975, A2 => n7974, ZN => n7973);
   U9110 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n790, A2 => n7976, ZN =>
                           n7975);
   U9111 : NAND2_X1 port map( A1 => n7978, A2 => n7977, ZN => n7976);
   U9112 : INV_X1 port map( A => DP_OP_751_130_5637_n733, ZN => n7977);
   U9113 : INV_X1 port map( A => DP_OP_751_130_5637_n791, ZN => n7978);
   U9114 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_17_port, B => 
                           n7828, ZN => DP_OP_751_130_5637_n1746);
   U9115 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1681, A2 => 
                           DP_OP_751_130_5637_n1637, ZN => n8131);
   U9116 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1579, B2 => 
                           DP_OP_751_130_5637_n1535, A => n8118, ZN => n8117);
   U9117 : XNOR2_X1 port map( A => n7987, B => n7985, ZN => 
                           DP_OP_751_130_5637_n1294);
   U9118 : XNOR2_X1 port map( A => n7986, B => DP_OP_751_130_5637_n1490, ZN => 
                           n7985);
   U9119 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1491, B => 
                           DP_OP_751_130_5637_n1440, ZN => n7986);
   U9120 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1393, B => 
                           DP_OP_751_130_5637_n1340, ZN => n7987);
   U9121 : XNOR2_X1 port map( A => n7988, B => n8068, ZN => 
                           DP_OP_751_130_5637_n1739);
   U9122 : OAI22_X1 port map( A1 => n8565, A2 => n8556, B1 => n8485, B2 => 
                           n10044, ZN => n7988);
   U9123 : NOR2_X1 port map( A1 => n8467, A2 => n7991, ZN => n8466);
   U9124 : NAND2_X1 port map( A1 => n7993, A2 => n7992, ZN => n7991);
   U9125 : INV_X1 port map( A => n10604, ZN => n7992);
   U9126 : NAND2_X1 port map( A1 => n10600, A2 => n10603, ZN => n7993);
   U9127 : BUF_X1 port map( A => n10700, Z => n7994);
   U9128 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1577, B2 => 
                           DP_OP_751_130_5637_n1534, A => 
                           DP_OP_751_130_5637_n1576, ZN => n8048);
   U9129 : XNOR2_X1 port map( A => n7996, B => n7828, ZN => 
                           DP_OP_751_130_5637_n1738);
   U9130 : OAI22_X1 port map( A1 => n8566, A2 => n8553, B1 => n9452, B2 => 
                           n10010, ZN => n7996);
   U9131 : XNOR2_X1 port map( A => n8002, B => n8001, ZN => 
                           DP_OP_751_130_5637_n1492);
   U9132 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1591, B => 
                           DP_OP_751_130_5637_n1541, ZN => n8002);
   U9133 : NAND2_X1 port map( A1 => n8004, A2 => n8003, ZN => 
                           DP_OP_751_130_5637_n1769);
   U9134 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1677, B2 => 
                           DP_OP_751_130_5637_n1635, A => 
                           DP_OP_751_130_5637_n1676, ZN => n8115);
   U9135 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n897, B => 
                           DP_OP_751_130_5637_n837, ZN => n8010);
   U9136 : XNOR2_X1 port map( A => n8010, B => DP_OP_751_130_5637_n896, ZN => 
                           DP_OP_751_130_5637_n798);
   U9137 : NAND2_X1 port map( A1 => n8006, A2 => n8005, ZN => 
                           DP_OP_751_130_5637_n797);
   U9138 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n896, A2 => n8007, ZN =>
                           n8006);
   U9139 : NAND2_X1 port map( A1 => n8009, A2 => n8008, ZN => n8007);
   U9140 : INV_X1 port map( A => DP_OP_751_130_5637_n837, ZN => n8008);
   U9141 : INV_X1 port map( A => DP_OP_751_130_5637_n897, ZN => n8009);
   U9142 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1685, B => 
                           DP_OP_751_130_5637_n1639, ZN => n8013);
   U9143 : XNOR2_X1 port map( A => n8014, B => n7828, ZN => 
                           DP_OP_751_130_5637_n1742);
   U9144 : OAI22_X1 port map( A1 => n8567, A2 => n10197, B1 => n9452, B2 => 
                           n10143, ZN => n8014);
   U9145 : XNOR2_X1 port map( A => n8017, B => n7979, ZN => 
                           DP_OP_751_130_5637_n1773);
   U9146 : BUF_X1 port map( A => n10658, Z => n8018);
   U9147 : INV_X1 port map( A => n8020, ZN => DP_OP_1090J1_126_7243_n20);
   U9148 : AOI21_X1 port map( B1 => DP_OP_1090J1_126_7243_n21, B2 => n8137, A 
                           => n8136, ZN => n8020);
   U9149 : OAI21_X1 port map( B1 => n8023, B2 => n8022, A => n8021, ZN => 
                           DP_OP_1090J1_126_7243_n21);
   U9150 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_11_port, ZN => n8021);
   U9151 : NOR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_11_port, ZN => n8022);
   U9152 : INV_X1 port map( A => DP_OP_1090J1_126_7243_n22, ZN => n8023);
   U9153 : NAND2_X1 port map( A1 => n8025, A2 => n8024, ZN => 
                           DP_OP_751_130_5637_n1093);
   U9154 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1192, A2 => n8026, ZN 
                           => n8025);
   U9155 : NAND2_X1 port map( A1 => n8028, A2 => n8027, ZN => n8026);
   U9156 : INV_X1 port map( A => DP_OP_751_130_5637_n1138, ZN => n8027);
   U9157 : INV_X1 port map( A => DP_OP_751_130_5637_n1193, ZN => n8028);
   U9158 : BUF_X1 port map( A => n9296, Z => n8029);
   U9159 : BUF_X1 port map( A => n10671, Z => n8031);
   U9160 : XNOR2_X1 port map( A => n8032, B => n8068, ZN => 
                           DP_OP_751_130_5637_n1740);
   U9161 : OAI22_X1 port map( A1 => n8565, A2 => n7795, B1 => n8485, B2 => 
                           n8556, ZN => n8032);
   U9162 : BUF_X1 port map( A => n9305, Z => n8034);
   U9163 : XNOR2_X1 port map( A => n8035, B => n7828, ZN => 
                           DP_OP_751_130_5637_n1736);
   U9164 : OAI22_X1 port map( A1 => n8563, A2 => n9979, B1 => n9452, B2 => 
                           n9944, ZN => n8035);
   U9165 : NAND2_X1 port map( A1 => n8037, A2 => n8036, ZN => 
                           DP_OP_1090J1_126_7243_n13);
   U9166 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n14, A2 => n8188, ZN 
                           => n8037);
   U9167 : NOR2_X1 port map( A1 => n8230, A2 => n8038, ZN => 
                           DP_OP_1090J1_126_7243_n14);
   U9168 : INV_X4 port map( A => n8676, ZN => DP_OP_751_130_5637_n1659);
   U9169 : NAND2_X1 port map( A1 => n8151, A2 => n8150, ZN => 
                           DP_OP_751_130_5637_n1389);
   U9170 : XNOR2_X1 port map( A => n8046, B => n8044, ZN => 
                           DP_OP_751_130_5637_n1180);
   U9171 : XNOR2_X1 port map( A => n8045, B => DP_OP_751_130_5637_n1376, ZN => 
                           n8044);
   U9172 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1377, B => 
                           DP_OP_751_130_5637_n1332, ZN => n8045);
   U9173 : XNOR2_X1 port map( A => n8052, B => n8050, ZN => 
                           DP_OP_751_130_5637_n1380);
   U9174 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1577, B => 
                           DP_OP_751_130_5637_n1534, ZN => n8051);
   U9175 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1479, B => 
                           DP_OP_751_130_5637_n1434, ZN => n8052);
   U9176 : BUF_X1 port map( A => DP_OP_751_130_5637_n107, Z => n8053);
   U9177 : NAND2_X1 port map( A1 => n7684, A2 => n7686, ZN => n10580);
   U9178 : XNOR2_X1 port map( A => n8054, B => DP_OP_751_130_5637_n1742, ZN => 
                           DP_OP_751_130_5637_n1688);
   U9179 : INV_X1 port map( A => DP_OP_751_130_5637_n1773, ZN => n8054);
   U9180 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1473, B => 
                           DP_OP_751_130_5637_n1431, ZN => n8178);
   U9181 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1472, B => n8178, ZN => 
                           DP_OP_751_130_5637_n1374);
   U9182 : XNOR2_X1 port map( A => n8055, B => n7979, ZN => 
                           DP_OP_751_130_5637_n1770);
   U9183 : OAI22_X1 port map( A1 => n7754, A2 => n10010, B1 => n7796, B2 => 
                           n9979, ZN => n8055);
   U9184 : AND2_X1 port map( A1 => n8705, A2 => n8703, ZN => n8111);
   U9185 : INV_X1 port map( A => DP_OP_751_130_5637_n1771, ZN => n8079);
   U9186 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1794, A2 => 
                           DP_OP_751_130_5637_n1761, ZN => n8095);
   U9187 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1533, B2 => 
                           DP_OP_751_130_5637_n1575, A => 
                           DP_OP_751_130_5637_n1574, ZN => n8060);
   U9188 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1739, B => n8057, ZN => 
                           DP_OP_751_130_5637_n1682);
   U9189 : INV_X1 port map( A => DP_OP_751_130_5637_n1770, ZN => n8057);
   U9190 : XNOR2_X1 port map( A => n8061, B => DP_OP_751_130_5637_n1574, ZN => 
                           DP_OP_751_130_5637_n1476);
   U9191 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1575, B => 
                           DP_OP_751_130_5637_n1533, ZN => n8061);
   U9192 : XNOR2_X1 port map( A => n8067, B => n8066, ZN => 
                           DP_OP_751_130_5637_n1376);
   U9193 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1475, B => 
                           DP_OP_751_130_5637_n1432, ZN => n8067);
   U9194 : NAND2_X1 port map( A1 => DataPath_ALUhw_MULT_mux_out_0_29_port, A2 
                           => n7979, ZN => n8085);
   U9195 : NAND3_X1 port map( A1 => n9016, A2 => n9015, A3 => n8069, ZN => 
                           n10453);
   U9196 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_20_port, B => 
                           n7828, ZN => DP_OP_751_130_5637_n1743);
   U9197 : XNOR2_X1 port map( A => n8073, B => n8072, ZN => 
                           DP_OP_751_130_5637_n1284);
   U9198 : XNOR2_X1 port map( A => n8074, B => n7828, ZN => 
                           DP_OP_751_130_5637_n1734);
   U9199 : OAI22_X1 port map( A1 => n8563, A2 => n10181, B1 => n8485, B2 => 
                           n9874, ZN => n8074);
   U9200 : BUF_X2 port map( A => n10466, Z => n8495);
   U9201 : XNOR2_X1 port map( A => n8075, B => n7828, ZN => 
                           DP_OP_751_130_5637_n1733);
   U9202 : OAI22_X1 port map( A1 => n8563, A2 => n9874, B1 => n8485, B2 => 
                           n10114, ZN => n8075);
   U9203 : BUF_X1 port map( A => DP_OP_751_130_5637_n1794, Z => n8076);
   U9204 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1581, B => 
                           DP_OP_751_130_5637_n1536, ZN => n8078);
   U9205 : NAND2_X1 port map( A1 => n8703, A2 => n8500, ZN => n9301);
   U9206 : NAND2_X1 port map( A1 => n9275, A2 => n10707, ZN => n8703);
   U9207 : OR2_X1 port map( A1 => DataPath_ALUhw_MULT_mux_out_0_29_port, A2 => 
                           n7979, ZN => n8086);
   U9208 : OAI22_X1 port map( A1 => n7754, A2 => n10114, B1 => n7796, B2 => 
                           n9817, ZN => DataPath_ALUhw_MULT_mux_out_0_29_port);
   U9209 : INV_X1 port map( A => n9563, ZN => n8081);
   U9210 : BUF_X1 port map( A => n10695, Z => n8082);
   U9211 : NAND2_X1 port map( A1 => n10516, A2 => n8687, ZN => n9028);
   U9212 : OAI211_X1 port map( C1 => n9108, C2 => n8428, A => n9026, B => n9025
                           , ZN => n10516);
   U9213 : NOR2_X1 port map( A1 => n8083, A2 => n8174, ZN => 
                           DP_OP_751_130_5637_n1673);
   U9214 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_28_port, B => 
                           n8263, ZN => n8174);
   U9215 : INV_X1 port map( A => n8175, ZN => n8083);
   U9216 : NAND2_X1 port map( A1 => n8086, A2 => n8085, ZN => 
                           DP_OP_751_130_5637_n1765);
   U9217 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_22_port, ZN => n8087);
   U9218 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n11, A2 => n8089, ZN 
                           => n8088);
   U9219 : OR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_22_port, ZN => n8089);
   U9220 : BUF_X2 port map( A => DP_OP_751_130_5637_n1659, Z => n8262);
   U9221 : NAND2_X1 port map( A1 => n8111, A2 => n8504, ZN => n9008);
   U9222 : NAND2_X1 port map( A1 => n10824, A2 => n10770, ZN => n8504);
   U9223 : NAND3_X1 port map( A1 => n9038, A2 => n9037, A3 => n8091, ZN => 
                           n10527);
   U9224 : OR2_X1 port map( A1 => n9036, A2 => i_RD1_1_port, ZN => n8140);
   U9225 : OAI21_X1 port map( B1 => n10517, B2 => n8685, A => n9024, ZN => 
                           n9036);
   U9226 : NAND2_X1 port map( A1 => n9035, A2 => n8092, ZN => n9042);
   U9227 : AND2_X1 port map( A1 => n9034, A2 => n8140, ZN => n8092);
   U9228 : NAND3_X1 port map( A1 => n9001, A2 => n8108, A3 => n9000, ZN => 
                           n10464);
   U9229 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1737, B => n8097, ZN => 
                           DP_OP_751_130_5637_n1678);
   U9230 : INV_X1 port map( A => DP_OP_751_130_5637_n1768, ZN => n8097);
   U9231 : INV_X1 port map( A => n8098, ZN => n8444);
   U9232 : OAI21_X1 port map( B1 => n8462, B2 => n8459, A => n8445, ZN => n8098
                           );
   U9233 : NAND2_X1 port map( A1 => n8131, A2 => DP_OP_751_130_5637_n1680, ZN 
                           => n8130);
   U9234 : NAND2_X1 port map( A1 => n9451, A2 => n7752, ZN => n8560);
   U9235 : NAND3_X1 port map( A1 => n9022, A2 => n9021, A3 => n8107, ZN => 
                           n10517);
   U9236 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1488, A2 => n8152, ZN 
                           => n8151);
   U9237 : XNOR2_X1 port map( A => n8109, B => DP_OP_751_130_5637_n1733, ZN => 
                           DP_OP_751_130_5637_n1670);
   U9238 : INV_X1 port map( A => DP_OP_751_130_5637_n1764, ZN => n8109);
   U9239 : AOI21_X1 port map( B1 => n10453, B2 => n8686, A => n9017, ZN => 
                           n9018);
   U9240 : OR2_X1 port map( A1 => n9018, A2 => i_RD1_7_port, ZN => n9054);
   U9241 : NAND2_X1 port map( A1 => n8112, A2 => n9306, ZN => n10658);
   U9242 : OAI21_X1 port map( B1 => n9305, B2 => n9304, A => n8113, ZN => n8112
                           );
   U9243 : NOR2_X1 port map( A1 => n7776, A2 => n9307, ZN => n8113);
   U9244 : XNOR2_X1 port map( A => n8120, B => n8118, ZN => 
                           DP_OP_751_130_5637_n1480);
   U9245 : XNOR2_X1 port map( A => n8119, B => DP_OP_751_130_5637_n1676, ZN => 
                           n8118);
   U9246 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1677, B => 
                           DP_OP_751_130_5637_n1635, ZN => n8119);
   U9247 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1579, B => 
                           DP_OP_751_130_5637_n1535, ZN => n8120);
   U9248 : NAND2_X1 port map( A1 => n8456, A2 => n8457, ZN => n10592);
   U9249 : NAND2_X1 port map( A1 => n8124, A2 => n8123, ZN => 
                           DP_OP_1090J1_126_7243_n28);
   U9250 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_4_port, ZN => n8123);
   U9251 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n29, A2 => n8125, ZN 
                           => n8124);
   U9252 : OR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_4_port, ZN => n8125);
   U9253 : NAND2_X1 port map( A1 => n9040, A2 => n9029, ZN => n9035);
   U9254 : NAND2_X1 port map( A1 => n9028, A2 => n9027, ZN => n9040);
   U9255 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n497, B => 
                           DP_OP_751_130_5637_n433, ZN => n8182);
   U9256 : XNOR2_X1 port map( A => n8182, B => n8181, ZN => 
                           DP_OP_751_130_5637_n398);
   U9257 : XNOR2_X1 port map( A => n8133, B => n8132, ZN => 
                           DP_OP_751_130_5637_n1484);
   U9258 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1583, B => 
                           DP_OP_751_130_5637_n1537, ZN => n8133);
   U9259 : NAND2_X1 port map( A1 => n8134, A2 => n8191, ZN => n9232);
   U9260 : OAI21_X1 port map( B1 => n8020, B2 => n8162, A => n8161, ZN => 
                           DP_OP_1090J1_126_7243_n19);
   U9261 : XNOR2_X1 port map( A => n8141, B => n7979, ZN => 
                           DP_OP_751_130_5637_n1764);
   U9262 : OAI21_X1 port map( B1 => n7755, B2 => n9817, A => n7750, ZN => n8141
                           );
   U9263 : NAND2_X1 port map( A1 => n8201, A2 => DP_OP_1090J1_126_7243_n30, ZN 
                           => n8200);
   U9264 : NAND2_X1 port map( A1 => n8143, A2 => n8142, ZN => 
                           DP_OP_1090J1_126_7243_n30);
   U9265 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_2_port, ZN => n8142);
   U9266 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n37, A2 => n8144, ZN 
                           => n8143);
   U9267 : OR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_2_port, ZN => n8144);
   U9268 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1489, B => 
                           DP_OP_751_130_5637_n1439, ZN => n8154);
   U9269 : NAND2_X1 port map( A1 => n8158, A2 => n9291, ZN => n9296);
   U9270 : OAI21_X1 port map( B1 => n10671, B2 => n10669, A => n8159, ZN => 
                           n8158);
   U9271 : NOR2_X1 port map( A1 => n9292, A2 => n7777, ZN => n8159);
   U9272 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_13_port, ZN => n8161);
   U9273 : NOR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_13_port, ZN => n8162);
   U9274 : NAND3_X1 port map( A1 => n9053, A2 => n9052, A3 => n8163, ZN => 
                           n9256);
   U9275 : INV_X1 port map( A => n10825, ZN => n10757);
   U9276 : OAI21_X1 port map( B1 => n7745, B2 => n8171, A => n8170, ZN => 
                           DP_OP_1090J1_126_7243_n17);
   U9277 : BUF_X1 port map( A => n9587, Z => n8167);
   U9278 : OAI21_X1 port map( B1 => n8169, B2 => n8176, A => n8172, ZN => 
                           DP_OP_1090J1_126_7243_n16);
   U9279 : INV_X1 port map( A => DP_OP_1090J1_126_7243_n17, ZN => n8169);
   U9280 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_15_port, ZN => n8170);
   U9281 : NOR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_15_port, ZN => n8171);
   U9282 : NOR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n16, A2 => n8232, ZN 
                           => n8230);
   U9283 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_16_port, ZN => n8172);
   U9284 : XNOR2_X1 port map( A => n8174, B => n8175, ZN => 
                           DP_OP_751_130_5637_n1674);
   U9285 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n497, A2 => 
                           DP_OP_751_130_5637_n433, ZN => n8180);
   U9286 : NAND2_X1 port map( A1 => n10796, A2 => n10823, ZN => n9315);
   U9287 : NAND2_X1 port map( A1 => n9270, A2 => n9269, ZN => n10796);
   U9288 : INV_X1 port map( A => DP_OP_1090J1_126_7243_n72, ZN => n8186);
   U9289 : NOR2_X1 port map( A1 => n8985, A2 => n9008, ZN => n9092);
   U9290 : AND2_X1 port map( A1 => C620_DATA2_29, A2 => n8379, ZN => n8482);
   U9291 : XNOR2_X1 port map( A => n8193, B => n8287, ZN => C620_DATA2_29);
   U9292 : NAND2_X1 port map( A1 => n8194, A2 => n8211, ZN => n8193);
   U9293 : NAND3_X1 port map( A1 => n8293, A2 => n8292, A3 => n8199, ZN => 
                           n8194);
   U9294 : NAND2_X1 port map( A1 => n8195, A2 => n8234, ZN => n8196);
   U9295 : NAND3_X1 port map( A1 => n8293, A2 => n8292, A3 => n8197, ZN => 
                           n8195);
   U9296 : AND2_X1 port map( A1 => C620_DATA2_31, A2 => n8379, ZN => n8480);
   U9297 : XNOR2_X1 port map( A => n8196, B => DP_OP_1090J1_126_7243_n1, ZN => 
                           C620_DATA2_31);
   U9298 : NOR2_X1 port map( A1 => n8198, A2 => n7766, ZN => n8197);
   U9299 : INV_X1 port map( A => n8244, ZN => n8198);
   U9300 : NOR2_X1 port map( A1 => n7791, A2 => n7766, ZN => n8199);
   U9301 : NAND2_X1 port map( A1 => n7935, A2 => DP_OP_1090J1_126_7243_n72, ZN 
                           => n8293);
   U9302 : NAND2_X1 port map( A1 => n7935, A2 => 
                           DataPath_WRF_CUhw_curr_addr_27_port, ZN => n8292);
   U9303 : NAND2_X1 port map( A1 => n8200, A2 => n8296, ZN => 
                           DP_OP_1090J1_126_7243_n29);
   U9304 : OR2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_27_port, ZN => n8204);
   U9305 : AOI21_X1 port map( B1 => n7935, B2 => n8209, A => n8206, ZN => n8205
                           );
   U9306 : AOI21_X1 port map( B1 => n7935, B2 => n8204, A => n7766, ZN => n8208
                           );
   U9307 : NAND2_X1 port map( A1 => n8212, A2 => n8213, ZN => n10628);
   U9308 : NAND2_X1 port map( A1 => n10645, A2 => n8215, ZN => n8212);
   U9309 : OAI21_X1 port map( B1 => n10649, B2 => n8222, A => n8219, ZN => 
                           n8456);
   U9310 : OR2_X1 port map( A1 => n10649, A2 => n10648, ZN => n10650);
   U9311 : NOR2_X1 port map( A1 => n8447, A2 => n7760, ZN => n8227);
   U9312 : OAI21_X1 port map( B1 => n10645, B2 => n10643, A => n10642, ZN => 
                           n8248);
   U9313 : OAI21_X1 port map( B1 => n8031, B2 => n10669, A => n10668, ZN => 
                           n8249);
   U9314 : AOI21_X1 port map( B1 => n9193, B2 => n9192, A => n9191, ZN => n8250
                           );
   U9315 : BUF_X1 port map( A => n10676, Z => n8251);
   U9316 : OAI21_X1 port map( B1 => n8034, B2 => n9304, A => n9303, ZN => n8252
                           );
   U9317 : AOI21_X1 port map( B1 => n8096, B2 => n10573, A => n10572, ZN => 
                           n8253);
   U9318 : AND2_X1 port map( A1 => C620_DATA2_29, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_29_port);
   U9319 : AND2_X1 port map( A1 => C620_DATA2_30, A2 => n8379, ZN => n8481);
   U9320 : AND2_X1 port map( A1 => C620_DATA2_30, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_30_port);
   U9321 : AOI222_X1 port map( A1 => DataPath_RF_c_win_1_port, A2 => n12041, B1
                           => DataPath_RF_c_win_2_port, B2 => n12042, C1 => 
                           DataPath_RF_c_win_0_port, C2 => n12043, ZN => n12038
                           );
   U9322 : AOI211_X1 port map( C1 => n9272, C2 => n9271, A => CU_I_i_FILL_delay
                           , B => n7768, ZN => n9273);
   U9323 : NOR2_X1 port map( A1 => n10876, A2 => n8723, ZN => n8976);
   U9324 : INV_X1 port map( A => n8102, ZN => n8254);
   U9325 : NOR2_X1 port map( A1 => n9272, A2 => n8720, ZN => n8256);
   U9326 : NOR2_X1 port map( A1 => n9272, A2 => n8720, ZN => n8977);
   U9327 : INV_X1 port map( A => DP_OP_751_130_5637_n119, ZN => 
                           DP_OP_751_130_5637_n117);
   U9328 : INV_X1 port map( A => DP_OP_751_130_5637_n127, ZN => 
                           DP_OP_751_130_5637_n125);
   U9329 : INV_X1 port map( A => DP_OP_751_130_5637_n139, ZN => 
                           DP_OP_751_130_5637_n137);
   U9330 : INV_X1 port map( A => DP_OP_751_130_5637_n147, ZN => 
                           DP_OP_751_130_5637_n145);
   U9331 : INV_X1 port map( A => DP_OP_751_130_5637_n155, ZN => 
                           DP_OP_751_130_5637_n153);
   U9332 : INV_X1 port map( A => DP_OP_751_130_5637_n169, ZN => 
                           DP_OP_751_130_5637_n167);
   U9333 : INV_X1 port map( A => DP_OP_751_130_5637_n177, ZN => 
                           DP_OP_751_130_5637_n175);
   U9334 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_31_port, ZN => 
                           DP_OP_751_130_5637_n1798);
   U9335 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_20_port, ZN => 
                           DP_OP_751_130_5637_n1809);
   U9336 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_19_port, ZN => 
                           DP_OP_751_130_5637_n1810);
   U9337 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_18_port, ZN => 
                           DP_OP_751_130_5637_n1811);
   U9338 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_17_port, ZN => 
                           DP_OP_751_130_5637_n1812);
   U9339 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_16_port, ZN => 
                           DP_OP_751_130_5637_n1813);
   U9340 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_15_port, ZN => 
                           DP_OP_751_130_5637_n1814);
   U9341 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_14_port, ZN => 
                           DP_OP_751_130_5637_n1815);
   U9342 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_13_port, ZN => 
                           DP_OP_751_130_5637_n1816);
   U9343 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_1_port, ZN => 
                           DP_OP_751_130_5637_n1828);
   U9344 : INV_X1 port map( A => DP_OP_751_130_5637_n191, ZN => 
                           DP_OP_751_130_5637_n189);
   U9345 : INV_X1 port map( A => DP_OP_751_130_5637_n198, ZN => 
                           DP_OP_751_130_5637_n196);
   U9346 : INV_X1 port map( A => DP_OP_751_130_5637_n71, ZN => 
                           DP_OP_751_130_5637_n201);
   U9347 : INV_X1 port map( A => DP_OP_751_130_5637_n91, ZN => 
                           DP_OP_751_130_5637_n206);
   U9348 : INV_X1 port map( A => DP_OP_751_130_5637_n105, ZN => 
                           DP_OP_751_130_5637_n209);
   U9349 : INV_X1 port map( A => DP_OP_751_130_5637_n113, ZN => 
                           DP_OP_751_130_5637_n211);
   U9350 : INV_X1 port map( A => DP_OP_751_130_5637_n121, ZN => 
                           DP_OP_751_130_5637_n213);
   U9351 : INV_X1 port map( A => DP_OP_751_130_5637_n129, ZN => 
                           DP_OP_751_130_5637_n215);
   U9352 : INV_X1 port map( A => DP_OP_751_130_5637_n133, ZN => 
                           DP_OP_751_130_5637_n216);
   U9353 : INV_X1 port map( A => DP_OP_751_130_5637_n141, ZN => 
                           DP_OP_751_130_5637_n218);
   U9354 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n171, B2 => 
                           DP_OP_751_130_5637_n173, A => 
                           DP_OP_751_130_5637_n172, ZN => 
                           DP_OP_751_130_5637_n170);
   U9355 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n163, B2 => 
                           DP_OP_751_130_5637_n165, A => 
                           DP_OP_751_130_5637_n164, ZN => 
                           DP_OP_751_130_5637_n162);
   U9356 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n141, B2 => 
                           DP_OP_751_130_5637_n143, A => 
                           DP_OP_751_130_5637_n142, ZN => 
                           DP_OP_751_130_5637_n140);
   U9357 : XOR2_X1 port map( A => DP_OP_751_130_5637_n8, B => n7748, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_57_port);
   U9358 : XOR2_X1 port map( A => DP_OP_751_130_5637_n20, B => 
                           DP_OP_751_130_5637_n143, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_45_port);
   U9359 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n7, B => n8056, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_58_port);
   U9360 : BUF_X1 port map( A => n7749, Z => n8265);
   U9361 : BUF_X1 port map( A => DP_OP_751_130_5637_n1455, Z => n8259);
   U9362 : BUF_X1 port map( A => DP_OP_751_130_5637_n1557, Z => n8260);
   U9363 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n502, A2 => 
                           DP_OP_751_130_5637_n600, ZN => n8271);
   U9364 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n908, A2 => 
                           DP_OP_751_130_5637_n909, ZN => n8275);
   U9365 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1010, A2 => 
                           DP_OP_751_130_5637_n1011, ZN => n8276);
   U9366 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1114, A2 => 
                           DP_OP_751_130_5637_n1212, ZN => n8277);
   U9367 : BUF_X1 port map( A => n7749, Z => n8264);
   U9368 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1216, A2 => 
                           DP_OP_751_130_5637_n1314, ZN => n8278);
   U9369 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1318, A2 => 
                           DP_OP_751_130_5637_n1416, ZN => n8279);
   U9370 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1418, A2 => 
                           DP_OP_751_130_5637_n1419, ZN => n8270);
   U9371 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1520, A2 => 
                           DP_OP_751_130_5637_n1521, ZN => n8280);
   U9372 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1622, A2 => 
                           DP_OP_751_130_5637_n1623, ZN => n8282);
   U9373 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1726, A2 => 
                           DP_OP_751_130_5637_n1792, ZN => n8281);
   U9374 : AND2_X1 port map( A1 => DP_OP_751_130_5637_n194, A2 => 
                           DP_OP_751_130_5637_n196, ZN => n8283);
   U9375 : BUF_X1 port map( A => DP_OP_751_130_5637_n843, Z => n8268);
   U9376 : BUF_X1 port map( A => DP_OP_751_130_5637_n1047, Z => n8266);
   U9377 : BUF_X1 port map( A => DP_OP_751_130_5637_n945, Z => n8267);
   U9378 : BUF_X1 port map( A => DP_OP_751_130_5637_n1353, Z => n8258);
   U9379 : BUF_X1 port map( A => DP_OP_751_130_5637_n1557, Z => n8261);
   U9380 : INV_X1 port map( A => DP_OP_1090J1_126_7243_n72, ZN => n8285);
   U9381 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_30_port, ZN => n8284);
   U9382 : XNOR2_X1 port map( A => DP_OP_1090J1_126_7243_n75, B => n8285, ZN =>
                           DP_OP_1090J1_126_7243_n37);
   U9383 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_29_port, ZN => n8286);
   U9384 : XOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_29_port, Z => n8287);
   U9385 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_28_port, ZN => n8288);
   U9386 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_27_port, ZN => n8291);
   U9387 : XOR2_X1 port map( A => n7935, B => n8294, Z => C620_DATA2_27);
   U9388 : XOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_27_port, Z => n8294);
   U9389 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_3_port, ZN => n8296);
   U9390 : XOR2_X1 port map( A => DP_OP_1090J1_126_7243_n30, B => n8297, Z => 
                           C620_DATA2_3);
   U9391 : XOR2_X1 port map( A => DP_OP_1090J1_126_7243_n72, B => 
                           DataPath_WRF_CUhw_curr_addr_3_port, Z => n8297);
   U9392 : NAND2_X1 port map( A1 => DP_OP_1090J1_126_7243_n72, A2 => 
                           DataPath_WRF_CUhw_curr_addr_24_port, ZN => n8298);
   U9393 : OR2_X1 port map( A1 => n7768, A2 => n10709, ZN => n8720);
   U9394 : OAI22_X2 port map( A1 => n9636, A2 => n8802, B1 => n577, B2 => 
                           n12094, ZN => n11418);
   U9395 : OAI22_X2 port map( A1 => n9641, A2 => n8802, B1 => n577, B2 => 
                           n12121, ZN => n11449);
   U9396 : INV_X2 port map( A => n12193, ZN => n8669);
   U9397 : INV_X2 port map( A => n12018, ZN => n8653);
   U9398 : INV_X2 port map( A => n11854, ZN => n8644);
   U9399 : OAI22_X2 port map( A1 => n9641, A2 => n8851, B1 => n11596, B2 => 
                           n12121, ZN => n11539);
   U9400 : OAI22_X2 port map( A1 => n9636, A2 => n8851, B1 => n11596, B2 => 
                           n12094, ZN => n11512);
   U9401 : OAI22_X2 port map( A1 => n9637, A2 => n8851, B1 => n11596, B2 => 
                           n12109, ZN => n11514);
   U9402 : NOR2_X1 port map( A1 => i_BUSY_WINDOW, A2 => CU_I_i_SPILL_delay, ZN 
                           => n8979);
   U9403 : BUF_X1 port map( A => n11660, Z => n8631);
   U9404 : BUF_X1 port map( A => n11653, Z => n8629);
   U9405 : BUF_X1 port map( A => n12154, Z => n8663);
   U9406 : BUF_X1 port map( A => n11696, Z => n8634);
   U9407 : AND2_X1 port map( A1 => n8696, A2 => n12107, ZN => n12106);
   U9408 : BUF_X1 port map( A => n11536, Z => n8621);
   U9409 : BUF_X1 port map( A => n11531, Z => n8619);
   U9410 : BUF_X1 port map( A => n11543, Z => n8623);
   U9411 : AND2_X1 port map( A1 => n8698, A2 => n11534, ZN => n11532);
   U9412 : BUF_X1 port map( A => n11585, Z => n8625);
   U9413 : AND2_X1 port map( A1 => n8690, A2 => n11418, ZN => n11420);
   U9414 : AND2_X1 port map( A1 => n8695, A2 => n11449, ZN => n11451);
   U9415 : INV_X1 port map( A => n8669, ZN => n8668);
   U9416 : INV_X1 port map( A => n8653, ZN => n8652);
   U9417 : AOI22_X1 port map( A1 => n8791, A2 => n3342, B1 => n11931, B2 => 
                           n8802, ZN => n11493);
   U9418 : INV_X1 port map( A => n8644, ZN => n8643);
   U9419 : NAND2_X1 port map( A1 => n8802, A2 => n8688, ZN => n8791);
   U9420 : INV_X2 port map( A => n8803, ZN => n8802);
   U9421 : INV_X1 port map( A => n8795, ZN => n9639);
   U9422 : OAI22_X1 port map( A1 => n9640, A2 => n8965, B1 => n12118, B2 => 
                           n8299, ZN => n11814);
   U9423 : OAI22_X1 port map( A1 => n9644, A2 => n8965, B1 => n12158, B2 => 
                           n8299, ZN => n11821);
   U9424 : INV_X1 port map( A => n8794, ZN => n9638);
   U9425 : NOR2_X1 port map( A1 => RST, A2 => n7804, ZN => n11819);
   U9426 : INV_X1 port map( A => n8680, ZN => n8679);
   U9427 : NAND2_X1 port map( A1 => n8256, A2 => n8976, ZN => n8724);
   U9428 : NOR2_X1 port map( A1 => n8702, A2 => n187, ZN => n10861);
   U9429 : INV_X1 port map( A => n8675, ZN => n8673);
   U9430 : INV_X1 port map( A => n8675, ZN => n8671);
   U9431 : AND2_X1 port map( A1 => n10877, A2 => n8688, ZN => n10857);
   U9432 : AND2_X1 port map( A1 => i_BUSY_WINDOW, A2 => n171, ZN => n9272);
   U9433 : NOR2_X1 port map( A1 => RST, A2 => n11816, ZN => n11818);
   U9434 : NOR2_X1 port map( A1 => RST, A2 => n7801, ZN => n11425);
   U9435 : OAI22_X1 port map( A1 => n9638, A2 => n8802, B1 => n577, B2 => 
                           n12112, ZN => n11426);
   U9436 : NOR2_X1 port map( A1 => RST, A2 => n8514, ZN => n11457);
   U9437 : NOR2_X1 port map( A1 => RST, A2 => n8513, ZN => n11454);
   U9438 : NOR2_X1 port map( A1 => RST, A2 => n8512, ZN => n11431);
   U9439 : NOR2_X1 port map( A1 => RST, A2 => n8511, ZN => n11423);
   U9440 : NOR2_X1 port map( A1 => RST, A2 => n8534, ZN => n11637);
   U9441 : NOR2_X1 port map( A1 => RST, A2 => n8536, ZN => n11661);
   U9442 : NOR2_X1 port map( A1 => RST, A2 => n8535, ZN => n11655);
   U9443 : NOR2_X1 port map( A1 => RST, A2 => n8533, ZN => n11635);
   U9444 : NOR2_X1 port map( A1 => RST, A2 => n8537, ZN => n11663);
   U9445 : NOR2_X1 port map( A1 => RST, A2 => n8666, ZN => n12176);
   U9446 : NOR2_X1 port map( A1 => RST, A2 => n8659, ZN => n12117);
   U9447 : NOR2_X1 port map( A1 => RST, A2 => n8655, ZN => n12111);
   U9448 : NOR2_X1 port map( A1 => RST, A2 => n8661, ZN => n12120);
   U9449 : NOR2_X1 port map( A1 => RST, A2 => n8523, ZN => n11538);
   U9450 : NOR2_X1 port map( A1 => RST, A2 => n8524, ZN => n11544);
   U9451 : NOR2_X1 port map( A1 => RST, A2 => n8521, ZN => n11513);
   U9452 : NOR2_X1 port map( A1 => RST, A2 => n8522, ZN => n11515);
   U9453 : INV_X1 port map( A => RST, ZN => n8698);
   U9454 : AND2_X1 port map( A1 => n8697, A2 => n11787, ZN => n11863);
   U9455 : AOI22_X1 port map( A1 => n8932, A2 => n3342, B1 => n11931, B2 => 
                           n8965, ZN => n11873);
   U9456 : NOR2_X1 port map( A1 => RST, A2 => n7805, ZN => n11815);
   U9457 : NOR2_X1 port map( A1 => RST, A2 => n7806, ZN => n11822);
   U9458 : AND2_X1 port map( A1 => n8697, A2 => n11795, ZN => n11872);
   U9459 : NOR2_X1 port map( A1 => RST, A2 => n7803, ZN => n11782);
   U9460 : OAI22_X1 port map( A1 => n9638, A2 => n8965, B1 => n8299, B2 => 
                           n12112, ZN => n11781);
   U9461 : NOR2_X1 port map( A1 => RST, A2 => n7802, ZN => n11766);
   U9462 : OAI22_X1 port map( A1 => n9636, A2 => n8965, B1 => n8299, B2 => 
                           n12094, ZN => n11765);
   U9463 : AND2_X1 port map( A1 => n8697, A2 => n11794, ZN => n11871);
   U9464 : AND2_X1 port map( A1 => n8697, A2 => n11790, ZN => n11867);
   U9465 : AND2_X1 port map( A1 => n8697, A2 => n11784, ZN => n11859);
   U9466 : AND2_X1 port map( A1 => n8697, A2 => n11789, ZN => n11866);
   U9467 : AND2_X1 port map( A1 => n8697, A2 => n11786, ZN => n11862);
   U9468 : AND2_X1 port map( A1 => n8697, A2 => n11783, ZN => n11858);
   U9469 : INV_X1 port map( A => RST, ZN => n8697);
   U9470 : OAI22_X1 port map( A1 => n9642, A2 => n8965, B1 => n12155, B2 => 
                           n8299, ZN => n11820);
   U9471 : NOR3_X1 port map( A1 => n11375, A2 => n10868, A3 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_15_port, ZN => 
                           n11377);
   U9472 : OAI211_X1 port map( C1 => n193, C2 => n8190, A => n8711, B => n8706,
                           ZN => i_ADD_WS1_0_port);
   U9473 : OAI211_X1 port map( C1 => n191, C2 => n8190, A => n8711, B => n8708,
                           ZN => i_ADD_WS1_2_port);
   U9474 : NOR2_X1 port map( A1 => n8702, A2 => n186, ZN => n10860);
   U9475 : INV_X1 port map( A => n8314, ZN => n8672);
   U9476 : INV_X1 port map( A => RST, ZN => n8696);
   U9477 : BUF_X1 port map( A => n12203, Z => n8670);
   U9478 : NOR2_X1 port map( A1 => RST, A2 => n12203, ZN => n12204);
   U9479 : NOR2_X1 port map( A1 => RST, A2 => n11796, ZN => n11813);
   U9480 : NOR2_X1 port map( A1 => RST, A2 => n11418, ZN => n11419);
   U9481 : NOR2_X1 port map( A1 => RST, A2 => n11774, ZN => n11780);
   U9482 : NOR2_X1 port map( A1 => RST, A2 => n11449, ZN => n11452);
   U9483 : AND2_X1 port map( A1 => n8698, A2 => n11667, ZN => n11719);
   U9484 : NOR2_X1 port map( A1 => RST, A2 => n11590, ZN => n11591);
   U9485 : AND2_X1 port map( A1 => n8688, A2 => n11436, ZN => n11482);
   U9486 : AND2_X1 port map( A1 => n8690, A2 => n11444, ZN => n11492);
   U9487 : AND2_X1 port map( A1 => n8689, A2 => n11450, ZN => n11510);
   U9488 : AND2_X1 port map( A1 => n8694, A2 => n11446, ZN => n11501);
   U9489 : AND2_X1 port map( A1 => n8691, A2 => n11437, ZN => n11483);
   U9490 : AND2_X1 port map( A1 => n8688, A2 => n11439, ZN => n11485);
   U9491 : AND2_X1 port map( A1 => n8690, A2 => n11433, ZN => n11479);
   U9492 : AND2_X1 port map( A1 => n8689, A2 => n11441, ZN => n11487);
   U9493 : AND2_X1 port map( A1 => n8689, A2 => n11421, ZN => n11506);
   U9494 : AND2_X1 port map( A1 => n8696, A2 => n11434, ZN => n11480);
   U9495 : AND2_X1 port map( A1 => n8691, A2 => n11448, ZN => n11504);
   U9496 : AND2_X1 port map( A1 => n8688, A2 => n11447, ZN => n11502);
   U9497 : AND2_X1 port map( A1 => n8690, A2 => n11435, ZN => n11481);
   U9498 : AND2_X1 port map( A1 => n8689, A2 => n11442, ZN => n11489);
   U9499 : AND2_X1 port map( A1 => n8698, A2 => n11445, ZN => n11496);
   U9500 : AND2_X1 port map( A1 => n8693, A2 => n11440, ZN => n11486);
   U9501 : AND2_X1 port map( A1 => n8691, A2 => n11438, ZN => n11484);
   U9502 : AND2_X1 port map( A1 => n8688, A2 => n11443, ZN => n11491);
   U9503 : AND2_X1 port map( A1 => n8690, A2 => n11432, ZN => n11478);
   U9504 : AND2_X1 port map( A1 => n8698, A2 => n11671, ZN => n11723);
   U9505 : AND2_X1 port map( A1 => n8696, A2 => n12126, ZN => n12181);
   U9506 : AND2_X1 port map( A1 => n8696, A2 => n12147, ZN => n12169);
   U9507 : AND2_X1 port map( A1 => n8696, A2 => n12123, ZN => n12178);
   U9508 : AND2_X1 port map( A1 => n8697, A2 => n11694, ZN => n11748);
   U9509 : AND2_X1 port map( A1 => n8698, A2 => n11687, ZN => n11739);
   U9510 : AND2_X1 port map( A1 => n8698, A2 => n11678, ZN => n11730);
   U9511 : AND2_X1 port map( A1 => n8698, A2 => n11690, ZN => n11742);
   U9512 : AND2_X1 port map( A1 => n8698, A2 => n11669, ZN => n11721);
   U9513 : AND2_X1 port map( A1 => n8698, A2 => n11688, ZN => n11740);
   U9514 : INV_X1 port map( A => n8854, ZN => n11716);
   U9515 : AND2_X1 port map( A1 => n8698, A2 => n11675, ZN => n11727);
   U9516 : AND2_X1 port map( A1 => n8698, A2 => n11668, ZN => n11720);
   U9517 : AND2_X1 port map( A1 => n8698, A2 => n11672, ZN => n11724);
   U9518 : AND2_X1 port map( A1 => n8696, A2 => n12144, ZN => n12167);
   U9519 : AND2_X1 port map( A1 => n8696, A2 => n12124, ZN => n12179);
   U9520 : AND2_X1 port map( A1 => n8696, A2 => n12125, ZN => n12180);
   U9521 : AND2_X1 port map( A1 => n8698, A2 => n11677, ZN => n11729);
   U9522 : AND2_X1 port map( A1 => n8698, A2 => n11666, ZN => n11718);
   U9523 : AND2_X1 port map( A1 => n8698, A2 => n11682, ZN => n11734);
   U9524 : AND2_X1 port map( A1 => n8698, A2 => n11670, ZN => n11722);
   U9525 : AND2_X1 port map( A1 => n8698, A2 => n11657, ZN => n11744);
   U9526 : AND2_X1 port map( A1 => n8698, A2 => n11665, ZN => n11717);
   U9527 : AND2_X1 port map( A1 => n8698, A2 => n11673, ZN => n11725);
   U9528 : AND2_X1 port map( A1 => n8698, A2 => n11575, ZN => n11620);
   U9529 : AND2_X1 port map( A1 => n8697, A2 => n11557, ZN => n11602);
   U9530 : AND2_X1 port map( A1 => n8698, A2 => n11576, ZN => n11621);
   U9531 : AND2_X1 port map( A1 => n8696, A2 => n12149, ZN => n12171);
   U9532 : INV_X1 port map( A => n8768, ZN => n12191);
   U9533 : AND2_X1 port map( A1 => n8696, A2 => n12127, ZN => n12182);
   U9534 : AND2_X1 port map( A1 => n8696, A2 => n12130, ZN => n12185);
   U9535 : INV_X1 port map( A => n8847, ZN => n11629);
   U9536 : AND2_X1 port map( A1 => n8696, A2 => n12138, ZN => n12161);
   U9537 : AND2_X1 port map( A1 => n8696, A2 => n12128, ZN => n12183);
   U9538 : AND2_X1 port map( A1 => n8696, A2 => n12131, ZN => n12186);
   U9539 : AND2_X1 port map( A1 => n8696, A2 => n12122, ZN => n12177);
   U9540 : AND2_X1 port map( A1 => n8696, A2 => n12133, ZN => n12188);
   U9541 : AND2_X1 port map( A1 => n8689, A2 => n12135, ZN => n12190);
   U9542 : AND2_X1 port map( A1 => n8696, A2 => n12129, ZN => n12184);
   U9543 : AND2_X1 port map( A1 => n8696, A2 => n12143, ZN => n12166);
   U9544 : AND2_X1 port map( A1 => n8690, A2 => n11555, ZN => n11600);
   U9545 : AND2_X1 port map( A1 => n8698, A2 => n11580, ZN => n11625);
   U9546 : AND2_X1 port map( A1 => n8696, A2 => n11565, ZN => n11610);
   U9547 : AND2_X1 port map( A1 => n8698, A2 => n11566, ZN => n11611);
   U9548 : AND2_X1 port map( A1 => n8698, A2 => n11570, ZN => n11615);
   U9549 : AND2_X1 port map( A1 => n8695, A2 => n11554, ZN => n11598);
   U9550 : AND2_X1 port map( A1 => n8697, A2 => n11558, ZN => n11603);
   U9551 : AND2_X1 port map( A1 => n8691, A2 => n11540, ZN => n11599);
   U9552 : AND2_X1 port map( A1 => n8697, A2 => n11561, ZN => n11606);
   U9553 : AND2_X1 port map( A1 => n8688, A2 => n11556, ZN => n11601);
   U9554 : AND2_X1 port map( A1 => n8690, A2 => n11553, ZN => n11597);
   U9555 : AND2_X1 port map( A1 => n8697, A2 => n11560, ZN => n11605);
   U9556 : AND2_X1 port map( A1 => n8697, A2 => n11563, ZN => n11608);
   U9557 : AND2_X1 port map( A1 => n8698, A2 => n11578, ZN => n11623);
   U9558 : AND2_X1 port map( A1 => n8696, A2 => n11806, ZN => n11884);
   U9559 : AND2_X1 port map( A1 => n8697, A2 => n11767, ZN => n11861);
   U9560 : AND2_X1 port map( A1 => n8697, A2 => n11804, ZN => n11882);
   U9561 : AND2_X1 port map( A1 => n8697, A2 => n11803, ZN => n11881);
   U9562 : AND2_X1 port map( A1 => n8697, A2 => n11788, ZN => n11864);
   U9563 : AND2_X1 port map( A1 => n8697, A2 => n11785, ZN => n11860);
   U9564 : AND2_X1 port map( A1 => n8697, A2 => n11811, ZN => n12017);
   U9565 : AND2_X1 port map( A1 => n8697, A2 => n11792, ZN => n11869);
   U9566 : AND2_X1 port map( A1 => n8697, A2 => n11808, ZN => n11886);
   U9567 : NOR2_X1 port map( A1 => n8700, A2 => n190, ZN => n10864);
   U9568 : NOR2_X1 port map( A1 => n8700, A2 => n193, ZN => n10867);
   U9569 : OR4_X1 port map( A1 => n9253, A2 => n9252, A3 => n9251, A4 => n9250,
                           ZN => n9257);
   U9570 : INV_X1 port map( A => n12087, ZN => n10115);
   U9571 : OR2_X1 port map( A1 => DataPath_RF_POP_ADDRGEN_curr_state_0_port, A2
                           => n851, ZN => n11375);
   U9572 : OAI21_X1 port map( B1 => i_DATAMEM_RM, B2 => i_DATAMEM_WM, A => 
                           CU_I_CW_MEM_2_port, ZN => n12194);
   U9573 : NOR2_X1 port map( A1 => n9005, A2 => n8978, ZN => n8712);
   U9574 : NOR2_X1 port map( A1 => RST, A2 => n11656, ZN => n11660);
   U9575 : NOR2_X1 port map( A1 => RST, A2 => n11638, ZN => n11653);
   U9576 : NOR2_X1 port map( A1 => RST, A2 => n12153, ZN => n12154);
   U9577 : NOR2_X1 port map( A1 => RST, A2 => n11692, ZN => n11696);
   U9578 : NOR2_X1 port map( A1 => RST, A2 => n12107, ZN => n12108);
   U9579 : NOR2_X1 port map( A1 => RST, A2 => n11537, ZN => n11536);
   U9580 : NOR2_X1 port map( A1 => RST, A2 => n11530, ZN => n11531);
   U9581 : NOR2_X1 port map( A1 => RST, A2 => n11542, ZN => n11543);
   U9582 : NOR2_X1 port map( A1 => RST, A2 => n11534, ZN => n11533);
   U9583 : NOR2_X1 port map( A1 => RST, A2 => n11584, ZN => n11585);
   U9584 : INV_X1 port map( A => n11589, ZN => n11844);
   U9585 : INV_X1 port map( A => n11552, ZN => n11835);
   U9586 : NOR2_X1 port map( A1 => i_ADD_WB_4_port, A2 => n11395, ZN => n11414)
                           ;
   U9587 : AND2_X1 port map( A1 => n8887, A2 => n8886, ZN => n11648);
   U9588 : AND2_X1 port map( A1 => n8881, A2 => n8880, ZN => n11646);
   U9589 : AND2_X1 port map( A1 => n8869, A2 => n8868, ZN => n11640);
   U9590 : AND2_X1 port map( A1 => n8740, A2 => n8739, ZN => n12145);
   U9591 : AND2_X1 port map( A1 => n8883, A2 => n8882, ZN => n11647);
   U9592 : AND2_X1 port map( A1 => n8877, A2 => n8876, ZN => n11644);
   U9593 : AND2_X1 port map( A1 => n8879, A2 => n8878, ZN => n11645);
   U9594 : AND2_X1 port map( A1 => n8873, A2 => n8872, ZN => n11641);
   U9595 : AND2_X1 port map( A1 => n8866, A2 => n8865, ZN => n11639);
   U9596 : AND2_X1 port map( A1 => n8890, A2 => n8889, ZN => n11649);
   U9597 : AND2_X1 port map( A1 => n8895, A2 => n8894, ZN => n11651);
   U9598 : AND2_X1 port map( A1 => n8893, A2 => n8892, ZN => n11650);
   U9599 : OAI22_X1 port map( A1 => n9644, A2 => n9643, B1 => n12158, B2 => 
                           n8441, ZN => n12174);
   U9600 : OAI22_X1 port map( A1 => n9639, A2 => n9643, B1 => n12115, B2 => 
                           n8441, ZN => n12116);
   U9601 : AND2_X1 port map( A1 => n8743, A2 => n8742, ZN => n12103);
   U9602 : OAI22_X1 port map( A1 => n9637, A2 => n9643, B1 => n12109, B2 => 
                           n8441, ZN => n12110);
   U9603 : AND2_X1 port map( A1 => n8736, A2 => n8735, ZN => n12102);
   U9604 : OAI22_X1 port map( A1 => n9640, A2 => n9643, B1 => n12118, B2 => 
                           n8441, ZN => n12119);
   U9605 : AND2_X1 port map( A1 => n8762, A2 => n8761, ZN => n12095);
   U9606 : AND2_X1 port map( A1 => n8748, A2 => n8747, ZN => n12105);
   U9607 : AND2_X1 port map( A1 => n8734, A2 => n8733, ZN => n12140);
   U9608 : AND2_X1 port map( A1 => n8732, A2 => n8731, ZN => n12100);
   U9609 : AND2_X1 port map( A1 => n8746, A2 => n8745, ZN => n12104);
   U9610 : AND2_X1 port map( A1 => n8765, A2 => n8764, ZN => n12096);
   U9611 : OAI22_X1 port map( A1 => n9638, A2 => n9643, B1 => n12112, B2 => 
                           n8441, ZN => n12113);
   U9612 : OAI22_X1 port map( A1 => n9642, A2 => n9643, B1 => n12155, B2 => 
                           n8441, ZN => n12156);
   U9613 : AND2_X1 port map( A1 => n8730, A2 => n8729, ZN => n12099);
   U9614 : AND2_X1 port map( A1 => n8697, A2 => n11559, ZN => n11604);
   U9615 : AND2_X1 port map( A1 => n8833, A2 => n8832, ZN => n11524);
   U9616 : AND2_X1 port map( A1 => n8925, A2 => n8924, ZN => n11769);
   U9617 : AND2_X1 port map( A1 => n8931, A2 => n8930, ZN => n11770);
   U9618 : AND2_X1 port map( A1 => n8940, A2 => n8939, ZN => n11801);
   U9619 : AND2_X1 port map( A1 => n8954, A2 => n8953, ZN => n11777);
   U9620 : AND2_X1 port map( A1 => n8946, A2 => n8945, ZN => n11775);
   U9621 : AND2_X1 port map( A1 => n8921, A2 => n8920, ZN => n11768);
   U9622 : AND2_X1 port map( A1 => n8934, A2 => n8933, ZN => n11772);
   U9623 : AND2_X1 port map( A1 => n8936, A2 => n8935, ZN => n11798);
   U9624 : AND2_X1 port map( A1 => n8956, A2 => n8955, ZN => n11778);
   U9625 : AND2_X1 port map( A1 => n8938, A2 => n8937, ZN => n11773);
   U9626 : AND2_X1 port map( A1 => n8950, A2 => n8949, ZN => n11776);
   U9627 : BUF_X1 port map( A => n8411, Z => n8680);
   U9628 : NAND2_X1 port map( A1 => n8693, A2 => n11950, ZN => n12206);
   U9629 : NOR2_X1 port map( A1 => n552, A2 => n11984, ZN => n11985);
   U9630 : NOR2_X1 port map( A1 => n550, A2 => n11981, ZN => n11982);
   U9631 : OAI211_X1 port map( C1 => n189, C2 => n8190, A => n8711, B => n8710,
                           ZN => i_ADD_WS1_4_port);
   U9632 : NAND3_X1 port map( A1 => n8701, A2 => i_RF2, A3 => n9004, ZN => 
                           n8700);
   U9633 : NOR2_X1 port map( A1 => n8702, A2 => n188, ZN => n10862);
   U9634 : NOR2_X1 port map( A1 => n8702, A2 => n184, ZN => n10858);
   U9635 : INV_X1 port map( A => n8705, ZN => n8997);
   U9636 : AND3_X1 port map( A1 => IR_26_port, A2 => n8312, A3 => n171, ZN => 
                           n10710);
   U9637 : INV_X1 port map( A => n10840, ZN => n10482);
   U9638 : AND2_X1 port map( A1 => n9532, A2 => n9531, ZN => n10458);
   U9639 : BUF_X1 port map( A => n9553, Z => n8488);
   U9640 : BUF_X1 port map( A => n9487, Z => n8576);
   U9641 : BUF_X1 port map( A => n10326, Z => n8493);
   U9642 : AND2_X1 port map( A1 => n10848, A2 => n8380, ZN => n10841);
   U9643 : NAND2_X1 port map( A1 => n8979, A2 => n8712, ZN => n8443);
   U9644 : BUF_X1 port map( A => n11892, Z => n8645);
   U9645 : BUF_X1 port map( A => n11948, Z => n8651);
   U9646 : BUF_X1 port map( A => n11912, Z => n8650);
   U9647 : BUF_X1 port map( A => n11904, Z => n8648);
   U9648 : BUF_X1 port map( A => n11908, Z => n8649);
   U9649 : BUF_X1 port map( A => n11896, Z => n8646);
   U9650 : BUF_X1 port map( A => n11900, Z => n8647);
   U9651 : INV_X1 port map( A => n11362, ZN => n11354);
   U9652 : INV_X1 port map( A => n11331, ZN => n11347);
   U9653 : INV_X1 port map( A => n11270, ZN => n11373);
   U9654 : OAI22_X1 port map( A1 => n9636, A2 => n9643, B1 => n12094, B2 => 
                           n8441, ZN => n12107);
   U9655 : OAI22_X1 port map( A1 => n9639, A2 => n8851, B1 => n11596, B2 => 
                           n12115, ZN => n11534);
   U9656 : OAI22_X1 port map( A1 => n9639, A2 => n8965, B1 => n8299, B2 => 
                           n12115, ZN => n11796);
   U9657 : OAI22_X1 port map( A1 => n9637, A2 => n8965, B1 => n8299, B2 => 
                           n12109, ZN => n11774);
   U9658 : NOR2_X1 port map( A1 => n8310, A2 => n11395, ZN => n11413);
   U9659 : NAND2_X1 port map( A1 => i_ADD_WB_3_port, A2 => i_WF, ZN => n11395);
   U9660 : NOR2_X1 port map( A1 => RST, A2 => n11527, ZN => n11626);
   U9661 : AND2_X1 port map( A1 => n8843, A2 => n8842, ZN => n11527);
   U9662 : NOR2_X1 port map( A1 => RST, A2 => n11522, ZN => n11617);
   U9663 : AND2_X1 port map( A1 => n8829, A2 => n8828, ZN => n11522);
   U9664 : NOR2_X1 port map( A1 => RST, A2 => n11521, ZN => n11616);
   U9665 : AND2_X1 port map( A1 => n8827, A2 => n8826, ZN => n11521);
   U9666 : NOR2_X1 port map( A1 => RST, A2 => n11519, ZN => n11613);
   U9667 : NOR2_X1 port map( A1 => RST, A2 => n11518, ZN => n11612);
   U9668 : AND2_X1 port map( A1 => n8822, A2 => n8821, ZN => n11518);
   U9669 : NOR2_X1 port map( A1 => RST, A2 => n11517, ZN => n11609);
   U9670 : AND2_X1 port map( A1 => n8818, A2 => n8817, ZN => n11517);
   U9671 : NOR2_X1 port map( A1 => RST, A2 => n11524, ZN => n11619);
   U9672 : NOR2_X1 port map( A1 => RST, A2 => n11523, ZN => n11618);
   U9673 : AND2_X1 port map( A1 => n8831, A2 => n8830, ZN => n11523);
   U9674 : NOR2_X1 port map( A1 => RST, A2 => n11520, ZN => n11614);
   U9675 : AND2_X1 port map( A1 => n8824, A2 => n8823, ZN => n11520);
   U9676 : NOR2_X1 port map( A1 => RST, A2 => n11516, ZN => n11607);
   U9677 : AND2_X1 port map( A1 => n8815, A2 => n8814, ZN => n11516);
   U9678 : NOR2_X1 port map( A1 => RST, A2 => n11525, ZN => n11622);
   U9679 : AND2_X1 port map( A1 => n8837, A2 => n8836, ZN => n11525);
   U9680 : AND2_X1 port map( A1 => n8845, A2 => n8844, ZN => n11528);
   U9681 : NOR2_X1 port map( A1 => RST, A2 => n11526, ZN => n11624);
   U9682 : AND2_X1 port map( A1 => n8840, A2 => n8839, ZN => n11526);
   U9683 : INV_X1 port map( A => n11921, ZN => n8912);
   U9684 : INV_X1 port map( A => n11942, ZN => n8947);
   U9685 : INV_X1 port map( A => n11919, ZN => n8908);
   U9686 : INV_X1 port map( A => n11930, ZN => n8928);
   U9687 : INV_X1 port map( A => n11940, ZN => n8943);
   U9688 : INV_X1 port map( A => n11929, ZN => n8926);
   U9689 : INV_X1 port map( A => n11939, ZN => n8941);
   U9690 : INV_X1 port map( A => n11922, ZN => n8914);
   U9691 : INV_X1 port map( A => n11925, ZN => n8918);
   U9692 : INV_X1 port map( A => n11918, ZN => n8906);
   U9693 : INV_X1 port map( A => n11917, ZN => n8904);
   U9694 : INV_X1 port map( A => n11924, ZN => n8916);
   U9695 : INV_X1 port map( A => n11949, ZN => n8957);
   U9696 : INV_X1 port map( A => n11920, ZN => n8910);
   U9697 : INV_X1 port map( A => n11927, ZN => n8922);
   U9698 : INV_X1 port map( A => n11916, ZN => n8902);
   U9699 : INV_X1 port map( A => n11944, ZN => n8951);
   U9700 : NOR2_X1 port map( A1 => n564, A2 => n12002, ZN => n12003);
   U9701 : NOR2_X1 port map( A1 => n562, A2 => n11999, ZN => n12000);
   U9702 : NOR2_X1 port map( A1 => n560, A2 => n11996, ZN => n11997);
   U9703 : NOR2_X1 port map( A1 => n558, A2 => n11993, ZN => n11994);
   U9704 : NOR2_X1 port map( A1 => n556, A2 => n11990, ZN => n11991);
   U9705 : NOR2_X1 port map( A1 => n554, A2 => n11987, ZN => n11988);
   U9706 : NOR2_X1 port map( A1 => n548, A2 => n11978, ZN => n11979);
   U9707 : NOR2_X1 port map( A1 => n546, A2 => n11975, ZN => n11976);
   U9708 : OAI211_X1 port map( C1 => n192, C2 => n8190, A => n8711, B => n8707,
                           ZN => i_ADD_WS1_1_port);
   U9709 : INV_X1 port map( A => n10444, ZN => n10493);
   U9710 : NOR2_X1 port map( A1 => n8700, A2 => n192, ZN => n10866);
   U9711 : NOR2_X1 port map( A1 => n10848, A2 => RST, ZN => n10847);
   U9712 : AND2_X1 port map( A1 => n9446, A2 => n9556, ZN => n10495);
   U9713 : AND2_X1 port map( A1 => n9532, A2 => i_ALU_OP_2_port, ZN => n10469);
   U9714 : AND2_X2 port map( A1 => n10857, A2 => CU_I_CW_EX_18, ZN => n10848);
   U9715 : NOR2_X1 port map( A1 => IR_26_port, A2 => n10771, ZN => n8699);
   U9716 : INV_X1 port map( A => n10744, ZN => n8455);
   U9717 : OR2_X1 port map( A1 => n476, A2 => n477, ZN => n8316);
   U9718 : NOR3_X2 port map( A1 => i_ADD_WB_4_port, A2 => i_ADD_WB_3_port, A3 
                           => n8409, ZN => n11913);
   U9719 : INV_X1 port map( A => n10851, ZN => n12032);
   U9720 : AND2_X1 port map( A1 => n8981, A2 => n8980, ZN => n12043);
   U9721 : INV_X2 port map( A => n11511, ZN => n11509);
   U9722 : BUF_X2 port map( A => n11511, Z => n8520);
   U9723 : INV_X2 port map( A => n11461, ZN => n11460);
   U9724 : BUF_X2 port map( A => n11461, Z => n8515);
   U9725 : AOI21_X1 port map( B1 => n8960, B2 => n8803, A => n8799, ZN => 
                           n11461);
   U9726 : INV_X2 port map( A => n11470, ZN => n11469);
   U9727 : BUF_X2 port map( A => n11470, Z => n8517);
   U9728 : AOI21_X1 port map( B1 => n8964, B2 => n8803, A => n8801, ZN => 
                           n11470);
   U9729 : INV_X2 port map( A => n11477, ZN => n11476);
   U9730 : BUF_X2 port map( A => n11477, Z => n8519);
   U9731 : INV_X2 port map( A => n11475, ZN => n11474);
   U9732 : BUF_X2 port map( A => n11475, Z => n8518);
   U9733 : INV_X2 port map( A => n11464, ZN => n11463);
   U9734 : BUF_X2 port map( A => n11464, Z => n8516);
   U9735 : AOI21_X1 port map( B1 => n8962, B2 => n8803, A => n8800, ZN => 
                           n11464);
   U9736 : BUF_X2 port map( A => n11429, Z => n8612);
   U9737 : NOR2_X1 port map( A1 => RST, A2 => n11427, ZN => n11429);
   U9738 : INV_X2 port map( A => n11593, ZN => n11592);
   U9739 : BUF_X2 port map( A => n11593, Z => n8528);
   U9740 : INV_X2 port map( A => n11551, ZN => n11550);
   U9741 : BUF_X2 port map( A => n11551, Z => n8526);
   U9742 : AOI21_X1 port map( B1 => n8962, B2 => n8852, A => n8849, ZN => 
                           n11551);
   U9743 : INV_X2 port map( A => n11548, ZN => n11547);
   U9744 : BUF_X2 port map( A => n11548, Z => n8525);
   U9745 : AOI21_X1 port map( B1 => n8960, B2 => n7761, A => n8848, ZN => 
                           n11548);
   U9746 : INV_X2 port map( A => n11588, ZN => n11587);
   U9747 : BUF_X2 port map( A => n11588, Z => n8527);
   U9748 : AOI21_X1 port map( B1 => n8964, B2 => n7761, A => n8850, ZN => 
                           n11588);
   U9749 : INV_X2 port map( A => n11595, ZN => n11594);
   U9750 : BUF_X2 port map( A => n11595, Z => n8529);
   U9751 : INV_X2 port map( A => n11630, ZN => n11628);
   U9752 : BUF_X2 port map( A => n11630, Z => n8530);
   U9753 : INV_X2 port map( A => n11405, ZN => n11404);
   U9754 : BUF_X2 port map( A => n11405, Z => n8507);
   U9755 : AOI21_X1 port map( B1 => n8964, B2 => n7762, A => n8769, ZN => 
                           n11405);
   U9756 : INV_X2 port map( A => n11410, ZN => n11409);
   U9757 : BUF_X2 port map( A => n11410, Z => n8508);
   U9758 : INV_X2 port map( A => n11412, ZN => n11411);
   U9759 : BUF_X2 port map( A => n11412, Z => n8509);
   U9760 : INV_X2 port map( A => n11416, ZN => n11415);
   U9761 : BUF_X2 port map( A => n11416, Z => n8510);
   U9762 : BUF_X2 port map( A => n11399, Z => n8506);
   U9763 : INV_X2 port map( A => n11749, ZN => n11747);
   U9764 : BUF_X2 port map( A => n11749, Z => n8543);
   U9765 : BUF_X2 port map( A => n11713, Z => n8541);
   U9766 : INV_X2 port map( A => n11699, ZN => n11698);
   U9767 : BUF_X2 port map( A => n11699, Z => n8538);
   U9768 : AOI21_X1 port map( B1 => n8960, B2 => n8531, A => n8897, ZN => 
                           n11699);
   U9769 : INV_X2 port map( A => n11715, ZN => n11714);
   U9770 : BUF_X2 port map( A => n11715, Z => n8542);
   U9771 : INV_X2 port map( A => n11702, ZN => n11701);
   U9772 : BUF_X2 port map( A => n11702, Z => n8539);
   U9773 : AOI21_X1 port map( B1 => n8962, B2 => n8901, A => n8898, ZN => 
                           n11702);
   U9774 : BUF_X2 port map( A => n11708, Z => n8540);
   U9775 : OAI22_X1 port map( A1 => n9641, A2 => n9643, B1 => n12121, B2 => 
                           n8441, ZN => n12153);
   U9776 : OAI22_X1 port map( A1 => n9640, A2 => n8851, B1 => n11596, B2 => 
                           n12118, ZN => n11537);
   U9777 : INV_X1 port map( A => n11521, ZN => n11571);
   U9778 : INV_X1 port map( A => n11520, ZN => n11569);
   U9779 : INV_X1 port map( A => n11518, ZN => n11567);
   U9780 : INV_X1 port map( A => n11516, ZN => n11562);
   U9781 : INV_X1 port map( A => n11517, ZN => n11564);
   U9782 : INV_X1 port map( A => n11527, ZN => n11581);
   U9783 : INV_X1 port map( A => n11519, ZN => n11568);
   U9784 : INV_X1 port map( A => n11525, ZN => n11577);
   U9785 : INV_X1 port map( A => n11523, ZN => n11573);
   U9786 : BUF_X2 port map( A => n11832, Z => n8546);
   U9787 : INV_X2 port map( A => n11841, ZN => n11840);
   U9788 : BUF_X2 port map( A => n11841, Z => n8547);
   U9789 : INV_X2 port map( A => n11850, ZN => n11849);
   U9790 : BUF_X2 port map( A => n11850, Z => n8548);
   U9791 : INV_X2 port map( A => n11827, ZN => n11826);
   U9792 : BUF_X2 port map( A => n11827, Z => n8545);
   U9793 : AOI21_X1 port map( B1 => n8960, B2 => n8544, A => n8959, ZN => 
                           n11827);
   U9794 : AOI21_X1 port map( B1 => n8960, B2 => n7762, A => n8725, ZN => 
                           n12193);
   U9795 : AOI21_X1 port map( B1 => n8972, B2 => n8971, A => n8970, ZN => 
                           n12018);
   U9796 : AOI21_X1 port map( B1 => n8969, B2 => n8544, A => n8968, ZN => 
                           n11854);
   U9797 : NOR3_X1 port map( A1 => n527, A2 => i_ADD_WB_0_port, A3 => 
                           i_ADD_WB_1_port, ZN => n11901);
   U9798 : NOR3_X1 port map( A1 => n526, A2 => i_ADD_WB_0_port, A3 => 
                           i_ADD_WB_2_port, ZN => n11909);
   U9799 : NOR3_X1 port map( A1 => n527, A2 => n526, A3 => i_ADD_WB_0_port, ZN 
                           => n11893);
   U9800 : NOR3_X1 port map( A1 => n525, A2 => n526, A3 => i_ADD_WB_2_port, ZN 
                           => n11905);
   U9801 : NOR3_X1 port map( A1 => n527, A2 => n525, A3 => i_ADD_WB_1_port, ZN 
                           => n11897);
   U9802 : NOR3_X1 port map( A1 => n525, A2 => i_ADD_WB_2_port, A3 => 
                           i_ADD_WB_1_port, ZN => n11914);
   U9803 : NAND2_X1 port map( A1 => n10857, A2 => CU_I_CW_ID_19, ZN => n12207);
   U9804 : INV_X1 port map( A => n10442, ZN => n10503);
   U9805 : INV_X1 port map( A => n10505, ZN => n10461);
   U9806 : INV_X1 port map( A => n10479, ZN => n10502);
   U9807 : INV_X1 port map( A => n10388, ZN => n10510);
   U9808 : AND4_X1 port map( A1 => n9804, A2 => n9803, A3 => n9802, A4 => n9801
                           , ZN => n8311);
   U9809 : INV_X1 port map( A => n10184, ZN => n10231);
   U9810 : OR2_X1 port map( A1 => n10021, A2 => n10115, ZN => n10184);
   U9811 : INV_X1 port map( A => n8094, ZN => n10229);
   U9812 : INV_X1 port map( A => n10182, ZN => n10232);
   U9813 : OR2_X1 port map( A1 => i_ALU_OP_0_port, A2 => i_ALU_OP_1_port, ZN =>
                           n10421);
   U9814 : NOR2_X1 port map( A1 => n8400, A2 => i_ALU_OP_1_port, ZN => n10492);
   U9815 : OR2_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_state_0_port, 
                           A2 => n838, ZN => n8713);
   U9816 : NOR2_X1 port map( A1 => n8455, A2 => n8308, ZN => n8454);
   U9817 : INV_X1 port map( A => RST, ZN => n8689);
   U9818 : INV_X1 port map( A => RST, ZN => n8690);
   U9819 : INV_X1 port map( A => RST, ZN => n8691);
   U9820 : OR2_X1 port map( A1 => RST, A2 => i_RF2, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3);
   U9821 : OR2_X1 port map( A1 => RST, A2 => i_RF1, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3);
   U9822 : INV_X1 port map( A => RST, ZN => n8694);
   U9823 : INV_X1 port map( A => RST, ZN => n8695);
   U9824 : OR2_X1 port map( A1 => n10921, A2 => n10920, ZN => n10926);
   U9825 : OR2_X1 port map( A1 => n10919, A2 => n10918, ZN => n10912);
   U9826 : NAND2_X1 port map( A1 => n10910, A2 => n10909, ZN => n10923);
   U9827 : OR2_X1 port map( A1 => n10740, A2 => n11391, ZN => n8716);
   U9828 : NAND3_X1 port map( A1 => n11889, A2 => n11913, A3 => n8692, ZN => 
                           n11892);
   U9829 : NAND3_X1 port map( A1 => n11914, A2 => n11913, A3 => n8692, ZN => 
                           n11948);
   U9830 : NAND3_X1 port map( A1 => n11909, A2 => n11913, A3 => n8692, ZN => 
                           n11912);
   U9831 : NAND3_X1 port map( A1 => n11901, A2 => n11913, A3 => n8692, ZN => 
                           n11904);
   U9832 : NAND3_X1 port map( A1 => n11905, A2 => n11913, A3 => n8692, ZN => 
                           n11908);
   U9833 : NAND3_X1 port map( A1 => n11893, A2 => n11913, A3 => n8692, ZN => 
                           n11896);
   U9834 : NAND3_X1 port map( A1 => n11897, A2 => n11913, A3 => n8692, ZN => 
                           n11900);
   U9835 : AND3_X1 port map( A1 => n10777, A2 => n10742, A3 => n10741, ZN => 
                           n10790);
   U9836 : OR3_X1 port map( A1 => n10759, A2 => IR_3_port, A3 => n8320, ZN => 
                           n10788);
   U9837 : NOR2_X2 port map( A1 => n10877, A2 => RST, ZN => n10851);
   U9838 : INV_X1 port map( A => n12058, ZN => n10846);
   U9839 : OR2_X1 port map( A1 => n11459, A2 => RST, ZN => n8799);
   U9840 : OR2_X1 port map( A1 => n11468, A2 => RST, ZN => n8801);
   U9841 : OR2_X1 port map( A1 => n11462, A2 => RST, ZN => n8800);
   U9842 : NOR2_X1 port map( A1 => n11329, A2 => n11348, ZN => n11357);
   U9843 : NOR2_X1 port map( A1 => n11305, A2 => n11325, ZN => n11329);
   U9844 : NOR2_X1 port map( A1 => DATA_SIZE_1_port, A2 => n11347, ZN => n11370
                           );
   U9845 : AOI21_X1 port map( B1 => n393, B2 => n8376, A => n11300, ZN => 
                           n11331);
   U9846 : INV_X1 port map( A => n11358, ZN => n11342);
   U9847 : NOR2_X1 port map( A1 => i_DATAMEM_RM, A2 => n11270, ZN => n11355);
   U9848 : NAND2_X1 port map( A1 => DATA_SIZE_1_port, A2 => n392, ZN => n11270)
                           ;
   U9849 : INV_X2 port map( A => i_DATAMEM_RM, ZN => n11305);
   U9850 : OR2_X1 port map( A1 => n11549, A2 => RST, ZN => n8849);
   U9851 : OR2_X1 port map( A1 => n11546, A2 => RST, ZN => n8848);
   U9852 : OR2_X1 port map( A1 => n11586, A2 => RST, ZN => n8850);
   U9853 : OR2_X1 port map( A1 => n11403, A2 => RST, ZN => n8769);
   U9854 : INV_X2 port map( A => n11399, ZN => n11398);
   U9855 : OR2_X1 port map( A1 => n11397, A2 => RST, ZN => n8751);
   U9856 : INV_X2 port map( A => n11713, ZN => n11712);
   U9857 : OR2_X1 port map( A1 => n11697, A2 => RST, ZN => n8897);
   U9858 : OR2_X1 port map( A1 => n11700, A2 => RST, ZN => n8898);
   U9859 : INV_X2 port map( A => n11708, ZN => n11707);
   U9860 : OR2_X1 port map( A1 => n11706, A2 => RST, ZN => n8899);
   U9861 : INV_X1 port map( A => n11526, ZN => n11579);
   U9862 : INV_X1 port map( A => n11522, ZN => n11572);
   U9863 : INV_X1 port map( A => n11524, ZN => n11574);
   U9864 : INV_X2 port map( A => n11832, ZN => n11831);
   U9865 : OR2_X1 port map( A1 => n11830, A2 => RST, ZN => n8961);
   U9866 : OR2_X1 port map( A1 => n11825, A2 => RST, ZN => n8959);
   U9867 : OR2_X1 port map( A1 => n11396, A2 => RST, ZN => n8725);
   U9868 : OR2_X1 port map( A1 => n11857, A2 => RST, ZN => n8970);
   U9869 : OR2_X1 port map( A1 => n11853, A2 => RST, ZN => n8968);
   U9870 : NAND2_X1 port map( A1 => n11456, A2 => n11893, ZN => n12109);
   U9871 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_12_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_12_port, B2 => n8680, ZN 
                           => n11928);
   U9872 : AOI22_X1 port map( A1 => n8679, A2 => 
                           DataPath_i_REG_LDSTR_OUT_16_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_16_port, B2 => n8680, ZN 
                           => n11932);
   U9873 : AOI22_X1 port map( A1 => n8679, A2 => 
                           DataPath_i_REG_LDSTR_OUT_18_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_18_port, B2 => n8680, ZN 
                           => n11934);
   U9874 : NOR3_X1 port map( A1 => n527, A2 => n525, A3 => n526, ZN => n11889);
   U9875 : AOI22_X1 port map( A1 => n8679, A2 => 
                           DataPath_i_REG_LDSTR_OUT_19_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_19_port, B2 => n8680, ZN 
                           => n11935);
   U9876 : AOI22_X1 port map( A1 => n8679, A2 => 
                           DataPath_i_REG_LDSTR_OUT_17_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_17_port, B2 => n8680, ZN 
                           => n11933);
   U9877 : INV_X1 port map( A => RST, ZN => n8692);
   U9878 : INV_X1 port map( A => RST, ZN => n8688);
   U9879 : INV_X1 port map( A => RST, ZN => n8693);
   U9880 : NOR2_X1 port map( A1 => n8700, A2 => n191, ZN => n10865);
   U9881 : AND2_X1 port map( A1 => n10746, A2 => n8062, ZN => n9276);
   U9882 : BUF_X1 port map( A => n8687, Z => n8686);
   U9883 : INV_X1 port map( A => n10498, ZN => n10376);
   U9884 : INV_X1 port map( A => n10495, ZN => n10462);
   U9885 : INV_X1 port map( A => n10507, ZN => n10476);
   U9886 : NAND2_X1 port map( A1 => i_ALU_OP_0_port, A2 => i_ALU_OP_1_port, ZN 
                           => n10452);
   U9887 : INV_X1 port map( A => n10421, ZN => n10450);
   U9888 : AND2_X1 port map( A1 => n7749, A2 => n7796, ZN => n9448);
   U9889 : AND2_X1 port map( A1 => n8673, A2 => DataPath_i_PIPLIN_A_31_port, ZN
                           => n9742);
   U9890 : INV_X1 port map( A => DP_OP_751_130_5637_n435, ZN => n9815);
   U9891 : AND2_X1 port map( A1 => n8673, A2 => DataPath_i_PIPLIN_A_29_port, ZN
                           => n9816);
   U9892 : BUF_X1 port map( A => n9721, Z => n8491);
   U9893 : INV_X1 port map( A => DP_OP_751_130_5637_n537, ZN => n9875);
   U9894 : INV_X1 port map( A => n9845, ZN => n10114);
   U9895 : AND2_X1 port map( A1 => n8673, A2 => DataPath_i_PIPLIN_A_28_port, ZN
                           => n9845);
   U9896 : BUF_X1 port map( A => n9494, Z => n8577);
   U9897 : INV_X1 port map( A => n10143, ZN => n8552);
   U9898 : BUF_X1 port map( A => n10466, Z => n8496);
   U9899 : OAI21_X1 port map( B1 => n9506, B2 => DP_OP_751_130_5637_n843, A => 
                           n9505, ZN => n9507);
   U9900 : INV_X1 port map( A => DP_OP_751_130_5637_n741, ZN => n10011);
   U9901 : AND2_X1 port map( A1 => n8674, A2 => DataPath_i_PIPLIN_A_26_port, ZN
                           => n9919);
   U9902 : OAI21_X1 port map( B1 => n8321, B2 => n8683, A => n9495, ZN => 
                           DP_OP_751_130_5637_n843);
   U9903 : AND2_X1 port map( A1 => n8674, A2 => DataPath_i_PIPLIN_A_25_port, ZN
                           => n9938);
   U9904 : INV_X1 port map( A => n9603, ZN => n9625);
   U9905 : INV_X1 port map( A => n10281, ZN => n9979);
   U9906 : AND2_X1 port map( A1 => n8674, A2 => DataPath_i_PIPLIN_A_24_port, ZN
                           => n10281);
   U9907 : OAI21_X2 port map( B1 => n7793, B2 => n10379, A => n9480, ZN => 
                           n9481);
   U9908 : BUF_X1 port map( A => n9454, Z => n8568);
   U9909 : OAI21_X2 port map( B1 => n7771, B2 => n10419, A => n9468, ZN => 
                           n9469);
   U9910 : OAI21_X1 port map( B1 => n8340, B2 => n8683, A => n9459, ZN => 
                           DP_OP_751_130_5637_n1455);
   U9911 : OAI21_X1 port map( B1 => n8341, B2 => n8138, A => n9460, ZN => 
                           n10446);
   U9912 : BUF_X1 port map( A => n9455, Z => n8569);
   U9913 : INV_X1 port map( A => n417, ZN => n8676);
   U9914 : OR2_X1 port map( A1 => DP_OP_751_130_5637_n1761, A2 => n10467, ZN =>
                           n10273);
   U9915 : INV_X2 port map( A => DRAMRF_READY, ZN => n10868);
   U9916 : AND2_X2 port map( A1 => n10856, A2 => n8413, ZN => n10855);
   U9917 : OAI22_X1 port map( A1 => n9644, A2 => n8900, B1 => n12158, B2 => 
                           n8442, ZN => n11692);
   U9918 : AOI211_X4 port map( C1 => n11844, C2 => DataPath_RF_c_win_3_port, A 
                           => RST, B => n11471, ZN => n11473);
   U9919 : AOI211_X4 port map( C1 => n11835, C2 => DataPath_RF_c_win_3_port, A 
                           => RST, B => n11465, ZN => n11467);
   U9920 : AOI211_X4 port map( C1 => DataPath_RF_c_win_4_port, C2 => n11844, A 
                           => RST, B => n11406, ZN => n11408);
   U9921 : AOI211_X4 port map( C1 => DataPath_RF_c_win_4_port, C2 => n11835, A 
                           => RST, B => n11400, ZN => n11402);
   U9922 : OAI222_X4 port map( A1 => n8851, A2 => n8966, B1 => n11596, B2 => 
                           n11589, C1 => n8442, C2 => n11842, ZN => n11590);
   U9923 : AOI211_X4 port map( C1 => DataPath_RF_c_win_1_port, C2 => n11844, A 
                           => RST, B => n11709, ZN => n11711);
   U9924 : AOI211_X4 port map( C1 => DataPath_RF_c_win_1_port, C2 => n11835, A 
                           => RST, B => n11703, ZN => n11705);
   U9925 : AOI211_X4 port map( C1 => DataPath_RF_c_win_0_port, C2 => n11844, A 
                           => RST, B => n11843, ZN => n11846);
   U9926 : AOI211_X4 port map( C1 => DataPath_RF_c_win_0_port, C2 => n11835, A 
                           => RST, B => n11834, ZN => n11837);
   U9927 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_15_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_15_port, B2 => n8411, ZN 
                           => n11931);
   U9928 : NOR3_X1 port map( A1 => i_ADD_WB_2_port, A2 => i_ADD_WB_0_port, A3 
                           => i_ADD_WB_1_port, ZN => n11455);
   U9929 : INV_X1 port map( A => i_NPC_SEL, ZN => n10577);
   U9930 : OR2_X2 port map( A1 => n8484, A2 => n9302, ZN => n10569);
   U9931 : OR2_X2 port map( A1 => n10638, A2 => n8101, ZN => n10571);
   U9932 : NOR2_X1 port map( A1 => n8503, A2 => n8502, ZN => n10707);
   U9933 : NOR2_X2 port map( A1 => n9427, A2 => n9561, ZN => n10498);
   U9934 : OAI21_X2 port map( B1 => n8322, B2 => n8683, A => n9509, ZN => 
                           DP_OP_751_130_5637_n639);
   U9935 : XNOR2_X2 port map( A => DP_OP_751_130_5637_n1251, B => n10379, ZN =>
                           n9482);
   U9936 : XNOR2_X2 port map( A => DP_OP_751_130_5637_n1353, B => n10337, ZN =>
                           n9475);
   U9937 : XNOR2_X2 port map( A => DP_OP_751_130_5637_n1455, B => n10419, ZN =>
                           n9470);
   U9938 : INV_X1 port map( A => n472, ZN => n8675);
   U9939 : XNOR2_X1 port map( A => n577, B => n823, ZN => n8721);
   U9940 : XNOR2_X1 port map( A => DataPath_RF_c_win_4_port, B => 
                           DataPath_RF_c_swin_4_port, ZN => n8722);
   U9941 : OAI221_X1 port map( B1 => DataPath_RF_c_swin_0_port, B2 => n8299, C1
                           => n8327, C2 => DataPath_RF_c_win_0_port, A => 
                           n10875, ZN => n10876);
   U9942 : MUX2_X1 port map( A => n5758, B => n8418, S => n10740, Z => n8795);
   U9943 : MUX2_X1 port map( A => n5830, B => n8416, S => n10740, Z => n8793);
   U9944 : MUX2_X1 port map( A => n5722, B => n8419, S => n10740, Z => n8796);
   U9945 : MUX2_X1 port map( A => n5614, B => n8422, S => n10740, Z => n8798);
   U9946 : MUX2_X1 port map( A => n5794, B => n8417, S => n10740, Z => n8794);
   U9947 : MUX2_X1 port map( A => n11417, B => n8410, S => n10740, Z => n8772);
   U9948 : MUX2_X1 port map( A => n5650, B => n8421, S => n10740, Z => n8797);
   U9949 : NOR2_X1 port map( A1 => n8440, A2 => n10795, ZN => CU_I_CW_IF_0);
   U9950 : OAI211_X1 port map( C1 => n8503, C2 => n10831, A => n10830, B => 
                           n10829, ZN => CU_I_CW_24_port);
   U9951 : NAND2_X1 port map( A1 => n10828, A2 => n10827, ZN => n10829);
   U9952 : AOI21_X1 port map( B1 => n10826, B2 => n8185, A => CU_I_CW_6_port, 
                           ZN => n10830);
   U9953 : AOI21_X1 port map( B1 => n8102, B2 => n10720, A => n10827, ZN => 
                           n10723);
   U9954 : NOR2_X1 port map( A1 => n10873, A2 => n10716, ZN => n10718);
   U9955 : NOR2_X1 port map( A1 => n10544, A2 => n10795, ZN => n10836);
   U9956 : AOI21_X1 port map( B1 => n10543, B2 => n8308, A => CU_I_CW_16_port, 
                           ZN => n10544);
   U9957 : NAND2_X1 port map( A1 => n8084, A2 => n8255, ZN => n9649);
   U9958 : OR2_X1 port map( A1 => n9648, A2 => n12022, ZN => n10542);
   U9959 : AOI21_X1 port map( B1 => n10826, B2 => n8080, A => n10768, ZN => 
                           n9648);
   U9960 : OAI211_X1 port map( C1 => n8973, C2 => n10721, A => n10715, B => 
                           n10714, ZN => CU_I_CW_22_port);
   U9961 : NAND4_X1 port map( A1 => n10873, A2 => n10744, A3 => n10720, A4 => 
                           n10713, ZN => n10714);
   U9962 : NAND2_X1 port map( A1 => n10712, A2 => n10711, ZN => n10721);
   U9963 : INV_X1 port map( A => n10710, ZN => n10712);
   U9964 : NAND2_X1 port map( A1 => n10709, A2 => n10708, ZN => CU_I_CW_21_port
                           );
   U9965 : NOR2_X1 port map( A1 => n12026, A2 => n10713, ZN => CU_I_CW_3_port);
   U9966 : NOR2_X1 port map( A1 => n10744, A2 => n10713, ZN => CU_I_CW_5_port);
   U9967 : OR2_X1 port map( A1 => n8084, A2 => n8080, ZN => n10713);
   U9968 : NOR2_X1 port map( A1 => n8453, A2 => n7773, ZN => 
                           DRAMRF_ADDRESS_31_port);
   U9969 : OAI21_X1 port map( B1 => n10740, B2 => n10736, A => n9645, ZN => 
                           DRAMRF_ISSUE);
   U9970 : INV_X1 port map( A => DRAMRF_READNOTWRITE_port, ZN => n9645);
   U9971 : OAI21_X1 port map( B1 => n10918, B2 => n8719, A => n8718, ZN => 
                           n10921);
   U9972 : AOI21_X1 port map( B1 => n10854, B2 => n10906, A => n8717, ZN => 
                           n10918);
   U9973 : INV_X1 port map( A => n10853, ZN => n8717);
   U9974 : INV_X1 port map( A => n10891, ZN => n10893);
   U9975 : INV_X1 port map( A => n10890, ZN => n10897);
   U9976 : INV_X1 port map( A => n10889, ZN => n10901);
   U9977 : INV_X1 port map( A => n10888, ZN => n10905);
   U9978 : NAND2_X1 port map( A1 => n8715, A2 => n8718, ZN => n10887);
   U9979 : AOI22_X1 port map( A1 => n8714, A2 => n12045, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, B2 => 
                           n8716, ZN => n8718);
   U9980 : INV_X1 port map( A => n8719, ZN => n8715);
   U9981 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, 
                           A2 => n10855, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, B2 => 
                           n8716, ZN => n10853);
   U9982 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, 
                           A2 => n10855, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, B2 => 
                           n8716, ZN => n10854);
   U9983 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port,
                           A2 => n10855, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, B2 => 
                           n8716, ZN => n10896);
   U9984 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port,
                           A2 => n10855, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, B2 => 
                           n8716, ZN => n10892);
   U9985 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, B2 => 
                           n8716, ZN => n10902);
   U9986 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, 
                           A2 => n10855, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, B2 => 
                           n8716, ZN => n10904);
   U9987 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, 
                           A2 => n10855, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, B2 => 
                           n8716, ZN => n10898);
   U9988 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, 
                           A2 => n10855, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, B2 => 
                           n8716, ZN => n10900);
   U9989 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, 
                           A2 => n10855, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, B2 => 
                           n8716, ZN => n10894);
   U9990 : OAI22_X1 port map( A1 => n8165, A2 => n12032, B1 => n10772, B2 => 
                           n12030, ZN => n7078);
   U9991 : OAI22_X1 port map( A1 => n12207, A2 => n10631, B1 => n12206, B2 => 
                           n8439, ZN => n6730);
   U9992 : AOI21_X1 port map( B1 => n10738, B2 => n10737, A => RST, ZN => n7068
                           );
   U9993 : NOR2_X1 port map( A1 => n10736, A2 => n12045, ZN => n10737);
   U9994 : INV_X1 port map( A => n12208, ZN => n10736);
   U9995 : NOR2_X1 port map( A1 => n10739, A2 => n12046, ZN => n7067);
   U9996 : INV_X1 port map( A => n10738, ZN => n10739);
   U9997 : NAND2_X1 port map( A1 => n8443, A2 => n838, ZN => n10738);
   U9998 : OAI211_X1 port map( C1 => n10763, C2 => n12026, A => n10762, B => 
                           n10761, ZN => n7084);
   U9999 : OAI22_X1 port map( A1 => n10781, A2 => n10788, B1 => n10766, B2 => 
                           n12029, ZN => n10760);
   U10000 : AOI21_X1 port map( B1 => i_ALU_OP_3_port, B2 => n10851, A => n10758
                           , ZN => n10762);
   U10001 : NOR3_X1 port map( A1 => n10772, A2 => n10757, A3 => n10756, ZN => 
                           n10758);
   U10002 : NOR2_X1 port map( A1 => n10740, A2 => RST, ZN => CU_I_N184);
   U10003 : NOR2_X1 port map( A1 => n10735, A2 => RST, ZN => 
                           DataPath_WRF_CUhw_N145);
   U10004 : AOI211_X1 port map( C1 => n10734, C2 => n8313, A => n10733, B => 
                           n10732, ZN => n10735);
   U10005 : OAI21_X1 port map( B1 => n10846, B2 => n8316, A => n10729, ZN => 
                           n10733);
   U10006 : OAI211_X1 port map( C1 => n235, C2 => n12032, A => n10793, B => 
                           n10792, ZN => n7080);
   U10007 : OAI211_X1 port map( C1 => n12032, C2 => n8438, A => n10755, B => 
                           n10754, ZN => n7082);
   U10008 : INV_X1 port map( A => n10751, ZN => n10753);
   U10009 : OAI21_X1 port map( B1 => IR_4_port, B2 => n210, A => n8315, ZN => 
                           n10750);
   U10010 : OAI211_X1 port map( C1 => n8380, C2 => n12032, A => n10745, B => 
                           n10747, ZN => n7079);
   U10011 : NAND2_X1 port map( A1 => IR_4_port, A2 => n12028, ZN => n10743);
   U10012 : OAI211_X1 port map( C1 => n8378, C2 => n12032, A => n10749, B => 
                           n10748, ZN => n7081);
   U10013 : NAND2_X1 port map( A1 => n10791, A2 => n8501, ZN => n10748);
   U10014 : NOR2_X1 port map( A1 => n10747, A2 => n10746, ZN => n10791);
   U10015 : OAI21_X1 port map( B1 => n10779, B2 => n210, A => n10778, ZN => 
                           n7085);
   U10016 : AOI211_X1 port map( C1 => n10777, C2 => n10776, A => n10775, B => 
                           n10774, ZN => n10778);
   U10017 : NOR3_X1 port map( A1 => n10773, A2 => n10772, A3 => n10771, ZN => 
                           n10774);
   U10018 : INV_X1 port map( A => n10716, ZN => n10768);
   U10019 : NOR2_X1 port map( A1 => n12032, A2 => n8681, ZN => n10775);
   U10020 : OAI22_X1 port map( A1 => n10767, A2 => n10788, B1 => n10766, B2 => 
                           n10765, ZN => n10776);
   U10021 : NAND2_X1 port map( A1 => n10764, A2 => n210, ZN => n10765);
   U10022 : INV_X1 port map( A => n10781, ZN => n10764);
   U10023 : INV_X1 port map( A => n10780, ZN => n10777);
   U10024 : INV_X1 port map( A => n10785, ZN => n10779);
   U10025 : NAND2_X1 port map( A1 => n10849, A2 => n10784, ZN => n7086);
   U10026 : AOI211_X1 port map( C1 => n10851, C2 => i_ALU_OP_1_port, A => 
                           n10783, B => n10782, ZN => n10784);
   U10027 : AOI211_X1 port map( C1 => n12025, C2 => n10781, A => n10788, B => 
                           n10780, ZN => n10782);
   U10028 : OAI21_X1 port map( B1 => n10788, B2 => n12027, A => n10787, ZN => 
                           n7083);
   U10029 : AOI211_X1 port map( C1 => n10850, C2 => n8501, A => n10786, B => 
                           n10785, ZN => n10787);
   U10030 : NOR2_X1 port map( A1 => n12032, A2 => n368, ZN => n10786);
   U10031 : INV_X1 port map( A => n10783, ZN => n10763);
   U10032 : INV_X1 port map( A => n10857, ZN => n10772);
   U10033 : AOI211_X1 port map( C1 => n8975, C2 => n10857, A => n8974, B => 
                           n10785, ZN => n10849);
   U10034 : NOR4_X1 port map( A1 => n10780, A2 => n12024, A3 => IR_1_port, A4 
                           => IR_2_port, ZN => n10785);
   U10035 : AOI211_X1 port map( C1 => n12029, C2 => n12025, A => n10766, B => 
                           n10780, ZN => n8974);
   U10036 : OR3_X1 port map( A1 => n10759, A2 => IR_3_port, A3 => IR_5_port, ZN
                           => n10766);
   U10037 : INV_X1 port map( A => n10715, ZN => n8975);
   U10038 : NAND2_X1 port map( A1 => n10857, A2 => n8997, ZN => n10780);
   U10039 : OR3_X1 port map( A1 => n10759, A2 => IR_5_port, A3 => n8318, ZN => 
                           n12024);
   U10040 : NAND2_X1 port map( A1 => n10742, A2 => n8317, ZN => n10759);
   U10041 : INV_X1 port map( A => n12043, ZN => n12037);
   U10042 : AOI21_X1 port map( B1 => n7695, B2 => IR_2_port, A => n10521, ZN =>
                           n2977);
   U10043 : OAI22_X1 port map( A1 => n12207, A2 => n10520, B1 => n12206, B2 => 
                           n8436, ZN => n10521);
   U10044 : NOR2_X1 port map( A1 => n10728, A2 => n8983, ZN => n10844);
   U10045 : INV_X1 port map( A => n12057, ZN => n8983);
   U10046 : NOR2_X1 port map( A1 => n8981, A2 => n8980, ZN => n12042);
   U10047 : AOI22_X1 port map( A1 => n7695, A2 => IR_1_port, B1 => 
                           DataPath_i_PIPLIN_IN1_1_port, B2 => n10871, ZN => 
                           n2981);
   U10048 : AOI22_X1 port map( A1 => n7695, A2 => n8427, B1 => 
                           DataPath_i_PIPLIN_IN1_0_port, B2 => n10871, ZN => 
                           n2982);
   U10049 : AOI22_X1 port map( A1 => n7695, A2 => n8391, B1 => 
                           DataPath_i_PIPLIN_IN1_14_port, B2 => n10871, ZN => 
                           n2965);
   U10050 : AOI22_X1 port map( A1 => n7695, A2 => IR_13_port, B1 => 
                           DataPath_i_PIPLIN_IN1_13_port, B2 => n10871, ZN => 
                           n2966);
   U10051 : AOI22_X1 port map( A1 => n7695, A2 => n8306, B1 => 
                           DataPath_i_PIPLIN_IN1_12_port, B2 => n10871, ZN => 
                           n2967);
   U10052 : AOI22_X1 port map( A1 => n7695, A2 => n8302, B1 => 
                           DataPath_i_PIPLIN_IN1_11_port, B2 => n10871, ZN => 
                           n2968);
   U10053 : AOI22_X1 port map( A1 => n7695, A2 => IR_10_port, B1 => 
                           DataPath_i_PIPLIN_IN1_10_port, B2 => n10871, ZN => 
                           n2969);
   U10054 : AOI22_X1 port map( A1 => n7695, A2 => IR_9_port, B1 => 
                           DataPath_i_PIPLIN_IN1_9_port, B2 => n10871, ZN => 
                           n2970);
   U10055 : AOI22_X1 port map( A1 => n7695, A2 => IR_8_port, B1 => 
                           DataPath_i_PIPLIN_IN1_8_port, B2 => n10871, ZN => 
                           n2971);
   U10056 : AOI22_X1 port map( A1 => n7695, A2 => IR_7_port, B1 => 
                           DataPath_i_PIPLIN_IN1_7_port, B2 => n10871, ZN => 
                           n2972);
   U10057 : AOI22_X1 port map( A1 => n7695, A2 => IR_6_port, B1 => 
                           DataPath_i_PIPLIN_IN1_6_port, B2 => n10871, ZN => 
                           n2973);
   U10058 : AOI22_X1 port map( A1 => n7695, A2 => n8304, B1 => 
                           DataPath_i_PIPLIN_IN1_15_port, B2 => n10871, ZN => 
                           n2963);
   U10059 : AOI22_X1 port map( A1 => n7695, A2 => IR_4_port, B1 => 
                           DataPath_i_PIPLIN_IN1_4_port, B2 => n10871, ZN => 
                           n2975);
   U10060 : AOI22_X1 port map( A1 => n7695, A2 => IR_3_port, B1 => 
                           DataPath_i_PIPLIN_IN1_3_port, B2 => n10871, ZN => 
                           n2976);
   U10061 : AOI22_X1 port map( A1 => n7695, A2 => IR_5_port, B1 => 
                           DataPath_i_PIPLIN_IN1_5_port, B2 => n10871, ZN => 
                           n2974);
   U10062 : OAI22_X1 port map( A1 => n10532, A2 => n12207, B1 => n12206, B2 => 
                           n8431, ZN => n7025);
   U10063 : INV_X1 port map( A => n10531, ZN => n10532);
   U10064 : OAI22_X1 port map( A1 => n10728, A2 => n8313, B1 => RST, B2 => 
                           n10727, ZN => n104);
   U10065 : AOI22_X1 port map( A1 => n10726, A2 => n10729, B1 => n477, B2 => 
                           n10868, ZN => n10727);
   U10066 : NAND2_X1 port map( A1 => n12208, A2 => n10725, ZN => n10729);
   U10067 : NAND2_X1 port map( A1 => n10724, A2 => n8313, ZN => n10726);
   U10068 : INV_X1 port map( A => n10845, ZN => n10728);
   U10069 : OAI22_X1 port map( A1 => n10538, A2 => n12207, B1 => n12206, B2 => 
                           n8432, ZN => n7022);
   U10070 : INV_X1 port map( A => n10537, ZN => n10538);
   U10071 : INV_X1 port map( A => n10515, ZN => n2491);
   U10072 : OAI22_X1 port map( A1 => n10514, A2 => n12207, B1 => n12206, B2 => 
                           n8435, ZN => n10515);
   U10073 : AND2_X1 port map( A1 => C620_DATA2_2, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_2_port);
   U10074 : AOI22_X1 port map( A1 => n10872, A2 => n10464, B1 => 
                           DataPath_i_PIPLIN_IN2_5_port, B2 => n10871, ZN => 
                           n2489);
   U10075 : AOI22_X1 port map( A1 => n10872, A2 => n10325, B1 => 
                           DataPath_i_PIPLIN_IN2_15_port, B2 => n10871, ZN => 
                           n2474);
   U10076 : AOI22_X1 port map( A1 => n10872, A2 => i_ADD_WS1_3_port, B1 => 
                           DataPath_i_PIPLIN_WRB1_3_port, B2 => n10871, ZN => 
                           n2987);
   U10077 : AOI22_X1 port map( A1 => n10872, A2 => n10391, B1 => 
                           DataPath_i_PIPLIN_IN2_11_port, B2 => n10871, ZN => 
                           n2480);
   U10078 : AOI22_X1 port map( A1 => n10872, A2 => n10438, B1 => 
                           DataPath_i_PIPLIN_IN2_9_port, B2 => n10871, ZN => 
                           n2483);
   U10079 : AOI22_X1 port map( A1 => n10872, A2 => i_ADD_WS1_4_port, B1 => 
                           DataPath_i_PIPLIN_WRB1_4_port, B2 => n10871, ZN => 
                           n2986);
   U10080 : AOI22_X1 port map( A1 => n10872, A2 => n9902, B1 => 
                           DataPath_i_PIPLIN_IN2_27_port, B2 => n10871, ZN => 
                           n2449);
   U10081 : AOI22_X1 port map( A1 => n10872, A2 => n10382, B1 => 
                           DataPath_i_PIPLIN_IN2_12_port, B2 => n10871, ZN => 
                           n2478);
   U10082 : AOI22_X1 port map( A1 => n10872, A2 => n10517, B1 => 
                           DataPath_i_PIPLIN_IN2_1_port, B2 => n10871, ZN => 
                           n2496);
   U10083 : AOI22_X1 port map( A1 => n10872, A2 => n10518, B1 => 
                           DataPath_i_PIPLIN_IN2_0_port, B2 => n10871, ZN => 
                           n2498);
   U10084 : AOI22_X1 port map( A1 => n10872, A2 => i_ADD_WS1_1_port, B1 => 
                           DataPath_i_PIPLIN_WRB1_1_port, B2 => n10871, ZN => 
                           n2989);
   U10085 : AOI22_X1 port map( A1 => n10872, A2 => i_ADD_WS1_0_port, B1 => 
                           DataPath_i_PIPLIN_WRB1_0_port, B2 => n10871, ZN => 
                           n2990);
   U10086 : AOI22_X1 port map( A1 => n10872, A2 => i_ADD_WS1_2_port, B1 => 
                           DataPath_i_PIPLIN_WRB1_2_port, B2 => n10871, ZN => 
                           n2988);
   U10087 : AOI22_X1 port map( A1 => n10872, A2 => n9812, B1 => 
                           DataPath_i_PIPLIN_IN2_30_port, B2 => n10871, ZN => 
                           n2443);
   U10088 : AOI22_X1 port map( A1 => n10872, A2 => n10070, B1 => 
                           DataPath_i_PIPLIN_IN2_22_port, B2 => n10871, ZN => 
                           n2459);
   U10089 : AOI22_X1 port map( A1 => n10872, A2 => n10248, B1 => 
                           DataPath_i_PIPLIN_IN2_17_port, B2 => n10871, ZN => 
                           n2469);
   U10090 : AOI22_X1 port map( A1 => n10872, A2 => n10212, B1 => 
                           DataPath_i_PIPLIN_IN2_18_port, B2 => n10871, ZN => 
                           n2467);
   U10091 : AOI22_X1 port map( A1 => n10872, A2 => n9790, B1 => 
                           DataPath_i_PIPLIN_IN2_31_port, B2 => n10871, ZN => 
                           n2441);
   U10092 : AOI22_X1 port map( A1 => n10872, A2 => n10000, B1 => 
                           DataPath_i_PIPLIN_IN2_24_port, B2 => n10871, ZN => 
                           n2455);
   U10093 : AOI22_X1 port map( A1 => n10872, A2 => n9836, B1 => 
                           DataPath_i_PIPLIN_IN2_29_port, B2 => n10871, ZN => 
                           n2445);
   U10094 : AOI22_X1 port map( A1 => n10872, A2 => n10135, B1 => 
                           DataPath_i_PIPLIN_IN2_20_port, B2 => n10871, ZN => 
                           n2463);
   U10095 : AOI22_X1 port map( A1 => n10872, A2 => n9931, B1 => 
                           DataPath_i_PIPLIN_IN2_26_port, B2 => n10871, ZN => 
                           n2451);
   U10096 : AOI22_X1 port map( A1 => n10872, A2 => n9864, B1 => 
                           DataPath_i_PIPLIN_IN2_28_port, B2 => n10871, ZN => 
                           n2447);
   U10097 : AOI22_X1 port map( A1 => n10872, A2 => n9963, B1 => 
                           DataPath_i_PIPLIN_IN2_25_port, B2 => n10871, ZN => 
                           n2453);
   U10098 : AOI22_X1 port map( A1 => n10872, A2 => n10102, B1 => 
                           DataPath_i_PIPLIN_IN2_21_port, B2 => n10871, ZN => 
                           n2461);
   U10099 : AOI22_X1 port map( A1 => n10872, A2 => n10037, B1 => 
                           DataPath_i_PIPLIN_IN2_23_port, B2 => n10871, ZN => 
                           n2457);
   U10100 : INV_X1 port map( A => n10530, ZN => n7026);
   U10101 : AOI22_X1 port map( A1 => n10872, A2 => n10173, B1 => 
                           DataPath_i_PIPLIN_IN2_19_port, B2 => n10871, ZN => 
                           n2465);
   U10102 : INV_X1 port map( A => n10534, ZN => n7024);
   U10103 : AOI22_X1 port map( A1 => n10872, A2 => n10533, B1 => 
                           DataPath_i_PIPLIN_IN2_10_port, B2 => n10871, ZN => 
                           n10534);
   U10104 : INV_X1 port map( A => n10528, ZN => n7027);
   U10105 : AOI22_X1 port map( A1 => n10872, A2 => n10527, B1 => 
                           DataPath_i_PIPLIN_IN2_3_port, B2 => n10871, ZN => 
                           n10528);
   U10106 : INV_X1 port map( A => n10536, ZN => n7023);
   U10107 : AOI22_X1 port map( A1 => n10872, A2 => n10535, B1 => 
                           DataPath_i_PIPLIN_IN2_13_port, B2 => n10871, ZN => 
                           n10536);
   U10108 : INV_X1 port map( A => n10540, ZN => n7021);
   U10109 : AOI22_X1 port map( A1 => n10872, A2 => n10539, B1 => 
                           DataPath_i_PIPLIN_IN2_16_port, B2 => n10871, ZN => 
                           n10540);
   U10110 : AND2_X1 port map( A1 => C620_DATA2_3, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_3_port);
   U10111 : AND2_X1 port map( A1 => C620_DATA2_4, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_4_port);
   U10112 : AND2_X1 port map( A1 => C620_DATA2_5, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_5_port);
   U10113 : OAI22_X1 port map( A1 => n9639, A2 => n8802, B1 => n577, B2 => 
                           n12115, ZN => n11427);
   U10114 : INV_X1 port map( A => n12140, ZN => n12141);
   U10115 : AND2_X1 port map( A1 => C620_DATA2_6, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_6_port);
   U10116 : INV_X1 port map( A => n11649, ZN => n11691);
   U10117 : INV_X1 port map( A => n11641, ZN => n11679);
   U10118 : INV_X1 port map( A => n11644, ZN => n11683);
   U10119 : INV_X1 port map( A => n11640, ZN => n11676);
   U10120 : INV_X1 port map( A => n11642, ZN => n11680);
   U10121 : INV_X1 port map( A => n11645, ZN => n11684);
   U10122 : INV_X1 port map( A => n11643, ZN => n11681);
   U10123 : INV_X1 port map( A => n11646, ZN => n11685);
   U10124 : INV_X1 port map( A => n11651, ZN => n11693);
   U10125 : INV_X1 port map( A => n11647, ZN => n11686);
   U10126 : INV_X1 port map( A => n11648, ZN => n11689);
   U10127 : INV_X1 port map( A => n11639, ZN => n11674);
   U10128 : INV_X1 port map( A => n11650, ZN => n11658);
   U10129 : OAI22_X1 port map( A1 => n9640, A2 => n8900, B1 => n12118, B2 => 
                           n8442, ZN => n11656);
   U10130 : OAI22_X1 port map( A1 => n9638, A2 => n8900, B1 => n12112, B2 => 
                           n8442, ZN => n11638);
   U10131 : INV_X1 port map( A => n12145, ZN => n12146);
   U10132 : INV_X1 port map( A => n12104, ZN => n12150);
   U10133 : INV_X1 port map( A => n12103, ZN => n12148);
   U10134 : INV_X1 port map( A => n12096, ZN => n12134);
   U10135 : INV_X1 port map( A => n12098, ZN => n12137);
   U10136 : INV_X1 port map( A => n12099, ZN => n12139);
   U10137 : INV_X1 port map( A => n12097, ZN => n12136);
   U10138 : INV_X1 port map( A => n12102, ZN => n12142);
   U10139 : INV_X1 port map( A => n12105, ZN => n12151);
   U10140 : INV_X1 port map( A => n12100, ZN => n12101);
   U10141 : INV_X1 port map( A => n12095, ZN => n12132);
   U10142 : OAI22_X1 port map( A1 => n9638, A2 => n8851, B1 => n11596, B2 => 
                           n12112, ZN => n11530);
   U10143 : INV_X1 port map( A => n11770, ZN => n11771);
   U10144 : OAI22_X1 port map( A1 => n9642, A2 => n8851, B1 => n11596, B2 => 
                           n12155, ZN => n11542);
   U10145 : INV_X1 port map( A => n11528, ZN => n11582);
   U10146 : INV_X1 port map( A => n11776, ZN => n11807);
   U10147 : INV_X1 port map( A => n11801, ZN => n11802);
   U10148 : INV_X1 port map( A => n11768, ZN => n11791);
   U10149 : OAI222_X1 port map( A1 => n8851, A2 => n8963, B1 => n11596, B2 => 
                           n11552, C1 => n8442, C2 => n11833, ZN => n11584);
   U10150 : INV_X1 port map( A => n11798, ZN => n11799);
   U10151 : INV_X1 port map( A => n11772, ZN => n11797);
   U10152 : INV_X1 port map( A => n11777, ZN => n11809);
   U10153 : INV_X1 port map( A => n11775, ZN => n11805);
   U10154 : INV_X1 port map( A => n11769, ZN => n11793);
   U10155 : INV_X1 port map( A => n11778, ZN => n11810);
   U10156 : INV_X1 port map( A => n11773, ZN => n11800);
   U10157 : OAI22_X1 port map( A1 => n8966, A2 => n8802, B1 => n11596, B2 => 
                           n11842, ZN => n11471);
   U10158 : OAI22_X1 port map( A1 => n8963, A2 => n8802, B1 => n11596, B2 => 
                           n11833, ZN => n11465);
   U10159 : OAI22_X1 port map( A1 => n8966, A2 => n9643, B1 => n577, B2 => 
                           n11842, ZN => n11406);
   U10160 : OAI22_X1 port map( A1 => n8963, A2 => n9643, B1 => n577, B2 => 
                           n11833, ZN => n11400);
   U10161 : INV_X1 port map( A => n12084, ZN => n10471);
   U10162 : AOI211_X1 port map( C1 => n10495, C2 => n10501, A => n9550, B => 
                           n9549, ZN => n12075);
   U10163 : OAI22_X1 port map( A1 => n10480, A2 => n10388, B1 => n10506, B2 => 
                           n10460, ZN => n9549);
   U10164 : OAI22_X1 port map( A1 => n10508, A2 => n10505, B1 => n10400, B2 => 
                           n10507, ZN => n9550);
   U10165 : AOI22_X1 port map( A1 => n10496, A2 => n10503, B1 => n10502, B2 => 
                           n10497, ZN => n12076);
   U10166 : AOI22_X1 port map( A1 => n10504, A2 => n10493, B1 => n10498, B2 => 
                           n10509, ZN => n12077);
   U10167 : OAI211_X1 port map( C1 => n9572, C2 => n9571, A => n9570, B => 
                           n9569, ZN => n12079);
   U10168 : AOI21_X1 port map( B1 => n9568, B2 => n10842, A => n9567, ZN => 
                           n9569);
   U10169 : OAI211_X1 port map( C1 => n9566, C2 => n10465, A => n9565, B => 
                           n9564, ZN => n9567);
   U10170 : XNOR2_X1 port map( A => n9561, B => n9560, ZN => n9566);
   U10171 : OAI21_X1 port map( B1 => n9573, B2 => n9559, A => n12080, ZN => 
                           n9568);
   U10172 : NAND2_X1 port map( A1 => DataPath_ALUhw_i_Q_EXTENDED_34_port, A2 =>
                           n8578, ZN => n9570);
   U10173 : XNOR2_X1 port map( A => n9558, B => n9573, ZN => n9571);
   U10174 : NOR2_X1 port map( A1 => n10491, A2 => n9557, ZN => n9558);
   U10175 : INV_X1 port map( A => n9591, ZN => n9557);
   U10176 : OAI211_X1 port map( C1 => n9419, C2 => n10181, A => n9359, B => 
                           n9358, ZN => n10504);
   U10177 : NAND2_X1 port map( A1 => n9374, A2 => n9562, ZN => n9358);
   U10178 : AOI21_X1 port map( B1 => n7785, B2 => n9544, A => n9357, ZN => 
                           n9359);
   U10179 : OAI211_X1 port map( C1 => n9379, C2 => n10183, A => n9356, B => 
                           n9355, ZN => n9357);
   U10180 : AOI22_X1 port map( A1 => n10288, A2 => n9542, B1 => n9983, B2 => 
                           n9917, ZN => n9356);
   U10181 : OAI21_X1 port map( B1 => n10511, B2 => n9372, A => n9344, ZN => 
                           n10494);
   U10182 : AOI211_X1 port map( C1 => n7785, C2 => n9535, A => n9343, B => 
                           n9342, ZN => n9344);
   U10183 : OAI21_X1 port map( B1 => n9579, B2 => n9951, A => n9341, ZN => 
                           n9342);
   U10184 : AOI22_X1 port map( A1 => n10288, A2 => n9534, B1 => n9983, B2 => 
                           n9953, ZN => n9341);
   U10185 : OAI21_X1 port map( B1 => n9952, B2 => n9434, A => n9338, ZN => 
                           n9343);
   U10186 : NAND2_X1 port map( A1 => n9433, A2 => n9730, ZN => n9338);
   U10187 : INV_X1 port map( A => n10490, ZN => n9572);
   U10188 : INV_X1 port map( A => n10842, ZN => n10484);
   U10189 : AOI21_X1 port map( B1 => n11959, B2 => n8901, A => n8857, ZN => 
                           n11667);
   U10190 : NOR2_X1 port map( A1 => n8531, A2 => n8908, ZN => n8857);
   U10191 : NAND4_X1 port map( A1 => n8408, A2 => n9426, A3 => n9425, A4 => 
                           n9424, ZN => n10501);
   U10192 : OR2_X1 port map( A1 => n9423, A2 => n8496, ZN => n9424);
   U10193 : AOI22_X1 port map( A1 => n9920, A2 => n10473, B1 => n9983, B2 => 
                           n10110, ZN => n9425);
   U10194 : NAND2_X1 port map( A1 => n9420, A2 => n9845, ZN => n9426);
   U10195 : NAND2_X1 port map( A1 => n9419, A2 => n10277, ZN => n9420);
   U10196 : NAND2_X1 port map( A1 => n10288, A2 => n9609, ZN => n9416);
   U10197 : NAND2_X1 port map( A1 => n9433, A2 => n9612, ZN => n9417);
   U10198 : NAND2_X1 port map( A1 => n9613, A2 => n10111, ZN => n9418);
   U10199 : OAI21_X1 port map( B1 => n9721, B2 => n9372, A => n9371, ZN => 
                           n10496);
   U10200 : AOI211_X1 port map( C1 => n7785, C2 => n9370, A => n9369, B => 
                           n9368, ZN => n9371);
   U10201 : OAI21_X1 port map( B1 => n9579, B2 => n9722, A => n9367, ZN => 
                           n9368);
   U10202 : AOI22_X1 port map( A1 => n10288, A2 => n9575, B1 => n9433, B2 => 
                           n9366, ZN => n9367);
   U10203 : OAI22_X1 port map( A1 => n9714, A2 => n9364, B1 => n9434, B2 => 
                           n10164, ZN => n9369);
   U10204 : INV_X1 port map( A => n9885, ZN => n9364);
   U10205 : INV_X1 port map( A => n9578, ZN => n9370);
   U10206 : INV_X1 port map( A => n9374, ZN => n9372);
   U10207 : NOR2_X1 port map( A1 => n10421, A2 => n7800, ZN => n10842);
   U10208 : NAND2_X1 port map( A1 => n9559, A2 => n9573, ZN => n12080);
   U10209 : OAI21_X1 port map( B1 => n10486, B2 => n10485, A => n9591, ZN => 
                           n9559);
   U10210 : NOR2_X1 port map( A1 => n9554, A2 => n8489, ZN => n10485);
   U10211 : NOR2_X1 port map( A1 => n10421, A2 => n8681, ZN => n10490);
   U10212 : AND2_X1 port map( A1 => n9595, A2 => n9592, ZN => n9573);
   U10213 : NOR2_X1 port map( A1 => n10486, A2 => n10483, ZN => n10491);
   U10214 : NAND2_X1 port map( A1 => n9554, A2 => n8488, ZN => n10483);
   U10215 : XNOR2_X1 port map( A => n8167, B => i_ALU_OP_2_port, ZN => n9554);
   U10216 : NAND2_X1 port map( A1 => n9591, A2 => n9590, ZN => n10486);
   U10217 : AND2_X1 port map( A1 => C620_DATA2_7, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_7_port);
   U10218 : OAI22_X1 port map( A1 => n8966, A2 => n8900, B1 => n8299, B2 => 
                           n11842, ZN => n11709);
   U10219 : OAI22_X1 port map( A1 => n8963, A2 => n8900, B1 => n8299, B2 => 
                           n11833, ZN => n11703);
   U10220 : OAI22_X1 port map( A1 => n9641, A2 => n8965, B1 => n8299, B2 => 
                           n12121, ZN => n11816);
   U10221 : OAI22_X1 port map( A1 => n8966, A2 => n8965, B1 => n11842, B2 => 
                           n8441, ZN => n11843);
   U10222 : OAI22_X1 port map( A1 => n8963, A2 => n8965, B1 => n11833, B2 => 
                           n8441, ZN => n11834);
   U10223 : AOI21_X1 port map( B1 => n11960, B2 => n8803, A => n8777, ZN => 
                           n11436);
   U10224 : NOR2_X1 port map( A1 => n8803, A2 => n8910, ZN => n8777);
   U10225 : AOI21_X1 port map( B1 => n11967, B2 => n8803, A => n8785, ZN => 
                           n11444);
   U10226 : NOR2_X1 port map( A1 => n8803, A2 => n8928, ZN => n8785);
   U10227 : AOI21_X1 port map( B1 => n11764, B2 => n8803, A => n8792, ZN => 
                           n11450);
   U10228 : NOR2_X1 port map( A1 => n8803, A2 => n8957, ZN => n8792);
   U10229 : AOI21_X1 port map( B1 => n11968, B2 => n8803, A => n8787, ZN => 
                           n11446);
   U10230 : NOR2_X1 port map( A1 => n8803, A2 => n8941, ZN => n8787);
   U10231 : AOI21_X1 port map( B1 => n11961, B2 => n8803, A => n8778, ZN => 
                           n11437);
   U10232 : NOR2_X1 port map( A1 => n8803, A2 => n8912, ZN => n8778);
   U10233 : AOI21_X1 port map( B1 => n11750, B2 => n8803, A => n8780, ZN => 
                           n11439);
   U10234 : NOR2_X1 port map( A1 => n8803, A2 => n8861, ZN => n8780);
   U10235 : AOI21_X1 port map( B1 => n11957, B2 => n8803, A => n8774, ZN => 
                           n11433);
   U10236 : NOR2_X1 port map( A1 => n8803, A2 => n8904, ZN => n8774);
   U10237 : AOI21_X1 port map( B1 => n11964, B2 => n8803, A => n8782, ZN => 
                           n11441);
   U10238 : NOR2_X1 port map( A1 => n8803, A2 => n8918, ZN => n8782);
   U10239 : AOI21_X1 port map( B1 => n11971, B2 => n8803, A => n8790, ZN => 
                           n11421);
   U10240 : NOR2_X1 port map( A1 => n8803, A2 => n8951, ZN => n8790);
   U10241 : AOI21_X1 port map( B1 => n11958, B2 => n8803, A => n8775, ZN => 
                           n11434);
   U10242 : NOR2_X1 port map( A1 => n8803, A2 => n8906, ZN => n8775);
   U10243 : AOI21_X1 port map( B1 => n11970, B2 => n8803, A => n8789, ZN => 
                           n11448);
   U10244 : NOR2_X1 port map( A1 => n8803, A2 => n8947, ZN => n8789);
   U10245 : AOI21_X1 port map( B1 => n11969, B2 => n8803, A => n8788, ZN => 
                           n11447);
   U10246 : NOR2_X1 port map( A1 => n8803, A2 => n8943, ZN => n8788);
   U10247 : AOI21_X1 port map( B1 => n11959, B2 => n8803, A => n8776, ZN => 
                           n11435);
   U10248 : NOR2_X1 port map( A1 => n8803, A2 => n8908, ZN => n8776);
   U10249 : AOI21_X1 port map( B1 => n11965, B2 => n8803, A => n8783, ZN => 
                           n11442);
   U10250 : NOR2_X1 port map( A1 => n8803, A2 => n8922, ZN => n8783);
   U10251 : INV_X1 port map( A => n12059, ZN => n8770);
   U10252 : AOI21_X1 port map( B1 => n11755, B2 => n8803, A => n8786, ZN => 
                           n11445);
   U10253 : NOR2_X1 port map( A1 => n8803, A2 => n8874, ZN => n8786);
   U10254 : AOI21_X1 port map( B1 => n11963, B2 => n8803, A => n8781, ZN => 
                           n11440);
   U10255 : NOR2_X1 port map( A1 => n8803, A2 => n8916, ZN => n8781);
   U10256 : AOI21_X1 port map( B1 => n11962, B2 => n8803, A => n8779, ZN => 
                           n11438);
   U10257 : NOR2_X1 port map( A1 => n8803, A2 => n8914, ZN => n8779);
   U10258 : AOI21_X1 port map( B1 => n11966, B2 => n8803, A => n8784, ZN => 
                           n11443);
   U10259 : NOR2_X1 port map( A1 => n8803, A2 => n8926, ZN => n8784);
   U10260 : AND2_X1 port map( A1 => C620_DATA2_8, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_8_port);
   U10261 : AOI21_X1 port map( B1 => n11956, B2 => n8803, A => n8773, ZN => 
                           n11432);
   U10262 : NOR2_X1 port map( A1 => n8803, A2 => n8902, ZN => n8773);
   U10263 : NAND2_X1 port map( A1 => n8531, A2 => n11760, ZN => n8886);
   U10264 : OR2_X1 port map( A1 => n8532, A2 => n11941, ZN => n8887);
   U10265 : NAND2_X1 port map( A1 => n8532, A2 => n11758, ZN => n8880);
   U10266 : OR2_X1 port map( A1 => n8901, A2 => n11937, ZN => n8881);
   U10267 : NAND2_X1 port map( A1 => n8531, A2 => n11752, ZN => n8868);
   U10268 : OR2_X1 port map( A1 => n8532, A2 => n11928, ZN => n8869);
   U10269 : AOI21_X1 port map( B1 => n11750, B2 => n8532, A => n8862, ZN => 
                           n11671);
   U10270 : NOR2_X1 port map( A1 => n8531, A2 => n8861, ZN => n8862);
   U10271 : AOI21_X1 port map( B1 => n11960, B2 => n7762, A => n8755, ZN => 
                           n12126);
   U10272 : NOR2_X1 port map( A1 => n7762, A2 => n8910, ZN => n8755);
   U10273 : NAND2_X1 port map( A1 => n8771, A2 => n11760, ZN => n8739);
   U10274 : OR2_X1 port map( A1 => n7762, A2 => n11941, ZN => n8740);
   U10275 : AOI21_X1 port map( B1 => n11970, B2 => n8771, A => n8741, ZN => 
                           n12147);
   U10276 : NOR2_X1 port map( A1 => n7762, A2 => n8947, ZN => n8741);
   U10277 : AOI21_X1 port map( B1 => n11957, B2 => n7762, A => n8752, ZN => 
                           n12123);
   U10278 : NOR2_X1 port map( A1 => n8771, A2 => n8904, ZN => n8752);
   U10279 : AOI21_X1 port map( B1 => n11764, B2 => n8532, A => n8896, ZN => 
                           n11694);
   U10280 : NOR2_X1 port map( A1 => n8532, A2 => n8957, ZN => n8896);
   U10281 : AOI21_X1 port map( B1 => n11968, B2 => n8901, A => n8884, ZN => 
                           n11687);
   U10282 : NOR2_X1 port map( A1 => n8532, A2 => n8941, ZN => n8884);
   U10283 : NAND2_X1 port map( A1 => n8532, A2 => n11759, ZN => n8882);
   U10284 : OR2_X1 port map( A1 => n8531, A2 => n11938, ZN => n8883);
   U10285 : AOI21_X1 port map( B1 => n11967, B2 => n8531, A => n8871, ZN => 
                           n11678);
   U10286 : NOR2_X1 port map( A1 => n8901, A2 => n8928, ZN => n8871);
   U10287 : AOI21_X1 port map( B1 => n11970, B2 => n8531, A => n8888, ZN => 
                           n11690);
   U10288 : NOR2_X1 port map( A1 => n8901, A2 => n8947, ZN => n8888);
   U10289 : AOI21_X1 port map( B1 => n11961, B2 => n8532, A => n8859, ZN => 
                           n11669);
   U10290 : NOR2_X1 port map( A1 => n8901, A2 => n8912, ZN => n8859);
   U10291 : AOI21_X1 port map( B1 => n11969, B2 => n8901, A => n8885, ZN => 
                           n11688);
   U10292 : NOR2_X1 port map( A1 => n8901, A2 => n8943, ZN => n8885);
   U10293 : NAND2_X1 port map( A1 => n8532, A2 => n11756, ZN => n8876);
   U10294 : OR2_X1 port map( A1 => n8532, A2 => n11935, ZN => n8877);
   U10295 : NAND2_X1 port map( A1 => n8531, A2 => n11757, ZN => n8878);
   U10296 : OR2_X1 port map( A1 => n8532, A2 => n11936, ZN => n8879);
   U10297 : OAI211_X1 port map( C1 => n8901, C2 => n8902, A => n8853, B => 
                           n8688, ZN => n8854);
   U10298 : NAND2_X1 port map( A1 => n8901, A2 => n11956, ZN => n8853);
   U10299 : AOI21_X1 port map( B1 => n11965, B2 => n8901, A => n8867, ZN => 
                           n11675);
   U10300 : NOR2_X1 port map( A1 => n8901, A2 => n8922, ZN => n8867);
   U10301 : AOI21_X1 port map( B1 => n11960, B2 => n8531, A => n8858, ZN => 
                           n11668);
   U10302 : NOR2_X1 port map( A1 => n8531, A2 => n8910, ZN => n8858);
   U10303 : NAND2_X1 port map( A1 => n8532, A2 => n11631, ZN => n8872);
   U10304 : OR2_X1 port map( A1 => n8901, A2 => n11931, ZN => n8873);
   U10305 : AOI21_X1 port map( B1 => n11963, B2 => n8901, A => n8863, ZN => 
                           n11672);
   U10306 : NOR2_X1 port map( A1 => n8532, A2 => n8916, ZN => n8863);
   U10307 : AOI21_X1 port map( B1 => n11969, B2 => n7762, A => n8738, ZN => 
                           n12144);
   U10308 : NOR2_X1 port map( A1 => n7762, A2 => n8943, ZN => n8738);
   U10309 : AOI21_X1 port map( B1 => n11958, B2 => n7762, A => n8753, ZN => 
                           n12124);
   U10310 : NOR2_X1 port map( A1 => n8771, A2 => n8906, ZN => n8753);
   U10311 : AOI21_X1 port map( B1 => n11959, B2 => n8771, A => n8754, ZN => 
                           n12125);
   U10312 : NOR2_X1 port map( A1 => n8771, A2 => n8908, ZN => n8754);
   U10313 : AOI21_X1 port map( B1 => n11966, B2 => n8532, A => n8870, ZN => 
                           n11677);
   U10314 : NOR2_X1 port map( A1 => n8901, A2 => n8926, ZN => n8870);
   U10315 : AOI21_X1 port map( B1 => n11958, B2 => n8531, A => n8856, ZN => 
                           n11666);
   U10316 : NOR2_X1 port map( A1 => n8901, A2 => n8906, ZN => n8856);
   U10317 : AOI21_X1 port map( B1 => n11755, B2 => n8531, A => n8875, ZN => 
                           n11682);
   U10318 : NOR2_X1 port map( A1 => n8532, A2 => n8874, ZN => n8875);
   U10319 : NAND2_X1 port map( A1 => n8532, A2 => n11751, ZN => n8865);
   U10320 : OR2_X1 port map( A1 => n8532, A2 => n11926, ZN => n8866);
   U10321 : NAND2_X1 port map( A1 => n8901, A2 => n11761, ZN => n8889);
   U10322 : OR2_X1 port map( A1 => n8531, A2 => n11943, ZN => n8890);
   U10323 : AOI21_X1 port map( B1 => n11962, B2 => n8531, A => n8860, ZN => 
                           n11670);
   U10324 : NOR2_X1 port map( A1 => n8531, A2 => n8914, ZN => n8860);
   U10325 : AOI21_X1 port map( B1 => n11971, B2 => n8901, A => n8891, ZN => 
                           n11657);
   U10326 : NOR2_X1 port map( A1 => n8901, A2 => n8951, ZN => n8891);
   U10327 : NAND2_X1 port map( A1 => n8901, A2 => n11763, ZN => n8894);
   U10328 : OR2_X1 port map( A1 => n8531, A2 => n11946, ZN => n8895);
   U10329 : NAND2_X1 port map( A1 => n8531, A2 => n11762, ZN => n8892);
   U10330 : OR2_X1 port map( A1 => n8532, A2 => n11945, ZN => n8893);
   U10331 : AOI21_X1 port map( B1 => n11957, B2 => n8532, A => n8855, ZN => 
                           n11665);
   U10332 : NOR2_X1 port map( A1 => n8901, A2 => n8904, ZN => n8855);
   U10333 : AOI21_X1 port map( B1 => n11964, B2 => n8901, A => n8864, ZN => 
                           n11673);
   U10334 : NOR2_X1 port map( A1 => n8532, A2 => n8918, ZN => n8864);
   U10335 : NAND2_X1 port map( A1 => n7761, A2 => n11762, ZN => n8842);
   U10336 : OR2_X1 port map( A1 => n7779, A2 => n11945, ZN => n8843);
   U10337 : NAND2_X1 port map( A1 => n7761, A2 => n11757, ZN => n8828);
   U10338 : OR2_X1 port map( A1 => n7761, A2 => n11936, ZN => n8829);
   U10339 : AOI21_X1 port map( B1 => n7779, B2 => n11968, A => n8834, ZN => 
                           n11575);
   U10340 : NOR2_X1 port map( A1 => n7761, A2 => n8941, ZN => n8834);
   U10341 : AOI21_X1 port map( B1 => n7779, B2 => n11961, A => n8809, ZN => 
                           n11557);
   U10342 : NOR2_X1 port map( A1 => n7779, A2 => n8912, ZN => n8809);
   U10343 : AOI21_X1 port map( B1 => n7779, B2 => n11969, A => n8835, ZN => 
                           n11576);
   U10344 : NOR2_X1 port map( A1 => n7761, A2 => n8943, ZN => n8835);
   U10345 : AOI21_X1 port map( B1 => n11971, B2 => n8771, A => n8744, ZN => 
                           n12149);
   U10346 : NOR2_X1 port map( A1 => n7762, A2 => n8951, ZN => n8744);
   U10347 : OAI211_X1 port map( C1 => n8771, C2 => n8928, A => n8767, B => 
                           n8688, ZN => n8768);
   U10348 : NAND2_X1 port map( A1 => n7762, A2 => n11967, ZN => n8767);
   U10349 : NAND2_X1 port map( A1 => n7762, A2 => n11761, ZN => n8742);
   U10350 : OR2_X1 port map( A1 => n8771, A2 => n11943, ZN => n8743);
   U10351 : NAND2_X1 port map( A1 => n7762, A2 => n11759, ZN => n8735);
   U10352 : OR2_X1 port map( A1 => n7762, A2 => n11938, ZN => n8736);
   U10353 : AOI21_X1 port map( B1 => n11961, B2 => n7762, A => n8756, ZN => 
                           n12127);
   U10354 : NOR2_X1 port map( A1 => n7762, A2 => n8912, ZN => n8756);
   U10355 : AOI21_X1 port map( B1 => n11963, B2 => n8771, A => n8759, ZN => 
                           n12130);
   U10356 : NOR2_X1 port map( A1 => n8771, A2 => n8916, ZN => n8759);
   U10357 : OAI211_X1 port map( C1 => n7779, C2 => n8957, A => n8846, B => 
                           n8688, ZN => n8847);
   U10358 : NAND2_X1 port map( A1 => n8852, A2 => n11764, ZN => n8846);
   U10359 : NAND2_X1 port map( A1 => n7762, A2 => n11751, ZN => n8761);
   U10360 : OR2_X1 port map( A1 => n7762, A2 => n11926, ZN => n8762);
   U10361 : AOI21_X1 port map( B1 => n11755, B2 => n8771, A => n8728, ZN => 
                           n12138);
   U10362 : NOR2_X1 port map( A1 => n7762, A2 => n8874, ZN => n8728);
   U10363 : NAND2_X1 port map( A1 => n7762, A2 => n11763, ZN => n8747);
   U10364 : OR2_X1 port map( A1 => n7762, A2 => n11946, ZN => n8748);
   U10365 : NAND2_X1 port map( A1 => n7762, A2 => n11758, ZN => n8733);
   U10366 : OR2_X1 port map( A1 => n7762, A2 => n11937, ZN => n8734);
   U10367 : NAND2_X1 port map( A1 => n8771, A2 => n11757, ZN => n8731);
   U10368 : OR2_X1 port map( A1 => n7762, A2 => n11936, ZN => n8732);
   U10369 : NAND2_X1 port map( A1 => n7762, A2 => n11762, ZN => n8745);
   U10370 : OR2_X1 port map( A1 => n7762, A2 => n11945, ZN => n8746);
   U10371 : NAND2_X1 port map( A1 => n7762, A2 => n11752, ZN => n8764);
   U10372 : OR2_X1 port map( A1 => n7762, A2 => n11928, ZN => n8765);
   U10373 : AOI21_X1 port map( B1 => n11962, B2 => n7762, A => n8757, ZN => 
                           n12128);
   U10374 : NOR2_X1 port map( A1 => n7762, A2 => n8914, ZN => n8757);
   U10375 : AOI21_X1 port map( B1 => n11964, B2 => n8771, A => n8760, ZN => 
                           n12131);
   U10376 : NOR2_X1 port map( A1 => n7762, A2 => n8918, ZN => n8760);
   U10377 : AOI21_X1 port map( B1 => n11956, B2 => n7762, A => n8750, ZN => 
                           n12122);
   U10378 : NOR2_X1 port map( A1 => n7762, A2 => n8902, ZN => n8750);
   U10379 : AOI21_X1 port map( B1 => n11965, B2 => n7762, A => n8763, ZN => 
                           n12133);
   U10380 : NOR2_X1 port map( A1 => n7762, A2 => n8922, ZN => n8763);
   U10381 : AOI21_X1 port map( B1 => n11966, B2 => n8771, A => n8766, ZN => 
                           n12135);
   U10382 : NOR2_X1 port map( A1 => n7762, A2 => n8926, ZN => n8766);
   U10383 : AOI21_X1 port map( B1 => n11750, B2 => n8771, A => n8758, ZN => 
                           n12129);
   U10384 : NOR2_X1 port map( A1 => n8771, A2 => n8861, ZN => n8758);
   U10385 : AOI21_X1 port map( B1 => n9643, B2 => n8688, A => n8726, ZN => 
                           n8727);
   U10386 : INV_X1 port map( A => n3341, ZN => n8726);
   U10387 : AOI21_X1 port map( B1 => n11968, B2 => n7762, A => n8737, ZN => 
                           n12143);
   U10388 : NOR2_X1 port map( A1 => n8771, A2 => n8941, ZN => n8737);
   U10389 : NAND2_X1 port map( A1 => n7762, A2 => n11756, ZN => n8729);
   U10390 : OR2_X1 port map( A1 => n7762, A2 => n11935, ZN => n8730);
   U10391 : NAND2_X1 port map( A1 => n7779, A2 => n11756, ZN => n8826);
   U10392 : OR2_X1 port map( A1 => n7761, A2 => n11935, ZN => n8827);
   U10393 : AOI21_X1 port map( B1 => n7779, B2 => n11750, A => n8811, ZN => 
                           n11559);
   U10394 : NOR2_X1 port map( A1 => n8852, A2 => n8861, ZN => n8811);
   U10395 : INV_X1 port map( A => n11923, ZN => n8861);
   U10396 : NAND2_X1 port map( A1 => n7761, A2 => n11631, ZN => n8821);
   U10397 : OR2_X1 port map( A1 => n7761, A2 => n11931, ZN => n8822);
   U10398 : AOI21_X1 port map( B1 => n7779, B2 => n11959, A => n8807, ZN => 
                           n11555);
   U10399 : NOR2_X1 port map( A1 => n7761, A2 => n8908, ZN => n8807);
   U10400 : AOI21_X1 port map( B1 => n7779, B2 => n11971, A => n8841, ZN => 
                           n11580);
   U10401 : NOR2_X1 port map( A1 => n7779, A2 => n8951, ZN => n8841);
   U10402 : NAND2_X1 port map( A1 => n7779, A2 => n11752, ZN => n8817);
   U10403 : OR2_X1 port map( A1 => n7779, A2 => n11928, ZN => n8818);
   U10404 : NAND2_X1 port map( A1 => n7761, A2 => n11759, ZN => n8832);
   U10405 : OR2_X1 port map( A1 => n8852, A2 => n11938, ZN => n8833);
   U10406 : NAND2_X1 port map( A1 => n7761, A2 => n11758, ZN => n8830);
   U10407 : OR2_X1 port map( A1 => n8852, A2 => n11937, ZN => n8831);
   U10408 : AOI21_X1 port map( B1 => n7761, B2 => n11966, A => n8819, ZN => 
                           n11565);
   U10409 : NOR2_X1 port map( A1 => n7779, A2 => n8926, ZN => n8819);
   U10410 : AOI21_X1 port map( B1 => n11967, B2 => n8852, A => n8820, ZN => 
                           n11566);
   U10411 : NOR2_X1 port map( A1 => n7761, A2 => n8928, ZN => n8820);
   U10412 : AOI21_X1 port map( B1 => n7761, B2 => n11755, A => n8825, ZN => 
                           n11570);
   U10413 : NOR2_X1 port map( A1 => n7779, A2 => n8874, ZN => n8825);
   U10414 : INV_X1 port map( A => n11934, ZN => n8874);
   U10415 : NAND2_X1 port map( A1 => n8852, A2 => n11633, ZN => n8823);
   U10416 : OR2_X1 port map( A1 => n7761, A2 => n11632, ZN => n8824);
   U10417 : NAND2_X1 port map( A1 => n7779, A2 => n11751, ZN => n8814);
   U10418 : OR2_X1 port map( A1 => n7761, A2 => n11926, ZN => n8815);
   U10419 : AOI21_X1 port map( B1 => n7779, B2 => n11957, A => n8805, ZN => 
                           n11554);
   U10420 : NOR2_X1 port map( A1 => n7779, A2 => n8904, ZN => n8805);
   U10421 : NAND2_X1 port map( A1 => n7761, A2 => n11760, ZN => n8836);
   U10422 : OR2_X1 port map( A1 => n8852, A2 => n11941, ZN => n8837);
   U10423 : AOI21_X1 port map( B1 => n8852, B2 => n11962, A => n8810, ZN => 
                           n11558);
   U10424 : NOR2_X1 port map( A1 => n7761, A2 => n8914, ZN => n8810);
   U10425 : AOI21_X1 port map( B1 => n7779, B2 => n11958, A => n8806, ZN => 
                           n11540);
   U10426 : NOR2_X1 port map( A1 => n7761, A2 => n8906, ZN => n8806);
   U10427 : AOI21_X1 port map( B1 => n8852, B2 => n11964, A => n8813, ZN => 
                           n11561);
   U10428 : NOR2_X1 port map( A1 => n8852, A2 => n8918, ZN => n8813);
   U10429 : AOI21_X1 port map( B1 => n7779, B2 => n11960, A => n8808, ZN => 
                           n11556);
   U10430 : NOR2_X1 port map( A1 => n7779, A2 => n8910, ZN => n8808);
   U10431 : AOI21_X1 port map( B1 => n11956, B2 => n8852, A => n8804, ZN => 
                           n11553);
   U10432 : NOR2_X1 port map( A1 => n7779, A2 => n8902, ZN => n8804);
   U10433 : AOI21_X1 port map( B1 => n7779, B2 => n11963, A => n8812, ZN => 
                           n11560);
   U10434 : NOR2_X1 port map( A1 => n8852, A2 => n8916, ZN => n8812);
   U10435 : NAND2_X1 port map( A1 => n8852, A2 => n11763, ZN => n8844);
   U10436 : OR2_X1 port map( A1 => n7779, A2 => n11946, ZN => n8845);
   U10437 : NAND2_X1 port map( A1 => n7761, A2 => n11761, ZN => n8839);
   U10438 : OR2_X1 port map( A1 => n8852, A2 => n11943, ZN => n8840);
   U10439 : AOI21_X1 port map( B1 => n7761, B2 => n11965, A => n8816, ZN => 
                           n11563);
   U10440 : NOR2_X1 port map( A1 => n7761, A2 => n8922, ZN => n8816);
   U10441 : AOI21_X1 port map( B1 => n7779, B2 => n11970, A => n8838, ZN => 
                           n11578);
   U10442 : NOR2_X1 port map( A1 => n7761, A2 => n8947, ZN => n8838);
   U10443 : AOI21_X1 port map( B1 => n11961, B2 => n8971, A => n8913, ZN => 
                           n11787);
   U10444 : NOR2_X1 port map( A1 => n8544, A2 => n8912, ZN => n8913);
   U10445 : AOI21_X1 port map( B1 => n11970, B2 => n8971, A => n8948, ZN => 
                           n11806);
   U10446 : NOR2_X1 port map( A1 => n8544, A2 => n8947, ZN => n8948);
   U10447 : NAND2_X1 port map( A1 => n8971, A2 => n11752, ZN => n8924);
   U10448 : OR2_X1 port map( A1 => n8971, A2 => n11928, ZN => n8925);
   U10449 : NAND2_X1 port map( A1 => n8544, A2 => n11754, ZN => n8930);
   U10450 : OR2_X1 port map( A1 => n8544, A2 => n11753, ZN => n8931);
   U10451 : NAND2_X1 port map( A1 => n8971, A2 => n11759, ZN => n8939);
   U10452 : OR2_X1 port map( A1 => n8971, A2 => n11938, ZN => n8940);
   U10453 : NAND2_X1 port map( A1 => n8544, A2 => n11762, ZN => n8953);
   U10454 : OR2_X1 port map( A1 => n8971, A2 => n11945, ZN => n8954);
   U10455 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_7_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_7_port, B2 => n8680, ZN =>
                           n11923);
   U10456 : AOI21_X1 port map( B1 => n11959, B2 => n8971, A => n8909, ZN => 
                           n11767);
   U10457 : NOR2_X1 port map( A1 => n8971, A2 => n8908, ZN => n8909);
   U10458 : NAND2_X1 port map( A1 => n8544, A2 => n11760, ZN => n8945);
   U10459 : OR2_X1 port map( A1 => n8544, A2 => n11941, ZN => n8946);
   U10460 : AOI21_X1 port map( B1 => n11967, B2 => n8544, A => n8929, ZN => 
                           n11795);
   U10461 : NOR2_X1 port map( A1 => n8544, A2 => n8928, ZN => n8929);
   U10462 : AOI21_X1 port map( B1 => n11969, B2 => n8971, A => n8944, ZN => 
                           n11804);
   U10463 : NOR2_X1 port map( A1 => n8971, A2 => n8943, ZN => n8944);
   U10464 : NAND2_X1 port map( A1 => n11375, A2 => n11374, ZN => n12057);
   U10465 : AOI21_X1 port map( B1 => n11966, B2 => n8971, A => n8927, ZN => 
                           n11794);
   U10466 : NOR2_X1 port map( A1 => n8544, A2 => n8926, ZN => n8927);
   U10467 : AOI21_X1 port map( B1 => n11968, B2 => n8544, A => n8942, ZN => 
                           n11803);
   U10468 : NOR2_X1 port map( A1 => n8971, A2 => n8941, ZN => n8942);
   U10469 : AOI21_X1 port map( B1 => n11962, B2 => n8971, A => n8915, ZN => 
                           n11788);
   U10470 : NOR2_X1 port map( A1 => n8971, A2 => n8914, ZN => n8915);
   U10471 : AOI21_X1 port map( B1 => n11964, B2 => n8544, A => n8919, ZN => 
                           n11790);
   U10472 : NOR2_X1 port map( A1 => n8971, A2 => n8918, ZN => n8919);
   U10473 : NAND2_X1 port map( A1 => n8971, A2 => n11751, ZN => n8920);
   U10474 : OR2_X1 port map( A1 => n8971, A2 => n11926, ZN => n8921);
   U10475 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_10_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_10_port, B2 => n8411, ZN 
                           => n11926);
   U10476 : AOI21_X1 port map( B1 => n11958, B2 => n8971, A => n8907, ZN => 
                           n11785);
   U10477 : NOR2_X1 port map( A1 => n8544, A2 => n8906, ZN => n8907);
   U10478 : NAND2_X1 port map( A1 => n8971, A2 => n11756, ZN => n8933);
   U10479 : OR2_X1 port map( A1 => n8544, A2 => n11935, ZN => n8934);
   U10480 : AOI21_X1 port map( B1 => n11957, B2 => n8544, A => n8905, ZN => 
                           n11784);
   U10481 : NOR2_X1 port map( A1 => n8971, A2 => n8904, ZN => n8905);
   U10482 : NAND2_X1 port map( A1 => n8544, A2 => n11757, ZN => n8935);
   U10483 : OR2_X1 port map( A1 => n8971, A2 => n11936, ZN => n8936);
   U10484 : AOI21_X1 port map( B1 => n11963, B2 => n8544, A => n8917, ZN => 
                           n11789);
   U10485 : NOR2_X1 port map( A1 => n8544, A2 => n8916, ZN => n8917);
   U10486 : AOI21_X1 port map( B1 => n11764, B2 => n8971, A => n8958, ZN => 
                           n11811);
   U10487 : NOR2_X1 port map( A1 => n8971, A2 => n8957, ZN => n8958);
   U10488 : AOI21_X1 port map( B1 => n11960, B2 => n8544, A => n8911, ZN => 
                           n11786);
   U10489 : NOR2_X1 port map( A1 => n8544, A2 => n8910, ZN => n8911);
   U10490 : AOI21_X1 port map( B1 => n11965, B2 => n8544, A => n8923, ZN => 
                           n11792);
   U10491 : NOR2_X1 port map( A1 => n8971, A2 => n8922, ZN => n8923);
   U10492 : NAND2_X1 port map( A1 => n8965, A2 => n8688, ZN => n8932);
   U10493 : AOI21_X1 port map( B1 => n11956, B2 => n8971, A => n8903, ZN => 
                           n11783);
   U10494 : NOR2_X1 port map( A1 => n8971, A2 => n8902, ZN => n8903);
   U10495 : NAND2_X1 port map( A1 => n8544, A2 => n11763, ZN => n8955);
   U10496 : OR2_X1 port map( A1 => n8971, A2 => n11946, ZN => n8956);
   U10497 : NAND2_X1 port map( A1 => n8971, A2 => n11758, ZN => n8937);
   U10498 : OR2_X1 port map( A1 => n8544, A2 => n11937, ZN => n8938);
   U10499 : AOI21_X1 port map( B1 => n11971, B2 => n8971, A => n8952, ZN => 
                           n11808);
   U10500 : NOR2_X1 port map( A1 => n8971, A2 => n8951, ZN => n8952);
   U10501 : INV_X1 port map( A => n11375, ZN => n10852);
   U10502 : NAND2_X1 port map( A1 => n8971, A2 => n11761, ZN => n8949);
   U10503 : OR2_X1 port map( A1 => n8544, A2 => n11943, ZN => n8950);
   U10504 : AOI22_X1 port map( A1 => n8679, A2 => 
                           DataPath_i_REG_LDSTR_OUT_27_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_27_port, B2 => n8411, ZN 
                           => n11943);
   U10505 : AND2_X1 port map( A1 => C620_DATA2_9, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_9_port);
   U10506 : NAND2_X1 port map( A1 => n9628, A2 => n8681, ZN => n9419);
   U10507 : INV_X1 port map( A => n9433, ZN => n9379);
   U10508 : NAND2_X1 port map( A1 => n9423, A2 => n9980, ZN => n9374);
   U10509 : INV_X1 port map( A => n10480, ZN => n10500);
   U10510 : NOR2_X1 port map( A1 => n9395, A2 => n9394, ZN => n10480);
   U10511 : NOR2_X1 port map( A1 => n9423, A2 => n9659, ZN => n9394);
   U10512 : NAND2_X1 port map( A1 => n9628, A2 => i_ALU_OP_2_port, ZN => n9423)
                           ;
   U10513 : NAND4_X1 port map( A1 => n9393, A2 => n9392, A3 => n9391, A4 => 
                           n9390, ZN => n9395);
   U10514 : NAND2_X1 port map( A1 => n9628, A2 => n9389, ZN => n9390);
   U10515 : INV_X1 port map( A => n12091, ZN => n9389);
   U10516 : AOI22_X1 port map( A1 => n9433, A2 => n9388, B1 => n10028, B2 => 
                           n9983, ZN => n9391);
   U10517 : INV_X1 port map( A => n9779, ZN => n9388);
   U10518 : INV_X1 port map( A => n9385, ZN => n9392);
   U10519 : OAI22_X1 port map( A1 => n9434, A2 => n9384, B1 => n9980, B2 => 
                           n9659, ZN => n9385);
   U10520 : INV_X1 port map( A => n10026, ZN => n9384);
   U10521 : OR2_X1 port map( A1 => n10284, A2 => n12085, ZN => n9434);
   U10522 : AOI22_X1 port map( A1 => n10288, A2 => n9630, B1 => n7785, B2 => 
                           n9742, ZN => n9393);
   U10523 : NAND2_X1 port map( A1 => n9653, A2 => n9634, ZN => n12083);
   U10524 : AND2_X1 port map( A1 => n9654, A2 => n10450, ZN => n10837);
   U10525 : OR2_X1 port map( A1 => n9654, A2 => n10421, ZN => n12084);
   U10526 : OAI21_X1 port map( B1 => n12206, B2 => n8386, A => n10525, ZN => 
                           n116);
   U10527 : INV_X1 port map( A => n10477, ZN => n10506);
   U10528 : NAND4_X1 port map( A1 => n9444, A2 => n9443, A3 => n9442, A4 => 
                           n9441, ZN => n10477);
   U10529 : NAND2_X1 port map( A1 => n9440, A2 => n10113, ZN => n9441);
   U10530 : OAI22_X1 port map( A1 => n10291, A2 => n12085, B1 => n12087, B2 => 
                           n9979, ZN => n9440);
   U10531 : NAND2_X1 port map( A1 => n9628, A2 => n9987, ZN => n9442);
   U10532 : INV_X1 port map( A => n9439, ZN => n9443);
   U10533 : OAI22_X1 port map( A1 => n8094, A2 => n10275, B1 => n10182, B2 => 
                           n10283, ZN => n9439);
   U10534 : AOI22_X1 port map( A1 => n10282, A2 => n7772, B1 => n7785, B2 => 
                           n10285, ZN => n9444);
   U10535 : INV_X1 port map( A => n10478, ZN => n10508);
   U10536 : AND2_X1 port map( A1 => C620_DATA2_10, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_10_port);
   U10537 : OAI22_X1 port map( A1 => n10526, A2 => n10525, B1 => n494, B2 => 
                           n12206, ZN => n7104);
   U10538 : NAND2_X1 port map( A1 => n10523, A2 => n10872, ZN => n10525);
   U10539 : OAI21_X1 port map( B1 => n10414, B2 => n10513, A => n10413, ZN => 
                           n7014);
   U10540 : AOI21_X1 port map( B1 => n10412, B2 => n10840, A => n10411, ZN => 
                           n10413);
   U10541 : OAI22_X1 port map( A1 => n10512, A2 => n10410, B1 => n8433, B2 => 
                           n12092, ZN => n10411);
   U10542 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1455, B => n8093, ZN =>
                           n10410);
   U10543 : INV_X1 port map( A => n10408, ZN => n10512);
   U10544 : NAND4_X1 port map( A1 => n10407, A2 => n10406, A3 => n10405, A4 => 
                           n10404, ZN => n10412);
   U10545 : AOI22_X1 port map( A1 => n10427, A2 => n10476, B1 => n10510, B2 => 
                           n10440, ZN => n10404);
   U10546 : AOI22_X1 port map( A1 => n10403, A2 => n10495, B1 => n10498, B2 => 
                           n10439, ZN => n10405);
   U10547 : INV_X1 port map( A => n10481, ZN => n10403);
   U10548 : AOI22_X1 port map( A1 => n10428, A2 => n10499, B1 => n10478, B2 => 
                           n10493, ZN => n10406);
   U10549 : NAND4_X1 port map( A1 => n9539, A2 => n9538, A3 => n9537, A4 => 
                           n9536, ZN => n10478);
   U10550 : OR2_X1 port map( A1 => n10277, A2 => n10237, ZN => n9536);
   U10551 : NAND2_X1 port map( A1 => n9628, A2 => n10228, ZN => n9537);
   U10552 : AOI22_X1 port map( A1 => n9920, A2 => n8093, B1 => n9983, B2 => 
                           n10487, ZN => n9538);
   U10553 : AOI22_X1 port map( A1 => n9535, A2 => n10113, B1 => n10232, B2 => 
                           n9534, ZN => n9539);
   U10554 : OR2_X1 port map( A1 => n9954, A2 => n9339, ZN => n9534);
   U10555 : NOR2_X1 port map( A1 => n9411, A2 => n8550, ZN => n9339);
   U10556 : OR2_X1 port map( A1 => n10230, A2 => n10233, ZN => n9535);
   U10557 : AOI21_X1 port map( B1 => n10402, B2 => n10461, A => n10401, ZN => 
                           n10407);
   U10558 : OAI22_X1 port map( A1 => n10431, A2 => n10479, B1 => n10400, B2 => 
                           n10442, ZN => n10401);
   U10559 : INV_X1 port map( A => n10474, ZN => n10400);
   U10560 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_41_port, B2 =>
                           n8578, A => n10399, ZN => n10414);
   U10561 : OAI211_X1 port map( C1 => n10398, C2 => n10421, A => n10397, B => 
                           n10396, ZN => n10399);
   U10562 : XNOR2_X1 port map( A => n10394, B => n10393, ZN => n10398);
   U10563 : XNOR2_X1 port map( A => n10392, B => n10395, ZN => n10393);
   U10564 : AOI21_X1 port map( B1 => n10451, B2 => n10448, A => n10449, ZN => 
                           n10394);
   U10565 : AND2_X1 port map( A1 => C620_DATA2_11, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_11_port);
   U10566 : OAI222_X1 port map( A1 => n12093, A2 => n10437, B1 => n10482, B2 =>
                           n10436, C1 => n12092, C2 => n500, ZN => n7013);
   U10567 : NOR3_X1 port map( A1 => n10435, A2 => n10434, A3 => n10433, ZN => 
                           n10436);
   U10568 : OAI22_X1 port map( A1 => n10481, A2 => n10442, B1 => n10459, B2 => 
                           n10479, ZN => n10433);
   U10569 : OAI22_X1 port map( A1 => n10432, A2 => n10507, B1 => n10431, B2 => 
                           n10462, ZN => n10434);
   U10570 : INV_X1 port map( A => n10475, ZN => n10431);
   U10571 : OAI211_X1 port map( C1 => n10441, C2 => n10460, A => n10430, B => 
                           n10429, ZN => n10435);
   U10572 : AOI22_X1 port map( A1 => n10428, A2 => n10510, B1 => n10493, B2 => 
                           n10474, ZN => n10429);
   U10573 : NAND4_X1 port map( A1 => n9548, A2 => n9547, A3 => n9546, A4 => 
                           n9545, ZN => n10474);
   U10574 : NAND2_X1 port map( A1 => n9544, A2 => n10113, ZN => n9545);
   U10575 : OAI22_X1 port map( A1 => n10183, A2 => n12085, B1 => n10181, B2 => 
                           n10286, ZN => n9544);
   U10576 : NAND2_X1 port map( A1 => n9628, A2 => n9543, ZN => n9546);
   U10577 : INV_X1 port map( A => n10185, ZN => n9543);
   U10578 : AOI22_X1 port map( A1 => n9542, A2 => n10232, B1 => n9541, B2 => 
                           n10229, ZN => n9547);
   U10579 : INV_X1 port map( A => n9921, ZN => n9541);
   U10580 : OR2_X1 port map( A1 => n10193, A2 => n10277, ZN => n9548);
   U10581 : AOI22_X1 port map( A1 => n10427, A2 => n10461, B1 => n10498, B2 => 
                           n10440, ZN => n10430);
   U10582 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_42_port, B2 =>
                           n10492, A => n10426, ZN => n10437);
   U10583 : OAI21_X1 port map( B1 => n10422, B2 => n10421, A => n10420, ZN => 
                           n10424);
   U10584 : INV_X1 port map( A => n10418, ZN => n10422);
   U10585 : OAI21_X1 port map( B1 => n10418, B2 => n10421, A => n10417, ZN => 
                           n10425);
   U10586 : XNOR2_X1 port map( A => n10416, B => n10415, ZN => n10418);
   U10587 : AND2_X1 port map( A1 => C620_DATA2_12, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_12_port);
   U10588 : NOR2_X1 port map( A1 => n9581, A2 => n9580, ZN => n10481);
   U10589 : OAI22_X1 port map( A1 => n9579, A2 => n10164, B1 => n9578, B2 => 
                           n10284, ZN => n9580);
   U10590 : AOI21_X1 port map( B1 => n9366, B2 => n12086, A => n10161, ZN => 
                           n9578);
   U10591 : INV_X1 port map( A => n10160, ZN => n9366);
   U10592 : INV_X1 port map( A => n9628, ZN => n9579);
   U10593 : OAI211_X1 port map( C1 => n10159, C2 => n10277, A => n9577, B => 
                           n9576, ZN => n9581);
   U10594 : NAND2_X1 port map( A1 => n9575, A2 => n10232, ZN => n9576);
   U10595 : AOI22_X1 port map( A1 => n9920, A2 => n8090, B1 => n9983, B2 => 
                           n8016, ZN => n9577);
   U10596 : AND2_X1 port map( A1 => C620_DATA2_13, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_13_port);
   U10597 : OAI22_X1 port map( A1 => n10342, A2 => n12093, B1 => n502, B2 => 
                           n12092, ZN => n7011);
   U10598 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_44_port, B2 =>
                           n10492, A => n10341, ZN => n10342);
   U10599 : OAI211_X1 port map( C1 => n10340, C2 => n10345, A => n10339, B => 
                           n10338, ZN => n10341);
   U10600 : NAND2_X1 port map( A1 => n10346, A2 => n10340, ZN => n10338);
   U10601 : AOI211_X1 port map( C1 => n10337, C2 => n10336, A => n10335, B => 
                           n10334, ZN => n10339);
   U10602 : NOR2_X1 port map( A1 => n10333, A2 => n10452, ZN => n10334);
   U10603 : NOR3_X1 port map( A1 => n10332, A2 => n10331, A3 => n10330, ZN => 
                           n10333);
   U10604 : OAI22_X1 port map( A1 => n10375, A2 => n10388, B1 => n10459, B2 => 
                           n10442, ZN => n10330);
   U10605 : INV_X1 port map( A => n10439, ZN => n10459);
   U10606 : OAI22_X1 port map( A1 => n10432, A2 => n10460, B1 => n10371, B2 => 
                           n10507, ZN => n10331);
   U10607 : OAI211_X1 port map( C1 => n10441, C2 => n10376, A => n10329, B => 
                           n10328, ZN => n10332);
   U10608 : AOI22_X1 port map( A1 => n10428, A2 => n10502, B1 => n10493, B2 => 
                           n10475, ZN => n10328);
   U10609 : NAND4_X1 port map( A1 => n9617, A2 => n9616, A3 => n9615, A4 => 
                           n9614, ZN => n10475);
   U10610 : NAND2_X1 port map( A1 => n9628, A2 => n10111, ZN => n9614);
   U10611 : OAI21_X1 port map( B1 => n10110, B2 => n10112, A => n7785, ZN => 
                           n9615);
   U10612 : AOI22_X1 port map( A1 => n9613, A2 => n9612, B1 => n10229, B2 => 
                           n10116, ZN => n9616);
   U10613 : INV_X1 port map( A => n10109, ZN => n9612);
   U10614 : NOR2_X1 port map( A1 => n10284, A2 => n12085, ZN => n9613);
   U10615 : AOI22_X1 port map( A1 => n10288, A2 => n9845, B1 => n10232, B2 => 
                           n9609, ZN => n9617);
   U10616 : OR2_X1 port map( A1 => n9414, A2 => n10112, ZN => n9609);
   U10617 : NOR2_X1 port map( A1 => n9411, A2 => n7795, ZN => n9414);
   U10618 : AOI22_X1 port map( A1 => n10387, A2 => n10461, B1 => n10495, B2 => 
                           n10440, ZN => n10329);
   U10619 : NOR2_X1 port map( A1 => n10327, A2 => n10337, ZN => n10335);
   U10620 : NOR2_X1 port map( A1 => n10343, A2 => n10350, ZN => n10340);
   U10621 : OAI21_X1 port map( B1 => n210, B2 => n10832, A => n10807, ZN => n48
                           );
   U10622 : NAND2_X1 port map( A1 => n8579, A2 => IRAM_DATA(0), ZN => n10807);
   U10623 : OAI21_X1 port map( B1 => n10832, B2 => n8428, A => n10805, ZN => 
                           n50);
   U10624 : NAND2_X1 port map( A1 => n8579, A2 => IRAM_DATA(2), ZN => n10805);
   U10625 : OAI21_X1 port map( B1 => n195, B2 => n10832, A => n10810, ZN => 
                           n7121);
   U10626 : NAND2_X1 port map( A1 => n8579, A2 => IRAM_DATA(14), ZN => n10810);
   U10627 : OAI21_X1 port map( B1 => n196, B2 => n10832, A => n10798, ZN => n57
                           );
   U10628 : NAND2_X1 port map( A1 => n8579, A2 => IRAM_DATA(12), ZN => n10798);
   U10629 : OAI21_X1 port map( B1 => n10832, B2 => n185, A => n10820, ZN => 
                           n7111);
   U10630 : NAND2_X1 port map( A1 => n8579, A2 => IRAM_DATA(24), ZN => n10820);
   U10631 : OAI211_X1 port map( C1 => n10367, C2 => n10513, A => n10366, B => 
                           n10365, ZN => n7010);
   U10632 : NAND2_X1 port map( A1 => n10364, A2 => n10840, ZN => n10365);
   U10633 : NAND4_X1 port map( A1 => n10363, A2 => n10362, A3 => n10361, A4 => 
                           n10360, ZN => n10364);
   U10634 : AOI21_X1 port map( B1 => n10402, B2 => n10502, A => n10359, ZN => 
                           n10360);
   U10635 : OAI22_X1 port map( A1 => n10443, A2 => n10462, B1 => n10371, B2 => 
                           n10505, ZN => n10359);
   U10636 : AOI22_X1 port map( A1 => n10427, A2 => n10498, B1 => n10476, B2 => 
                           n10358, ZN => n10361);
   U10637 : AOI22_X1 port map( A1 => n10389, A2 => n10510, B1 => n10493, B2 => 
                           n10439, ZN => n10362);
   U10638 : NAND4_X1 port map( A1 => n9624, A2 => n9623, A3 => n9622, A4 => 
                           n9621, ZN => n10439);
   U10639 : OAI21_X1 port map( B1 => n10090, B2 => n10087, A => n7785, ZN => 
                           n9621);
   U10640 : AOI22_X1 port map( A1 => n10232, A2 => n9620, B1 => n10091, B2 => 
                           n10229, ZN => n9622);
   U10641 : OR2_X1 port map( A1 => n9402, A2 => n10087, ZN => n9620);
   U10642 : NOR2_X1 port map( A1 => n9411, A2 => n8556, ZN => n9402);
   U10643 : NAND2_X1 port map( A1 => n9628, A2 => n10089, ZN => n9623);
   U10644 : OAI21_X1 port map( B1 => n10085, B2 => n9618, A => n10113, ZN => 
                           n9624);
   U10645 : INV_X1 port map( A => n10088, ZN => n9618);
   U10646 : AOI22_X1 port map( A1 => n10387, A2 => n10499, B1 => n10503, B2 => 
                           n10440, ZN => n10363);
   U10647 : AOI22_X1 port map( A1 => n10408, A2 => n10357, B1 => n7764, B2 => 
                           DRAM_ADDRESS_13_port, ZN => n10366);
   U10648 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1251, B => n8555, ZN =>
                           n10357);
   U10649 : AOI211_X1 port map( C1 => DataPath_ALUhw_i_Q_EXTENDED_45_port, C2 
                           => n8578, A => n10356, B => n10355, ZN => n10367);
   U10650 : OAI211_X1 port map( C1 => n10381, C2 => n10354, A => n10353, B => 
                           n10352, ZN => n10355);
   U10651 : AOI21_X1 port map( B1 => n10350, B2 => n10349, A => n10348, ZN => 
                           n10354);
   U10652 : INV_X1 port map( A => n10347, ZN => n10348);
   U10653 : NOR2_X1 port map( A1 => n10345, A2 => n10344, ZN => n10356);
   U10654 : XNOR2_X1 port map( A => n10349, B => n10343, ZN => n10344);
   U10655 : INV_X1 port map( A => n10380, ZN => n10345);
   U10656 : AND2_X1 port map( A1 => C620_DATA2_14, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_14_port);
   U10657 : AOI22_X1 port map( A1 => n9105, A2 => n8399, B1 => n8997, B2 => 
                           n8304, ZN => n8710);
   U10658 : AOI22_X1 port map( A1 => n9105, A2 => n8305, B1 => n8997, B2 => 
                           n8391, ZN => n8709);
   U10659 : AOI22_X1 port map( A1 => n9105, A2 => n8395, B1 => n8997, B2 => 
                           n8302, ZN => n8706);
   U10660 : AOI22_X1 port map( A1 => n9105, A2 => n8397, B1 => n8997, B2 => 
                           IR_13_port, ZN => n8708);
   U10661 : AOI22_X1 port map( A1 => n9105, A2 => n8396, B1 => n8997, B2 => 
                           n8306, ZN => n8707);
   U10662 : OAI211_X1 port map( C1 => n10277, C2 => n10058, A => n9608, B => 
                           n9607, ZN => n10440);
   U10663 : AOI22_X1 port map( A1 => n10229, A2 => n9606, B1 => n10232, B2 => 
                           n9605, ZN => n9607);
   U10664 : OAI211_X1 port map( C1 => n8553, C2 => n9411, A => n9377, B => 
                           n9376, ZN => n9605);
   U10665 : NAND2_X1 port map( A1 => n9603, A2 => n12082, ZN => n9376);
   U10666 : INV_X1 port map( A => n9375, ZN => n9377);
   U10667 : INV_X1 port map( A => n9797, ZN => n9606);
   U10668 : AOI22_X1 port map( A1 => n9628, A2 => n9799, B1 => n9602, B2 => 
                           n10113, ZN => n9608);
   U10669 : OAI22_X1 port map( A1 => n10059, A2 => n12085, B1 => n12087, B2 => 
                           n9761, ZN => n9602);
   U10670 : INV_X1 port map( A => n10428, ZN => n10443);
   U10671 : INV_X1 port map( A => n10346, ZN => n10381);
   U10672 : AND2_X1 port map( A1 => C620_DATA2_15, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_15_port);
   U10673 : AOI22_X1 port map( A1 => n8580, A2 => IRAM_DATA(10), B1 => 
                           IR_10_port, B2 => n10808, ZN => n3009);
   U10674 : AOI22_X1 port map( A1 => n8580, A2 => IRAM_DATA(13), B1 => 
                           IR_13_port, B2 => n10808, ZN => n3006);
   U10675 : AOI22_X1 port map( A1 => n8580, A2 => IRAM_DATA(8), B1 => IR_8_port
                           , B2 => n10808, ZN => n3010);
   U10676 : AOI22_X1 port map( A1 => n8580, A2 => n12019, B1 => n8501, B2 => 
                           n10795, ZN => n7109);
   U10677 : INV_X1 port map( A => n10823, ZN => n10795);
   U10678 : NAND2_X1 port map( A1 => n8580, A2 => IRAM_DATA(27), ZN => n10822);
   U10679 : AOI22_X1 port map( A1 => n8580, A2 => n12021, B1 => n8308, B2 => 
                           n10808, ZN => n7105);
   U10680 : OAI21_X1 port map( B1 => n194, B2 => n10832, A => n10811, ZN => 
                           n7120);
   U10681 : NAND2_X1 port map( A1 => n8580, A2 => IRAM_DATA(15), ZN => n10811);
   U10682 : INV_X1 port map( A => n10803, ZN => n52);
   U10683 : AOI22_X1 port map( A1 => n8580, A2 => IRAM_DATA(4), B1 => IR_4_port
                           , B2 => n10808, ZN => n10803);
   U10684 : INV_X1 port map( A => n10806, ZN => n49);
   U10685 : AOI22_X1 port map( A1 => n8580, A2 => IRAM_DATA(1), B1 => IR_1_port
                           , B2 => n10808, ZN => n10806);
   U10686 : INV_X1 port map( A => n10809, ZN => n7122);
   U10687 : AOI22_X1 port map( A1 => n8580, A2 => IRAM_DATA(9), B1 => IR_9_port
                           , B2 => n10808, ZN => n10809);
   U10688 : INV_X1 port map( A => n10804, ZN => n51);
   U10689 : AOI22_X1 port map( A1 => n8580, A2 => IRAM_DATA(3), B1 => IR_3_port
                           , B2 => n10808, ZN => n10804);
   U10690 : INV_X1 port map( A => n10800, ZN => n55);
   U10691 : AOI22_X1 port map( A1 => n8580, A2 => IRAM_DATA(7), B1 => IR_7_port
                           , B2 => n10808, ZN => n10800);
   U10692 : INV_X1 port map( A => n10801, ZN => n54);
   U10693 : AOI22_X1 port map( A1 => n8580, A2 => IRAM_DATA(6), B1 => IR_6_port
                           , B2 => n10808, ZN => n10801);
   U10694 : INV_X1 port map( A => n10802, ZN => n53);
   U10695 : AOI22_X1 port map( A1 => n8580, A2 => IRAM_DATA(5), B1 => IR_5_port
                           , B2 => n10808, ZN => n10802);
   U10696 : OAI21_X1 port map( B1 => n10832, B2 => n186, A => n10819, ZN => 
                           n7112);
   U10697 : NAND2_X1 port map( A1 => n8580, A2 => IRAM_DATA(23), ZN => n10819);
   U10698 : OAI21_X1 port map( B1 => n10832, B2 => n192, A => n10813, ZN => 
                           n7118);
   U10699 : NAND2_X1 port map( A1 => n8580, A2 => IRAM_DATA(17), ZN => n10813);
   U10700 : OAI21_X1 port map( B1 => n10832, B2 => n191, A => n10814, ZN => 
                           n7117);
   U10701 : NAND2_X1 port map( A1 => n8580, A2 => IRAM_DATA(18), ZN => n10814);
   U10702 : OAI21_X1 port map( B1 => n10832, B2 => n190, A => n10815, ZN => 
                           n7116);
   U10703 : NAND2_X1 port map( A1 => n8580, A2 => IRAM_DATA(19), ZN => n10815);
   U10704 : OAI21_X1 port map( B1 => n10832, B2 => n189, A => n10816, ZN => 
                           n7115);
   U10705 : NAND2_X1 port map( A1 => n8580, A2 => IRAM_DATA(20), ZN => n10816);
   U10706 : OAI21_X1 port map( B1 => n10832, B2 => n187, A => n10818, ZN => 
                           n7113);
   U10707 : NAND2_X1 port map( A1 => n8580, A2 => IRAM_DATA(22), ZN => n10818);
   U10708 : OAI21_X1 port map( B1 => n10832, B2 => n193, A => n10812, ZN => 
                           n7119);
   U10709 : NAND2_X1 port map( A1 => n8580, A2 => IRAM_DATA(16), ZN => n10812);
   U10710 : OAI21_X1 port map( B1 => n10832, B2 => n188, A => n10817, ZN => 
                           n7114);
   U10711 : NAND2_X1 port map( A1 => n8580, A2 => IRAM_DATA(21), ZN => n10817);
   U10712 : OAI21_X1 port map( B1 => n197, B2 => n10832, A => n10799, ZN => n56
                           );
   U10713 : NAND2_X1 port map( A1 => n8580, A2 => IRAM_DATA(11), ZN => n10799);
   U10714 : OAI21_X1 port map( B1 => n10832, B2 => n184, A => n10821, ZN => 
                           n7110);
   U10715 : NAND2_X1 port map( A1 => n8580, A2 => IRAM_DATA(25), ZN => n10821);
   U10716 : OAI222_X1 port map( A1 => n12093, A2 => n10301, B1 => n10482, B2 =>
                           n10300, C1 => n12092, C2 => n504, ZN => n7008);
   U10717 : NOR3_X1 port map( A1 => n10299, A2 => n10298, A3 => n10297, ZN => 
                           n10300);
   U10718 : OAI22_X1 port map( A1 => n10375, A2 => n10462, B1 => n10374, B2 => 
                           n10460, ZN => n10297);
   U10719 : INV_X1 port map( A => n10358, ZN => n10374);
   U10720 : OAI22_X1 port map( A1 => n10432, A2 => n10479, B1 => n10371, B2 => 
                           n10388, ZN => n10298);
   U10721 : INV_X1 port map( A => n10389, ZN => n10432);
   U10722 : OAI211_X1 port map( C1 => n10441, C2 => n10442, A => n10296, B => 
                           n10295, ZN => n10299);
   U10723 : AOI22_X1 port map( A1 => n10428, A2 => n10493, B1 => n10476, B2 => 
                           n10294, ZN => n10295);
   U10724 : OAI21_X1 port map( B1 => n10028, B2 => n10027, A => n7785, ZN => 
                           n9631);
   U10725 : AOI22_X1 port map( A1 => n10232, A2 => n9630, B1 => n9743, B2 => 
                           n10229, ZN => n9632);
   U10726 : OR2_X1 port map( A1 => n9381, A2 => n10027, ZN => n9630);
   U10727 : NOR2_X1 port map( A1 => n9411, A2 => n10010, ZN => n9381);
   U10728 : OR2_X1 port map( A1 => n7800, A2 => n12074, ZN => n9411);
   U10729 : AOI22_X1 port map( A1 => n9628, A2 => n10026, B1 => n9627, B2 => 
                           n10022, ZN => n9633);
   U10730 : AOI21_X1 port map( B1 => n10115, B2 => n10024, A => n10284, ZN => 
                           n9627);
   U10731 : NOR2_X1 port map( A1 => n10184, A2 => n368, ZN => n9628);
   U10732 : AOI22_X1 port map( A1 => n10498, A2 => n10387, B1 => n10293, B2 => 
                           n10461, ZN => n10296);
   U10733 : INV_X1 port map( A => n10402, ZN => n10441);
   U10734 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_47_port, B2 =>
                           n8578, A => n10272, ZN => n10301);
   U10735 : OAI211_X1 port map( C1 => n10271, C2 => n10270, A => n10269, B => 
                           n10268, ZN => n10272);
   U10736 : INV_X1 port map( A => n10265, ZN => n10267);
   U10737 : AOI211_X1 port map( C1 => n10264, C2 => n10468, A => n10263, B => 
                           n10262, ZN => n10269);
   U10738 : NOR3_X1 port map( A1 => n10489, A2 => n8554, A3 => n7794, ZN => 
                           n10262);
   U10739 : INV_X1 port map( A => n10458, ZN => n10489);
   U10740 : NOR3_X1 port map( A1 => n10488, A2 => n10261, A3 => 
                           DP_OP_751_130_5637_n1149, ZN => n10263);
   U10741 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1149, B => n8554, ZN =>
                           n10264);
   U10742 : OAI21_X1 port map( B1 => n10369, B2 => n10370, A => n10258, ZN => 
                           n10259);
   U10743 : NAND2_X1 port map( A1 => n10258, A2 => n10257, ZN => n10370);
   U10744 : AOI21_X1 port map( B1 => n10256, B2 => n10255, A => n10254, ZN => 
                           n10369);
   U10745 : INV_X1 port map( A => n10253, ZN => n10254);
   U10746 : INV_X1 port map( A => n10343, ZN => n10256);
   U10747 : INV_X1 port map( A => n10266, ZN => n10260);
   U10748 : AND2_X1 port map( A1 => n10252, A2 => n10251, ZN => n10266);
   U10749 : AOI21_X1 port map( B1 => n10346, B2 => n10265, A => n10380, ZN => 
                           n10271);
   U10750 : NOR2_X1 port map( A1 => n10250, A2 => n10421, ZN => n10380);
   U10751 : INV_X1 port map( A => n10249, ZN => n10250);
   U10752 : NOR2_X1 port map( A1 => n10249, A2 => n10421, ZN => n10346);
   U10753 : OAI22_X1 port map( A1 => n10324, A2 => n12093, B1 => n505, B2 => 
                           n12092, ZN => n7007);
   U10754 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_48_port, B2 =>
                           n10492, A => n10323, ZN => n10324);
   U10755 : OAI211_X1 port map( C1 => n10322, C2 => n10321, A => n10320, B => 
                           n10319, ZN => n10323);
   U10756 : NAND2_X1 port map( A1 => n10318, A2 => n10321, ZN => n10319);
   U10757 : AOI21_X1 port map( B1 => n10317, B2 => n10390, A => n10316, ZN => 
                           n10320);
   U10758 : AOI22_X1 port map( A1 => n10308, A2 => n10476, B1 => n10358, B2 => 
                           n10510, ZN => n10309);
   U10759 : AOI22_X1 port map( A1 => n10427, A2 => n10503, B1 => n10389, B2 => 
                           n10495, ZN => n10310);
   U10760 : AOI211_X1 port map( C1 => n10493, C2 => n10402, A => n10307, B => 
                           n10306, ZN => n10311);
   U10761 : OAI22_X1 port map( A1 => n10373, A2 => n10479, B1 => n10372, B2 => 
                           n10460, ZN => n10306);
   U10762 : OAI22_X1 port map( A1 => n10371, A2 => n10376, B1 => n10305, B2 => 
                           n10505, ZN => n10307);
   U10763 : OAI211_X1 port map( C1 => n10292, C2 => n10291, A => n10290, B => 
                           n10289, ZN => n10402);
   U10764 : OAI22_X1 port map( A1 => n10288, A2 => n10287, B1 => n10286, B2 => 
                           n10285, ZN => n10289);
   U10765 : NOR2_X1 port map( A1 => n10284, A2 => n10283, ZN => n10287);
   U10766 : AOI211_X1 port map( C1 => n10282, C2 => n10281, A => n10280, B => 
                           n10279, ZN => n10290);
   U10767 : NOR2_X1 port map( A1 => n10278, A2 => n10277, ZN => n10279);
   U10768 : INV_X1 port map( A => n10276, ZN => n10278);
   U10769 : OAI22_X1 port map( A1 => n10180, A2 => n10275, B1 => n10274, B2 => 
                           n8094, ZN => n10280);
   U10770 : INV_X1 port map( A => n9987, ZN => n10274);
   U10771 : NOR2_X1 port map( A1 => n10304, A2 => n10303, ZN => n10321);
   U10772 : INV_X1 port map( A => n10302, ZN => n10322);
   U10773 : OAI211_X1 port map( C1 => n10247, C2 => n10513, A => n10246, B => 
                           n10245, ZN => n7006);
   U10774 : NAND2_X1 port map( A1 => n10244, A2 => n10840, ZN => n10245);
   U10775 : AOI22_X1 port map( A1 => n10308, A2 => n10461, B1 => n10358, B2 => 
                           n10498, ZN => n10241);
   U10776 : AOI22_X1 port map( A1 => n10427, A2 => n10493, B1 => n10389, B2 => 
                           n10503, ZN => n10242);
   U10777 : INV_X1 port map( A => n10375, ZN => n10427);
   U10778 : AOI21_X1 port map( B1 => n7785, B2 => n10239, A => n10238, ZN => 
                           n10375);
   U10779 : OAI211_X1 port map( C1 => n10237, C2 => n10284, A => n10236, B => 
                           n10235, ZN => n10238);
   U10780 : OAI21_X1 port map( B1 => n10234, B2 => n10233, A => n10232, ZN => 
                           n10235);
   U10781 : NOR2_X1 port map( A1 => n9951, A2 => n12074, ZN => n10233);
   U10782 : AOI22_X1 port map( A1 => n10231, A2 => n10230, B1 => n10229, B2 => 
                           n10228, ZN => n10236);
   U10783 : AND2_X1 port map( A1 => n9730, A2 => n12086, ZN => n10230);
   U10784 : AOI21_X1 port map( B1 => n10115, B2 => n9953, A => n9954, ZN => 
                           n10237);
   U10785 : AOI211_X1 port map( C1 => n10476, C2 => n10227, A => n10226, B => 
                           n10225, ZN => n10243);
   U10786 : OAI22_X1 port map( A1 => n10373, A2 => n10462, B1 => n10372, B2 => 
                           n10388, ZN => n10225);
   U10787 : OAI22_X1 port map( A1 => n10371, A2 => n10479, B1 => n10305, B2 => 
                           n10460, ZN => n10226);
   U10788 : AOI22_X1 port map( A1 => n10408, A2 => n10224, B1 => n7764, B2 => 
                           DRAM_ADDRESS_17_port, ZN => n10246);
   U10789 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1047, B => n8550, ZN =>
                           n10224);
   U10790 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_49_port, B2 =>
                           n10492, A => n10222, ZN => n10247);
   U10791 : NAND4_X1 port map( A1 => n10221, A2 => n10220, A3 => n10219, A4 => 
                           n10218, ZN => n10222);
   U10792 : OAI211_X1 port map( C1 => n10304, C2 => n10216, A => n10318, B => 
                           n10215, ZN => n10220);
   U10793 : NAND2_X1 port map( A1 => n10302, A2 => n10214, ZN => n10221);
   U10794 : OAI21_X1 port map( B1 => n10303, B2 => n10216, A => n10213, ZN => 
                           n10214);
   U10795 : OAI222_X1 port map( A1 => n10691, A2 => n7759, B1 => n8549, B2 => 
                           n9045, C1 => n8326, C2 => n10702, ZN => n7056);
   U10796 : XNOR2_X1 port map( A => n10690, B => n10689, ZN => n10691);
   U10797 : NOR2_X1 port map( A1 => n10688, A2 => n10687, ZN => n10689);
   U10798 : INV_X1 port map( A => n10686, ZN => n10688);
   U10799 : OAI222_X1 port map( A1 => n7759, A2 => n10697, B1 => n10702, B2 => 
                           intadd_1_A_1_port, C1 => n8549, C2 => n9029, ZN => 
                           n7057);
   U10800 : NAND2_X1 port map( A1 => n10694, A2 => n10693, ZN => n10696);
   U10801 : INV_X1 port map( A => n10692, ZN => n10694);
   U10802 : OAI222_X1 port map( A1 => n7759, A2 => n10703, B1 => n10702, B2 => 
                           intadd_1_A_0_port, C1 => n8549, C2 => n12060, ZN => 
                           n7058);
   U10803 : NAND2_X1 port map( A1 => n10698, A2 => n10699, ZN => n10701);
   U10804 : OAI222_X1 port map( A1 => n10685, A2 => n7759, B1 => n8549, B2 => 
                           n9047, C1 => n8325, C2 => n10702, ZN => n7055);
   U10805 : XNOR2_X1 port map( A => n10684, B => n10683, ZN => n10685);
   U10806 : NAND2_X1 port map( A1 => n10682, A2 => n10681, ZN => n10683);
   U10807 : INV_X1 port map( A => n10680, ZN => n10682);
   U10808 : OAI222_X1 port map( A1 => n10679, A2 => n7759, B1 => n10702, B2 => 
                           n226, C1 => n8549, C2 => n10678, ZN => n7054);
   U10809 : NAND2_X1 port map( A1 => n10675, A2 => n10674, ZN => n10677);
   U10810 : OAI21_X1 port map( B1 => n10673, B2 => n7759, A => n10672, ZN => 
                           n7053);
   U10811 : AOI22_X1 port map( A1 => n12070, A2 => i_RD1_6_port, B1 => 
                           IRAM_ADDRESS_6_port, B2 => n10835, ZN => n10672);
   U10812 : XNOR2_X1 port map( A => n8031, B => n10670, ZN => n10673);
   U10813 : NOR2_X1 port map( A1 => n7777, A2 => n10669, ZN => n10670);
   U10814 : OAI21_X1 port map( B1 => n9240, B2 => n8549, A => n10706, ZN => 
                           n7059);
   U10815 : NAND2_X1 port map( A1 => n10705, A2 => n8549, ZN => n10706);
   U10816 : OAI21_X1 port map( B1 => n10667, B2 => n7759, A => n10666, ZN => 
                           n7052);
   U10817 : AOI22_X1 port map( A1 => n12070, A2 => i_RD1_7_port, B1 => 
                           IRAM_ADDRESS_7_port, B2 => n10835, ZN => n10666);
   U10818 : XNOR2_X1 port map( A => n10664, B => IRAM_ADDRESS_7_port, ZN => 
                           n10665);
   U10819 : OAI22_X1 port map( A1 => n10211, A2 => n12093, B1 => n506, B2 => 
                           n12092, ZN => n7005);
   U10820 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_50_port, B2 =>
                           n10492, A => n10210, ZN => n10211);
   U10821 : NAND4_X1 port map( A1 => n10209, A2 => n10208, A3 => n10207, A4 => 
                           n10206, ZN => n10210);
   U10822 : AOI21_X1 port map( B1 => n10202, B2 => n10390, A => n10201, ZN => 
                           n10208);
   U10823 : AOI22_X1 port map( A1 => n10293, A2 => n10498, B1 => n10499, B2 => 
                           n10308, ZN => n10194);
   U10824 : AOI22_X1 port map( A1 => n10389, A2 => n10493, B1 => n10502, B2 => 
                           n10358, ZN => n10195);
   U10825 : OAI211_X1 port map( C1 => n10193, C2 => n10284, A => n10192, B => 
                           n10191, ZN => n10389);
   U10826 : NAND2_X1 port map( A1 => n10190, A2 => n7785, ZN => n10191);
   U10827 : AOI211_X1 port map( C1 => n10189, C2 => n10188, A => n10187, B => 
                           n10186, ZN => n10192);
   U10828 : NOR2_X1 port map( A1 => n8094, A2 => n10185, ZN => n10186);
   U10829 : NOR3_X1 port map( A1 => n10184, A2 => n12085, A3 => n10183, ZN => 
                           n10187);
   U10830 : OAI21_X1 port map( B1 => n10182, B2 => n10181, A => n10180, ZN => 
                           n10189);
   U10831 : AOI21_X1 port map( B1 => n10115, B2 => n9917, A => n9918, ZN => 
                           n10193);
   U10832 : AOI211_X1 port map( C1 => n10461, C2 => n10227, A => n10179, B => 
                           n10178, ZN => n10196);
   U10833 : OAI22_X1 port map( A1 => n10373, A2 => n10442, B1 => n10177, B2 => 
                           n10507, ZN => n10178);
   U10834 : OAI22_X1 port map( A1 => n10371, A2 => n10462, B1 => n10305, B2 => 
                           n10388, ZN => n10179);
   U10835 : OAI211_X1 port map( C1 => n10205, C2 => n10176, A => n10302, B => 
                           n10175, ZN => n10209);
   U10836 : INV_X1 port map( A => n10174, ZN => n10176);
   U10837 : AOI22_X1 port map( A1 => n9294, A2 => n8303, B1 => 
                           IRAM_ADDRESS_8_port, B2 => n10835, ZN => n12061);
   U10838 : XNOR2_X1 port map( A => n9295, B => IRAM_ADDRESS_8_port, ZN => 
                           n9293);
   U10839 : OAI222_X1 port map( A1 => n12093, A2 => n10172, B1 => n10482, B2 =>
                           n10171, C1 => n12092, C2 => n507, ZN => n7004);
   U10840 : AND3_X1 port map( A1 => n10170, A2 => n10169, A3 => n10168, ZN => 
                           n10171);
   U10841 : AOI22_X1 port map( A1 => n10493, A2 => n10387, B1 => n10293, B2 => 
                           n10502, ZN => n10168);
   U10842 : INV_X1 port map( A => n10373, ZN => n10387);
   U10843 : AOI211_X1 port map( C1 => n7785, C2 => n10167, A => n10166, B => 
                           n10165, ZN => n10373);
   U10844 : OAI21_X1 port map( B1 => n10164, B2 => n8094, A => n10163, ZN => 
                           n10165);
   U10845 : OAI21_X1 port map( B1 => n10162, B2 => n10161, A => n10232, ZN => 
                           n10163);
   U10846 : AND2_X1 port map( A1 => n9886, A2 => n10870, ZN => n10161);
   U10847 : OAI22_X1 port map( A1 => n10292, A2 => n10160, B1 => n10159, B2 => 
                           n10284, ZN => n10166);
   U10848 : AOI21_X1 port map( B1 => n10115, B2 => n9885, A => n9574, ZN => 
                           n10159);
   U10849 : INV_X1 port map( A => n9889, ZN => n9574);
   U10850 : AOI22_X1 port map( A1 => n10308, A2 => n10510, B1 => n10358, B2 => 
                           n10495, ZN => n10169);
   U10851 : AOI211_X1 port map( C1 => n10461, C2 => n10158, A => n10157, B => 
                           n10156, ZN => n10170);
   U10852 : OAI22_X1 port map( A1 => n10155, A2 => n10507, B1 => n10154, B2 => 
                           n10460, ZN => n10156);
   U10853 : OAI22_X1 port map( A1 => n10371, A2 => n10442, B1 => n10305, B2 => 
                           n10376, ZN => n10157);
   U10854 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_51_port, B2 =>
                           n10492, A => n10153, ZN => n10172);
   U10855 : OAI21_X1 port map( B1 => n10152, B2 => n10151, A => n10150, ZN => 
                           n10153);
   U10856 : AOI21_X1 port map( B1 => n10302, B2 => n10149, A => n10148, ZN => 
                           n10150);
   U10857 : OAI211_X1 port map( C1 => n10147, C2 => n10465, A => n10146, B => 
                           n10145, ZN => n10148);
   U10858 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n945, B => n8552, ZN => 
                           n10147);
   U10859 : XNOR2_X1 port map( A => n10142, B => n10141, ZN => n10149);
   U10860 : NOR2_X1 port map( A1 => n10140, A2 => n10421, ZN => n10302);
   U10861 : INV_X1 port map( A => n10139, ZN => n10140);
   U10862 : INV_X1 port map( A => n10318, ZN => n10151);
   U10863 : NOR2_X1 port map( A1 => n10139, A2 => n10421, ZN => n10318);
   U10864 : NAND2_X1 port map( A1 => n10137, A2 => n10136, ZN => n10141);
   U10865 : AOI22_X1 port map( A1 => n12070, A2 => i_RD1_9_port, B1 => n10835, 
                           B2 => IRAM_ADDRESS_9_port, ZN => n12063);
   U10866 : XNOR2_X1 port map( A => n8034, B => n9300, ZN => n12064);
   U10867 : NOR2_X1 port map( A1 => n7776, A2 => n9304, ZN => n9300);
   U10868 : AND2_X1 port map( A1 => C620_DATA2_20, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_20_port);
   U10869 : OAI22_X1 port map( A1 => n10134, A2 => n12093, B1 => n508, B2 => 
                           n12092, ZN => n7003);
   U10870 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_52_port, B2 =>
                           n10492, A => n10133, ZN => n10134);
   U10871 : OAI211_X1 port map( C1 => n10132, C2 => n10131, A => n10130, B => 
                           n10129, ZN => n10133);
   U10872 : AOI21_X1 port map( B1 => n10128, B2 => n10390, A => n10127, ZN => 
                           n10129);
   U10873 : INV_X1 port map( A => n10452, ZN => n10390);
   U10874 : NAND4_X1 port map( A1 => n10121, A2 => n10120, A3 => n10119, A4 => 
                           n10118, ZN => n10128);
   U10875 : AOI21_X1 port map( B1 => n10499, B2 => n10158, A => n10117, ZN => 
                           n10118);
   U10876 : OAI22_X1 port map( A1 => n10371, A2 => n10444, B1 => n10305, B2 => 
                           n10479, ZN => n10117);
   U10877 : INV_X1 port map( A => n10294, ZN => n10305);
   U10878 : AOI22_X1 port map( A1 => n10293, A2 => n10495, B1 => n10476, B2 => 
                           n10107, ZN => n10119);
   U10879 : AOI22_X1 port map( A1 => n10308, A2 => n10498, B1 => n10358, B2 => 
                           n10503, ZN => n10120);
   U10880 : AOI22_X1 port map( A1 => n10106, A2 => n10461, B1 => n10510, B2 => 
                           n10227, ZN => n10121);
   U10881 : NAND2_X1 port map( A1 => n10105, A2 => n10132, ZN => n10130);
   U10882 : AND2_X1 port map( A1 => n10104, A2 => n10103, ZN => n10132);
   U10883 : OAI222_X1 port map( A1 => n10663, A2 => n7759, B1 => n8549, B2 => 
                           n9077, C1 => n8429, C2 => n10702, ZN => n7049);
   U10884 : XNOR2_X1 port map( A => n10661, B => IRAM_ADDRESS_10_port, ZN => 
                           n10662);
   U10885 : OAI222_X1 port map( A1 => n8549, A2 => n10660, B1 => n7759, B2 => 
                           n10659, C1 => n8383, C2 => n10702, ZN => n7048);
   U10886 : XNOR2_X1 port map( A => n10656, B => IRAM_ADDRESS_11_port, ZN => 
                           n10657);
   U10887 : INV_X1 port map( A => i_RD1_11_port, ZN => n10660);
   U10888 : AND2_X1 port map( A1 => C620_DATA2_21, A2 => n10730, ZN => 
                           DRAMRF_ADDRESS_21_port);
   U10889 : OAI211_X1 port map( C1 => n10101, C2 => n10513, A => n10100, B => 
                           n10099, ZN => n7002);
   U10890 : OAI21_X1 port map( B1 => n10098, B2 => n10097, A => n10840, ZN => 
                           n10099);
   U10891 : NAND2_X1 port map( A1 => n10096, A2 => n10095, ZN => n10097);
   U10892 : AOI22_X1 port map( A1 => n10107, A2 => n10461, B1 => n10476, B2 => 
                           n10094, ZN => n10095);
   U10893 : AOI22_X1 port map( A1 => n10293, A2 => n10503, B1 => n10502, B2 => 
                           n10308, ZN => n10096);
   U10894 : INV_X1 port map( A => n10372, ZN => n10293);
   U10895 : OAI211_X1 port map( C1 => n10154, C2 => n10376, A => n10093, B => 
                           n10092, ZN => n10098);
   U10896 : AOI22_X1 port map( A1 => n10358, A2 => n10493, B1 => n10294, B2 => 
                           n10495, ZN => n10092);
   U10897 : NAND2_X1 port map( A1 => n9816, A2 => n10115, ZN => n10088);
   U10898 : NOR2_X1 port map( A1 => n9747, A2 => n12085, ZN => n10085);
   U10899 : AOI22_X1 port map( A1 => n10106, A2 => n10499, B1 => n10510, B2 => 
                           n10158, ZN => n10093);
   U10900 : INV_X1 port map( A => n10227, ZN => n10154);
   U10901 : AOI22_X1 port map( A1 => n10408, A2 => n10083, B1 => n7764, B2 => 
                           DRAM_ADDRESS_21_port, ZN => n10100);
   U10902 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n843, B => n8556, ZN => 
                           n10083);
   U10903 : AOI211_X1 port map( C1 => DataPath_ALUhw_i_Q_EXTENDED_53_port, C2 
                           => n8578, A => n10081, B => n10080, ZN => n10101);
   U10904 : OAI211_X1 port map( C1 => n10131, C2 => n10079, A => n10078, B => 
                           n10077, ZN => n10080);
   U10905 : INV_X1 port map( A => DP_OP_751_130_5637_n843, ZN => n10076);
   U10906 : AOI21_X1 port map( B1 => n10075, B2 => n10104, A => n10074, ZN => 
                           n10079);
   U10907 : INV_X1 port map( A => n10073, ZN => n10074);
   U10908 : NOR2_X1 port map( A1 => n10072, A2 => n10071, ZN => n10081);
   U10909 : XNOR2_X1 port map( A => n10075, B => n10103, ZN => n10071);
   U10910 : INV_X1 port map( A => n10105, ZN => n10072);
   U10911 : OAI222_X1 port map( A1 => n10655, A2 => n7759, B1 => n10702, B2 => 
                           n222, C1 => n8549, C2 => n10654, ZN => n7047);
   U10912 : INV_X1 port map( A => i_RD1_12_port, ZN => n10654);
   U10913 : XNOR2_X1 port map( A => n10651, B => n222, ZN => n10652);
   U10914 : OAI222_X1 port map( A1 => n12093, A2 => n10069, B1 => n10482, B2 =>
                           n10068, C1 => n12092, C2 => n509, ZN => n7001);
   U10915 : NOR3_X1 port map( A1 => n10067, A2 => n10066, A3 => n10065, ZN => 
                           n10068);
   U10916 : OAI22_X1 port map( A1 => n10064, A2 => n10460, B1 => n10177, B2 => 
                           n10376, ZN => n10065);
   U10917 : OAI22_X1 port map( A1 => n10372, A2 => n10444, B1 => n10063, B2 => 
                           n10505, ZN => n10066);
   U10918 : AOI211_X1 port map( C1 => n7785, C2 => n10062, A => n10061, B => 
                           n10060, ZN => n10372);
   U10919 : OAI22_X1 port map( A1 => n10292, A2 => n10059, B1 => n10284, B2 => 
                           n10058, ZN => n10060);
   U10920 : INV_X1 port map( A => n9796, ZN => n10058);
   U10921 : NAND2_X1 port map( A1 => n10231, A2 => n12086, ZN => n10292);
   U10922 : OAI21_X1 port map( B1 => n10057, B2 => n8094, A => n10056, ZN => 
                           n10061);
   U10923 : OAI211_X1 port map( C1 => n12087, C2 => n7792, A => n10055, B => 
                           n10232, ZN => n10056);
   U10924 : INV_X1 port map( A => n9799, ZN => n10057);
   U10925 : OAI211_X1 port map( C1 => n8311, C2 => n10507, A => n10054, B => 
                           n10053, ZN => n10067);
   U10926 : AOI22_X1 port map( A1 => n10308, A2 => n10495, B1 => n10294, B2 => 
                           n10503, ZN => n10053);
   U10927 : AOI22_X1 port map( A1 => n10106, A2 => n10510, B1 => n10502, B2 => 
                           n10227, ZN => n10054);
   U10928 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_54_port, B2 =>
                           n10492, A => n10052, ZN => n10069);
   U10929 : OAI211_X1 port map( C1 => n10051, C2 => n10131, A => n10050, B => 
                           n10049, ZN => n10052);
   U10930 : AOI21_X1 port map( B1 => n10458, B2 => n7769, A => n10045, ZN => 
                           n10047);
   U10931 : NOR2_X1 port map( A1 => n10465, A2 => n7769, ZN => n10045);
   U10932 : NAND2_X1 port map( A1 => n10105, A2 => n10043, ZN => n10050);
   U10933 : OAI21_X1 port map( B1 => n10042, B2 => n10041, A => n10040, ZN => 
                           n10043);
   U10934 : XNOR2_X1 port map( A => n10039, B => n10038, ZN => n10051);
   U10935 : OAI222_X1 port map( A1 => n12093, A2 => n10036, B1 => n10482, B2 =>
                           n10035, C1 => n12092, C2 => n510, ZN => n7000);
   U10936 : NOR3_X1 port map( A1 => n10034, A2 => n10033, A3 => n10032, ZN => 
                           n10035);
   U10937 : OAI22_X1 port map( A1 => n10063, A2 => n10460, B1 => n10177, B2 => 
                           n10479, ZN => n10032);
   U10938 : OAI22_X1 port map( A1 => n10031, A2 => n10507, B1 => n10064, B2 => 
                           n10388, ZN => n10033);
   U10939 : OAI211_X1 port map( C1 => n8311, C2 => n10505, A => n10030, B => 
                           n10029, ZN => n10034);
   U10940 : AOI22_X1 port map( A1 => n10308, A2 => n10503, B1 => n10294, B2 => 
                           n10493, ZN => n10029);
   U10941 : OAI21_X1 port map( B1 => n9779, B2 => n368, A => n10286, ZN => 
                           n10022);
   U10942 : INV_X1 port map( A => n10021, ZN => n10084);
   U10943 : AOI22_X1 port map( A1 => n10106, A2 => n10498, B1 => n10495, B2 => 
                           n10227, ZN => n10030);
   U10944 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_55_port, B2 =>
                           n10492, A => n10020, ZN => n10036);
   U10945 : OAI21_X1 port map( B1 => n10019, B2 => n10131, A => n10018, ZN => 
                           n10020);
   U10946 : AOI21_X1 port map( B1 => n10105, B2 => n10017, A => n10016, ZN => 
                           n10018);
   U10947 : OAI211_X1 port map( C1 => n10015, C2 => n10465, A => n10014, B => 
                           n10013, ZN => n10016);
   U10948 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n741, B => n10012, ZN =>
                           n10015);
   U10949 : XNOR2_X1 port map( A => n10009, B => n10008, ZN => n10017);
   U10950 : NAND2_X1 port map( A1 => n10007, A2 => n10040, ZN => n10009);
   U10951 : NAND2_X1 port map( A1 => n10041, A2 => n10042, ZN => n10040);
   U10952 : NAND2_X1 port map( A1 => n10006, A2 => n10005, ZN => n10042);
   U10953 : INV_X1 port map( A => n10038, ZN => n10041);
   U10954 : NOR2_X1 port map( A1 => n10004, A2 => n10421, ZN => n10105);
   U10955 : NAND2_X1 port map( A1 => n10004, A2 => n10450, ZN => n10131);
   U10956 : XNOR2_X1 port map( A => n10007, B => n10008, ZN => n10019);
   U10957 : NOR2_X1 port map( A1 => n10003, A2 => n10002, ZN => n10008);
   U10958 : INV_X1 port map( A => n10001, ZN => n10003);
   U10959 : OAI222_X1 port map( A1 => n8549, A2 => n10647, B1 => n7759, B2 => 
                           n10646, C1 => n8384, C2 => n10702, ZN => n7045);
   U10960 : XNOR2_X1 port map( A => n10645, B => n10644, ZN => n10646);
   U10961 : NOR2_X1 port map( A1 => n7760, A2 => n10643, ZN => n10644);
   U10962 : OAI222_X1 port map( A1 => n12093, A2 => n9999, B1 => n10482, B2 => 
                           n9998, C1 => n12092, C2 => n511, ZN => n6999);
   U10963 : NOR3_X1 port map( A1 => n9997, A2 => n9996, A3 => n9995, ZN => 
                           n9998);
   U10964 : OAI22_X1 port map( A1 => n10155, A2 => n10479, B1 => n10177, B2 => 
                           n10462, ZN => n9995);
   U10965 : OAI22_X1 port map( A1 => n10063, A2 => n10388, B1 => n10064, B2 => 
                           n10376, ZN => n9996);
   U10966 : OAI211_X1 port map( C1 => n8311, C2 => n10460, A => n9994, B => 
                           n9993, ZN => n9997);
   U10967 : AOI22_X1 port map( A1 => n10461, A2 => n9992, B1 => n10308, B2 => 
                           n10493, ZN => n9993);
   U10968 : NAND4_X1 port map( A1 => n9991, A2 => n9990, A3 => n9989, A4 => 
                           n9988, ZN => n10308);
   U10969 : NAND2_X1 port map( A1 => n10276, A2 => n10288, ZN => n9988);
   U10970 : OAI211_X1 port map( C1 => n10115, C2 => n9987, A => n10232, B => 
                           n9986, ZN => n9989);
   U10971 : OR2_X1 port map( A1 => n10285, A2 => n12087, ZN => n9986);
   U10972 : AOI22_X1 port map( A1 => n9985, A2 => n9984, B1 => n7772, B2 => 
                           n9983, ZN => n9990);
   U10973 : INV_X1 port map( A => n10275, ZN => n9984);
   U10974 : NOR2_X1 port map( A1 => n9982, A2 => n9981, ZN => n9991);
   U10975 : OAI22_X1 port map( A1 => n9980, A2 => n9979, B1 => n10184, B2 => 
                           n10283, ZN => n9981);
   U10976 : AOI22_X1 port map( A1 => n9533, A2 => n12082, B1 => n10281, B2 => 
                           n12071, ZN => n10283);
   U10977 : AND2_X1 port map( A1 => n9978, A2 => n7785, ZN => n9982);
   U10978 : AOI22_X1 port map( A1 => n9977, A2 => n10476, B1 => n10503, B2 => 
                           n10227, ZN => n9994);
   U10979 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_56_port, B2 =>
                           n8578, A => n9976, ZN => n9999);
   U10980 : OAI211_X1 port map( C1 => n9975, C2 => n9974, A => n9973, B => 
                           n9972, ZN => n9976);
   U10981 : AOI21_X1 port map( B1 => n10458, B2 => n10281, A => n9968, ZN => 
                           n9970);
   U10982 : NOR2_X1 port map( A1 => n10465, A2 => n10281, ZN => n9968);
   U10983 : NAND2_X1 port map( A1 => n9967, A2 => n9975, ZN => n9973);
   U10984 : NOR2_X1 port map( A1 => n9966, A2 => n9965, ZN => n9975);
   U10985 : INV_X1 port map( A => n9964, ZN => n9966);
   U10986 : OAI211_X1 port map( C1 => n9962, C2 => n10513, A => n9961, B => 
                           n9960, ZN => n6998);
   U10987 : NAND2_X1 port map( A1 => n9959, A2 => n10840, ZN => n9960);
   U10988 : AOI22_X1 port map( A1 => n10106, A2 => n10495, B1 => n10493, B2 => 
                           n10227, ZN => n9956);
   U10989 : INV_X1 port map( A => n10228, ZN => n9952);
   U10990 : INV_X1 port map( A => n10155, ZN => n10106);
   U10991 : AOI22_X1 port map( A1 => n10094, A2 => n10498, B1 => n10158, B2 => 
                           n10503, ZN => n9957);
   U10992 : AOI211_X1 port map( C1 => n10476, C2 => n9949, A => n9948, B => 
                           n9947, ZN => n9958);
   U10993 : OAI22_X1 port map( A1 => n9946, A2 => n10505, B1 => n8311, B2 => 
                           n10388, ZN => n9947);
   U10994 : OAI22_X1 port map( A1 => n10031, A2 => n10460, B1 => n10064, B2 => 
                           n10479, ZN => n9948);
   U10995 : AOI22_X1 port map( A1 => n10408, A2 => n9945, B1 => n7764, B2 => 
                           DRAM_ADDRESS_25_port, ZN => n9961);
   U10996 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n639, B => n9944, ZN => 
                           n9945);
   U10997 : AOI211_X1 port map( C1 => DataPath_ALUhw_i_Q_EXTENDED_57_port, C2 
                           => n8578, A => n9943, B => n9942, ZN => n9962);
   U10998 : OAI211_X1 port map( C1 => n9974, C2 => n9941, A => n9940, B => 
                           n9939, ZN => n9942);
   U10999 : AOI21_X1 port map( B1 => n9937, B2 => n9964, A => n9936, ZN => 
                           n9941);
   U11000 : INV_X1 port map( A => n9935, ZN => n9936);
   U11001 : NOR2_X1 port map( A1 => n9934, A2 => n9933, ZN => n9943);
   U11002 : XNOR2_X1 port map( A => n9932, B => n9937, ZN => n9933);
   U11003 : INV_X1 port map( A => n9967, ZN => n9934);
   U11004 : OAI222_X1 port map( A1 => n8549, A2 => n10641, B1 => n10702, B2 => 
                           n8381, C1 => n7759, C2 => n10640, ZN => n7044);
   U11005 : XNOR2_X1 port map( A => n10638, B => n8381, ZN => n10639);
   U11006 : OAI222_X1 port map( A1 => n12093, A2 => n9930, B1 => n10482, B2 => 
                           n9929, C1 => n12092, C2 => n512, ZN => n6997);
   U11007 : NOR4_X1 port map( A1 => n9928, A2 => n9927, A3 => n9926, A4 => 
                           n9925, ZN => n9929);
   U11008 : OAI21_X1 port map( B1 => n9924, B2 => n10505, A => n9923, ZN => 
                           n9925);
   U11009 : AOI22_X1 port map( A1 => n10094, A2 => n10502, B1 => n9992, B2 => 
                           n10510, ZN => n9923);
   U11010 : OAI22_X1 port map( A1 => n10064, A2 => n10462, B1 => n10177, B2 => 
                           n10444, ZN => n9926);
   U11011 : INV_X1 port map( A => n10158, ZN => n10177);
   U11012 : NAND2_X1 port map( A1 => n9921, A2 => n10286, ZN => n10188);
   U11013 : OAI21_X1 port map( B1 => n9560, B2 => n12081, A => n9352, ZN => 
                           n9918);
   U11014 : OAI22_X1 port map( A1 => n9946, A2 => n10460, B1 => n8311, B2 => 
                           n10376, ZN => n9927);
   U11015 : OAI22_X1 port map( A1 => n10155, A2 => n10442, B1 => n9916, B2 => 
                           n10507, ZN => n9928);
   U11016 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_58_port, B2 =>
                           n8578, A => n9915, ZN => n9930);
   U11017 : OAI211_X1 port map( C1 => n9974, C2 => n9914, A => n9913, B => 
                           n9912, ZN => n9915);
   U11018 : AOI21_X1 port map( B1 => n10458, B2 => n9919, A => n9908, ZN => 
                           n9910);
   U11019 : NOR2_X1 port map( A1 => n10465, A2 => n9919, ZN => n9908);
   U11020 : AOI21_X1 port map( B1 => n10469, B2 => n10181, A => n9907, ZN => 
                           n9911);
   U11021 : NOR2_X1 port map( A1 => n10465, A2 => n10181, ZN => n9907);
   U11022 : NAND2_X1 port map( A1 => n9967, A2 => n9906, ZN => n9913);
   U11023 : XNOR2_X1 port map( A => n9903, B => n9905, ZN => n9914);
   U11024 : OAI21_X1 port map( B1 => n10594, B2 => n7759, A => n10593, ZN => 
                           n7034);
   U11025 : AOI22_X1 port map( A1 => n12070, A2 => i_RD1_25_port, B1 => 
                           IRAM_ADDRESS_25_port, B2 => n10835, ZN => n10593);
   U11026 : XNOR2_X1 port map( A => n10590, B => IRAM_ADDRESS_25_port, ZN => 
                           n10591);
   U11027 : OAI211_X1 port map( C1 => n220, C2 => n10702, A => n10637, B => 
                           n10636, ZN => n7043);
   U11028 : OR2_X1 port map( A1 => n8549, A2 => n10635, ZN => n10636);
   U11029 : INV_X1 port map( A => i_RD1_16_port, ZN => n10635);
   U11030 : OAI21_X1 port map( B1 => n8248, B2 => n9317, A => n8451, ZN => 
                           n10633);
   U11031 : OAI21_X1 port map( B1 => n10589, B2 => n7759, A => n10588, ZN => 
                           n7033);
   U11032 : AOI22_X1 port map( A1 => n12070, A2 => i_RD1_26_port, B1 => 
                           IRAM_ADDRESS_26_port, B2 => n10835, ZN => n10588);
   U11033 : AOI22_X1 port map( A1 => n12070, A2 => i_RD1_18_port, B1 => 
                           IRAM_ADDRESS_18_port, B2 => n10835, ZN => n12066);
   U11034 : NAND2_X1 port map( A1 => n10554, A2 => n9330, ZN => n9326);
   U11035 : NAND2_X1 port map( A1 => n10545, A2 => n9329, ZN => n9327);
   U11036 : OAI222_X1 port map( A1 => n12093, A2 => n9901, B1 => n10482, B2 => 
                           n9900, C1 => n12092, C2 => n513, ZN => n6996);
   U11037 : NOR4_X1 port map( A1 => n9899, A2 => n9898, A3 => n9897, A4 => 
                           n9896, ZN => n9900);
   U11038 : OAI22_X1 port map( A1 => n9895, A2 => n10507, B1 => n9924, B2 => 
                           n10460, ZN => n9896);
   U11039 : OAI21_X1 port map( B1 => n8311, B2 => n10479, A => n9894, ZN => 
                           n9897);
   U11040 : AOI22_X1 port map( A1 => n10094, A2 => n10495, B1 => n9992, B2 => 
                           n10498, ZN => n9894);
   U11041 : OAI22_X1 port map( A1 => n9916, A2 => n10505, B1 => n10064, B2 => 
                           n10442, ZN => n9898);
   U11042 : OAI22_X1 port map( A1 => n10155, A2 => n10444, B1 => n9946, B2 => 
                           n10388, ZN => n9899);
   U11043 : AOI211_X1 port map( C1 => n7785, C2 => n9893, A => n9892, B => 
                           n9891, ZN => n10155);
   U11044 : NOR2_X1 port map( A1 => n9890, A2 => n10284, ZN => n9891);
   U11045 : OAI211_X1 port map( C1 => n9889, C2 => n10184, A => n9888, B => 
                           n9887, ZN => n9892);
   U11046 : AOI22_X1 port map( A1 => n9983, A2 => n8552, B1 => n10229, B2 => 
                           n9886, ZN => n9887);
   U11047 : OAI21_X1 port map( B1 => n10286, B2 => n9885, A => n9884, ZN => 
                           n9888);
   U11048 : AOI21_X1 port map( B1 => n12087, B2 => n10164, A => n10182, ZN => 
                           n9884);
   U11049 : AOI21_X1 port map( B1 => n12082, B2 => n8016, A => n9365, ZN => 
                           n9889);
   U11050 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_59_port, B2 =>
                           n8578, A => n9883, ZN => n9901);
   U11051 : OAI21_X1 port map( B1 => n9882, B2 => n9974, A => n9881, ZN => 
                           n9883);
   U11052 : AOI21_X1 port map( B1 => n9967, B2 => n9880, A => n9879, ZN => 
                           n9881);
   U11053 : OAI211_X1 port map( C1 => n9878, C2 => n10465, A => n9877, B => 
                           n9876, ZN => n9879);
   U11054 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n537, B => n7797, ZN => 
                           n9878);
   U11055 : XNOR2_X1 port map( A => n9873, B => n9872, ZN => n9880);
   U11056 : OAI21_X1 port map( B1 => n9904, B2 => n9905, A => n9871, ZN => 
                           n9873);
   U11057 : OAI21_X1 port map( B1 => n9870, B2 => n9965, A => n9869, ZN => 
                           n9904);
   U11058 : NOR2_X1 port map( A1 => n9868, A2 => n10421, ZN => n9967);
   U11059 : NAND2_X1 port map( A1 => n9868, A2 => n10450, ZN => n9974);
   U11060 : NAND2_X1 port map( A1 => n9866, A2 => n9865, ZN => n9872);
   U11061 : OAI21_X1 port map( B1 => n10586, B2 => n7759, A => n10585, ZN => 
                           n7032);
   U11062 : AOI22_X1 port map( A1 => n12070, A2 => i_RD1_27_port, B1 => 
                           IRAM_ADDRESS_27_port, B2 => n10835, ZN => n10585);
   U11063 : XNOR2_X1 port map( A => n10584, B => n10583, ZN => n10586);
   U11064 : XNOR2_X1 port map( A => n10590, B => IRAM_ADDRESS_27_port, ZN => 
                           n10583);
   U11065 : AOI22_X1 port map( A1 => n12070, A2 => i_RD1_19_port, B1 => 
                           IRAM_ADDRESS_19_port, B2 => n10835, ZN => n12068);
   U11066 : OAI21_X1 port map( B1 => n9331, B2 => n10551, A => n10545, ZN => 
                           n9332);
   U11067 : INV_X1 port map( A => n10554, ZN => n9331);
   U11068 : OAI22_X1 port map( A1 => n9863, A2 => n12093, B1 => n514, B2 => 
                           n12092, ZN => n6995);
   U11069 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_60_port, B2 =>
                           n8578, A => n9862, ZN => n9863);
   U11070 : OAI21_X1 port map( B1 => n9861, B2 => n10114, A => n9860, ZN => 
                           n9862);
   U11071 : AOI211_X1 port map( C1 => n10114, C2 => n9859, A => n9858, B => 
                           n9857, ZN => n9860);
   U11072 : AOI21_X1 port map( B1 => n9856, B2 => n9855, A => n9854, ZN => 
                           n9857);
   U11073 : NOR2_X1 port map( A1 => n9853, A2 => n10452, ZN => n9858);
   U11074 : NOR3_X1 port map( A1 => n9852, A2 => n9851, A3 => n9850, ZN => 
                           n9853);
   U11075 : OAI22_X1 port map( A1 => n9849, A2 => n10507, B1 => n10063, B2 => 
                           n10442, ZN => n9850);
   U11076 : INV_X1 port map( A => n10094, ZN => n10063);
   U11077 : OAI211_X1 port map( C1 => n8311, C2 => n10462, A => n9848, B => 
                           n9847, ZN => n9851);
   U11078 : AOI22_X1 port map( A1 => n10107, A2 => n10493, B1 => n10502, B2 => 
                           n9992, ZN => n9847);
   U11079 : INV_X1 port map( A => n10064, ZN => n10107);
   U11080 : NAND2_X1 port map( A1 => n9413, A2 => n9421, ZN => n10112);
   U11081 : NAND2_X1 port map( A1 => n10473, A2 => n12082, ZN => n9413);
   U11082 : AOI22_X1 port map( A1 => n9843, A2 => n10461, B1 => n9949, B2 => 
                           n10510, ZN => n9848);
   U11083 : OAI22_X1 port map( A1 => n9946, A2 => n10376, B1 => n9916, B2 => 
                           n10460, ZN => n9852);
   U11084 : OAI21_X1 port map( B1 => n9842, B2 => n9841, A => n9840, ZN => 
                           n9859);
   U11085 : INV_X1 port map( A => n10469, ZN => n10488);
   U11086 : AOI21_X1 port map( B1 => n9838, B2 => n9841, A => n9837, ZN => 
                           n9861);
   U11087 : OAI222_X1 port map( A1 => n8549, A2 => n10599, B1 => n7759, B2 => 
                           n10598, C1 => n8377, C2 => n10702, ZN => n7035);
   U11088 : XNOR2_X1 port map( A => n10595, B => n8377, ZN => n10596);
   U11089 : NAND2_X1 port map( A1 => n8466, A2 => n8458, ZN => n10597);
   U11090 : NAND2_X1 port map( A1 => n10554, A2 => n8469, ZN => n8458);
   U11091 : INV_X1 port map( A => i_RD1_24_port, ZN => n10599);
   U11092 : OAI222_X1 port map( A1 => n10631, A2 => n8549, B1 => n10702, B2 => 
                           intadd_0_A_0_port, C1 => n7759, C2 => n10630, ZN => 
                           n7039);
   U11093 : NAND2_X1 port map( A1 => n10627, A2 => n10626, ZN => n10629);
   U11094 : INV_X1 port map( A => i_RD1_20_port, ZN => n10631);
   U11095 : OAI222_X1 port map( A1 => n8549, A2 => n10582, B1 => n10702, B2 => 
                           n8156, C1 => n7759, C2 => n10581, ZN => n7031);
   U11096 : INV_X1 port map( A => i_RD1_28_port, ZN => n10582);
   U11097 : OAI222_X1 port map( A1 => n8549, A2 => n10625, B1 => n10702, B2 => 
                           n8387, C1 => n7759, C2 => n10624, ZN => n7038);
   U11098 : XNOR2_X1 port map( A => n10623, B => n10622, ZN => n10624);
   U11099 : NAND2_X1 port map( A1 => n10621, A2 => n10620, ZN => n10622);
   U11100 : INV_X1 port map( A => n10627, ZN => n10619);
   U11101 : INV_X1 port map( A => i_RD1_21_port, ZN => n10625);
   U11102 : OAI222_X1 port map( A1 => n8549, A2 => n10618, B1 => n10702, B2 => 
                           n8390, C1 => n7759, C2 => n10617, ZN => n7037);
   U11103 : XNOR2_X1 port map( A => n10616, B => n10615, ZN => n10617);
   U11104 : NAND2_X1 port map( A1 => n10614, A2 => n10613, ZN => n10615);
   U11105 : INV_X1 port map( A => n10610, ZN => n10611);
   U11106 : INV_X1 port map( A => i_RD1_22_port, ZN => n10618);
   U11107 : OAI222_X1 port map( A1 => n8549, A2 => n10609, B1 => n10702, B2 => 
                           n8394, C1 => n7759, C2 => n10608, ZN => n7036);
   U11108 : XNOR2_X1 port map( A => n10607, B => n10606, ZN => n10608);
   U11109 : NOR2_X1 port map( A1 => n10605, A2 => n10604, ZN => n10606);
   U11110 : INV_X1 port map( A => n10603, ZN => n10605);
   U11111 : AOI21_X1 port map( B1 => n10602, B2 => n10601, A => n10600, ZN => 
                           n10607);
   U11112 : OAI21_X1 port map( B1 => n9833, B2 => n9832, A => n10840, ZN => 
                           n9834);
   U11113 : OAI211_X1 port map( C1 => n8311, C2 => n10442, A => n9831, B => 
                           n9830, ZN => n9832);
   U11114 : AOI22_X1 port map( A1 => n9829, A2 => n10476, B1 => n9992, B2 => 
                           n10495, ZN => n9830);
   U11115 : AOI22_X1 port map( A1 => n9843, A2 => n10499, B1 => n9949, B2 => 
                           n10498, ZN => n9831);
   U11116 : OAI211_X1 port map( C1 => n9849, C2 => n10505, A => n9828, B => 
                           n9827, ZN => n9833);
   U11117 : NAND2_X1 port map( A1 => n10094, A2 => n10493, ZN => n9827);
   U11118 : NAND4_X1 port map( A1 => n9826, A2 => n9825, A3 => n9824, A4 => 
                           n9823, ZN => n10094);
   U11119 : NAND2_X1 port map( A1 => n9822, A2 => n7785, ZN => n9823);
   U11120 : INV_X1 port map( A => n9821, ZN => n9822);
   U11121 : AOI22_X1 port map( A1 => n9985, A2 => n10091, B1 => n10229, B2 => 
                           n9820, ZN => n9824);
   U11122 : NOR2_X1 port map( A1 => n10284, A2 => n10115, ZN => n9985);
   U11123 : AOI22_X1 port map( A1 => n10282, A2 => n10090, B1 => n10231, B2 => 
                           n10087, ZN => n9825);
   U11124 : NAND2_X1 port map( A1 => n9401, A2 => n9403, ZN => n10087);
   U11125 : NAND2_X1 port map( A1 => n7818, A2 => n12082, ZN => n9401);
   U11126 : AOI22_X1 port map( A1 => n10089, A2 => n9844, B1 => n10086, B2 => 
                           n10288, ZN => n9826);
   U11127 : AOI22_X1 port map( A1 => n10502, A2 => n9977, B1 => n9819, B2 => 
                           n10510, ZN => n9828);
   U11128 : INV_X1 port map( A => n9916, ZN => n9819);
   U11129 : INV_X1 port map( A => n9946, ZN => n9977);
   U11130 : AOI22_X1 port map( A1 => n10408, A2 => n9818, B1 => n7782, B2 => 
                           DRAM_ADDRESS_29_port, ZN => n9835);
   U11131 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n435, B => n9817, ZN => 
                           n9818);
   U11132 : NOR2_X1 port map( A1 => n10513, A2 => n10465, ZN => n10408);
   U11133 : NAND2_X1 port map( A1 => n10841, A2 => n10452, ZN => n10513);
   U11134 : AOI21_X1 port map( B1 => n8471, B2 => n8303, A => n8470, ZN => 
                           n8477);
   U11135 : INV_X1 port map( A => n10575, ZN => n8470);
   U11136 : AOI22_X1 port map( A1 => n12070, A2 => i_RD1_30_port, B1 => 
                           IRAM_ADDRESS_30_port, B2 => n10835, ZN => n10575);
   U11137 : XNOR2_X1 port map( A => n8472, B => IRAM_ADDRESS_30_port, ZN => 
                           n8471);
   U11138 : NOR2_X1 port map( A1 => n10834, A2 => n10833, ZN => n8472);
   U11139 : NAND2_X1 port map( A1 => n9276, A2 => n8110, ZN => n9277);
   U11140 : NAND2_X1 port map( A1 => n10833, A2 => IRAM_ADDRESS_30_port, ZN => 
                           n8473);
   U11141 : NOR2_X1 port map( A1 => n10576, A2 => IRAM_ADDRESS_29_port, ZN => 
                           n10834);
   U11142 : OAI21_X1 port map( B1 => IRAM_ADDRESS_26_port, B2 => 
                           IRAM_ADDRESS_27_port, A => n10590, ZN => n10574);
   U11143 : XNOR2_X1 port map( A => n10590, B => IRAM_ADDRESS_26_port, ZN => 
                           n10587);
   U11144 : NOR2_X1 port map( A1 => n10590, A2 => IRAM_ADDRESS_25_port, ZN => 
                           n10572);
   U11145 : NAND2_X1 port map( A1 => n10590, A2 => IRAM_ADDRESS_25_port, ZN => 
                           n10573);
   U11146 : OR2_X1 port map( A1 => n10569, A2 => n184, ZN => n10570);
   U11147 : NAND2_X1 port map( A1 => n8446, A2 => n7775, ZN => n8445);
   U11148 : NAND2_X1 port map( A1 => n8448, A2 => n8450, ZN => n8447);
   U11149 : XNOR2_X1 port map( A => n12065, B => IRAM_ADDRESS_17_port, ZN => 
                           n9321);
   U11150 : AND2_X1 port map( A1 => n10638, A2 => n8381, ZN => n9317);
   U11151 : AND2_X1 port map( A1 => n9324, A2 => n9320, ZN => n10634);
   U11152 : NAND2_X1 port map( A1 => n9316, A2 => n8384, ZN => n10642);
   U11153 : NOR2_X1 port map( A1 => n9316, A2 => n8384, ZN => n10643);
   U11154 : NAND2_X1 port map( A1 => n9313, A2 => IRAM_ADDRESS_13_port, ZN => 
                           n9314);
   U11155 : INV_X1 port map( A => n9312, ZN => n9313);
   U11156 : XNOR2_X1 port map( A => n9312, B => n8398, ZN => n10648);
   U11157 : NOR2_X1 port map( A1 => n10656, A2 => n8383, ZN => n9308);
   U11158 : NAND2_X1 port map( A1 => n10656, A2 => n8383, ZN => n9309);
   U11159 : NAND2_X1 port map( A1 => n10661, A2 => IRAM_ADDRESS_10_port, ZN => 
                           n9306);
   U11160 : NOR2_X1 port map( A1 => n10661, A2 => IRAM_ADDRESS_10_port, ZN => 
                           n9307);
   U11161 : NAND2_X1 port map( A1 => n9299, A2 => n224, ZN => n9303);
   U11162 : NOR2_X1 port map( A1 => n9299, A2 => n224, ZN => n9304);
   U11163 : NAND2_X1 port map( A1 => n9298, A2 => n9297, ZN => n9305);
   U11164 : NAND2_X1 port map( A1 => n10664, A2 => IRAM_ADDRESS_7_port, ZN => 
                           n9291);
   U11165 : NOR2_X1 port map( A1 => n10664, A2 => IRAM_ADDRESS_7_port, ZN => 
                           n9292);
   U11166 : NAND2_X1 port map( A1 => IRAM_ADDRESS_6_port, A2 => IR_6_port, ZN 
                           => n9290);
   U11167 : NAND2_X1 port map( A1 => n9289, A2 => n10675, ZN => n10671);
   U11168 : NAND2_X1 port map( A1 => n9288, A2 => IRAM_ADDRESS_5_port, ZN => 
                           n10675);
   U11169 : INV_X1 port map( A => n9287, ZN => n9288);
   U11170 : AOI21_X1 port map( B1 => n10684, B2 => n10681, A => n10680, ZN => 
                           n10676);
   U11171 : AND2_X1 port map( A1 => n9286, A2 => n8325, ZN => n10680);
   U11172 : NAND2_X1 port map( A1 => n9285, A2 => IRAM_ADDRESS_4_port, ZN => 
                           n10681);
   U11173 : INV_X1 port map( A => n9286, ZN => n9285);
   U11174 : AOI21_X1 port map( B1 => n10692, B2 => n10686, A => n10687, ZN => 
                           n9283);
   U11175 : NAND2_X1 port map( A1 => n9281, A2 => IRAM_ADDRESS_2_port, ZN => 
                           n10693);
   U11176 : NAND2_X1 port map( A1 => n9279, A2 => intadd_1_A_0_port, ZN => 
                           n10698);
   U11177 : AOI22_X1 port map( A1 => n8462, A2 => n8465, B1 => n8459, B2 => 
                           n8461, ZN => n8457);
   U11178 : INV_X1 port map( A => n8466, ZN => n8461);
   U11179 : AOI21_X1 port map( B1 => n8466, B2 => n8460, A => 
                           IRAM_ADDRESS_24_port, ZN => n8459);
   U11180 : INV_X1 port map( A => n8469, ZN => n8460);
   U11181 : NAND2_X1 port map( A1 => n8466, A2 => IRAM_ADDRESS_24_port, ZN => 
                           n8465);
   U11182 : AOI21_X1 port map( B1 => n8466, B2 => n8464, A => n8463, ZN => 
                           n8462);
   U11183 : INV_X1 port map( A => n10595, ZN => n8463);
   U11184 : AND2_X1 port map( A1 => n10571, A2 => n10568, ZN => n10595);
   U11185 : OR2_X1 port map( A1 => n10569, A2 => n185, ZN => n10568);
   U11186 : AND2_X1 port map( A1 => n10566, A2 => n8394, ZN => n10604);
   U11187 : NAND2_X1 port map( A1 => n10565, A2 => n10613, ZN => n10600);
   U11188 : NAND2_X1 port map( A1 => n10564, A2 => n8390, ZN => n10613);
   U11189 : NAND2_X1 port map( A1 => n10610, A2 => n10614, ZN => n10565);
   U11190 : OAI21_X1 port map( B1 => n10563, B2 => n10626, A => n10620, ZN => 
                           n10610);
   U11191 : NAND2_X1 port map( A1 => n10562, A2 => n8387, ZN => n10620);
   U11192 : NAND2_X1 port map( A1 => n10561, A2 => intadd_0_A_0_port, ZN => 
                           n10626);
   U11193 : NOR2_X1 port map( A1 => n8468, A2 => n10567, ZN => n8467);
   U11194 : NAND2_X1 port map( A1 => n10552, A2 => n10553, ZN => n8468);
   U11195 : NAND2_X1 port map( A1 => n10546, A2 => n10545, ZN => n10553);
   U11196 : INV_X1 port map( A => n10548, ZN => n10545);
   U11197 : XNOR2_X1 port map( A => n10549, B => n8392, ZN => n10546);
   U11198 : NOR2_X1 port map( A1 => n8469, A2 => n8377, ZN => n8464);
   U11199 : NOR2_X1 port map( A1 => n7758, A2 => n10567, ZN => n8469);
   U11200 : NAND2_X1 port map( A1 => n10601, A2 => n10603, ZN => n10567);
   U11201 : OR2_X1 port map( A1 => n10566, A2 => n8394, ZN => n10603);
   U11202 : NAND2_X1 port map( A1 => n10560, A2 => n10559, ZN => n10566);
   U11203 : NAND2_X1 port map( A1 => n10571, A2 => n186, ZN => n10559);
   U11204 : NOR2_X1 port map( A1 => n10612, A2 => n10558, ZN => n10601);
   U11205 : INV_X1 port map( A => n10614, ZN => n10558);
   U11206 : OR2_X1 port map( A1 => n10564, A2 => n8390, ZN => n10614);
   U11207 : NAND2_X1 port map( A1 => n10560, A2 => n10557, ZN => n10564);
   U11208 : NAND2_X1 port map( A1 => n10571, A2 => n187, ZN => n10557);
   U11209 : NAND2_X1 port map( A1 => n10627, A2 => n10621, ZN => n10612);
   U11210 : INV_X1 port map( A => n10563, ZN => n10621);
   U11211 : NOR2_X1 port map( A1 => n10562, A2 => n8387, ZN => n10563);
   U11212 : NAND2_X1 port map( A1 => n10560, A2 => n10556, ZN => n10562);
   U11213 : NAND2_X1 port map( A1 => n10571, A2 => n188, ZN => n10556);
   U11214 : OR2_X1 port map( A1 => n10561, A2 => intadd_0_A_0_port, ZN => 
                           n10627);
   U11215 : NAND2_X1 port map( A1 => n10560, A2 => n10555, ZN => n10561);
   U11216 : NAND2_X1 port map( A1 => n10571, A2 => n189, ZN => n10555);
   U11217 : NAND2_X1 port map( A1 => n10571, A2 => n10569, ZN => n10560);
   U11218 : NOR2_X1 port map( A1 => n10548, A2 => n10547, ZN => n10550);
   U11219 : NOR2_X1 port map( A1 => n10549, A2 => IRAM_ADDRESS_19_port, ZN => 
                           n10547);
   U11220 : NAND2_X1 port map( A1 => n10571, A2 => n9328, ZN => n10549);
   U11221 : OR2_X1 port map( A1 => n10569, A2 => n190, ZN => n9328);
   U11222 : NOR2_X1 port map( A1 => n9323, A2 => IRAM_ADDRESS_18_port, ZN => 
                           n10548);
   U11223 : NAND2_X1 port map( A1 => n9330, A2 => n9329, ZN => n10551);
   U11224 : NAND2_X1 port map( A1 => n9323, A2 => IRAM_ADDRESS_18_port, ZN => 
                           n9329);
   U11225 : NAND2_X1 port map( A1 => n10571, A2 => n9322, ZN => n9323);
   U11226 : OR2_X1 port map( A1 => n10569, A2 => n191, ZN => n9322);
   U11227 : AOI21_X1 port map( B1 => n9325, B2 => n8367, A => n8309, ZN => 
                           n9330);
   U11228 : INV_X1 port map( A => n9324, ZN => n9325);
   U11229 : NAND2_X1 port map( A1 => n9318, A2 => IRAM_ADDRESS_16_port, ZN => 
                           n9324);
   U11230 : NAND2_X1 port map( A1 => n10571, A2 => n9319, ZN => n9318);
   U11231 : OR2_X1 port map( A1 => n10569, A2 => n193, ZN => n9319);
   U11232 : INV_X1 port map( A => n8101, ZN => n9302);
   U11233 : NAND2_X1 port map( A1 => n10740, A2 => n9273, ZN => n9274);
   U11234 : AOI21_X1 port map( B1 => n10828, B2 => n9268, A => n9267, ZN => 
                           n9269);
   U11235 : OAI21_X1 port map( B1 => n10523, B2 => n9266, A => n10719, ZN => 
                           n9267);
   U11236 : NAND2_X1 port map( A1 => n9265, A2 => n9264, ZN => n9268);
   U11237 : NOR2_X1 port map( A1 => n10720, A2 => n8102, ZN => n10827);
   U11238 : INV_X1 port map( A => n10711, ZN => n10828);
   U11239 : AND2_X1 port map( A1 => n9259, A2 => n9258, ZN => n9260);
   U11240 : INV_X1 port map( A => n9246, ZN => n9248);
   U11241 : NAND2_X1 port map( A1 => n9242, A2 => n9241, ZN => n9243);
   U11242 : AOI21_X1 port map( B1 => n8685, B2 => i_RD2_0_port, A => n9240, ZN 
                           => n9241);
   U11243 : NAND2_X1 port map( A1 => n10518, A2 => n8687, ZN => n9242);
   U11244 : NAND4_X1 port map( A1 => n9236, A2 => n9235, A3 => n9234, A4 => 
                           n9233, ZN => n9253);
   U11245 : INV_X1 port map( A => n7689, ZN => n9259);
   U11246 : INV_X1 port map( A => n9223, ZN => n9224);
   U11247 : OAI22_X1 port map( A1 => n9222, A2 => n9221, B1 => n9220, B2 => 
                           n10578, ZN => n9225);
   U11248 : INV_X1 port map( A => i_RD1_29_port, ZN => n10578);
   U11249 : NAND2_X1 port map( A1 => n9219, A2 => i_RD1_28_port, ZN => n9221);
   U11250 : INV_X1 port map( A => n9218, ZN => n9219);
   U11251 : INV_X1 port map( A => n9217, ZN => n9222);
   U11252 : NOR2_X1 port map( A1 => n9216, A2 => n9215, ZN => n9226);
   U11253 : INV_X1 port map( A => n9214, ZN => n9216);
   U11254 : NAND4_X1 port map( A1 => n9212, A2 => n9211, A3 => n9214, A4 => 
                           n9217, ZN => n9255);
   U11255 : XNOR2_X1 port map( A => n9220, B => i_RD1_29_port, ZN => n9217);
   U11256 : NAND2_X1 port map( A1 => n9210, A2 => n9209, ZN => n9220);
   U11257 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_29_port, ZN => 
                           n9209);
   U11258 : NAND2_X1 port map( A1 => n9836, A2 => n8687, ZN => n9210);
   U11259 : OAI211_X1 port map( C1 => n8106, C2 => n8334, A => n7698, B => 
                           n9206, ZN => n9836);
   U11260 : NAND2_X1 port map( A1 => n7690, A2 => IRAM_ADDRESS_29_port, ZN => 
                           n9206);
   U11261 : XNOR2_X1 port map( A => n9205, B => i_RD1_30_port, ZN => n9214);
   U11262 : XNOR2_X1 port map( A => n9218, B => i_RD1_28_port, ZN => n9211);
   U11263 : NAND2_X1 port map( A1 => n9204, A2 => n9203, ZN => n9218);
   U11264 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_28_port, ZN => 
                           n9203);
   U11265 : NAND2_X1 port map( A1 => n9864, A2 => n8687, ZN => n9204);
   U11266 : OAI211_X1 port map( C1 => n571, C2 => n8106, A => n7697, B => n9202
                           , ZN => n9864);
   U11267 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_28_port, ZN => 
                           n9202);
   U11268 : NAND2_X1 port map( A1 => n9199, A2 => n9198, ZN => n9201);
   U11269 : OAI21_X1 port map( B1 => n9197, B2 => n9196, A => n9195, ZN => 
                           n9199);
   U11270 : INV_X1 port map( A => n9194, ZN => n9197);
   U11271 : AND2_X1 port map( A1 => n9200, A2 => n9196, ZN => n9189);
   U11272 : NAND2_X1 port map( A1 => n9188, A2 => i_RD1_24_port, ZN => n9196);
   U11273 : NAND2_X1 port map( A1 => n9187, A2 => i_RD1_27_port, ZN => n9200);
   U11274 : INV_X1 port map( A => n9186, ZN => n9187);
   U11275 : AOI22_X1 port map( A1 => n9186, A2 => n9185, B1 => n9184, B2 => 
                           n9183, ZN => n9198);
   U11276 : INV_X1 port map( A => i_RD1_26_port, ZN => n9183);
   U11277 : INV_X1 port map( A => n9182, ZN => n9184);
   U11278 : INV_X1 port map( A => i_RD1_27_port, ZN => n9185);
   U11279 : NAND2_X1 port map( A1 => n7699, A2 => IRAM_ADDRESS_27_port, ZN => 
                           n9181);
   U11280 : INV_X1 port map( A => n9180, ZN => n9190);
   U11281 : OAI21_X1 port map( B1 => i_RD1_24_port, B2 => n9188, A => n9194, ZN
                           => n9180);
   U11282 : NAND2_X1 port map( A1 => n9179, A2 => n9178, ZN => n9194);
   U11283 : INV_X1 port map( A => i_RD1_25_port, ZN => n9178);
   U11284 : AOI21_X1 port map( B1 => n10000, B2 => n8686, A => n9177, ZN => 
                           n9188);
   U11285 : AND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_24_port, ZN => 
                           n9177);
   U11286 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_24_port, ZN => 
                           n9176);
   U11287 : AOI22_X1 port map( A1 => n9182, A2 => i_RD1_26_port, B1 => n9175, 
                           B2 => i_RD1_25_port, ZN => n9195);
   U11288 : INV_X1 port map( A => n9179, ZN => n9175);
   U11289 : NAND2_X1 port map( A1 => n9174, A2 => n9173, ZN => n9179);
   U11290 : NAND2_X1 port map( A1 => n8685, A2 => i_RD2_25_port, ZN => n9173);
   U11291 : NAND2_X1 port map( A1 => n9963, A2 => n8686, ZN => n9174);
   U11292 : OAI211_X1 port map( C1 => n568, C2 => n8106, A => n7698, B => n9172
                           , ZN => n9963);
   U11293 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_25_port, ZN => 
                           n9172);
   U11294 : AOI21_X1 port map( B1 => n9931, B2 => n8686, A => n9171, ZN => 
                           n9182);
   U11295 : AND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_26_port, ZN => 
                           n9171);
   U11296 : OAI211_X1 port map( C1 => n8106, C2 => n8370, A => n7697, B => 
                           n9170, ZN => n9931);
   U11297 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_26_port, ZN => 
                           n9170);
   U11298 : NAND2_X1 port map( A1 => n9169, A2 => n9168, ZN => n9192);
   U11299 : NAND2_X1 port map( A1 => n9167, A2 => n9166, ZN => n9169);
   U11300 : NAND2_X1 port map( A1 => n9165, A2 => i_RD1_22_port, ZN => n9166);
   U11301 : INV_X1 port map( A => n9164, ZN => n9165);
   U11302 : NOR2_X1 port map( A1 => n9254, A2 => n9162, ZN => n9163);
   U11303 : NOR2_X1 port map( A1 => n9161, A2 => i_RD1_21_port, ZN => n9162);
   U11304 : NAND2_X1 port map( A1 => n9159, A2 => n10609, ZN => n9168);
   U11305 : INV_X1 port map( A => i_RD1_23_port, ZN => n10609);
   U11306 : INV_X1 port map( A => n9158, ZN => n9159);
   U11307 : NAND2_X1 port map( A1 => n9158, A2 => i_RD1_23_port, ZN => n9167);
   U11308 : AOI21_X1 port map( B1 => n10037, B2 => n8686, A => n9157, ZN => 
                           n9158);
   U11309 : AND2_X1 port map( A1 => n8685, A2 => i_RD2_23_port, ZN => n9157);
   U11310 : OAI211_X1 port map( C1 => n566, C2 => n8106, A => n7698, B => n9156
                           , ZN => n10037);
   U11311 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_23_port, ZN => 
                           n9156);
   U11312 : XNOR2_X1 port map( A => n9164, B => i_RD1_22_port, ZN => n9160);
   U11313 : NAND2_X1 port map( A1 => n9155, A2 => n9154, ZN => n9164);
   U11314 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_22_port, ZN => 
                           n9154);
   U11315 : NAND2_X1 port map( A1 => n10070, A2 => n8687, ZN => n9155);
   U11316 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_22_port, ZN => 
                           n9153);
   U11317 : NAND2_X1 port map( A1 => n9152, A2 => n9151, ZN => n9237);
   U11318 : NAND2_X1 port map( A1 => n9150, A2 => i_RD1_20_port, ZN => n9151);
   U11319 : NAND2_X1 port map( A1 => n9161, A2 => i_RD1_21_port, ZN => n9152);
   U11320 : AOI21_X1 port map( B1 => n10102, B2 => n8686, A => n9149, ZN => 
                           n9161);
   U11321 : AND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_21_port, ZN => 
                           n9149);
   U11322 : OAI211_X1 port map( C1 => n564, C2 => n8106, A => n7697, B => n9148
                           , ZN => n10102);
   U11323 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_21_port, ZN => 
                           n9148);
   U11324 : AOI21_X1 port map( B1 => n10135, B2 => n8687, A => n9145, ZN => 
                           n9150);
   U11325 : AND2_X1 port map( A1 => n8685, A2 => i_RD2_20_port, ZN => n9145);
   U11326 : OAI211_X1 port map( C1 => n8106, C2 => n8369, A => n7698, B => 
                           n9144, ZN => n10135);
   U11327 : NAND2_X1 port map( A1 => n7690, A2 => IRAM_ADDRESS_20_port, ZN => 
                           n9144);
   U11328 : AOI21_X1 port map( B1 => n9143, B2 => n9142, A => n9141, ZN => 
                           n9147);
   U11329 : INV_X1 port map( A => n9140, ZN => n9142);
   U11330 : OAI211_X1 port map( C1 => n9139, C2 => n9138, A => n9137, B => 
                           n9136, ZN => n9143);
   U11331 : NAND2_X1 port map( A1 => n9135, A2 => i_RD1_17_port, ZN => n9136);
   U11332 : INV_X1 port map( A => n9134, ZN => n9135);
   U11333 : INV_X1 port map( A => n9133, ZN => n9137);
   U11334 : NAND2_X1 port map( A1 => n9132, A2 => i_RD1_16_port, ZN => n9138);
   U11335 : AOI21_X1 port map( B1 => n10173, B2 => n8687, A => n9129, ZN => 
                           n9141);
   U11336 : OAI21_X1 port map( B1 => n8687, B2 => n9128, A => i_RD1_19_port, ZN
                           => n9129);
   U11337 : AND2_X1 port map( A1 => n9127, A2 => i_RD1_18_port, ZN => n9133);
   U11338 : OAI21_X1 port map( B1 => n9127, B2 => i_RD1_18_port, A => n9126, ZN
                           => n9140);
   U11339 : OAI21_X1 port map( B1 => n10173, B2 => n8685, A => n9125, ZN => 
                           n9126);
   U11340 : AOI21_X1 port map( B1 => n8685, B2 => n9128, A => i_RD1_19_port, ZN
                           => n9125);
   U11341 : INV_X1 port map( A => i_RD2_19_port, ZN => n9128);
   U11342 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_19_port, ZN => 
                           n9124);
   U11343 : OAI21_X1 port map( B1 => n10212, B2 => n8685, A => n9123, ZN => 
                           n9127);
   U11344 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => n9122, ZN => n9123);
   U11345 : INV_X1 port map( A => i_RD2_18_port, ZN => n9122);
   U11346 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_18_port, ZN => 
                           n9121);
   U11347 : XNOR2_X1 port map( A => n9132, B => i_RD1_16_port, ZN => n9131);
   U11348 : AOI21_X1 port map( B1 => n10539, B2 => n8687, A => n9120, ZN => 
                           n9132);
   U11349 : AND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_16_port, ZN => 
                           n9120);
   U11350 : OAI211_X1 port map( C1 => n8106, C2 => n8368, A => n7698, B => 
                           n9119, ZN => n10539);
   U11351 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_16_port, ZN => 
                           n9119);
   U11352 : XNOR2_X1 port map( A => n9134, B => n9118, ZN => n9139);
   U11353 : INV_X1 port map( A => i_RD1_17_port, ZN => n9118);
   U11354 : NAND2_X1 port map( A1 => n9117, A2 => n9116, ZN => n9134);
   U11355 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_17_port, ZN => 
                           n9116);
   U11356 : NAND2_X1 port map( A1 => n10248, A2 => n8687, ZN => n9117);
   U11357 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_17_port, ZN => 
                           n9115);
   U11358 : INV_X1 port map( A => n9112, ZN => n9113);
   U11359 : AOI22_X1 port map( A1 => n9111, A2 => n10647, B1 => n9112, B2 => 
                           n10641, ZN => n9114);
   U11360 : INV_X1 port map( A => i_RD1_15_port, ZN => n10641);
   U11361 : NAND2_X1 port map( A1 => n9110, A2 => n9109, ZN => n9112);
   U11362 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_15_port, ZN => 
                           n9109);
   U11363 : NAND2_X1 port map( A1 => n10325, A2 => n8686, ZN => n9110);
   U11364 : NAND2_X1 port map( A1 => n9105, A2 => n8331, ZN => n9106);
   U11365 : NAND2_X1 port map( A1 => n7756, A2 => IRAM_ADDRESS_15_port, ZN => 
                           n9107);
   U11366 : INV_X1 port map( A => i_RD1_14_port, ZN => n10647);
   U11367 : INV_X1 port map( A => n9104, ZN => n9111);
   U11368 : NAND2_X1 port map( A1 => n9102, A2 => i_RD1_13_port, ZN => n9234);
   U11369 : NAND2_X1 port map( A1 => n9104, A2 => i_RD1_14_port, ZN => n9239);
   U11370 : OAI21_X1 port map( B1 => n10537, B2 => n8685, A => n9101, ZN => 
                           n9104);
   U11371 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => n9100, ZN => n9101);
   U11372 : INV_X1 port map( A => i_RD2_14_port, ZN => n9100);
   U11373 : NAND2_X1 port map( A1 => n9105, A2 => 
                           DECODEhw_i_tickcounter_14_port, ZN => n9098);
   U11374 : NAND2_X1 port map( A1 => n7756, A2 => IRAM_ADDRESS_14_port, ZN => 
                           n9099);
   U11375 : OAI21_X1 port map( B1 => n10535, B2 => n8685, A => n9096, ZN => 
                           n9102);
   U11376 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => n9095, ZN => n9096);
   U11377 : INV_X1 port map( A => i_RD2_13_port, ZN => n9095);
   U11378 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_13_port, ZN => 
                           n9094);
   U11379 : OAI211_X1 port map( C1 => n9249, C2 => n9088, A => n9235, B => 
                           n9233, ZN => n9089);
   U11380 : NAND2_X1 port map( A1 => n9097, A2 => i_RD1_12_port, ZN => n9233);
   U11381 : OAI21_X1 port map( B1 => n10382, B2 => n8685, A => n9087, ZN => 
                           n9097);
   U11382 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => n9086, ZN => n9087);
   U11383 : INV_X1 port map( A => i_RD2_12_port, ZN => n9086);
   U11384 : NAND2_X1 port map( A1 => n9105, A2 => 
                           DECODEhw_i_tickcounter_12_port, ZN => n9084);
   U11385 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_12_port, ZN => 
                           n9085);
   U11386 : NAND2_X1 port map( A1 => n9083, A2 => i_RD1_11_port, ZN => n9235);
   U11387 : AOI22_X1 port map( A1 => n9082, A2 => i_RD1_9_port, B1 => n9081, B2
                           => i_RD1_10_port, ZN => n9249);
   U11388 : NOR2_X1 port map( A1 => n9080, A2 => n9088, ZN => n9090);
   U11389 : OAI21_X1 port map( B1 => n9083, B2 => i_RD1_11_port, A => n9079, ZN
                           => n9088);
   U11390 : NAND2_X1 port map( A1 => n9078, A2 => n9077, ZN => n9079);
   U11391 : INV_X1 port map( A => n9081, ZN => n9078);
   U11392 : AOI21_X1 port map( B1 => n10533, B2 => n8687, A => n9076, ZN => 
                           n9081);
   U11393 : AND2_X1 port map( A1 => n8685, A2 => i_RD2_10_port, ZN => n9076);
   U11394 : NAND2_X1 port map( A1 => n9105, A2 => 
                           DECODEhw_i_tickcounter_10_port, ZN => n9074);
   U11395 : NAND2_X1 port map( A1 => n7699, A2 => IRAM_ADDRESS_10_port, ZN => 
                           n9075);
   U11396 : OAI21_X1 port map( B1 => n10391, B2 => n8685, A => n9073, ZN => 
                           n9083);
   U11397 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => n9072, ZN => n9073);
   U11398 : INV_X1 port map( A => i_RD2_11_port, ZN => n9072);
   U11399 : NAND2_X1 port map( A1 => n9105, A2 => n8330, ZN => n9070);
   U11400 : NAND2_X1 port map( A1 => n7756, A2 => IRAM_ADDRESS_11_port, ZN => 
                           n9071);
   U11401 : OAI22_X1 port map( A1 => n9082, A2 => i_RD1_9_port, B1 => n9069, B2
                           => i_RD1_8_port, ZN => n9080);
   U11402 : AOI21_X1 port map( B1 => n10438, B2 => n8687, A => n9068, ZN => 
                           n9082);
   U11403 : AND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_9_port, ZN => n9068
                           );
   U11404 : OAI211_X1 port map( C1 => n552, C2 => n9208, A => n9067, B => n9066
                           , ZN => n10438);
   U11405 : NAND2_X1 port map( A1 => n7756, A2 => IRAM_ADDRESS_9_port, ZN => 
                           n9067);
   U11406 : INV_X1 port map( A => n9062, ZN => n9063);
   U11407 : OAI211_X1 port map( C1 => n9061, C2 => n9060, A => n9059, B => 
                           n9236, ZN => n9062);
   U11408 : NAND2_X1 port map( A1 => n9069, A2 => i_RD1_8_port, ZN => n9236);
   U11409 : OAI21_X1 port map( B1 => n10531, B2 => n8685, A => n9058, ZN => 
                           n9069);
   U11410 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => n9057, ZN => n9058);
   U11411 : INV_X1 port map( A => i_RD2_8_port, ZN => n9057);
   U11412 : NAND2_X1 port map( A1 => n9105, A2 => DECODEhw_i_tickcounter_8_port
                           , ZN => n9055);
   U11413 : NAND2_X1 port map( A1 => n7756, A2 => IRAM_ADDRESS_8_port, ZN => 
                           n9056);
   U11414 : INV_X1 port map( A => n9054, ZN => n9061);
   U11415 : XNOR2_X1 port map( A => n9049, B => i_RD1_5_port, ZN => n9050);
   U11416 : AOI22_X1 port map( A1 => n9048, A2 => n9047, B1 => n9046, B2 => 
                           n9045, ZN => n9051);
   U11417 : INV_X1 port map( A => n9044, ZN => n9046);
   U11418 : INV_X1 port map( A => n9064, ZN => n9052);
   U11419 : NAND4_X1 port map( A1 => n9042, A2 => n9043, A3 => n9247, A4 => 
                           n9245, ZN => n9053);
   U11420 : NAND2_X1 port map( A1 => n9041, A2 => i_RD1_2_port, ZN => n9245);
   U11421 : INV_X1 port map( A => n9040, ZN => n9041);
   U11422 : NAND2_X1 port map( A1 => n9044, A2 => i_RD1_3_port, ZN => n9247);
   U11423 : AOI21_X1 port map( B1 => n10527, B2 => n8687, A => n9039, ZN => 
                           n9044);
   U11424 : AND2_X1 port map( A1 => n8685, A2 => i_RD2_3_port, ZN => n9039);
   U11425 : NAND2_X1 port map( A1 => n7699, A2 => IRAM_ADDRESS_3_port, ZN => 
                           n9038);
   U11426 : OAI21_X1 port map( B1 => n10518, B2 => n8685, A => n9033, ZN => 
                           n9034);
   U11427 : AOI21_X1 port map( B1 => n8685, B2 => n9032, A => i_RD1_0_port, ZN 
                           => n9033);
   U11428 : INV_X1 port map( A => i_RD2_0_port, ZN => n9032);
   U11429 : NAND2_X1 port map( A1 => n9105, A2 => n8328, ZN => n9030);
   U11430 : NAND2_X1 port map( A1 => n7756, A2 => IRAM_ADDRESS_0_port, ZN => 
                           n9031);
   U11431 : NAND2_X1 port map( A1 => n9035, A2 => n9246, ZN => n9043);
   U11432 : NAND2_X1 port map( A1 => n9105, A2 => DECODEhw_i_tickcounter_2_port
                           , ZN => n9025);
   U11433 : NAND2_X1 port map( A1 => n7696, A2 => IRAM_ADDRESS_2_port, ZN => 
                           n9026);
   U11434 : AND2_X1 port map( A1 => n9036, A2 => i_RD1_1_port, ZN => n9246);
   U11435 : NAND2_X1 port map( A1 => n8685, A2 => n9023, ZN => n9024);
   U11436 : INV_X1 port map( A => i_RD2_1_port, ZN => n9023);
   U11437 : NAND2_X1 port map( A1 => n7696, A2 => IRAM_ADDRESS_1_port, ZN => 
                           n9022);
   U11438 : NAND4_X1 port map( A1 => n9020, A2 => n9059, A3 => n9054, A4 => 
                           n9060, ZN => n9064);
   U11439 : NAND2_X1 port map( A1 => n9018, A2 => i_RD1_7_port, ZN => n9059);
   U11440 : AND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_7_port, ZN => n9017
                           );
   U11441 : NAND2_X1 port map( A1 => n7699, A2 => IRAM_ADDRESS_7_port, ZN => 
                           n9016);
   U11442 : AND2_X1 port map( A1 => n8685, A2 => i_RD2_6_port, ZN => n9014);
   U11443 : NAND2_X1 port map( A1 => n9105, A2 => DECODEhw_i_tickcounter_6_port
                           , ZN => n9012);
   U11444 : NAND2_X1 port map( A1 => n7699, A2 => IRAM_ADDRESS_6_port, ZN => 
                           n9013);
   U11445 : NAND2_X1 port map( A1 => n9011, A2 => i_RD1_4_port, ZN => n9244);
   U11446 : INV_X1 port map( A => n9048, ZN => n9011);
   U11447 : AOI21_X1 port map( B1 => n10514, B2 => n8687, A => n9010, ZN => 
                           n9048);
   U11448 : NOR2_X1 port map( A1 => i_RD2_4_port, A2 => n8686, ZN => n9010);
   U11449 : NAND2_X1 port map( A1 => n9105, A2 => DECODEhw_i_tickcounter_4_port
                           , ZN => n9006);
   U11450 : INV_X1 port map( A => i_RD1_5_port, ZN => n10678);
   U11451 : NAND2_X1 port map( A1 => n9003, A2 => n9002, ZN => n9049);
   U11452 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_5_port, ZN => 
                           n9002);
   U11453 : NAND2_X1 port map( A1 => n10464, A2 => n8687, ZN => n9003);
   U11454 : NAND2_X1 port map( A1 => n7696, A2 => IRAM_ADDRESS_5_port, ZN => 
                           n9001);
   U11455 : OAI21_X1 port map( B1 => n9215, B2 => n8999, A => n9230, ZN => 
                           n9231);
   U11456 : NAND2_X1 port map( A1 => n9215, A2 => n8998, ZN => n9230);
   U11457 : AOI21_X1 port map( B1 => n8329, B2 => n8997, A => CU_I_CW_ID_22, ZN
                           => n8998);
   U11458 : AND2_X1 port map( A1 => IR_3_port, A2 => IR_5_port, ZN => n10741);
   U11459 : NAND2_X1 port map( A1 => n10781, A2 => n10767, ZN => n10789);
   U11460 : NAND2_X1 port map( A1 => n8428, A2 => IR_1_port, ZN => n10767);
   U11461 : NAND2_X1 port map( A1 => n8315, A2 => IR_2_port, ZN => n10781);
   U11462 : NAND2_X1 port map( A1 => n8996, A2 => i_RD1_30_port, ZN => n8999);
   U11463 : INV_X1 port map( A => n9205, ZN => n8996);
   U11464 : NAND2_X1 port map( A1 => n8995, A2 => n8994, ZN => n9205);
   U11465 : NAND2_X1 port map( A1 => n8685, A2 => i_RD2_30_port, ZN => n8994);
   U11466 : NAND2_X1 port map( A1 => n9812, A2 => n8687, ZN => n8995);
   U11467 : NAND2_X1 port map( A1 => n7757, A2 => IRAM_ADDRESS_30_port, ZN => 
                           n8993);
   U11468 : NAND2_X1 port map( A1 => n8991, A2 => n8990, ZN => n8992);
   U11469 : INV_X1 port map( A => i_RD1_31_port, ZN => n8990);
   U11470 : INV_X1 port map( A => n8989, ZN => n8991);
   U11471 : NAND2_X1 port map( A1 => n8989, A2 => i_RD1_31_port, ZN => n9223);
   U11472 : AOI21_X1 port map( B1 => n9790, B2 => n8686, A => n8988, ZN => 
                           n8989);
   U11473 : AND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_31_port, ZN => 
                           n8988);
   U11474 : NAND2_X1 port map( A1 => n7699, A2 => IRAM_ADDRESS_31_port, ZN => 
                           n8987);
   U11475 : NAND2_X1 port map( A1 => n8308, A2 => n8704, ZN => n10720);
   U11476 : NOR2_X1 port map( A1 => n194, A2 => CU_I_CW_ID_22, ZN => n8986);
   U11477 : NAND2_X1 port map( A1 => n10543, A2 => n9275, ZN => n8705);
   U11478 : NAND2_X1 port map( A1 => n10843, A2 => n171, ZN => n10519);
   U11479 : NOR2_X1 port map( A1 => n10756, A2 => n8984, ZN => n10843);
   U11480 : AND2_X1 port map( A1 => n8454, A2 => n8255, ZN => n9271);
   U11481 : NOR2_X1 port map( A1 => n9264, A2 => n8501, ZN => n10826);
   U11482 : INV_X1 port map( A => n10707, ZN => n9264);
   U11483 : NOR3_X1 port map( A1 => n9810, A2 => n9809, A3 => n9808, ZN => 
                           n9811);
   U11484 : OAI22_X1 port map( A1 => n9916, A2 => n10376, B1 => n9849, B2 => 
                           n10460, ZN => n9808);
   U11485 : OAI22_X1 port map( A1 => n9946, A2 => n10462, B1 => n9807, B2 => 
                           n10507, ZN => n9809);
   U11486 : OAI211_X1 port map( C1 => n8311, C2 => n10444, A => n9806, B => 
                           n9805, ZN => n9810);
   U11487 : AOI22_X1 port map( A1 => n9829, A2 => n10461, B1 => n9992, B2 => 
                           n10503, ZN => n9805);
   U11488 : AOI22_X1 port map( A1 => n9843, A2 => n10510, B1 => n9949, B2 => 
                           n10502, ZN => n9806);
   U11489 : OAI22_X1 port map( A1 => n7781, A2 => n9800, B1 => n9799, B2 => 
                           n10115, ZN => n9801);
   U11490 : NOR2_X1 port map( A1 => n9798, A2 => n10182, ZN => n9800);
   U11491 : AOI22_X1 port map( A1 => n7769, A2 => n9983, B1 => n9920, B2 => 
                           n7792, ZN => n9802);
   U11492 : INV_X1 port map( A => n9980, ZN => n9920);
   U11493 : OAI211_X1 port map( C1 => n10062, C2 => n10286, A => n10113, B => 
                           n10055, ZN => n9803);
   U11494 : NAND2_X1 port map( A1 => n9797, A2 => n10286, ZN => n10055);
   U11495 : AOI22_X1 port map( A1 => n9796, A2 => n10231, B1 => n9795, B2 => 
                           n7785, ZN => n9804);
   U11496 : AOI21_X1 port map( B1 => n9798, B2 => n12081, A => n9601, ZN => 
                           n9796);
   U11497 : NOR2_X1 port map( A1 => n9603, A2 => n12081, ZN => n9601);
   U11498 : INV_X1 port map( A => n10465, ZN => n10468);
   U11499 : NOR3_X1 port map( A1 => n9788, A2 => n9787, A3 => n9786, ZN => 
                           n9789);
   U11500 : OAI22_X1 port map( A1 => n9849, A2 => n10388, B1 => n10031, B2 => 
                           n10444, ZN => n9786);
   U11501 : NAND2_X1 port map( A1 => n9448, A2 => n9428, ZN => n10444);
   U11502 : NOR2_X1 port map( A1 => n8099, A2 => n7800, ZN => n9428);
   U11503 : INV_X1 port map( A => n9992, ZN => n10031);
   U11504 : NAND4_X1 port map( A1 => n9785, A2 => n9784, A3 => n9783, A4 => 
                           n9782, ZN => n9992);
   U11505 : NAND2_X1 port map( A1 => n9844, A2 => n10026, ZN => n9782);
   U11506 : OAI21_X1 port map( B1 => n10277, B2 => n10869, A => n10180, ZN => 
                           n9844);
   U11507 : NAND2_X1 port map( A1 => n9781, A2 => n10286, ZN => n10025);
   U11508 : OAI211_X1 port map( C1 => n9780, C2 => n9779, A => n9778, B => 
                           n10115, ZN => n10023);
   U11509 : NAND2_X1 port map( A1 => n9629, A2 => n9386, ZN => n9779);
   U11510 : NAND2_X1 port map( A1 => n7800, A2 => n10010, ZN => n9386);
   U11511 : AOI22_X1 port map( A1 => n10012, A2 => n9983, B1 => n10231, B2 => 
                           n10027, ZN => n9784);
   U11512 : NOR2_X1 port map( A1 => n9777, A2 => n9776, ZN => n9785);
   U11513 : NOR2_X1 port map( A1 => n9778, A2 => n10277, ZN => n9776);
   U11514 : INV_X1 port map( A => n10240, ZN => n10277);
   U11515 : OAI22_X1 port map( A1 => n9775, A2 => n9774, B1 => n8094, B2 => 
                           n12091, ZN => n9777);
   U11516 : INV_X1 port map( A => n10282, ZN => n9775);
   U11517 : NOR2_X1 port map( A1 => n10182, A2 => n12087, ZN => n10282);
   U11518 : AOI21_X1 port map( B1 => n9845, B2 => n9773, A => n9772, ZN => 
                           n9849);
   U11519 : OAI211_X1 port map( C1 => n9771, C2 => n9770, A => n9769, B => 
                           n9768, ZN => n9772);
   U11520 : AOI22_X1 port map( A1 => n9767, A2 => n10111, B1 => n10231, B2 => 
                           n10116, ZN => n9768);
   U11521 : AND2_X1 port map( A1 => n9611, A2 => n9610, ZN => n10116);
   U11522 : OR2_X1 port map( A1 => n10473, A2 => n8681, ZN => n9610);
   U11523 : NAND2_X1 port map( A1 => n9409, A2 => n9408, ZN => n10111);
   U11524 : NAND2_X1 port map( A1 => n8681, A2 => n10122, ZN => n9408);
   U11525 : NAND2_X1 port map( A1 => n9669, A2 => i_ALU_OP_2_port, ZN => n9409)
                           ;
   U11526 : AOI22_X1 port map( A1 => n9766, A2 => n10122, B1 => n10232, B2 => 
                           n10108, ZN => n9769);
   U11527 : OAI21_X1 port map( B1 => n9780, B2 => n10109, A => n9846, ZN => 
                           n10108);
   U11528 : NAND2_X1 port map( A1 => n10110, A2 => n9765, ZN => n9846);
   U11529 : NAND2_X1 port map( A1 => n9611, A2 => n9410, ZN => n10109);
   U11530 : NAND2_X1 port map( A1 => n7795, A2 => n7800, ZN => n9410);
   U11531 : OR2_X1 port map( A1 => n9669, A2 => n7800, ZN => n9611);
   U11532 : INV_X1 port map( A => n10110, ZN => n9770);
   U11533 : NAND2_X1 port map( A1 => n9845, A2 => n12071, ZN => n9421);
   U11534 : NAND2_X1 port map( A1 => n10473, A2 => n12089, ZN => n9422);
   U11535 : INV_X1 port map( A => n9764, ZN => n9773);
   U11536 : OAI22_X1 port map( A1 => n9916, A2 => n10479, B1 => n9807, B2 => 
                           n10505, ZN => n9787);
   U11537 : NAND2_X1 port map( A1 => n9396, A2 => n9552, ZN => n10505);
   U11538 : NOR2_X1 port map( A1 => n9556, A2 => n7796, ZN => n9396);
   U11539 : AOI211_X1 port map( C1 => n10232, C2 => n10062, A => n9763, B => 
                           n9762, ZN => n9807);
   U11540 : OAI21_X1 port map( B1 => n9764, B2 => n9761, A => n9760, ZN => 
                           n9762);
   U11541 : AOI22_X1 port map( A1 => n9766, A2 => n7769, B1 => n10113, B2 => 
                           n9795, ZN => n9760);
   U11542 : NAND2_X1 port map( A1 => n9759, A2 => n9758, ZN => n9795);
   U11543 : NAND2_X1 port map( A1 => n9799, A2 => n12088, ZN => n9758);
   U11544 : OAI22_X1 port map( A1 => n9771, A2 => n9798, B1 => n9797, B2 => 
                           n10184, ZN => n9763);
   U11545 : OAI21_X1 port map( B1 => n10059, B2 => n9780, A => n9759, ZN => 
                           n10062);
   U11546 : NAND2_X1 port map( A1 => n9757, A2 => n9765, ZN => n9759);
   U11547 : INV_X1 port map( A => n9798, ZN => n9757);
   U11548 : NOR2_X1 port map( A1 => n9761, A2 => n12073, ZN => n9375);
   U11549 : NAND2_X1 port map( A1 => n9604, A2 => n9378, ZN => n10059);
   U11550 : NAND2_X1 port map( A1 => n7800, A2 => n8553, ZN => n9378);
   U11551 : NAND2_X1 port map( A1 => n7789, A2 => n8681, ZN => n9604);
   U11552 : NAND3_X1 port map( A1 => n8486, A2 => n9552, A3 => n8167, ZN => 
                           n10479);
   U11553 : AOI211_X1 port map( C1 => n10232, C2 => n10190, A => n9756, B => 
                           n9755, ZN => n9916);
   U11554 : OAI21_X1 port map( B1 => n9764, B2 => n10181, A => n9754, ZN => 
                           n9755);
   U11555 : OAI21_X1 port map( B1 => n9664, B2 => n8681, A => n9354, ZN => 
                           n10185);
   U11556 : NAND2_X1 port map( A1 => n8681, A2 => n10197, ZN => n9354);
   U11557 : OAI22_X1 port map( A1 => n9771, A2 => n9752, B1 => n9921, B2 => 
                           n10184, ZN => n9756);
   U11558 : INV_X1 port map( A => n9917, ZN => n9752);
   U11559 : OAI21_X1 port map( B1 => n9780, B2 => n10183, A => n9753, ZN => 
                           n10190);
   U11560 : NAND2_X1 port map( A1 => n9917, A2 => n9765, ZN => n9753);
   U11561 : NAND2_X1 port map( A1 => n9919, A2 => n12071, ZN => n9352);
   U11562 : NAND2_X1 port map( A1 => n9562, A2 => n12089, ZN => n9353);
   U11563 : NAND2_X1 port map( A1 => n9540, A2 => n9349, ZN => n10183);
   U11564 : NAND2_X1 port map( A1 => n7800, A2 => n10197, ZN => n9349);
   U11565 : OR2_X1 port map( A1 => n9664, A2 => n7800, ZN => n9540);
   U11566 : OAI211_X1 port map( C1 => n9946, C2 => n10442, A => n9751, B => 
                           n9750, ZN => n9788);
   U11567 : AOI22_X1 port map( A1 => n10476, A2 => n9749, B1 => n9829, B2 => 
                           n10499, ZN => n9750);
   U11568 : INV_X1 port map( A => n10460, ZN => n10499);
   U11569 : NAND2_X1 port map( A1 => n9446, A2 => n9555, ZN => n10460);
   U11570 : AOI21_X1 port map( B1 => n8555, B2 => i_ALU_OP_2_port, A => n9399, 
                           ZN => n10089);
   U11571 : NOR2_X1 port map( A1 => n10082, A2 => n7800, ZN => n9399);
   U11572 : OAI21_X1 port map( B1 => n9747, B2 => n9780, A => n9821, ZN => 
                           n10086);
   U11573 : NAND2_X1 port map( A1 => n10090, A2 => n9765, ZN => n9821);
   U11574 : NAND2_X1 port map( A1 => n9816, A2 => n12071, ZN => n9403);
   U11575 : NAND2_X1 port map( A1 => n7818, A2 => n12089, ZN => n9404);
   U11576 : NAND2_X1 port map( A1 => n9619, A2 => n9405, ZN => n9747);
   U11577 : NAND2_X1 port map( A1 => n7800, A2 => n8556, ZN => n9405);
   U11578 : NAND2_X1 port map( A1 => n8555, A2 => n8681, ZN => n9619);
   U11579 : OAI21_X1 port map( B1 => n7800, B2 => n9817, A => n9406, ZN => 
                           n9820);
   U11580 : NAND2_X1 port map( A1 => n10082, A2 => n7800, ZN => n9406);
   U11581 : OAI211_X1 port map( C1 => n7780, C2 => n10010, A => n9746, B => 
                           n9745, ZN => n9749);
   U11582 : AOI22_X1 port map( A1 => n10113, A2 => n9744, B1 => n10231, B2 => 
                           n9743, ZN => n9745);
   U11583 : INV_X1 port map( A => n9781, ZN => n9743);
   U11584 : OR2_X1 port map( A1 => n10261, A2 => i_ALU_OP_2_port, ZN => n9629);
   U11585 : INV_X1 port map( A => n9778, ZN => n9744);
   U11586 : NAND2_X1 port map( A1 => n10028, A2 => n9765, ZN => n9778);
   U11587 : INV_X1 port map( A => n9774, ZN => n10028);
   U11588 : NOR2_X1 port map( A1 => n10024, A2 => n12073, ZN => n9387);
   U11589 : AOI22_X1 port map( A1 => n9767, A2 => n10026, B1 => n10229, B2 => 
                           n9742, ZN => n9746);
   U11590 : NAND2_X1 port map( A1 => n9383, A2 => n9382, ZN => n10026);
   U11591 : NAND2_X1 port map( A1 => n8681, A2 => n10012, ZN => n9382);
   U11592 : NAND2_X1 port map( A1 => n10261, A2 => n7800, ZN => n9383);
   U11593 : NOR2_X1 port map( A1 => n10284, A2 => n10869, ZN => n9767);
   U11594 : NAND2_X1 port map( A1 => n9448, A2 => n9445, ZN => n10507);
   U11595 : NOR2_X1 port map( A1 => n8099, A2 => n8681, ZN => n9445);
   U11596 : AOI22_X1 port map( A1 => n9843, A2 => n10498, B1 => n9949, B2 => 
                           n10495, ZN => n9751);
   U11597 : INV_X1 port map( A => n9924, ZN => n9949);
   U11598 : AOI21_X1 port map( B1 => n10231, B2 => n9950, A => n9741, ZN => 
                           n9924);
   U11599 : OAI211_X1 port map( C1 => n9740, C2 => n10182, A => n9739, B => 
                           n9738, ZN => n9741);
   U11600 : NAND2_X1 port map( A1 => n9955, A2 => n10113, ZN => n9738);
   U11601 : NAND2_X1 port map( A1 => n9737, A2 => n9736, ZN => n9955);
   U11602 : NAND2_X1 port map( A1 => n10228, A2 => n12088, ZN => n9736);
   U11603 : NAND2_X1 port map( A1 => n9336, A2 => n9335, ZN => n10228);
   U11604 : NAND2_X1 port map( A1 => n8681, A2 => n7767, ZN => n9335);
   U11605 : NAND2_X1 port map( A1 => n8093, A2 => n7800, ZN => n9336);
   U11606 : AOI22_X1 port map( A1 => n9938, A2 => n9748, B1 => n9735, B2 => 
                           n9953, ZN => n9739);
   U11607 : AOI21_X1 port map( B1 => n10286, B2 => n9734, A => n10239, ZN => 
                           n9740);
   U11608 : OAI21_X1 port map( B1 => n8551, B2 => n8681, A => n9951, ZN => 
                           n9734);
   U11609 : NAND2_X1 port map( A1 => n8681, A2 => n9938, ZN => n9951);
   U11610 : OR2_X1 port map( A1 => n10239, A2 => n10234, ZN => n9950);
   U11611 : NOR2_X1 port map( A1 => n9733, A2 => n9732, ZN => n10234);
   U11612 : NOR2_X1 port map( A1 => n10487, A2 => n8681, ZN => n9732);
   U11613 : OAI21_X1 port map( B1 => n8093, B2 => n7800, A => n10286, ZN => 
                           n9733);
   U11614 : NAND2_X1 port map( A1 => n9737, A2 => n9731, ZN => n10239);
   U11615 : NAND2_X1 port map( A1 => n9730, A2 => n12089, ZN => n9731);
   U11616 : NAND2_X1 port map( A1 => n9953, A2 => n9765, ZN => n9737);
   U11617 : NOR2_X1 port map( A1 => n9944, A2 => n12073, ZN => n9340);
   U11618 : INV_X1 port map( A => n8099, ZN => n9561);
   U11619 : INV_X1 port map( A => n9448, ZN => n9427);
   U11620 : INV_X1 port map( A => n9895, ZN => n9843);
   U11621 : AOI21_X1 port map( B1 => n10231, B2 => n9729, A => n9728, ZN => 
                           n9895);
   U11622 : OAI211_X1 port map( C1 => n9727, C2 => n10182, A => n9726, B => 
                           n9725, ZN => n9728);
   U11623 : NAND2_X1 port map( A1 => n9893, A2 => n10113, ZN => n9725);
   U11624 : OAI21_X1 port map( B1 => n10164, B2 => n10869, A => n9724, ZN => 
                           n9893);
   U11625 : AOI21_X1 port map( B1 => n7800, B2 => n8090, A => n9363, ZN => 
                           n10164);
   U11626 : NOR2_X1 port map( A1 => n7800, A2 => n10143, ZN => n9363);
   U11627 : AOI22_X1 port map( A1 => n7797, A2 => n9748, B1 => n9735, B2 => 
                           n9885, ZN => n9726);
   U11628 : INV_X1 port map( A => n9771, ZN => n9735);
   U11629 : AOI21_X1 port map( B1 => n10286, B2 => n9723, A => n10167, ZN => 
                           n9727);
   U11630 : OAI21_X1 port map( B1 => n8681, B2 => n10143, A => n9722, ZN => 
                           n9723);
   U11631 : INV_X1 port map( A => n9886, ZN => n9722);
   U11632 : NOR2_X1 port map( A1 => n7800, A2 => n9874, ZN => n9886);
   U11633 : INV_X1 port map( A => n10115, ZN => n10286);
   U11634 : INV_X1 port map( A => n9890, ZN => n9729);
   U11635 : NOR2_X1 port map( A1 => n10162, A2 => n10167, ZN => n9890);
   U11636 : OAI21_X1 port map( B1 => n10160, B2 => n9780, A => n9724, ZN => 
                           n10167);
   U11637 : NAND2_X1 port map( A1 => n9885, A2 => n9765, ZN => n9724);
   U11638 : NOR2_X1 port map( A1 => n9874, A2 => n12073, ZN => n9365);
   U11639 : AOI211_X1 port map( C1 => n8491, C2 => i_ALU_OP_2_port, A => n10115
                           , B => n9720, ZN => n10162);
   U11640 : NOR2_X1 port map( A1 => n8090, A2 => n7800, ZN => n9720);
   U11641 : NAND2_X1 port map( A1 => n9347, A2 => n9551, ZN => n10442);
   U11642 : NOR2_X1 port map( A1 => n9555, A2 => n7796, ZN => n9347);
   U11643 : OAI21_X1 port map( B1 => n9764, B2 => n9979, A => n9717, ZN => 
                           n9718);
   U11644 : AOI22_X1 port map( A1 => n9766, A2 => n7772, B1 => n10113, B2 => 
                           n9978, ZN => n9717);
   U11645 : NAND2_X1 port map( A1 => n9716, A2 => n9715, ZN => n9978);
   U11646 : NAND2_X1 port map( A1 => n9987, A2 => n12088, ZN => n9715);
   U11647 : INV_X1 port map( A => n10284, ZN => n10113);
   U11648 : NAND2_X1 port map( A1 => n7828, A2 => n8015, ZN => n10284);
   U11649 : NOR2_X1 port map( A1 => n10180, A2 => n8681, ZN => n9766);
   U11650 : AOI21_X1 port map( B1 => n7781, B2 => n8681, A => n9748, ZN => 
                           n9764);
   U11651 : INV_X1 port map( A => n9983, ZN => n9714);
   U11652 : OR2_X1 port map( A1 => n10182, A2 => n10115, ZN => n10180);
   U11653 : OAI22_X1 port map( A1 => n9771, A2 => n9713, B1 => n10275, B2 => 
                           n10184, ZN => n9719);
   U11654 : NAND2_X1 port map( A1 => n9438, A2 => n9437, ZN => n10275);
   U11655 : OR2_X1 port map( A1 => n9533, A2 => n8681, ZN => n9437);
   U11656 : INV_X1 port map( A => n10285, ZN => n9713);
   U11657 : AND2_X1 port map( A1 => n9980, A2 => n12090, ZN => n9771);
   U11658 : NAND2_X1 port map( A1 => n10229, A2 => n8300, ZN => n9980);
   U11659 : OAI21_X1 port map( B1 => n10291, B2 => n9780, A => n9716, ZN => 
                           n10276);
   U11660 : NAND2_X1 port map( A1 => n10285, A2 => n9765, ZN => n9716);
   U11661 : INV_X1 port map( A => n12090, ZN => n9765);
   U11662 : INV_X1 port map( A => n12088, ZN => n10869);
   U11663 : NAND2_X1 port map( A1 => n9436, A2 => n9435, ZN => n10285);
   U11664 : INV_X1 port map( A => n12072, ZN => n9435);
   U11665 : NAND2_X1 port map( A1 => n9533, A2 => n12089, ZN => n9436);
   U11666 : INV_X1 port map( A => n12089, ZN => n9780);
   U11667 : NAND2_X1 port map( A1 => n9438, A2 => n9432, ZN => n10291);
   U11668 : NAND2_X1 port map( A1 => n7800, A2 => n8557, ZN => n9432);
   U11669 : NAND2_X1 port map( A1 => n8559, A2 => n8681, ZN => n9438);
   U11670 : NAND2_X1 port map( A1 => n9337, A2 => n8263, ZN => n10182);
   U11671 : INV_X1 port map( A => n8015, ZN => n9337);
   U11672 : NOR2_X1 port map( A1 => n9527, A2 => i_ALU_OP_0_port, ZN => n9532);
   U11673 : NAND2_X1 port map( A1 => i_ALU_OP_1_port, A2 => n10870, ZN => n9527
                           );
   U11674 : INV_X1 port map( A => n12074, ZN => n10870);
   U11675 : NAND2_X1 port map( A1 => n9529, A2 => n9528, ZN => n10465);
   U11676 : AOI21_X1 port map( B1 => i_ALU_OP_3_port, B2 => n12088, A => n8412,
                           ZN => n9528);
   U11677 : NAND2_X1 port map( A1 => n9531, A2 => n8319, ZN => n9529);
   U11678 : XNOR2_X1 port map( A => i_ALU_OP_2_port, B => n8385, ZN => n9531);
   U11679 : OAI22_X1 port map( A1 => n9814, A2 => n9855, B1 => n9711, B2 => 
                           n9817, ZN => n9793);
   U11680 : NAND2_X1 port map( A1 => n9710, A2 => n9845, ZN => n9855);
   U11681 : INV_X1 port map( A => n9841, ZN => n9710);
   U11682 : INV_X1 port map( A => n9842, ZN => n9838);
   U11683 : NAND2_X1 port map( A1 => n9709, A2 => n10450, ZN => n9842);
   U11684 : INV_X1 port map( A => n9708, ZN => n9709);
   U11685 : NAND2_X1 port map( A1 => n9708, A2 => n10450, ZN => n9854);
   U11686 : AOI21_X1 port map( B1 => n9707, B2 => n9865, A => n9706, ZN => 
                           n9708);
   U11687 : INV_X1 port map( A => n9866, ZN => n9706);
   U11688 : NAND2_X1 port map( A1 => n9705, A2 => n9874, ZN => n9866);
   U11689 : NAND2_X1 port map( A1 => n9704, A2 => n7797, ZN => n9865);
   U11690 : INV_X1 port map( A => n9705, ZN => n9704);
   U11691 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n537, B => 
                           i_ALU_OP_2_port, ZN => n9705);
   U11692 : OAI21_X1 port map( B1 => n9868, B2 => n9703, A => n9867, ZN => 
                           n9707);
   U11693 : OAI21_X1 port map( B1 => n9903, B2 => n9905, A => n9871, ZN => 
                           n9867);
   U11694 : NAND2_X1 port map( A1 => n9935, A2 => n9869, ZN => n9903);
   U11695 : OR2_X1 port map( A1 => n9937, A2 => n9964, ZN => n9935);
   U11696 : NAND2_X1 port map( A1 => n9701, A2 => n9979, ZN => n9964);
   U11697 : INV_X1 port map( A => n9700, ZN => n9701);
   U11698 : NAND2_X1 port map( A1 => n9869, A2 => n9699, ZN => n9937);
   U11699 : NAND2_X1 port map( A1 => n9698, A2 => n9944, ZN => n9869);
   U11700 : INV_X1 port map( A => n9697, ZN => n9698);
   U11701 : NAND2_X1 port map( A1 => n9702, A2 => n9919, ZN => n9871);
   U11702 : XNOR2_X1 port map( A => n9909, B => n8681, ZN => n9702);
   U11703 : INV_X1 port map( A => n9965, ZN => n9932);
   U11704 : AND2_X1 port map( A1 => n9700, A2 => n10281, ZN => n9965);
   U11705 : XNOR2_X1 port map( A => n9969, B => n8681, ZN => n9700);
   U11706 : INV_X1 port map( A => n9870, ZN => n9699);
   U11707 : AND2_X1 port map( A1 => n9697, A2 => n9938, ZN => n9870);
   U11708 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n639, B => n8681, ZN => 
                           n9697);
   U11709 : AND2_X1 port map( A1 => n9696, A2 => n10010, ZN => n10002);
   U11710 : NAND2_X1 port map( A1 => n9695, A2 => n10012, ZN => n10001);
   U11711 : INV_X1 port map( A => n9696, ZN => n9695);
   U11712 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n741, B => 
                           i_ALU_OP_2_port, ZN => n9696);
   U11713 : OAI21_X1 port map( B1 => n10039, B2 => n10038, A => n9694, ZN => 
                           n10007);
   U11714 : XNOR2_X1 port map( A => n9693, B => n8553, ZN => n10038);
   U11715 : NAND2_X1 port map( A1 => n10073, A2 => n10005, ZN => n10039);
   U11716 : OR2_X1 port map( A1 => n10075, A2 => n10104, ZN => n10073);
   U11717 : NAND2_X1 port map( A1 => n9692, A2 => n10123, ZN => n10104);
   U11718 : NAND2_X1 port map( A1 => n10005, A2 => n9691, ZN => n10075);
   U11719 : NAND2_X1 port map( A1 => n9690, A2 => n8556, ZN => n10005);
   U11720 : NAND2_X1 port map( A1 => n9689, A2 => n7769, ZN => n9694);
   U11721 : INV_X1 port map( A => n9693, ZN => n9689);
   U11722 : XNOR2_X1 port map( A => n10046, B => i_ALU_OP_2_port, ZN => n9693);
   U11723 : NAND2_X1 port map( A1 => n9691, A2 => n10103, ZN => n10006);
   U11724 : NAND2_X1 port map( A1 => n9688, A2 => n10122, ZN => n10103);
   U11725 : INV_X1 port map( A => n9692, ZN => n9688);
   U11726 : XNOR2_X1 port map( A => n10124, B => i_ALU_OP_2_port, ZN => n9692);
   U11727 : NAND2_X1 port map( A1 => n9687, A2 => n10082, ZN => n9691);
   U11728 : INV_X1 port map( A => n9690, ZN => n9687);
   U11729 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n843, B => 
                           i_ALU_OP_2_port, ZN => n9690);
   U11730 : NAND2_X1 port map( A1 => n9686, A2 => n10137, ZN => n10004);
   U11731 : NAND2_X1 port map( A1 => n9685, A2 => n8552, ZN => n10137);
   U11732 : INV_X1 port map( A => n9684, ZN => n9685);
   U11733 : OAI211_X1 port map( C1 => n10139, C2 => n10138, A => n10136, B => 
                           n10142, ZN => n9686);
   U11734 : NAND2_X1 port map( A1 => n10175, A2 => n9683, ZN => n10142);
   U11735 : OR2_X1 port map( A1 => n10174, A2 => n9682, ZN => n10175);
   U11736 : NAND2_X1 port map( A1 => n10216, A2 => n10303, ZN => n10213);
   U11737 : AND2_X1 port map( A1 => n9680, A2 => n8557, ZN => n10303);
   U11738 : NAND2_X1 port map( A1 => n9684, A2 => n10143, ZN => n10136);
   U11739 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n945, B => 
                           i_ALU_OP_2_port, ZN => n9684);
   U11740 : NAND2_X1 port map( A1 => n10204, A2 => n9683, ZN => n10138);
   U11741 : NAND2_X1 port map( A1 => n10203, A2 => n10205, ZN => n10204);
   U11742 : INV_X1 port map( A => n9682, ZN => n10205);
   U11743 : XNOR2_X1 port map( A => n10198, B => n8681, ZN => n9679);
   U11744 : NAND2_X1 port map( A1 => n10215, A2 => n9678, ZN => n10203);
   U11745 : NAND2_X1 port map( A1 => n9681, A2 => n7767, ZN => n9678);
   U11746 : NAND2_X1 port map( A1 => n10216, A2 => n10304, ZN => n10215);
   U11747 : XNOR2_X1 port map( A => n10313, B => i_ALU_OP_2_port, ZN => n9680);
   U11748 : XNOR2_X1 port map( A => n9681, B => n8551, ZN => n10216);
   U11749 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1047, B => n8300, ZN =>
                           n9681);
   U11750 : OAI21_X1 port map( B1 => n9677, B2 => n9676, A => n10252, ZN => 
                           n10139);
   U11751 : NAND2_X1 port map( A1 => n9675, A2 => n10261, ZN => n10252);
   U11752 : INV_X1 port map( A => n8554, ZN => n10261);
   U11753 : INV_X1 port map( A => n9674, ZN => n9675);
   U11754 : NAND2_X1 port map( A1 => n10251, A2 => n10257, ZN => n9676);
   U11755 : NAND2_X1 port map( A1 => n9673, A2 => n8494, ZN => n10257);
   U11756 : INV_X1 port map( A => n9672, ZN => n9673);
   U11757 : NAND2_X1 port map( A1 => n9674, A2 => n8554, ZN => n10251);
   U11758 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1149, B => 
                           i_ALU_OP_2_port, ZN => n9674);
   U11759 : AOI21_X1 port map( B1 => n10249, B2 => n9671, A => n10265, ZN => 
                           n9677);
   U11760 : NAND2_X1 port map( A1 => n10368, A2 => n10258, ZN => n10265);
   U11761 : NAND2_X1 port map( A1 => n9672, A2 => n10377, ZN => n10258);
   U11762 : XNOR2_X1 port map( A => n10379, B => n8681, ZN => n9672);
   U11763 : NAND2_X1 port map( A1 => n10347, A2 => n10255, ZN => n10368);
   U11764 : OR2_X1 port map( A1 => n10349, A2 => n10350, ZN => n10347);
   U11765 : AND2_X1 port map( A1 => n9670, A2 => n9669, ZN => n10350);
   U11766 : NOR2_X1 port map( A1 => n10349, A2 => n10343, ZN => n9671);
   U11767 : XNOR2_X1 port map( A => n10337, B => n8300, ZN => n9670);
   U11768 : NAND2_X1 port map( A1 => n10255, A2 => n10253, ZN => n10349);
   U11769 : NAND2_X1 port map( A1 => n9668, A2 => n10351, ZN => n10253);
   U11770 : INV_X1 port map( A => n8555, ZN => n10351);
   U11771 : INV_X1 port map( A => n9667, ZN => n9668);
   U11772 : NAND2_X1 port map( A1 => n9667, A2 => n8555, ZN => n10255);
   U11773 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1251, B => 
                           i_ALU_OP_2_port, ZN => n9667);
   U11774 : AOI21_X1 port map( B1 => n10384, B2 => n9666, A => n9665, ZN => 
                           n10249);
   U11775 : NOR2_X1 port map( A1 => n10383, A2 => n8090, ZN => n9665);
   U11776 : NAND2_X1 port map( A1 => n10383, A2 => n8090, ZN => n9666);
   U11777 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1353, B => n8300, ZN =>
                           n10383);
   U11778 : XNOR2_X1 port map( A => n10419, B => n8300, ZN => n10415);
   U11779 : NAND2_X1 port map( A1 => n9663, A2 => n10445, ZN => n10448);
   U11780 : INV_X1 port map( A => n8559, ZN => n10445);
   U11781 : INV_X1 port map( A => n10447, ZN => n9663);
   U11782 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1455, B => n8300, ZN =>
                           n10392);
   U11783 : AND2_X1 port map( A1 => n10447, A2 => n8559, ZN => n10449);
   U11784 : XNOR2_X1 port map( A => n10446, B => i_ALU_OP_2_port, ZN => n10447)
                           ;
   U11785 : NAND2_X1 port map( A1 => n9662, A2 => n9661, ZN => n10451);
   U11786 : NAND2_X1 port map( A1 => n9660, A2 => n9659, ZN => n9661);
   U11787 : INV_X1 port map( A => n9658, ZN => n9660);
   U11788 : NAND4_X1 port map( A1 => n9654, A2 => n9653, A3 => n9652, A4 => 
                           n10472, ZN => n9655);
   U11789 : OR2_X1 port map( A1 => n10470, A2 => n10473, ZN => n10472);
   U11790 : AOI21_X1 port map( B1 => n9600, B2 => n9599, A => n9598, ZN => 
                           n9654);
   U11791 : NOR2_X1 port map( A1 => n9597, A2 => n8016, ZN => n9598);
   U11792 : AND2_X1 port map( A1 => n9595, A2 => n9594, ZN => n9599);
   U11793 : NAND2_X1 port map( A1 => n9597, A2 => n8016, ZN => n9594);
   U11794 : XNOR2_X1 port map( A => n8263, B => n8300, ZN => n9597);
   U11795 : NAND2_X1 port map( A1 => n9555, A2 => n9562, ZN => n9595);
   U11796 : INV_X1 port map( A => n9560, ZN => n9562);
   U11797 : INV_X1 port map( A => n9556, ZN => n9555);
   U11798 : NAND2_X1 port map( A1 => n9551, A2 => n10511, ZN => n9591);
   U11799 : INV_X1 port map( A => n9552, ZN => n9551);
   U11800 : NAND2_X1 port map( A1 => n9556, A2 => n9560, ZN => n9592);
   U11801 : XNOR2_X1 port map( A => n8099, B => i_ALU_OP_2_port, ZN => n9556);
   U11802 : NAND2_X1 port map( A1 => n9590, A2 => n9589, ZN => n9593);
   U11803 : NOR2_X1 port map( A1 => DataPath_ALUhw_MULT_mux_out_0_0_port, A2 =>
                           n9588, ZN => n9589);
   U11804 : NOR2_X1 port map( A1 => n8167, A2 => n8681, ZN => n9588);
   U11805 : NAND2_X1 port map( A1 => n9552, A2 => n10487, ZN => n9590);
   U11806 : XNOR2_X1 port map( A => n7979, B => i_ALU_OP_2_port, ZN => n9552);
   U11807 : NAND2_X1 port map( A1 => n9658, A2 => n8011, ZN => n9656);
   U11808 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1557, B => n8300, ZN =>
                           n9658);
   U11809 : NAND2_X1 port map( A1 => n9635, A2 => n9653, ZN => n9657);
   U11810 : NAND2_X1 port map( A1 => n9582, A2 => n7787, ZN => n9653);
   U11811 : INV_X1 port map( A => n9583, ZN => n9582);
   U11812 : NAND2_X1 port map( A1 => n10838, A2 => n9634, ZN => n9635);
   U11813 : NAND2_X1 port map( A1 => n9583, A2 => n9603, ZN => n9634);
   U11814 : XNOR2_X1 port map( A => n9626, B => n8300, ZN => n9583);
   U11815 : AND2_X1 port map( A1 => n10455, A2 => n9586, ZN => n10838);
   U11816 : OR2_X1 port map( A1 => n10456, A2 => n10454, ZN => n10455);
   U11817 : NAND2_X1 port map( A1 => n10470, A2 => n10473, ZN => n10454);
   U11818 : XNOR2_X1 port map( A => n8015, B => n8300, ZN => n10470);
   U11819 : NAND2_X1 port map( A1 => n9586, A2 => n9652, ZN => n10456);
   U11820 : NAND2_X1 port map( A1 => n9584, A2 => n10457, ZN => n9652);
   U11821 : INV_X1 port map( A => n9585, ZN => n9584);
   U11822 : NAND2_X1 port map( A1 => n9585, A2 => n7818, ZN => n9586);
   U11823 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1659, B => n8300, ZN =>
                           n9585);
   U11824 : XNOR2_X1 port map( A => n9650, B => n7792, ZN => n9792);
   U11825 : XNOR2_X1 port map( A => n9794, B => i_ALU_OP_2_port, ZN => n9650);
   U11826 : AOI21_X1 port map( B1 => n9711, B2 => n9817, A => n9813, ZN => 
                           n9791);
   U11827 : NOR2_X1 port map( A1 => n9814, A2 => n9856, ZN => n9813);
   U11828 : NAND2_X1 port map( A1 => n9841, A2 => n10114, ZN => n9856);
   U11829 : XNOR2_X1 port map( A => n9839, B => i_ALU_OP_2_port, ZN => n9841);
   U11830 : XNOR2_X1 port map( A => n9711, B => n9817, ZN => n9814);
   U11831 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n435, B => 
                           i_ALU_OP_2_port, ZN => n9711);
   U11832 : NAND2_X1 port map( A1 => n8681, A2 => n9742, ZN => n12091);
   U11833 : AND2_X1 port map( A1 => n8167, A2 => n9533, ZN => 
                           DataPath_ALUhw_MULT_mux_out_0_0_port);
   U11834 : AOI211_X1 port map( C1 => n10511, C2 => n8167, A => n9449, B => 
                           n9448, ZN => DataPath_ALUhw_MULT_mux_out_0_1_port);
   U11835 : NOR2_X1 port map( A1 => n8167, A2 => n9533, ZN => n9449);
   U11836 : OAI22_X1 port map( A1 => n8489, A2 => n8566, B1 => n9452, B2 => 
                           n10511, ZN => DataPath_ALUhw_MULT_mux_out_1_3_port);
   U11837 : NOR2_X1 port map( A1 => n8485, A2 => n9553, ZN => 
                           DataPath_ALUhw_MULT_mux_out_1_2_port);
   U11838 : OAI22_X1 port map( A1 => n8568, A2 => n8488, B1 => n10511, B2 => 
                           n7786, ZN => DataPath_ALUhw_MULT_mux_out_2_5_port);
   U11839 : OAI22_X1 port map( A1 => n8573, A2 => n8488, B1 => n10511, B2 => 
                           n9458, ZN => DataPath_ALUhw_MULT_mux_out_3_7_port);
   U11840 : OAI22_X1 port map( A1 => n7788, A2 => n10511, B1 => n9560, B2 => 
                           n8570, ZN => DataPath_ALUhw_MULT_mux_out_2_6_port);
   U11841 : OAI22_X1 port map( A1 => n8574, A2 => n8488, B1 => n10511, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_9_port);
   U11842 : OAI22_X1 port map( A1 => n8573, A2 => n10511, B1 => n9560, B2 => 
                           n7700, ZN => DataPath_ALUhw_MULT_mux_out_3_8_port);
   U11843 : OAI22_X1 port map( A1 => n7788, A2 => n9560, B1 => n9721, B2 => 
                           n7786, ZN => DataPath_ALUhw_MULT_mux_out_2_7_port);
   U11844 : OAI22_X1 port map( A1 => n9721, A2 => n8563, B1 => n8485, B2 => 
                           n8495, ZN => DataPath_ALUhw_MULT_mux_out_1_6_port);
   U11845 : NOR2_X1 port map( A1 => n9470, A2 => n8488, ZN => 
                           DataPath_ALUhw_MULT_mux_out_5_10_port);
   U11846 : OAI22_X1 port map( A1 => n9469, A2 => n8488, B1 => n10511, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_11_port);
   U11847 : OAI22_X1 port map( A1 => n8574, A2 => n10511, B1 => n9560, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_10_port);
   U11848 : OAI22_X1 port map( A1 => n8572, A2 => n9560, B1 => n9721, B2 => 
                           n7700, ZN => DataPath_ALUhw_MULT_mux_out_3_9_port);
   U11849 : OAI22_X1 port map( A1 => n7788, A2 => n9721, B1 => n8496, B2 => 
                           n8569, ZN => DataPath_ALUhw_MULT_mux_out_2_8_port);
   U11850 : OAI22_X1 port map( A1 => n8496, A2 => n8563, B1 => n8485, B2 => 
                           n10457, ZN => DataPath_ALUhw_MULT_mux_out_1_7_port);
   U11851 : OAI22_X1 port map( A1 => n7763, A2 => n8488, B1 => n10511, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_13_port);
   U11852 : OAI22_X1 port map( A1 => n9469, A2 => n10511, B1 => n9560, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_12_port);
   U11853 : OAI22_X1 port map( A1 => n8574, A2 => n9560, B1 => n9721, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_11_port);
   U11854 : OAI22_X1 port map( A1 => n8573, A2 => n9721, B1 => n8496, B2 => 
                           n9458, ZN => DataPath_ALUhw_MULT_mux_out_3_10_port);
   U11855 : OAI22_X1 port map( A1 => n8568, A2 => n8495, B1 => n10457, B2 => 
                           n8569, ZN => DataPath_ALUhw_MULT_mux_out_2_9_port);
   U11856 : OAI22_X1 port map( A1 => n10457, A2 => n8563, B1 => n8485, B2 => 
                           n8490, ZN => DataPath_ALUhw_MULT_mux_out_1_8_port);
   U11857 : OAI22_X1 port map( A1 => n9481, A2 => n8488, B1 => n10511, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_15_port);
   U11858 : OAI22_X1 port map( A1 => n7763, A2 => n10511, B1 => n9560, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_14_port);
   U11859 : OAI22_X1 port map( A1 => n9469, A2 => n9560, B1 => n9721, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_13_port);
   U11860 : OAI22_X1 port map( A1 => n8574, A2 => n9721, B1 => n8495, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_12_port);
   U11861 : OAI22_X1 port map( A1 => n7783, A2 => n8495, B1 => n10457, B2 => 
                           n7700, ZN => DataPath_ALUhw_MULT_mux_out_3_11_port);
   U11862 : OAI22_X1 port map( A1 => n7788, A2 => n10457, B1 => n8490, B2 => 
                           n8570, ZN => DataPath_ALUhw_MULT_mux_out_2_10_port);
   U11863 : NOR2_X1 port map( A1 => n9487, A2 => n8488, ZN => 
                           DataPath_ALUhw_MULT_mux_out_8_16_port);
   U11864 : OAI22_X1 port map( A1 => n9486, A2 => n8488, B1 => n10511, B2 => 
                           n8576, ZN => DataPath_ALUhw_MULT_mux_out_8_17_port);
   U11865 : OAI22_X1 port map( A1 => n9481, A2 => n10511, B1 => n9560, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_16_port);
   U11866 : OAI22_X1 port map( A1 => n7763, A2 => n9560, B1 => n8491, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_15_port);
   U11867 : OAI22_X1 port map( A1 => n9469, A2 => n9721, B1 => n8495, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_14_port);
   U11868 : OAI22_X1 port map( A1 => n8574, A2 => n8495, B1 => n10457, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_13_port);
   U11869 : OAI22_X1 port map( A1 => n7783, A2 => n10457, B1 => n8490, B2 => 
                           n7701, ZN => DataPath_ALUhw_MULT_mux_out_3_12_port);
   U11870 : OAI22_X1 port map( A1 => n7788, A2 => n7787, B1 => n9659, B2 => 
                           n8570, ZN => DataPath_ALUhw_MULT_mux_out_2_11_port);
   U11871 : OAI22_X1 port map( A1 => n7754, A2 => n10395, B1 => n8487, B2 => 
                           n10423, ZN => DataPath_ALUhw_MULT_mux_out_0_10_port)
                           ;
   U11872 : OAI22_X1 port map( A1 => n9493, A2 => n8488, B1 => n10511, B2 => 
                           n8577, ZN => DataPath_ALUhw_MULT_mux_out_9_19_port);
   U11873 : OAI22_X1 port map( A1 => n9486, A2 => n10511, B1 => n9560, B2 => 
                           n8576, ZN => DataPath_ALUhw_MULT_mux_out_8_18_port);
   U11874 : OAI22_X1 port map( A1 => n9481, A2 => n9560, B1 => n8491, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_17_port);
   U11875 : OAI22_X1 port map( A1 => n7763, A2 => n9721, B1 => n8495, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_16_port);
   U11876 : OAI22_X1 port map( A1 => n9469, A2 => n8495, B1 => n10457, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_15_port);
   U11877 : OAI22_X1 port map( A1 => n8574, A2 => n10457, B1 => n8490, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_14_port);
   U11878 : OAI22_X1 port map( A1 => n7783, A2 => n8490, B1 => n9659, B2 => 
                           n9458, ZN => DataPath_ALUhw_MULT_mux_out_3_13_port);
   U11879 : OAI22_X1 port map( A1 => n8568, A2 => n9659, B1 => n8559, B2 => 
                           n7786, ZN => DataPath_ALUhw_MULT_mux_out_2_12_port);
   U11880 : OAI22_X1 port map( A1 => n7754, A2 => n10423, B1 => n8487, B2 => 
                           n10386, ZN => DataPath_ALUhw_MULT_mux_out_0_11_port)
                           ;
   U11881 : NOR2_X1 port map( A1 => n9501, A2 => n8488, ZN => 
                           DataPath_ALUhw_MULT_mux_out_10_20_port);
   U11882 : OAI22_X1 port map( A1 => n9500, A2 => n8488, B1 => n10511, B2 => 
                           n9501, ZN => DataPath_ALUhw_MULT_mux_out_10_21_port)
                           ;
   U11883 : OAI22_X1 port map( A1 => n9493, A2 => n10511, B1 => n9560, B2 => 
                           n8577, ZN => DataPath_ALUhw_MULT_mux_out_9_20_port);
   U11884 : OAI22_X1 port map( A1 => n9486, A2 => n9560, B1 => n8491, B2 => 
                           n8576, ZN => DataPath_ALUhw_MULT_mux_out_8_19_port);
   U11885 : OAI22_X1 port map( A1 => n9481, A2 => n9721, B1 => n8495, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_18_port);
   U11886 : OAI22_X1 port map( A1 => n7763, A2 => n8495, B1 => n10457, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_17_port);
   U11887 : OAI22_X1 port map( A1 => n9469, A2 => n10457, B1 => n8490, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_16_port);
   U11888 : OAI22_X1 port map( A1 => n8574, A2 => n7787, B1 => n9659, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_15_port);
   U11889 : OAI22_X1 port map( A1 => n7784, A2 => n9659, B1 => n8559, B2 => 
                           n7700, ZN => DataPath_ALUhw_MULT_mux_out_3_14_port);
   U11890 : OAI22_X1 port map( A1 => n7788, A2 => n8559, B1 => n10395, B2 => 
                           n8570, ZN => DataPath_ALUhw_MULT_mux_out_2_13_port);
   U11891 : OAI22_X1 port map( A1 => n10395, A2 => n8562, B1 => n9452, B2 => 
                           n10423, ZN => DataPath_ALUhw_MULT_mux_out_1_12_port)
                           ;
   U11892 : NOR2_X1 port map( A1 => n9508, A2 => n8488, ZN => 
                           DataPath_ALUhw_MULT_mux_out_11_22_port);
   U11893 : OAI22_X1 port map( A1 => n9507, A2 => n8488, B1 => n10511, B2 => 
                           n9508, ZN => DataPath_ALUhw_MULT_mux_out_11_23_port)
                           ;
   U11894 : OAI22_X1 port map( A1 => n9500, A2 => n10511, B1 => n9560, B2 => 
                           n9501, ZN => DataPath_ALUhw_MULT_mux_out_10_22_port)
                           ;
   U11895 : OAI22_X1 port map( A1 => n9493, A2 => n9560, B1 => n8491, B2 => 
                           n8577, ZN => DataPath_ALUhw_MULT_mux_out_9_21_port);
   U11896 : OAI22_X1 port map( A1 => n9486, A2 => n9721, B1 => n8495, B2 => 
                           n8576, ZN => DataPath_ALUhw_MULT_mux_out_8_20_port);
   U11897 : OAI22_X1 port map( A1 => n9481, A2 => n8495, B1 => n10457, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_19_port);
   U11898 : OAI22_X1 port map( A1 => n7763, A2 => n10457, B1 => n8490, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_18_port);
   U11899 : OAI22_X1 port map( A1 => n9469, A2 => n7787, B1 => n9659, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_17_port);
   U11900 : OAI22_X1 port map( A1 => n8574, A2 => n9659, B1 => n8559, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_16_port);
   U11901 : OAI22_X1 port map( A1 => n7784, A2 => n8559, B1 => n10395, B2 => 
                           n7700, ZN => DataPath_ALUhw_MULT_mux_out_3_15_port);
   U11902 : OAI22_X1 port map( A1 => n7788, A2 => n10395, B1 => n10423, B2 => 
                           n7786, ZN => DataPath_ALUhw_MULT_mux_out_2_14_port);
   U11903 : OAI22_X1 port map( A1 => n7755, A2 => n8492, B1 => n8487, B2 => 
                           n8555, ZN => DataPath_ALUhw_MULT_mux_out_0_13_port);
   U11904 : OAI22_X1 port map( A1 => n10423, A2 => n8567, B1 => n9452, B2 => 
                           n10386, ZN => DataPath_ALUhw_MULT_mux_out_1_13_port)
                           ;
   U11905 : NOR2_X1 port map( A1 => n9512, A2 => n8488, ZN => 
                           DataPath_ALUhw_MULT_mux_out_12_24_port);
   U11906 : OAI22_X1 port map( A1 => n9511, A2 => n8488, B1 => n10511, B2 => 
                           n9512, ZN => DataPath_ALUhw_MULT_mux_out_12_25_port)
                           ;
   U11907 : OAI22_X1 port map( A1 => n9507, A2 => n10511, B1 => n9560, B2 => 
                           n9508, ZN => DataPath_ALUhw_MULT_mux_out_11_24_port)
                           ;
   U11908 : OAI22_X1 port map( A1 => n9500, A2 => n9560, B1 => n8491, B2 => 
                           n9501, ZN => DataPath_ALUhw_MULT_mux_out_10_23_port)
                           ;
   U11909 : OAI22_X1 port map( A1 => n9493, A2 => n9721, B1 => n8495, B2 => 
                           n8577, ZN => DataPath_ALUhw_MULT_mux_out_9_22_port);
   U11910 : OAI22_X1 port map( A1 => n9486, A2 => n8495, B1 => n10457, B2 => 
                           n9487, ZN => DataPath_ALUhw_MULT_mux_out_8_21_port);
   U11911 : OAI22_X1 port map( A1 => n9481, A2 => n10457, B1 => n8490, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_20_port);
   U11912 : OAI22_X1 port map( A1 => n7763, A2 => n7787, B1 => n9659, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_19_port);
   U11913 : OAI22_X1 port map( A1 => n9469, A2 => n9659, B1 => n8559, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_18_port);
   U11914 : OAI22_X1 port map( A1 => n8574, A2 => n8559, B1 => n10395, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_17_port);
   U11915 : OAI22_X1 port map( A1 => n7784, A2 => n10395, B1 => n10423, B2 => 
                           n9458, ZN => DataPath_ALUhw_MULT_mux_out_3_16_port);
   U11916 : OAI22_X1 port map( A1 => n8568, A2 => n10423, B1 => n10386, B2 => 
                           n8570, ZN => DataPath_ALUhw_MULT_mux_out_2_15_port);
   U11917 : OAI22_X1 port map( A1 => n7754, A2 => n8555, B1 => n8487, B2 => 
                           n8494, ZN => DataPath_ALUhw_MULT_mux_out_0_14_port);
   U11918 : OAI22_X1 port map( A1 => n10386, A2 => n8567, B1 => n8485, B2 => 
                           n8492, ZN => DataPath_ALUhw_MULT_mux_out_1_14_port);
   U11919 : NOR2_X1 port map( A1 => n9519, A2 => n8488, ZN => 
                           DataPath_ALUhw_MULT_mux_out_13_26_port);
   U11920 : OAI22_X1 port map( A1 => n9518, A2 => n8488, B1 => n10511, B2 => 
                           n9519, ZN => DataPath_ALUhw_MULT_mux_out_13_27_port)
                           ;
   U11921 : OAI22_X1 port map( A1 => n9511, A2 => n10511, B1 => n9560, B2 => 
                           n9512, ZN => DataPath_ALUhw_MULT_mux_out_12_26_port)
                           ;
   U11922 : OAI22_X1 port map( A1 => n9507, A2 => n9560, B1 => n8491, B2 => 
                           n9508, ZN => DataPath_ALUhw_MULT_mux_out_11_25_port)
                           ;
   U11923 : OAI22_X1 port map( A1 => n9500, A2 => n8491, B1 => n8495, B2 => 
                           n9501, ZN => DataPath_ALUhw_MULT_mux_out_10_24_port)
                           ;
   U11924 : OAI22_X1 port map( A1 => n9493, A2 => n8495, B1 => n10457, B2 => 
                           n8577, ZN => DataPath_ALUhw_MULT_mux_out_9_23_port);
   U11925 : OAI22_X1 port map( A1 => n9486, A2 => n10457, B1 => n8490, B2 => 
                           n8576, ZN => DataPath_ALUhw_MULT_mux_out_8_22_port);
   U11926 : OAI22_X1 port map( A1 => n9481, A2 => n7787, B1 => n9659, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_21_port);
   U11927 : OAI22_X1 port map( A1 => n7763, A2 => n9659, B1 => n8559, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_20_port);
   U11928 : OAI22_X1 port map( A1 => n9469, A2 => n8559, B1 => n10395, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_19_port);
   U11929 : OAI22_X1 port map( A1 => n8574, A2 => n10395, B1 => n10423, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_18_port);
   U11930 : OAI22_X1 port map( A1 => n7784, A2 => n10423, B1 => n10386, B2 => 
                           n7701, ZN => DataPath_ALUhw_MULT_mux_out_3_17_port);
   U11931 : OAI22_X1 port map( A1 => n7788, A2 => n10386, B1 => n8492, B2 => 
                           n7786, ZN => DataPath_ALUhw_MULT_mux_out_2_16_port);
   U11932 : OAI22_X1 port map( A1 => n7755, A2 => n8494, B1 => n8554, B2 => 
                           n7796, ZN => DataPath_ALUhw_MULT_mux_out_0_15_port);
   U11933 : OAI22_X1 port map( A1 => n8493, A2 => n8567, B1 => n8485, B2 => 
                           n8555, ZN => DataPath_ALUhw_MULT_mux_out_1_15_port);
   U11934 : NOR2_X1 port map( A1 => n9523, A2 => n8489, ZN => 
                           DataPath_ALUhw_MULT_mux_out_14_28_port);
   U11935 : OAI22_X1 port map( A1 => n9522, A2 => n8488, B1 => n10511, B2 => 
                           n9523, ZN => DataPath_ALUhw_MULT_mux_out_14_29_port)
                           ;
   U11936 : OAI22_X1 port map( A1 => n9518, A2 => n10511, B1 => n9560, B2 => 
                           n9519, ZN => DataPath_ALUhw_MULT_mux_out_13_28_port)
                           ;
   U11937 : OAI22_X1 port map( A1 => n9511, A2 => n9560, B1 => n8491, B2 => 
                           n9512, ZN => DataPath_ALUhw_MULT_mux_out_12_27_port)
                           ;
   U11938 : OAI22_X1 port map( A1 => n9507, A2 => n9721, B1 => n8495, B2 => 
                           n9508, ZN => DataPath_ALUhw_MULT_mux_out_11_26_port)
                           ;
   U11939 : OAI22_X1 port map( A1 => n9500, A2 => n8495, B1 => n10457, B2 => 
                           n9501, ZN => DataPath_ALUhw_MULT_mux_out_10_25_port)
                           ;
   U11940 : OAI22_X1 port map( A1 => n9493, A2 => n10457, B1 => n8490, B2 => 
                           n8577, ZN => DataPath_ALUhw_MULT_mux_out_9_24_port);
   U11941 : OAI22_X1 port map( A1 => n9486, A2 => n8490, B1 => n9659, B2 => 
                           n8576, ZN => DataPath_ALUhw_MULT_mux_out_8_23_port);
   U11942 : OAI22_X1 port map( A1 => n9481, A2 => n9659, B1 => n8559, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_22_port);
   U11943 : OAI22_X1 port map( A1 => n7763, A2 => n8559, B1 => n10395, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_21_port);
   U11944 : OAI22_X1 port map( A1 => n9469, A2 => n10395, B1 => n10423, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_20_port);
   U11945 : OAI22_X1 port map( A1 => n8574, A2 => n10423, B1 => n10386, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_19_port);
   U11946 : OAI22_X1 port map( A1 => n8572, A2 => n10386, B1 => n8493, B2 => 
                           n7701, ZN => DataPath_ALUhw_MULT_mux_out_3_18_port);
   U11947 : OAI22_X1 port map( A1 => n7788, A2 => n8492, B1 => n8555, B2 => 
                           n7786, ZN => DataPath_ALUhw_MULT_mux_out_2_17_port);
   U11948 : OAI22_X1 port map( A1 => n7754, A2 => n8554, B1 => n8487, B2 => 
                           n10312, ZN => DataPath_ALUhw_MULT_mux_out_0_16_port)
                           ;
   U11949 : OAI22_X1 port map( A1 => n8555, A2 => n8565, B1 => n9452, B2 => 
                           n8494, ZN => DataPath_ALUhw_MULT_mux_out_1_16_port);
   U11950 : NOR2_X1 port map( A1 => n9526, A2 => n8489, ZN => 
                           DataPath_ALUhw_MULT_mux_out_15_30_port);
   U11951 : BUF_X1 port map( A => n9553, Z => n8489);
   U11952 : OAI22_X1 port map( A1 => n7755, A2 => n9761, B1 => n7796, B2 => 
                           n10024, ZN => DataPath_ALUhw_MULT_mux_out_0_31_port)
                           ;
   U11953 : OAI22_X1 port map( A1 => n10114, A2 => n8563, B1 => n9452, B2 => 
                           n9817, ZN => DataPath_ALUhw_MULT_mux_out_1_31_port);
   U11954 : OAI22_X1 port map( A1 => n8568, A2 => n10181, B1 => n9874, B2 => 
                           n8570, ZN => DataPath_ALUhw_MULT_mux_out_2_31_port);
   U11955 : OAI22_X1 port map( A1 => n7784, A2 => n9979, B1 => n9944, B2 => 
                           n7701, ZN => DataPath_ALUhw_MULT_mux_out_3_31_port);
   U11956 : OAI22_X1 port map( A1 => n8574, A2 => n8553, B1 => n10010, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_31_port);
   U11957 : OAI22_X1 port map( A1 => n9469, A2 => n7795, B1 => n8556, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_31_port);
   U11958 : OAI22_X1 port map( A1 => n7763, A2 => n10197, B1 => n10143, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_31_port);
   U11959 : OAI22_X1 port map( A1 => n9481, A2 => n8557, B1 => n8550, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_31_port);
   U11960 : OAI22_X1 port map( A1 => n9486, A2 => n8494, B1 => n8554, B2 => 
                           n8576, ZN => DataPath_ALUhw_MULT_mux_out_8_31_port);
   U11961 : OAI22_X1 port map( A1 => n9493, A2 => n8492, B1 => n8555, B2 => 
                           n8577, ZN => DataPath_ALUhw_MULT_mux_out_9_31_port);
   U11962 : OAI22_X1 port map( A1 => n9500, A2 => n10423, B1 => n10386, B2 => 
                           n9501, ZN => DataPath_ALUhw_MULT_mux_out_10_31_port)
                           ;
   U11963 : OAI22_X1 port map( A1 => n9507, A2 => n8559, B1 => n10395, B2 => 
                           n9508, ZN => DataPath_ALUhw_MULT_mux_out_11_31_port)
                           ;
   U11964 : OAI22_X1 port map( A1 => n9511, A2 => n7787, B1 => n9659, B2 => 
                           n9512, ZN => DataPath_ALUhw_MULT_mux_out_12_31_port)
                           ;
   U11965 : OAI22_X1 port map( A1 => n9518, A2 => n8495, B1 => n10457, B2 => 
                           n9519, ZN => DataPath_ALUhw_MULT_mux_out_13_31_port)
                           ;
   U11966 : OAI22_X1 port map( A1 => n9522, A2 => n9560, B1 => n8491, B2 => 
                           n9523, ZN => DataPath_ALUhw_MULT_mux_out_14_31_port)
                           ;
   U11967 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n435, B => n9794, ZN => 
                           n9526);
   U11968 : OAI21_X1 port map( B1 => n8365, B2 => n8673, A => n9429, ZN => 
                           n9533);
   U11969 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_0_port, A2 => n8671, 
                           ZN => n9429);
   U11970 : OAI21_X1 port map( B1 => n8404, B2 => n8683, A => n9524, ZN => 
                           DP_OP_751_130_5637_n333);
   U11971 : NAND2_X1 port map( A1 => n8682, A2 => DataPath_i_PIPLIN_IN2_31_port
                           , ZN => n9524);
   U11972 : OAI21_X1 port map( B1 => n8405, B2 => n8683, A => n9525, ZN => 
                           n9794);
   U11973 : NAND2_X1 port map( A1 => n8682, A2 => DataPath_i_PIPLIN_IN2_30_port
                           , ZN => n9525);
   U11974 : OAI22_X1 port map( A1 => n7788, A2 => n9944, B1 => n10181, B2 => 
                           n8569, ZN => DataPath_ALUhw_MULT_mux_out_2_30_port);
   U11975 : OAI22_X1 port map( A1 => n7784, A2 => n10010, B1 => n9979, B2 => 
                           n7701, ZN => DataPath_ALUhw_MULT_mux_out_3_30_port);
   U11976 : OAI22_X1 port map( A1 => n8574, A2 => n8556, B1 => n8553, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_30_port);
   U11977 : OAI22_X1 port map( A1 => n9469, A2 => n10143, B1 => n7795, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_30_port);
   U11978 : OAI22_X1 port map( A1 => n7763, A2 => n8550, B1 => n10197, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_30_port);
   U11979 : OAI22_X1 port map( A1 => n9481, A2 => n8554, B1 => n9482, B2 => 
                           n8558, ZN => DataPath_ALUhw_MULT_mux_out_7_30_port);
   U11980 : OAI22_X1 port map( A1 => n9486, A2 => n8555, B1 => n7789, B2 => 
                           n9487, ZN => DataPath_ALUhw_MULT_mux_out_8_30_port);
   U11981 : OAI22_X1 port map( A1 => n9493, A2 => n10386, B1 => n8493, B2 => 
                           n8577, ZN => DataPath_ALUhw_MULT_mux_out_9_30_port);
   U11982 : OAI22_X1 port map( A1 => n9500, A2 => n10395, B1 => n10423, B2 => 
                           n9501, ZN => DataPath_ALUhw_MULT_mux_out_10_30_port)
                           ;
   U11983 : OAI22_X1 port map( A1 => n9507, A2 => n9659, B1 => n8559, B2 => 
                           n9508, ZN => DataPath_ALUhw_MULT_mux_out_11_30_port)
                           ;
   U11984 : OAI22_X1 port map( A1 => n9511, A2 => n10457, B1 => n7787, B2 => 
                           n9512, ZN => DataPath_ALUhw_MULT_mux_out_12_30_port)
                           ;
   U11985 : OAI22_X1 port map( A1 => n9518, A2 => n9721, B1 => n8495, B2 => 
                           n9519, ZN => DataPath_ALUhw_MULT_mux_out_13_30_port)
                           ;
   U11986 : OAI22_X1 port map( A1 => n9522, A2 => n10511, B1 => n9560, B2 => 
                           n9523, ZN => DataPath_ALUhw_MULT_mux_out_14_30_port)
                           ;
   U11987 : NAND2_X1 port map( A1 => n8682, A2 => DataPath_i_PIPLIN_IN2_29_port
                           , ZN => n9520);
   U11988 : OAI21_X1 port map( B1 => n8403, B2 => n8683, A => n9521, ZN => 
                           n9839);
   U11989 : NAND2_X1 port map( A1 => n8682, A2 => DataPath_i_PIPLIN_IN2_28_port
                           , ZN => n9521);
   U11990 : OAI22_X1 port map( A1 => n8568, A2 => n9979, B1 => n9944, B2 => 
                           n7786, ZN => DataPath_ALUhw_MULT_mux_out_2_29_port);
   U11991 : OAI22_X1 port map( A1 => n7784, A2 => n8553, B1 => n10010, B2 => 
                           n9458, ZN => DataPath_ALUhw_MULT_mux_out_3_29_port);
   U11992 : OAI22_X1 port map( A1 => n8574, A2 => n7795, B1 => n8556, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_29_port);
   U11993 : OAI22_X1 port map( A1 => n9469, A2 => n10197, B1 => n10143, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_29_port);
   U11994 : OAI22_X1 port map( A1 => n7763, A2 => n8557, B1 => n8551, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_29_port);
   U11995 : OAI22_X1 port map( A1 => n9481, A2 => n8494, B1 => n8554, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_29_port);
   U11996 : OAI22_X1 port map( A1 => n9486, A2 => n8492, B1 => n8555, B2 => 
                           n8576, ZN => DataPath_ALUhw_MULT_mux_out_8_29_port);
   U11997 : OAI22_X1 port map( A1 => n9493, A2 => n10423, B1 => n10386, B2 => 
                           n8577, ZN => DataPath_ALUhw_MULT_mux_out_9_29_port);
   U11998 : OAI22_X1 port map( A1 => n9500, A2 => n8559, B1 => n10395, B2 => 
                           n9501, ZN => DataPath_ALUhw_MULT_mux_out_10_29_port)
                           ;
   U11999 : OAI22_X1 port map( A1 => n9507, A2 => n7787, B1 => n9659, B2 => 
                           n9508, ZN => DataPath_ALUhw_MULT_mux_out_11_29_port)
                           ;
   U12000 : OAI22_X1 port map( A1 => n9511, A2 => n8496, B1 => n10457, B2 => 
                           n9512, ZN => DataPath_ALUhw_MULT_mux_out_12_29_port)
                           ;
   U12001 : OAI22_X1 port map( A1 => n9518, A2 => n9560, B1 => n8491, B2 => 
                           n9519, ZN => DataPath_ALUhw_MULT_mux_out_13_29_port)
                           ;
   U12002 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_2_port, A2 => n8671, 
                           ZN => n9350);
   U12003 : NAND2_X1 port map( A1 => n8314, A2 => DataPath_i_PIPLIN_IN1_2_port,
                           ZN => n9351);
   U12004 : OAI21_X1 port map( B1 => n9875, B2 => DP_OP_751_130_5637_n639, A =>
                           n9515, ZN => n9516);
   U12005 : NAND2_X1 port map( A1 => n9875, A2 => n9909, ZN => n9515);
   U12006 : NAND2_X1 port map( A1 => n8682, A2 => DataPath_i_PIPLIN_IN2_27_port
                           , ZN => n9513);
   U12007 : INV_X1 port map( A => n9909, ZN => n9517);
   U12008 : OAI21_X1 port map( B1 => n8356, B2 => n8683, A => n9514, ZN => 
                           n9909);
   U12009 : NAND2_X1 port map( A1 => n8682, A2 => DataPath_i_PIPLIN_IN2_26_port
                           , ZN => n9514);
   U12010 : OAI22_X1 port map( A1 => n9944, A2 => n8560, B1 => n9452, B2 => 
                           n10181, ZN => DataPath_ALUhw_MULT_mux_out_1_28_port)
                           ;
   U12011 : OAI22_X1 port map( A1 => n8568, A2 => n10010, B1 => n9979, B2 => 
                           n8570, ZN => DataPath_ALUhw_MULT_mux_out_2_28_port);
   U12012 : OAI22_X1 port map( A1 => n7784, A2 => n8556, B1 => n8553, B2 => 
                           n7700, ZN => DataPath_ALUhw_MULT_mux_out_3_28_port);
   U12013 : OAI22_X1 port map( A1 => n8574, A2 => n10143, B1 => n7795, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_28_port);
   U12014 : OAI22_X1 port map( A1 => n9469, A2 => n8551, B1 => n10197, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_28_port);
   U12015 : INV_X1 port map( A => n7767, ZN => n8550);
   U12016 : OAI22_X1 port map( A1 => n7763, A2 => n8554, B1 => n9475, B2 => 
                           n8558, ZN => DataPath_ALUhw_MULT_mux_out_6_28_port);
   U12017 : OAI22_X1 port map( A1 => n9481, A2 => n8555, B1 => n7789, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_28_port);
   U12018 : OAI22_X1 port map( A1 => n9486, A2 => n10386, B1 => n8493, B2 => 
                           n9487, ZN => DataPath_ALUhw_MULT_mux_out_8_28_port);
   U12019 : OAI22_X1 port map( A1 => n9493, A2 => n10395, B1 => n10423, B2 => 
                           n8577, ZN => DataPath_ALUhw_MULT_mux_out_9_28_port);
   U12020 : OAI22_X1 port map( A1 => n9500, A2 => n9659, B1 => n8559, B2 => 
                           n9501, ZN => DataPath_ALUhw_MULT_mux_out_10_28_port)
                           ;
   U12021 : OAI22_X1 port map( A1 => n9507, A2 => n10457, B1 => n7787, B2 => 
                           n9508, ZN => DataPath_ALUhw_MULT_mux_out_11_28_port)
                           ;
   U12022 : OAI22_X1 port map( A1 => n9511, A2 => n9721, B1 => n8495, B2 => 
                           n9512, ZN => DataPath_ALUhw_MULT_mux_out_12_28_port)
                           ;
   U12023 : NAND2_X1 port map( A1 => n9361, A2 => n9360, ZN => n9596);
   U12024 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_3_port, A2 => n8671, 
                           ZN => n9360);
   U12025 : NAND2_X1 port map( A1 => n8314, A2 => DataPath_i_PIPLIN_IN1_3_port,
                           ZN => n9361);
   U12026 : OAI21_X1 port map( B1 => n8354, B2 => n8683, A => n9510, ZN => 
                           n9969);
   U12027 : NAND2_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_24_port
                           , ZN => n9510);
   U12028 : NAND2_X1 port map( A1 => n8682, A2 => DataPath_i_PIPLIN_IN2_25_port
                           , ZN => n9509);
   U12029 : OAI22_X1 port map( A1 => n7754, A2 => n10181, B1 => n7796, B2 => 
                           n9874, ZN => DataPath_ALUhw_MULT_mux_out_0_27_port);
   U12030 : OAI22_X1 port map( A1 => n8568, A2 => n8553, B1 => n10010, B2 => 
                           n7786, ZN => DataPath_ALUhw_MULT_mux_out_2_27_port);
   U12031 : OAI22_X1 port map( A1 => n7783, A2 => n7795, B1 => n8556, B2 => 
                           n7700, ZN => DataPath_ALUhw_MULT_mux_out_3_27_port);
   U12032 : OAI22_X1 port map( A1 => n8574, A2 => n10197, B1 => n10143, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_27_port);
   U12033 : OAI22_X1 port map( A1 => n9469, A2 => n8557, B1 => n8550, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_27_port);
   U12034 : OAI22_X1 port map( A1 => n7763, A2 => n8494, B1 => n8554, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_27_port);
   U12035 : OAI22_X1 port map( A1 => n9481, A2 => n8492, B1 => n8555, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_27_port);
   U12036 : OAI22_X1 port map( A1 => n9486, A2 => n10423, B1 => n10386, B2 => 
                           n8576, ZN => DataPath_ALUhw_MULT_mux_out_8_27_port);
   U12037 : OAI22_X1 port map( A1 => n9493, A2 => n8559, B1 => n10395, B2 => 
                           n9494, ZN => DataPath_ALUhw_MULT_mux_out_9_27_port);
   U12038 : OAI22_X1 port map( A1 => n9500, A2 => n7787, B1 => n9659, B2 => 
                           n9501, ZN => DataPath_ALUhw_MULT_mux_out_10_27_port)
                           ;
   U12039 : OAI22_X1 port map( A1 => n9507, A2 => n8496, B1 => n10457, B2 => 
                           n9508, ZN => DataPath_ALUhw_MULT_mux_out_11_27_port)
                           ;
   U12040 : OAI21_X1 port map( B1 => n8364, B2 => n8673, A => n9412, ZN => 
                           n10473);
   U12041 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_4_port, A2 => n8671, 
                           ZN => n9412);
   U12042 : OAI21_X1 port map( B1 => n10011, B2 => DP_OP_751_130_5637_n843, A 
                           => n9504, ZN => n9505);
   U12043 : NAND2_X1 port map( A1 => n10011, A2 => n10046, ZN => n9504);
   U12044 : NAND2_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_23_port
                           , ZN => n9502);
   U12045 : INV_X1 port map( A => n10046, ZN => n9506);
   U12046 : OAI21_X1 port map( B1 => n8353, B2 => n8682, A => n9503, ZN => 
                           n10046);
   U12047 : NAND2_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_22_port
                           , ZN => n9503);
   U12048 : OAI22_X1 port map( A1 => n10010, A2 => n8567, B1 => n8485, B2 => 
                           n9979, ZN => DataPath_ALUhw_MULT_mux_out_1_26_port);
   U12049 : OAI22_X1 port map( A1 => n7788, A2 => n8556, B1 => n8553, B2 => 
                           n8570, ZN => DataPath_ALUhw_MULT_mux_out_2_26_port);
   U12050 : OAI22_X1 port map( A1 => n7783, A2 => n10143, B1 => n7795, B2 => 
                           n9458, ZN => DataPath_ALUhw_MULT_mux_out_3_26_port);
   U12051 : OAI22_X1 port map( A1 => n8574, A2 => n8550, B1 => n10197, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_26_port);
   U12052 : OAI22_X1 port map( A1 => n9469, A2 => n8554, B1 => n9470, B2 => 
                           n8558, ZN => DataPath_ALUhw_MULT_mux_out_5_26_port);
   U12053 : OAI22_X1 port map( A1 => n7763, A2 => n8555, B1 => n7789, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_26_port);
   U12054 : OAI22_X1 port map( A1 => n9481, A2 => n10386, B1 => n8493, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_26_port);
   U12055 : OAI22_X1 port map( A1 => n9486, A2 => n10395, B1 => n10423, B2 => 
                           n8576, ZN => DataPath_ALUhw_MULT_mux_out_8_26_port);
   U12056 : OAI22_X1 port map( A1 => n9493, A2 => n9659, B1 => n8559, B2 => 
                           n9494, ZN => DataPath_ALUhw_MULT_mux_out_9_26_port);
   U12057 : OAI22_X1 port map( A1 => n9500, A2 => n10457, B1 => n8490, B2 => 
                           n9501, ZN => DataPath_ALUhw_MULT_mux_out_10_26_port)
                           ;
   U12058 : OAI21_X1 port map( B1 => n8362, B2 => n8673, A => n9400, ZN => 
                           n10463);
   U12059 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_5_port, A2 => n8672, 
                           ZN => n9400);
   U12060 : OAI21_X1 port map( B1 => n10144, B2 => DP_OP_751_130_5637_n843, A 
                           => n9498, ZN => n9499);
   U12061 : NAND2_X1 port map( A1 => n9497, A2 => DP_OP_751_130_5637_n843, ZN 
                           => n9498);
   U12062 : INV_X1 port map( A => n10124, ZN => n9497);
   U12063 : NAND2_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_21_port
                           , ZN => n9495);
   U12064 : OAI21_X1 port map( B1 => n8351, B2 => n8682, A => n9496, ZN => 
                           n10124);
   U12065 : NAND2_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_20_port
                           , ZN => n9496);
   U12066 : INV_X1 port map( A => DP_OP_751_130_5637_n945, ZN => n10144);
   U12067 : OAI22_X1 port map( A1 => n8574, A2 => n8557, B1 => n8551, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_25_port);
   U12068 : OAI22_X1 port map( A1 => n9469, A2 => n8494, B1 => n8554, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_25_port);
   U12069 : OAI22_X1 port map( A1 => n7763, A2 => n8492, B1 => n8555, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_25_port);
   U12070 : OAI22_X1 port map( A1 => n9481, A2 => n10423, B1 => n10386, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_25_port);
   U12071 : OAI22_X1 port map( A1 => n9486, A2 => n8559, B1 => n10395, B2 => 
                           n8576, ZN => DataPath_ALUhw_MULT_mux_out_8_25_port);
   U12072 : OAI22_X1 port map( A1 => n9493, A2 => n7787, B1 => n9659, B2 => 
                           n9494, ZN => DataPath_ALUhw_MULT_mux_out_9_25_port);
   U12073 : OAI21_X1 port map( B1 => n8360, B2 => n8673, A => n9373, ZN => 
                           n9603);
   U12074 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_6_port, A2 => n8674, 
                           ZN => n9373);
   U12075 : OAI21_X1 port map( B1 => n10217, B2 => DP_OP_751_130_5637_n945, A 
                           => n9491, ZN => n9492);
   U12076 : NAND2_X1 port map( A1 => n9490, A2 => DP_OP_751_130_5637_n945, ZN 
                           => n9491);
   U12077 : INV_X1 port map( A => n10198, ZN => n9490);
   U12078 : OAI21_X1 port map( B1 => n8349, B2 => n8682, A => n9488, ZN => 
                           DP_OP_751_130_5637_n945);
   U12079 : NAND2_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_19_port
                           , ZN => n9488);
   U12080 : OAI21_X1 port map( B1 => n8350, B2 => n8682, A => n9489, ZN => 
                           n10198);
   U12081 : NAND2_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_18_port
                           , ZN => n9489);
   U12082 : OAI22_X1 port map( A1 => n7784, A2 => n8550, B1 => n10197, B2 => 
                           n7701, ZN => DataPath_ALUhw_MULT_mux_out_3_24_port);
   U12083 : OAI22_X1 port map( A1 => n8574, A2 => n8554, B1 => n7694, B2 => 
                           n8557, ZN => DataPath_ALUhw_MULT_mux_out_4_24_port);
   U12084 : OAI22_X1 port map( A1 => n9469, A2 => n8555, B1 => n7789, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_24_port);
   U12085 : OAI22_X1 port map( A1 => n7763, A2 => n10386, B1 => n8493, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_24_port);
   U12086 : OAI22_X1 port map( A1 => n9481, A2 => n10395, B1 => n10423, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_24_port);
   U12087 : OAI22_X1 port map( A1 => n9486, A2 => n9659, B1 => n8559, B2 => 
                           n8576, ZN => DataPath_ALUhw_MULT_mux_out_8_24_port);
   U12088 : OAI21_X1 port map( B1 => n8361, B2 => n8673, A => n9380, ZN => 
                           n9651);
   U12089 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_7_port, A2 => n8674, 
                           ZN => n9380);
   U12090 : AOI21_X1 port map( B1 => n7794, B2 => n10313, A => n9484, ZN => 
                           n9485);
   U12091 : NOR2_X1 port map( A1 => n7794, A2 => n10217, ZN => n9484);
   U12092 : INV_X1 port map( A => DP_OP_751_130_5637_n1047, ZN => n10217);
   U12093 : OAI21_X1 port map( B1 => n8348, B2 => n8683, A => n9483, ZN => 
                           DP_OP_751_130_5637_n1047);
   U12094 : NAND2_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_17_port
                           , ZN => n9483);
   U12095 : OAI22_X1 port map( A1 => n7788, A2 => n10197, B1 => n10143, B2 => 
                           n8570, ZN => DataPath_ALUhw_MULT_mux_out_2_23_port);
   U12096 : OAI22_X1 port map( A1 => n7784, A2 => n8557, B1 => n8550, B2 => 
                           n9458, ZN => DataPath_ALUhw_MULT_mux_out_3_23_port);
   U12097 : OAI22_X1 port map( A1 => n8574, A2 => n8494, B1 => n8554, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_23_port);
   U12098 : OAI22_X1 port map( A1 => n9469, A2 => n8492, B1 => n8555, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_23_port);
   U12099 : OAI22_X1 port map( A1 => n7763, A2 => n10423, B1 => n10386, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_23_port);
   U12100 : OAI22_X1 port map( A1 => n9481, A2 => n8559, B1 => n10395, B2 => 
                           n9482, ZN => DataPath_ALUhw_MULT_mux_out_7_23_port);
   U12101 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_8_port, A2 => n8671, 
                           ZN => n9430);
   U12102 : NAND2_X1 port map( A1 => n8314, A2 => DataPath_i_PIPLIN_IN1_8_port,
                           ZN => n9431);
   U12103 : OAI21_X1 port map( B1 => n7793, B2 => DP_OP_751_130_5637_n1149, A 
                           => n9479, ZN => n9480);
   U12104 : NAND2_X1 port map( A1 => n9478, A2 => DP_OP_751_130_5637_n1149, ZN 
                           => n9479);
   U12105 : INV_X1 port map( A => n10379, ZN => n9478);
   U12106 : OAI21_X1 port map( B1 => n8346, B2 => n8683, A => n9476, ZN => 
                           DP_OP_751_130_5637_n1149);
   U12107 : NAND2_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_15_port
                           , ZN => n9476);
   U12108 : OAI21_X1 port map( B1 => n8347, B2 => n8683, A => n9477, ZN => 
                           n10379);
   U12109 : NAND2_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_14_port
                           , ZN => n9477);
   U12110 : OAI22_X1 port map( A1 => n8568, A2 => n8551, B1 => n10197, B2 => 
                           n8569, ZN => DataPath_ALUhw_MULT_mux_out_2_22_port);
   U12111 : OAI22_X1 port map( A1 => n7784, A2 => n8554, B1 => n7701, B2 => 
                           n8557, ZN => DataPath_ALUhw_MULT_mux_out_3_22_port);
   U12112 : OAI22_X1 port map( A1 => n8574, A2 => n8555, B1 => n8494, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_22_port);
   U12113 : OAI22_X1 port map( A1 => n9469, A2 => n10386, B1 => n8493, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_22_port);
   U12114 : OAI22_X1 port map( A1 => n7763, A2 => n10395, B1 => n10423, B2 => 
                           n9475, ZN => DataPath_ALUhw_MULT_mux_out_6_22_port);
   U12115 : OAI21_X1 port map( B1 => n8357, B2 => n8673, A => n9334, ZN => 
                           n10409);
   U12116 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_9_port, A2 => n8671, 
                           ZN => n9334);
   U12117 : OAI211_X1 port map( C1 => DP_OP_751_130_5637_n1251, C2 => n10337, A
                           => n9473, B => n9472, ZN => n9474);
   U12118 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1353, A2 => 
                           DP_OP_751_130_5637_n1251, ZN => n9472);
   U12119 : NAND2_X1 port map( A1 => n8677, A2 => n10337, ZN => n9473);
   U12120 : OAI21_X1 port map( B1 => n8345, B2 => n8683, A => n9471, ZN => 
                           n10337);
   U12121 : NAND2_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_12_port
                           , ZN => n9471);
   U12122 : OAI22_X1 port map( A1 => n8568, A2 => n8557, B1 => n8550, B2 => 
                           n8569, ZN => DataPath_ALUhw_MULT_mux_out_2_21_port);
   U12123 : OAI22_X1 port map( A1 => n8573, A2 => n8494, B1 => n8554, B2 => 
                           n7700, ZN => DataPath_ALUhw_MULT_mux_out_3_21_port);
   U12124 : OAI21_X1 port map( B1 => DP_OP_751_130_5637_n1659, B2 => 
                           DP_OP_751_130_5637_n1557, A => n9457, ZN => n8572);
   U12125 : OAI22_X1 port map( A1 => n8574, A2 => n8492, B1 => n8555, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_21_port);
   U12126 : OAI22_X1 port map( A1 => n9469, A2 => n10423, B1 => n10386, B2 => 
                           n9470, ZN => DataPath_ALUhw_MULT_mux_out_5_21_port);
   U12127 : OAI21_X1 port map( B1 => n8358, B2 => n8673, A => n9348, ZN => 
                           n9664);
   U12128 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_10_port, A2 => n8671, 
                           ZN => n9348);
   U12129 : OAI21_X1 port map( B1 => n7771, B2 => DP_OP_751_130_5637_n1353, A 
                           => n9467, ZN => n9468);
   U12130 : NAND2_X1 port map( A1 => n9466, A2 => DP_OP_751_130_5637_n1353, ZN 
                           => n9467);
   U12131 : INV_X1 port map( A => n10419, ZN => n9466);
   U12132 : INV_X1 port map( A => n411, ZN => n8677);
   U12133 : OAI21_X1 port map( B1 => n8342, B2 => n8683, A => n9464, ZN => n411
                           );
   U12134 : NAND2_X1 port map( A1 => n8682, A2 => DataPath_i_PIPLIN_IN2_11_port
                           , ZN => n9464);
   U12135 : OAI21_X1 port map( B1 => n8343, B2 => n8683, A => n9465, ZN => 
                           n10419);
   U12136 : NAND2_X1 port map( A1 => n8682, A2 => DataPath_i_PIPLIN_IN2_10_port
                           , ZN => n9465);
   U12137 : OAI22_X1 port map( A1 => n7754, A2 => n10143, B1 => n8487, B2 => 
                           n7795, ZN => DataPath_ALUhw_MULT_mux_out_0_20_port);
   U12138 : OAI22_X1 port map( A1 => n10223, A2 => n8560, B1 => n9452, B2 => 
                           n10197, ZN => DataPath_ALUhw_MULT_mux_out_1_20_port)
                           ;
   U12139 : OAI22_X1 port map( A1 => n8568, A2 => n8554, B1 => n8570, B2 => 
                           n8558, ZN => DataPath_ALUhw_MULT_mux_out_2_20_port);
   U12140 : BUF_X1 port map( A => n9455, Z => n8570);
   U12141 : OAI22_X1 port map( A1 => n7784, A2 => n8555, B1 => n7789, B2 => 
                           n7700, ZN => DataPath_ALUhw_MULT_mux_out_3_20_port);
   U12142 : XNOR2_X1 port map( A => n9626, B => DP_OP_751_130_5637_n1659, ZN =>
                           n8571);
   U12143 : OAI22_X1 port map( A1 => n8574, A2 => n10386, B1 => n8493, B2 => 
                           n7694, ZN => DataPath_ALUhw_MULT_mux_out_4_20_port);
   U12144 : OAI21_X1 port map( B1 => n8359, B2 => n8673, A => n9362, ZN => 
                           n10385);
   U12145 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_11_port, A2 => n8671, 
                           ZN => n9362);
   U12146 : OAI21_X1 port map( B1 => n415, B2 => DP_OP_751_130_5637_n1455, A =>
                           n9462, ZN => n9463);
   U12147 : NAND2_X1 port map( A1 => n9461, A2 => DP_OP_751_130_5637_n1455, ZN 
                           => n9462);
   U12148 : INV_X1 port map( A => n10446, ZN => n9461);
   U12149 : NAND2_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_9_port,
                           ZN => n9459);
   U12150 : NAND2_X1 port map( A1 => n8683, A2 => DataPath_i_PIPLIN_IN2_8_port,
                           ZN => n9460);
   U12151 : OAI22_X1 port map( A1 => n9447, A2 => n10197, B1 => n8487, B2 => 
                           n10143, ZN => DataPath_ALUhw_MULT_mux_out_0_19_port)
                           ;
   U12152 : OAI22_X1 port map( A1 => n8557, A2 => n8566, B1 => n9452, B2 => 
                           n10223, ZN => DataPath_ALUhw_MULT_mux_out_1_19_port)
                           ;
   U12153 : OAI22_X1 port map( A1 => n8568, A2 => n8494, B1 => n8554, B2 => 
                           n7786, ZN => DataPath_ALUhw_MULT_mux_out_2_19_port);
   U12154 : OAI22_X1 port map( A1 => n7784, A2 => n8492, B1 => n8555, B2 => 
                           n9458, ZN => DataPath_ALUhw_MULT_mux_out_3_19_port);
   U12155 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_12_port, A2 => n8672, 
                           ZN => n9407);
   U12156 : NAND2_X1 port map( A1 => n8682, A2 => DataPath_i_PIPLIN_IN2_7_port,
                           ZN => n9456);
   U12157 : OAI22_X1 port map( A1 => n9447, A2 => n10223, B1 => n8487, B2 => 
                           n10197, ZN => DataPath_ALUhw_MULT_mux_out_0_18_port)
                           ;
   U12158 : OAI22_X1 port map( A1 => n8554, A2 => n8566, B1 => n9452, B2 => 
                           n8558, ZN => DataPath_ALUhw_MULT_mux_out_1_18_port);
   U12159 : OAI22_X1 port map( A1 => n7788, A2 => n8555, B1 => n7789, B2 => 
                           n8569, ZN => DataPath_ALUhw_MULT_mux_out_2_18_port);
   U12160 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_13_port, A2 => n8672, 
                           ZN => n9397);
   U12161 : NAND2_X1 port map( A1 => n8314, A2 => DataPath_i_PIPLIN_IN1_13_port
                           , ZN => n9398);
   U12162 : OAI21_X1 port map( B1 => n8338, B2 => n8138, A => n9453, ZN => n417
                           );
   U12163 : NAND2_X1 port map( A1 => i_S2, A2 => DataPath_i_PIPLIN_IN2_5_port, 
                           ZN => n9453);
   U12164 : NAND2_X1 port map( A1 => DP_OP_751_130_5637_n1761, A2 => n10467, ZN
                           => n10021);
   U12165 : OAI21_X1 port map( B1 => n8335, B2 => n8138, A => n9333, ZN => 
                           n10467);
   U12166 : NAND2_X1 port map( A1 => i_S2, A2 => DataPath_i_PIPLIN_IN2_4_port, 
                           ZN => n9333);
   U12167 : OAI22_X1 port map( A1 => n9447, A2 => n10312, B1 => n8487, B2 => 
                           n10223, ZN => DataPath_ALUhw_MULT_mux_out_0_17_port)
                           ;
   U12168 : INV_X1 port map( A => n9587, ZN => n9530);
   U12169 : OAI21_X1 port map( B1 => n8337, B2 => i_S2, A => n9346, ZN => n9587
                           );
   U12170 : NAND2_X1 port map( A1 => i_S2, A2 => DataPath_i_PIPLIN_IN2_0_port, 
                           ZN => n9346);
   U12171 : OAI22_X1 port map( A1 => n7789, A2 => n8567, B1 => n9452, B2 => 
                           n8554, ZN => DataPath_ALUhw_MULT_mux_out_1_17_port);
   U12172 : OAI21_X1 port map( B1 => n8336, B2 => i_S2, A => n9345, ZN => n9563
                           );
   U12173 : NAND2_X1 port map( A1 => i_S2, A2 => DataPath_i_PIPLIN_IN2_2_port, 
                           ZN => n9345);
   U12174 : INV_X1 port map( A => DP_OP_751_130_5637_I2, ZN => 
                           DP_OP_751_130_5637_n1794);
   U12175 : INV_X1 port map( A => n10377, ZN => n10378);
   U12176 : NAND4_X1 port map( A1 => n8443, A2 => DP_OP_1090J1_126_7243_n72, A3
                           => DRAMRF_READY, A4 => n8713, ZN => n9646);
   U12177 : NAND2_X1 port map( A1 => n10856, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_15_port, ZN => 
                           n12208);
   U12178 : NOR3_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_state_0_port,
                           A2 => n838, A3 => n10868, ZN => n10856);
   U12179 : NAND2_X1 port map( A1 => n8722, A2 => n8721, ZN => n8723);
   U12180 : INV_X1 port map( A => n10473, ZN => n10466);
   U12181 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n639, B => n9909, ZN => 
                           n9519);
   U12182 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n843, B => n10046, ZN =>
                           n9508);
   U12183 : INV_X1 port map( A => n9742, ZN => n10024);
   U12184 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n537, B => n9839, ZN => 
                           n9523);
   U12185 : INV_X1 port map( A => n10010, ZN => n10012);
   U12186 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_20_port, A2 => n8671, 
                           ZN => n10123);
   U12187 : INV_X1 port map( A => n10123, ZN => n10122);
   U12188 : INV_X1 port map( A => n9669, ZN => n10326);
   U12189 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n945, B => n10124, ZN =>
                           n9501);
   U12190 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n1047, B => n10198, ZN 
                           => n9494);
   U12191 : XNOR2_X1 port map( A => DP_OP_751_130_5637_n741, B => n9969, ZN => 
                           n9512);
   U12192 : XNOR2_X1 port map( A => n10313, B => DP_OP_751_130_5637_n1149, ZN 
                           => n9487);
   U12193 : AND2_X1 port map( A1 => IRAM_ADDRESS_17_port, A2 => n12065, ZN => 
                           n8309);
   U12194 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_17_port, A2 => n8671, 
                           ZN => n10223);
   U12195 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_16_port, A2 => n8671, 
                           ZN => n10312);
   U12196 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_22_port, A2 => n8672, 
                           ZN => n10044);
   U12197 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_30_port, A2 => n8674, 
                           ZN => n9761);
   U12198 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_27_port, A2 => n8672, 
                           ZN => n9874);
   U12199 : INV_X1 port map( A => i_RD1_4_port, ZN => n9047);
   U12200 : NAND2_X1 port map( A1 => n8681, A2 => n10870, ZN => n12087);
   U12201 : INV_X1 port map( A => n9533, ZN => n9553);
   U12202 : OAI21_X1 port map( B1 => n9517, B2 => DP_OP_751_130_5637_n639, A =>
                           n9516, ZN => n9518);
   U12203 : NAND2_X1 port map( A1 => n10273, A2 => n10021, ZN => n9455);
   U12204 : AND4_X1 port map( A1 => n10789, A2 => n10742, A3 => IR_4_port, A4 
                           => n10741, ZN => n8329);
   U12205 : OR2_X1 port map( A1 => IRAM_ADDRESS_17_port, A2 => n12065, ZN => 
                           n8367);
   U12206 : AND3_X1 port map( A1 => n12208, A2 => n10725, A3 => DRAMRF_READY, 
                           ZN => n8371);
   U12207 : INV_X1 port map( A => n8447, ZN => n8446);
   U12208 : AOI21_X1 port map( B1 => n8962, B2 => n8771, A => n8751, ZN => 
                           n11399);
   U12209 : AOI21_X1 port map( B1 => n8964, B2 => n8901, A => n8899, ZN => 
                           n11708);
   U12210 : AOI21_X1 port map( B1 => n8962, B2 => n8971, A => n8961, ZN => 
                           n11832);
   U12211 : AND2_X1 port map( A1 => n10730, A2 => n8696, ZN => n8379);
   U12212 : NOR2_X1 port map( A1 => n10021, A2 => n12087, ZN => n10240);
   U12213 : AND4_X1 port map( A1 => n9418, A2 => n9417, A3 => n9416, A4 => 
                           n9415, ZN => n8408);
   U12214 : NAND2_X1 port map( A1 => n8400, A2 => i_ALU_OP_1_port, ZN => n8412)
                           ;
   U12215 : INV_X1 port map( A => n12022, ZN => n8973);
   U12216 : INV_X1 port map( A => i_RD1_2_port, ZN => n9029);
   U12217 : INV_X1 port map( A => i_RD1_10_port, ZN => n9077);
   U12218 : INV_X1 port map( A => i_RD1_3_port, ZN => n9045);
   U12219 : INV_X1 port map( A => i_RD1_0_port, ZN => n9240);
   U12220 : NAND3_X1 port map( A1 => n9647, A2 => n8452, A3 => n9646, ZN => 
                           DP_OP_1090J1_126_7243_n75);
   U12221 : AND2_X1 port map( A1 => n10634, A2 => n8449, ZN => n8448);
   U12222 : NAND2_X1 port map( A1 => n9317, A2 => n8451, ZN => n8449);
   U12223 : INV_X1 port map( A => n9321, ZN => n8450);
   U12224 : OR2_X1 port map( A1 => n10638, A2 => n8381, ZN => n8451);
   U12225 : INV_X1 port map( A => C620_DATA2_31, ZN => n8453);
   U12226 : NAND3_X1 port map( A1 => n8454, A2 => n8699, A3 => n8255, ZN => 
                           n9005);
   U12227 : AOI21_X1 port map( B1 => n10529, B2 => n8687, A => n9014, ZN => 
                           n9019);
   U12228 : INV_X1 port map( A => n8443, ZN => n8714);
   U12229 : AOI22_X1 port map( A1 => n10872, A2 => n10453, B1 => 
                           DataPath_i_PIPLIN_IN2_7_port, B2 => n10871, ZN => 
                           n2486);
   U12230 : BUF_X1 port map( A => n9315, Z => n8483);
   U12231 : INV_X1 port map( A => n8485, ZN => n8486);
   U12232 : XNOR2_X1 port map( A => DP_OP_751_130_5637_I2, B => n9563, ZN => 
                           n9450);
   U12233 : NAND2_X1 port map( A1 => n8977, A2 => n8976, ZN => n8498);
   U12234 : NAND2_X1 port map( A1 => n8498, A2 => n8499, ZN => n9647);
   U12235 : AND2_X1 port map( A1 => n8371, A2 => n11375, ZN => n8499);
   U12236 : INV_X1 port map( A => n10740, ZN => n10724);
   U12237 : NAND2_X1 port map( A1 => n9271, A2 => n8699, ZN => n8500);
   U12238 : INV_X1 port map( A => n10824, ZN => n10831);
   U12239 : NAND2_X1 port map( A1 => n9283, A2 => n9284, ZN => n10684);
   U12240 : NAND2_X1 port map( A1 => n9282, A2 => IRAM_ADDRESS_3_port, ZN => 
                           n10686);
   U12241 : OAI21_X1 port map( B1 => n9263, B2 => n9262, A => n10824, ZN => 
                           n9270);
   U12242 : NAND2_X1 port map( A1 => n9019, A2 => i_RD1_6_port, ZN => n9060);
   U12243 : OAI22_X1 port map( A1 => n8062, A2 => n10719, B1 => n10718, B2 => 
                           n10717, ZN => CU_I_CW_23_port);
   U12244 : INV_X1 port map( A => n10770, ZN => n10722);
   U12245 : NOR2_X1 port map( A1 => n8062, A2 => n10713, ZN => CU_I_CW_4_port);
   U12246 : NAND2_X1 port map( A1 => n10791, A2 => n8062, ZN => n10792);
   U12247 : XNOR2_X1 port map( A => n8252, B => n10662, ZN => n10663);
   U12248 : XNOR2_X1 port map( A => n10696, B => n8082, ZN => n10697);
   U12249 : AOI21_X1 port map( B1 => n8082, B2 => n10693, A => n10692, ZN => 
                           n10690);
   U12250 : AOI21_X1 port map( B1 => n10770, B2 => n8185, A => n10769, ZN => 
                           n10773);
   U12251 : NAND2_X1 port map( A1 => n10770, A2 => n8110, ZN => n9266);
   U12252 : NAND2_X1 port map( A1 => n10717, A2 => n9649, ZN => n10541);
   U12253 : OAI21_X1 port map( B1 => n8254, B2 => n10823, A => n10822, ZN => 
                           n7108);
   U12254 : NOR2_X1 port map( A1 => n10763, A2 => n8254, ZN => n10850);
   U12255 : AOI22_X1 port map( A1 => n10872, A2 => n10516, B1 => 
                           DataPath_i_PIPLIN_IN2_2_port, B2 => n10871, ZN => 
                           n2494);
   U12256 : NOR3_X1 port map( A1 => n8177, A2 => IRAM_DATA(28), A3 => n12020, 
                           ZN => n10797);
   U12257 : XNOR2_X1 port map( A => n8096, B => n10591, ZN => n10594);
   U12258 : NAND2_X1 port map( A1 => n9280, A2 => n10698, ZN => n10695);
   U12259 : OAI211_X1 port map( C1 => n8139, C2 => n8373, A => n7697, B => 
                           n9176, ZN => n10000);
   U12260 : OAI211_X1 port map( C1 => n8139, C2 => n8372, A => n7698, B => 
                           n8987, ZN => n9790);
   U12261 : OAI211_X1 port map( C1 => n572, C2 => n8139, A => n7697, B => n8993
                           , ZN => n9812);
   U12262 : OAI211_X1 port map( C1 => n570, C2 => n8139, A => n7698, B => n9181
                           , ZN => n9902);
   U12263 : OAI211_X1 port map( C1 => n8139, C2 => n8374, A => n7697, B => 
                           n9153, ZN => n10070);
   U12264 : OAI211_X1 port map( C1 => n560, C2 => n8139, A => n7697, B => n9115
                           , ZN => n10248);
   U12265 : OAI211_X1 port map( C1 => n556, C2 => n8139, A => n9094, B => n9093
                           , ZN => n10535);
   U12266 : OAI211_X1 port map( C1 => n562, C2 => n8139, A => n7698, B => n9124
                           , ZN => n10173);
   U12267 : OAI211_X1 port map( C1 => n8139, C2 => n8375, A => n7697, B => 
                           n9121, ZN => n10212);
   U12268 : OAI22_X1 port map( A1 => n10797, A2 => n10808, B1 => n181, B2 => 
                           n10823, ZN => n7107);
   U12269 : OR2_X1 port map( A1 => n10751, A2 => n8255, ZN => n10747);
   U12270 : AND2_X1 port map( A1 => n8502, A2 => n181, ZN => n10746);
   U12271 : NAND2_X1 port map( A1 => IR_26_port, A2 => n181, ZN => n8704);
   U12272 : NAND2_X1 port map( A1 => n8255, A2 => IR_26_port, ZN => n10756);
   U12273 : NOR2_X1 port map( A1 => n8313, A2 => n477, ZN => n10725);
   U12274 : NOR2_X1 port map( A1 => n10731, A2 => n10846, ZN => 
                           DRAMRF_READNOTWRITE_port);
   U12275 : NOR3_X1 port map( A1 => n10731, A2 => n7773, A3 => 
                           DP_OP_1090J1_126_7243_n72, ZN => n10732);
   U12276 : NOR2_X1 port map( A1 => n10731, A2 => RST, ZN => n10845);
   U12277 : XNOR2_X1 port map( A => n10701, B => n7994, ZN => n10703);
   U12278 : XNOR2_X1 port map( A => n8018, B => n10657, ZN => n10659);
   U12279 : NAND2_X1 port map( A1 => n9311, A2 => n9310, ZN => n10649);
   U12280 : NAND2_X1 port map( A1 => n10700, A2 => n10699, ZN => n9280);
   U12281 : NOR4_X1 port map( A1 => n9257, A2 => n9254, A3 => n9255, A4 => 
                           n9256, ZN => n9258);
   U12282 : OAI211_X1 port map( C1 => n9065, C2 => n9064, A => n9256, B => 
                           n9063, ZN => n9091);
   U12283 : INV_X1 port map( A => n9271, ZN => n10719);
   U12284 : INV_X1 port map( A => n8982, ZN => n10731);
   U12285 : XNOR2_X1 port map( A => n8249, B => n10665, ZN => n10667);
   U12286 : XNOR2_X1 port map( A => n8248, B => n10639, ZN => n10640);
   U12287 : XNOR2_X1 port map( A => n10580, B => n10579, ZN => n10581);
   U12288 : OAI211_X1 port map( C1 => n190, C2 => n8190, A => n8711, B => n8709
                           , ZN => i_ADD_WS1_3_port);
   U12289 : NAND2_X1 port map( A1 => n10676, A2 => n10674, ZN => n9289);
   U12290 : INV_X1 port map( A => n9278, ZN => n9279);
   U12291 : NAND2_X1 port map( A1 => n9278, A2 => IRAM_ADDRESS_1_port, ZN => 
                           n10699);
   U12292 : NAND2_X1 port map( A1 => n9228, A2 => n9227, ZN => n9229);
   U12293 : NAND2_X1 port map( A1 => n7692, A2 => IR_13_port, ZN => n9093);
   U12294 : NAND2_X1 port map( A1 => n7692, A2 => IR_9_port, ZN => n9066);
   U12295 : NAND2_X1 port map( A1 => n7693, A2 => IR_5_port, ZN => n9000);
   U12296 : NAND2_X1 port map( A1 => n7693, A2 => IR_3_port, ZN => n9037);
   U12297 : OAI211_X1 port map( C1 => n8190, C2 => n9007, A => n10519, B => 
                           n9006, ZN => n9009);
   U12298 : NAND2_X1 port map( A1 => n7693, A2 => IR_1_port, ZN => n9021);
   U12299 : NAND2_X1 port map( A1 => n7693, A2 => IR_7_port, ZN => n9015);
   U12300 : AOI22_X1 port map( A1 => n10872, A2 => n10529, B1 => 
                           DataPath_i_PIPLIN_IN2_6_port, B2 => n10871, ZN => 
                           n10530);
   U12301 : XNOR2_X1 port map( A => n10597, B => n10596, ZN => n10598);
   U12302 : OAI21_X1 port map( B1 => n10653, B2 => n222, A => n10651, ZN => 
                           n9311);
   U12303 : OR2_X1 port map( A1 => n8484, A2 => n8406, ZN => n9312);
   U12304 : OR2_X1 port map( A1 => n8484, A2 => n196, ZN => n10651);
   U12305 : OR2_X1 port map( A1 => n8192, A2 => n197, ZN => n10656);
   U12306 : NAND2_X1 port map( A1 => n9296, A2 => IRAM_ADDRESS_8_port, ZN => 
                           n9297);
   U12307 : OAI21_X1 port map( B1 => n9296, B2 => IRAM_ADDRESS_8_port, A => 
                           n9295, ZN => n9298);
   U12308 : OR2_X1 port map( A1 => n8484, A2 => n8407, ZN => n9299);
   U12309 : NOR2_X1 port map( A1 => n8192, A2 => n8324, ZN => n9295);
   U12310 : NOR2_X1 port map( A1 => n8484, A2 => n8332, ZN => n10664);
   U12311 : NOR2_X1 port map( A1 => n8484, A2 => n9290, ZN => n10669);
   U12312 : OAI21_X1 port map( B1 => n8192, B2 => n8307, A => n8366, ZN => 
                           n10668);
   U12313 : OR2_X1 port map( A1 => n8192, A2 => n8320, ZN => n9287);
   U12314 : OR2_X1 port map( A1 => n8484, A2 => n8317, ZN => n9286);
   U12315 : NAND2_X1 port map( A1 => n10704, A2 => IRAM_ADDRESS_0_port, ZN => 
                           n10700);
   U12316 : OR2_X1 port map( A1 => n8484, A2 => IR_2_port, ZN => n9281);
   U12317 : NOR2_X1 port map( A1 => n8484, A2 => n8318, ZN => n9282);
   U12318 : NOR2_X1 port map( A1 => n8483, A2 => n8315, ZN => n9278);
   U12319 : NOR2_X1 port map( A1 => n8483, A2 => n210, ZN => n10704);
   U12320 : NAND2_X1 port map( A1 => n10524, A2 => n10523, ZN => n9261);
   U12321 : OAI211_X1 port map( C1 => n195, C2 => n9108, A => n9099, B => n9098
                           , ZN => n10537);
   U12322 : OAI211_X1 port map( C1 => n194, C2 => n9108, A => n9107, B => n9106
                           , ZN => n10325);
   U12323 : OAI211_X1 port map( C1 => n196, C2 => n9108, A => n9085, B => n9084
                           , ZN => n10382);
   U12324 : OAI211_X1 port map( C1 => n197, C2 => n9108, A => n9071, B => n9070
                           , ZN => n10391);
   U12325 : OAI211_X1 port map( C1 => n9108, C2 => n8324, A => n9056, B => 
                           n9055, ZN => n10531);
   U12326 : OAI211_X1 port map( C1 => n9108, C2 => n8323, A => n9075, B => 
                           n9074, ZN => n10533);
   U12327 : OAI211_X1 port map( C1 => n210, C2 => n9108, A => n9031, B => n9030
                           , ZN => n10518);
   U12328 : OAI211_X1 port map( C1 => n9108, C2 => n8307, A => n9013, B => 
                           n9012, ZN => n10529);
   U12329 : NOR2_X1 port map( A1 => n10713, A2 => n176, ZN => CU_I_CW_6_port);
   U12330 : NAND2_X1 port map( A1 => n10713, A2 => n8455, ZN => n10717);
   U12331 : INV_X1 port map( A => n10524, ZN => n10526);
   U12332 : OAI211_X1 port map( C1 => n10634, C2 => n10633, A => n10632, B => 
                           n8303, ZN => n10637);
   U12333 : XNOR2_X1 port map( A => n8040, B => n10652, ZN => n10655);
   U12334 : XNOR2_X1 port map( A => n10704, B => n230, ZN => n10705);
   U12335 : XNOR2_X1 port map( A => n8029, B => n9293, ZN => n9294);
   U12336 : OAI22_X1 port map( A1 => n8253, A2 => n10587, B1 => 
                           IRAM_ADDRESS_26_port, B2 => n10590, ZN => n10584);
   U12337 : OAI21_X1 port map( B1 => n10628, B2 => n10619, A => n10626, ZN => 
                           n10623);
   U12338 : OAI21_X1 port map( B1 => n10628, B2 => n10612, A => n10611, ZN => 
                           n10616);
   U12339 : INV_X1 port map( A => n10628, ZN => n10602);
   U12340 : NOR3_X1 port map( A1 => n10772, A2 => n8455, A3 => n8973, ZN => 
                           n10783);
   U12341 : NOR4_X1 port map( A1 => n10768, A2 => n8084, A3 => n8455, A4 => 
                           n8254, ZN => n10769);
   U12342 : OR2_X1 port map( A1 => n8484, A2 => n195, ZN => n9316);
   U12343 : NAND2_X1 port map( A1 => n10653, A2 => n222, ZN => n9310);
   U12344 : NOR2_X1 port map( A1 => n8192, A2 => n8323, ZN => n10661);
   U12345 : OR2_X1 port map( A1 => n8084, A2 => n176, ZN => n8984);
   U12346 : INV_X1 port map( A => n7767, ZN => n8551);
   U12347 : INV_X1 port map( A => n7769, ZN => n8553);
   U12348 : INV_X1 port map( A => n7772, ZN => n8557);
   U12349 : INV_X1 port map( A => n7772, ZN => n8558);
   U12350 : INV_X1 port map( A => n8560, ZN => n8561);
   U12351 : INV_X1 port map( A => n8561, ZN => n8562);
   U12352 : INV_X1 port map( A => n8564, ZN => n8565);
   U12353 : INV_X1 port map( A => n8564, ZN => n8566);
   U12354 : NOR2_X1 port map( A1 => n10927, A2 => n10913, ZN => n8582);
   U12355 : NOR2_X1 port map( A1 => n10927, A2 => n10912, ZN => n8585);
   U12356 : NOR2_X1 port map( A1 => n10927, A2 => n10912, ZN => n8586);
   U12357 : NOR2_X1 port map( A1 => n10922, A2 => n10912, ZN => n8587);
   U12358 : NOR2_X1 port map( A1 => n10922, A2 => n10912, ZN => n8588);
   U12359 : NOR2_X1 port map( A1 => n10923, A2 => n10913, ZN => n8589);
   U12360 : NOR2_X1 port map( A1 => n10923, A2 => n10913, ZN => n8590);
   U12361 : NOR2_X1 port map( A1 => n10925, A2 => n10913, ZN => n8592);
   U12362 : NOR2_X1 port map( A1 => n10925, A2 => n10913, ZN => n8593);
   U12363 : NOR2_X1 port map( A1 => n10926, A2 => n10922, ZN => n8596);
   U12364 : NOR2_X1 port map( A1 => n10924, A2 => n10925, ZN => n8599);
   U12365 : NOR2_X1 port map( A1 => n10924, A2 => n10925, ZN => n8600);
   U12366 : NOR2_X1 port map( A1 => n10926, A2 => n10923, ZN => n8601);
   U12367 : NOR2_X1 port map( A1 => n10926, A2 => n10923, ZN => n8602);
   U12368 : NOR2_X1 port map( A1 => n10924, A2 => n10923, ZN => n8603);
   U12369 : NOR2_X1 port map( A1 => n10924, A2 => n10923, ZN => n8604);
   U12370 : NOR2_X1 port map( A1 => n10926, A2 => n10925, ZN => n8605);
   U12371 : NOR2_X1 port map( A1 => n10926, A2 => n10925, ZN => n8606);
   U12372 : NOR2_X1 port map( A1 => n10927, A2 => n10926, ZN => n8607);
   U12373 : NOR2_X1 port map( A1 => n10927, A2 => n10926, ZN => n8608);
   U12374 : INV_X1 port map( A => n8675, ZN => n8674);
   U12375 : MUX2_X1 port map( A => n6146, B => n8423, S => n10740, Z => n8960);
   U12376 : NAND3_X1 port map( A1 => n9643, A2 => n8692, A3 => n8957, ZN => 
                           n8749);
   U12377 : MUX2_X1 port map( A => n6126, B => n8424, S => n10740, Z => n8962);
   U12378 : MUX2_X1 port map( A => n6052, B => n8425, S => n10740, Z => n8964);
   U12379 : MUX2_X1 port map( A => n5978, B => n8426, S => n10740, Z => n8967);
   U12380 : MUX2_X1 port map( A => n5941, B => n8401, S => n10740, Z => n8969);
   U12381 : MUX2_X1 port map( A => n8770, B => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_15_port, S => 
                           n10740, Z => n8972);
   U12382 : NAND3_X1 port map( A1 => n7685, A2 => n10519, A3 => n9004, ZN => 
                           n8985);
   U12383 : NAND3_X1 port map( A1 => n7685, A2 => IR_4_port, A3 => n9004, ZN =>
                           n9007);
   U12384 : FA_X1 port map( A => n9049, B => n10678, CI => n9244, CO => n9065, 
                           S => n_3950);
   U12385 : NAND3_X1 port map( A1 => n9160, A2 => n9167, A3 => n9168, ZN => 
                           n9254);
   U12386 : MUX2_X1 port map( A => i_RD2_27_port, B => n9902, S => n8686, Z => 
                           n9186);
   U12387 : MUX2_X1 port map( A => n9231, B => n9230, S => n9229, Z => n10524);
   U12388 : NAND3_X1 port map( A1 => n7778, A2 => n9238, A3 => n9239, ZN => 
                           n9252);
   U12389 : NAND3_X1 port map( A1 => n9245, A2 => n9244, A3 => n9243, ZN => 
                           n9251);
   U12390 : NAND3_X1 port map( A1 => n9249, A2 => n9248, A3 => n9247, ZN => 
                           n9250);
   U12391 : MUX2_X1 port map( A => n10543, B => n10826, S => n9261, Z => n9263)
                           ;
   U12392 : MUX2_X1 port map( A => n10707, B => n9276, S => n10524, Z => n9262)
                           ;
   U12393 : NAND3_X1 port map( A1 => n10523, A2 => n8062, A3 => n10827, ZN => 
                           n9265);
   U12394 : NAND3_X1 port map( A1 => n10695, A2 => n10686, A3 => n10693, ZN => 
                           n9284);
   U12395 : NAND3_X1 port map( A1 => n10571, A2 => n9319, A3 => n220, ZN => 
                           n9320);
   U12396 : XOR2_X1 port map( A => n9327, B => n9326, Z => n12067);
   U12397 : XOR2_X1 port map( A => n10546, B => n9332, Z => n12069);
   U12398 : NAND3_X1 port map( A1 => n9353, A2 => n9435, A3 => n9352, ZN => 
                           n9917);
   U12399 : NAND3_X1 port map( A1 => n9613, A2 => n9543, A3 => n8385, ZN => 
                           n9355);
   U12400 : NAND3_X1 port map( A1 => n9404, A2 => n9435, A3 => n9403, ZN => 
                           n10090);
   U12401 : NAND3_X1 port map( A1 => n9551, A2 => n8486, A3 => n8167, ZN => 
                           n10388);
   U12402 : NAND3_X1 port map( A1 => n7785, A2 => n9612, A3 => n12086, ZN => 
                           n9415);
   U12403 : NAND3_X1 port map( A1 => n9422, A2 => n9435, A3 => n9421, ZN => 
                           n10110);
   U12404 : MUX2_X1 port map( A => n10273, B => n10021, S => n8676, Z => n9454)
                           ;
   U12405 : MUX2_X1 port map( A => n8676, B => n415, S => n9626, Z => n9457);
   U12406 : NAND3_X1 port map( A1 => n10469, A2 => n9561, A3 => n9560, ZN => 
                           n9565);
   U12407 : NAND3_X1 port map( A1 => n10458, A2 => n8099, A3 => n9562, ZN => 
                           n9564);
   U12408 : NAND3_X1 port map( A1 => n9593, A2 => n9592, A3 => n9591, ZN => 
                           n9600);
   U12409 : NAND3_X1 port map( A1 => n9633, A2 => n9632, A3 => n9631, ZN => 
                           n10428);
   U12410 : NAND3_X1 port map( A1 => n9657, A2 => n9656, A3 => n9655, ZN => 
                           n9662);
   U12411 : NAND3_X1 port map( A1 => n9699, A2 => n9932, A3 => n9871, ZN => 
                           n9703);
   U12412 : NAND3_X1 port map( A1 => n10023, A2 => n10113, A3 => n10025, ZN => 
                           n9783);
   U12413 : MUX2_X1 port map( A => n10468, B => n10458, S => n9839, Z => n9837)
                           ;
   U12414 : MUX2_X1 port map( A => n10488, B => n10465, S => n9839, Z => n9840)
                           ;
   U12415 : XOR2_X1 port map( A => n9872, B => n9867, Z => n9882);
   U12416 : NAND3_X1 port map( A1 => n10469, A2 => n9875, A3 => n9874, ZN => 
                           n9877);
   U12417 : NAND3_X1 port map( A1 => n10458, A2 => n7797, A3 => 
                           DP_OP_751_130_5637_n537, ZN => n9876);
   U12418 : XOR2_X1 port map( A => n9905, B => n9904, Z => n9906);
   U12419 : MUX2_X1 port map( A => n9911, B => n9910, S => n9909, Z => n9912);
   U12420 : NAND3_X1 port map( A1 => n10469, A2 => n7790, A3 => n9944, ZN => 
                           n9940);
   U12421 : NAND3_X1 port map( A1 => n10458, A2 => n9938, A3 => 
                           DP_OP_751_130_5637_n639, ZN => n9939);
   U12422 : NAND3_X1 port map( A1 => n9958, A2 => n9957, A3 => n9956, ZN => 
                           n9959);
   U12423 : MUX2_X1 port map( A => n10465, B => n10488, S => n9979, Z => n9971)
                           ;
   U12424 : MUX2_X1 port map( A => n9971, B => n9970, S => n9969, Z => n9972);
   U12425 : NAND3_X1 port map( A1 => n10469, A2 => n10011, A3 => n10010, ZN => 
                           n10014);
   U12426 : NAND3_X1 port map( A1 => n10458, A2 => n10012, A3 => 
                           DP_OP_751_130_5637_n741, ZN => n10013);
   U12427 : MUX2_X1 port map( A => n10465, B => n10488, S => n8553, Z => n10048
                           );
   U12428 : MUX2_X1 port map( A => n10048, B => n10047, S => n10046, Z => 
                           n10049);
   U12429 : NAND3_X1 port map( A1 => n10469, A2 => n10076, A3 => n8556, ZN => 
                           n10078);
   U12430 : NAND3_X1 port map( A1 => n10458, A2 => n10082, A3 => 
                           DP_OP_751_130_5637_n843, ZN => n10077);
   U12431 : MUX2_X1 port map( A => n10469, B => n10468, S => n10122, Z => 
                           n10126);
   U12432 : MUX2_X1 port map( A => n10458, B => n10468, S => n10123, Z => 
                           n10125);
   U12433 : MUX2_X1 port map( A => n10126, B => n10125, S => n10124, Z => 
                           n10127);
   U12434 : XOR2_X1 port map( A => n10141, B => n10138, Z => n10152);
   U12435 : NAND3_X1 port map( A1 => n10469, A2 => n10144, A3 => n10143, ZN => 
                           n10146);
   U12436 : NAND3_X1 port map( A1 => n10458, A2 => n8552, A3 => 
                           DP_OP_751_130_5637_n945, ZN => n10145);
   U12437 : NAND3_X1 port map( A1 => n10196, A2 => n10195, A3 => n10194, ZN => 
                           n10202);
   U12438 : MUX2_X1 port map( A => n10468, B => n10469, S => n10197, Z => 
                           n10200);
   U12439 : MUX2_X1 port map( A => n10200, B => n10199, S => n10198, Z => 
                           n10201);
   U12440 : NAND3_X1 port map( A1 => n10318, A2 => n10203, A3 => n10204, ZN => 
                           n10207);
   U12441 : NAND3_X1 port map( A1 => n10318, A2 => n10205, A3 => n10204, ZN => 
                           n10206);
   U12442 : NAND3_X1 port map( A1 => n10469, A2 => n10217, A3 => n8550, ZN => 
                           n10219);
   U12443 : NAND3_X1 port map( A1 => n10458, A2 => n7767, A3 => 
                           DP_OP_751_130_5637_n1047, ZN => n10218);
   U12444 : NAND3_X1 port map( A1 => n10243, A2 => n10242, A3 => n10241, ZN => 
                           n10244);
   U12445 : XOR2_X1 port map( A => n10260, B => n10259, Z => n10270);
   U12446 : NAND3_X1 port map( A1 => n10346, A2 => n10267, A3 => n10266, ZN => 
                           n10268);
   U12447 : NAND3_X1 port map( A1 => n10311, A2 => n10310, A3 => n10309, ZN => 
                           n10317);
   U12448 : MUX2_X1 port map( A => n10469, B => n10468, S => n7772, Z => n10315
                           );
   U12449 : MUX2_X1 port map( A => n10458, B => n10468, S => n8557, Z => n10314
                           );
   U12450 : MUX2_X1 port map( A => n10315, B => n10314, S => n10313, Z => 
                           n10316);
   U12451 : MUX2_X1 port map( A => n10458, B => n10468, S => n8493, Z => n10336
                           );
   U12452 : MUX2_X1 port map( A => n10465, B => n10488, S => n8493, Z => n10327
                           );
   U12453 : NAND3_X1 port map( A1 => n10469, A2 => n8555, A3 => n7793, ZN => 
                           n10353);
   U12454 : NAND3_X1 port map( A1 => n10458, A2 => n10351, A3 => 
                           DP_OP_751_130_5637_n1251, ZN => n10352);
   U12455 : NAND3_X1 port map( A1 => n10469, A2 => n10395, A3 => n7771, ZN => 
                           n10397);
   U12456 : NAND3_X1 port map( A1 => n10458, A2 => n8093, A3 => 
                           DP_OP_751_130_5637_n1455, ZN => n10396);
   U12457 : MUX2_X1 port map( A => n10465, B => n10489, S => n10419, Z => 
                           n10417);
   U12458 : MUX2_X1 port map( A => n10488, B => n10465, S => n10419, Z => 
                           n10420);
   U12459 : MUX2_X1 port map( A => n10425, B => n10424, S => n10423, Z => 
                           n10426);
   U12460 : XOR2_X1 port map( A => IRAM_ADDRESS_28_port, B => n10590, Z => 
                           n10579);
   U12461 : XOR2_X1 port map( A => n10587, B => n8253, Z => n10589);
   U12462 : XOR2_X1 port map( A => n10629, B => n10628, Z => n10630);
   U12463 : XOR2_X1 port map( A => n10677, B => n8251, Z => n10679);
   U12464 : NAND3_X1 port map( A1 => n8185, A2 => n10707, A3 => n8080, ZN => 
                           n10708);
   U12465 : NAND3_X1 port map( A1 => n10723, A2 => n10722, A3 => n10721, ZN => 
                           CU_I_CW_25_port);
   U12466 : NAND3_X1 port map( A1 => n10790, A2 => n12029, A3 => n10743, ZN => 
                           n10745);
   U12467 : NAND3_X1 port map( A1 => n10790, A2 => n210, A3 => n10789, ZN => 
                           n10749);
   U12468 : NAND3_X1 port map( A1 => n10790, A2 => n8428, A3 => n10750, ZN => 
                           n10755);
   U12469 : NAND3_X1 port map( A1 => n10752, A2 => n181, A3 => n10753, ZN => 
                           n10754);
   U12470 : NAND3_X1 port map( A1 => n10760, A2 => n10777, A3 => n8427, ZN => 
                           n10761);
   U12471 : NAND3_X1 port map( A1 => n10790, A2 => n10789, A3 => n8427, ZN => 
                           n10793);
   DataPath_RF_bus_complete_win_data_0_port <= '0';
   U12473 : NOR2_X1 port map( A1 => n8084, A2 => n181, ZN => n12022);
   U12474 : NAND2_X1 port map( A1 => n8084, A2 => n8080, ZN => n10873);
   U12475 : NAND2_X1 port map( A1 => n8254, A2 => n8062, ZN => n12026);
   U12476 : AND2_X1 port map( A1 => n10857, A2 => CU_I_CW_MEM_0_port, ZN => 
                           CU_I_N170);
   U12477 : AND2_X1 port map( A1 => n10857, A2 => CU_I_CW_MEM_1_port, ZN => 
                           CU_I_N171);
   U12478 : OAI22_X1 port map( A1 => n821, A2 => DataPath_RF_c_win_1_port, B1 
                           => DataPath_RF_c_win_2_port, B2 => n822, ZN => 
                           n10874);
   U12479 : AOI221_X1 port map( B1 => n821, B2 => DataPath_RF_c_win_1_port, C1 
                           => n822, C2 => DataPath_RF_c_win_2_port, A => n10874
                           , ZN => n10875);
   U12480 : NAND2_X1 port map( A1 => CU_I_CW_ID_19, A2 => n10877, ZN => n11950)
                           ;
   U12481 : NOR2_X1 port map( A1 => n473, A2 => n11950, ZN => DECODEhw_i_WR1);
   U12482 : XOR2_X1 port map( A => n838, B => 
                           DataPath_RF_PUSH_ADDRGEN_curr_state_0_port, Z => 
                           n12045);
   U12483 : NAND2_X1 port map( A1 => n10890, A2 => n10894, ZN => n10882);
   U12484 : NAND2_X1 port map( A1 => n10900, A2 => n10889, ZN => n10883);
   U12485 : NOR2_X1 port map( A1 => n10882, A2 => n10883, ZN => n10879);
   U12486 : NAND2_X1 port map( A1 => n10898, A2 => n10904, ZN => n10886);
   U12487 : INV_X1 port map( A => n10886, ZN => n10878);
   U12488 : AND2_X1 port map( A1 => n10888, A2 => n10902, ZN => n10885);
   U12489 : NAND2_X1 port map( A1 => n10878, A2 => n10885, ZN => n10909);
   U12490 : NAND2_X1 port map( A1 => n10854, A2 => n10853, ZN => n10880);
   U12491 : NOR2_X1 port map( A1 => n10880, A2 => n10887, ZN => n10910);
   U12492 : AOI21_X1 port map( B1 => n10856, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_14_port, A => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_15_port, ZN => 
                           n11394);
   U12493 : NAND2_X1 port map( A1 => n11394, A2 => n10891, ZN => n10881);
   U12494 : NAND2_X1 port map( A1 => n10892, A2 => n10896, ZN => n10884);
   U12495 : INV_X1 port map( A => n10879, ZN => n10907);
   U12496 : NOR2_X1 port map( A1 => n10909, A2 => n10911, ZN => n10908);
   U12497 : NAND2_X1 port map( A1 => n10879, A2 => n10908, ZN => n10927);
   U12498 : OAI21_X1 port map( B1 => n11394, B2 => n10893, A => n10892, ZN => 
                           n10895);
   U12499 : OAI221_X1 port map( B1 => n10897, B2 => n10896, C1 => n10897, C2 =>
                           n10895, A => n10894, ZN => n10899);
   U12500 : OAI221_X1 port map( B1 => n10901, B2 => n10900, C1 => n10901, C2 =>
                           n10899, A => n10898, ZN => n10903);
   U12501 : OAI221_X1 port map( B1 => n10905, B2 => n10904, C1 => n10905, C2 =>
                           n10903, A => n10902, ZN => n10906);
   U12502 : NAND2_X1 port map( A1 => n10920, A2 => n10918, ZN => n10913);
   U12503 : NOR2_X1 port map( A1 => n10927, A2 => n10913, ZN => n11235);
   U12504 : NAND2_X1 port map( A1 => n10908, A2 => n10907, ZN => n10922);
   U12505 : AOI22_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_480_port, B1 => 
                           n11239, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_352_port, ZN => 
                           n10917);
   U12506 : INV_X1 port map( A => n10920, ZN => n10919);
   U12507 : NOR2_X1 port map( A1 => n10927, A2 => n10912, ZN => n11237);
   U12508 : AOI22_X1 port map( A1 => n8584, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_192_port, B1 => 
                           n8585, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_448_port, ZN => 
                           n10916);
   U12509 : NOR2_X1 port map( A1 => n10922, A2 => n10912, ZN => n11240);
   U12510 : NOR2_X1 port map( A1 => n10923, A2 => n10913, ZN => n11238);
   U12511 : AOI22_X1 port map( A1 => n8587, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_320_port, B1 => 
                           n8590, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_224_port, ZN => 
                           n10915);
   U12512 : NAND2_X1 port map( A1 => n10911, A2 => n10923, ZN => n10925);
   U12513 : NOR2_X1 port map( A1 => n10925, A2 => n10913, ZN => n11234);
   U12514 : AOI22_X1 port map( A1 => n8591, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_64_port, B1 => 
                           n8593, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_96_port, ZN => 
                           n10914);
   U12515 : NAND4_X1 port map( A1 => n10917, A2 => n10916, A3 => n10915, A4 => 
                           n10914, ZN => n10933);
   U12516 : NAND2_X1 port map( A1 => n10919, A2 => n10921, ZN => n10924);
   U12517 : NOR2_X1 port map( A1 => n10926, A2 => n10922, ZN => n11246);
   U12518 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_384_port, B1 => 
                           n8596, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_288_port, ZN => 
                           n10931);
   U12519 : NOR2_X1 port map( A1 => n10924, A2 => n10922, ZN => n11249);
   U12520 : NOR2_X1 port map( A1 => n10924, A2 => n10925, ZN => n11253);
   U12521 : AOI22_X1 port map( A1 => n8597, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_256_port, B1 => 
                           n8599, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_0_port, ZN => 
                           n10930);
   U12522 : NOR2_X1 port map( A1 => n10926, A2 => n10923, ZN => n11252);
   U12523 : NOR2_X1 port map( A1 => n10924, A2 => n10923, ZN => n11248);
   U12524 : AOI22_X1 port map( A1 => n8601, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_160_port, B1 => 
                           n8604, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_128_port, ZN => 
                           n10929);
   U12525 : NOR2_X1 port map( A1 => n10926, A2 => n10925, ZN => n11251);
   U12526 : NOR2_X1 port map( A1 => n10927, A2 => n10926, ZN => n11250);
   U12527 : AOI22_X1 port map( A1 => n8605, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_32_port, B1 => 
                           n8607, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_416_port, ZN => 
                           n10928);
   U12528 : NAND4_X1 port map( A1 => n10931, A2 => n10930, A3 => n10929, A4 => 
                           n10928, ZN => n10932);
   U12529 : OR2_X1 port map( A1 => n10933, A2 => n10932, ZN => 
                           DRAMRF_DATA_OUT(0));
   U12530 : AOI22_X1 port map( A1 => n11235, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_490_port, B1 => 
                           n8587, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_330_port, ZN => 
                           n10937);
   U12531 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_362_port, B1 => 
                           n11238, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_234_port, ZN => 
                           n10936);
   U12532 : AOI22_X1 port map( A1 => n8585, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_458_port, B1 => 
                           n11234, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_106_port, ZN => 
                           n10935);
   U12533 : AOI22_X1 port map( A1 => n8584, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_202_port, B1 => 
                           n8591, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_74_port, ZN => 
                           n10934);
   U12534 : NAND4_X1 port map( A1 => n10937, A2 => n10936, A3 => n10935, A4 => 
                           n10934, ZN => n10943);
   U12535 : AOI22_X1 port map( A1 => n11249, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_266_port, B1 => 
                           n8605, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_42_port, ZN => 
                           n10941);
   U12536 : AOI22_X1 port map( A1 => n11246, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_298_port, B1 => 
                           n11248, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_138_port, ZN => 
                           n10940);
   U12537 : AOI22_X1 port map( A1 => n8607, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_426_port, B1 => 
                           n8601, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_170_port, ZN => 
                           n10939);
   U12538 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_394_port, B1 => 
                           n8600, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_10_port, ZN => 
                           n10938);
   U12539 : NAND4_X1 port map( A1 => n10941, A2 => n10940, A3 => n10939, A4 => 
                           n10938, ZN => n10942);
   U12540 : OR2_X1 port map( A1 => n10943, A2 => n10942, ZN => 
                           DRAMRF_DATA_OUT(10));
   U12541 : AOI22_X1 port map( A1 => n11236, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_75_port, B1 => 
                           n8592, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_107_port, ZN => 
                           n10947);
   U12542 : AOI22_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_491_port, B1 => 
                           n11241, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_203_port, ZN => 
                           n10946);
   U12543 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_363_port, B1 => 
                           n8586, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_459_port, ZN => 
                           n10945);
   U12544 : AOI22_X1 port map( A1 => n8588, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_331_port, B1 => 
                           n11238, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_235_port, ZN => 
                           n10944);
   U12545 : NAND4_X1 port map( A1 => n10947, A2 => n10946, A3 => n10945, A4 => 
                           n10944, ZN => n10953);
   U12546 : AOI22_X1 port map( A1 => n8608, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_427_port, B1 => 
                           n8603, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_139_port, ZN => 
                           n10951);
   U12547 : AOI22_X1 port map( A1 => n8597, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_267_port, B1 => 
                           n8606, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_43_port, ZN => 
                           n10950);
   U12548 : AOI22_X1 port map( A1 => n8595, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_299_port, B1 => 
                           n11253, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_11_port, ZN => 
                           n10949);
   U12549 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_395_port, B1 => 
                           n8602, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_171_port, ZN => 
                           n10948);
   U12550 : NAND4_X1 port map( A1 => n10951, A2 => n10950, A3 => n10949, A4 => 
                           n10948, ZN => n10952);
   U12551 : OR2_X1 port map( A1 => n10953, A2 => n10952, ZN => 
                           DRAMRF_DATA_OUT(11));
   U12552 : AOI22_X1 port map( A1 => n8586, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_460_port, B1 => 
                           n8588, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_332_port, ZN => 
                           n10957);
   U12553 : AOI22_X1 port map( A1 => n11238, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_236_port, B1 => 
                           n8592, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_108_port, ZN => 
                           n10956);
   U12554 : AOI22_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_492_port, B1 => 
                           n11236, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_76_port, ZN => 
                           n10955);
   U12555 : AOI22_X1 port map( A1 => n11239, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_364_port, B1 => 
                           n11241, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_204_port, ZN => 
                           n10954);
   U12556 : NAND4_X1 port map( A1 => n10957, A2 => n10956, A3 => n10955, A4 => 
                           n10954, ZN => n10963);
   U12557 : AOI22_X1 port map( A1 => n11250, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_428_port, B1 => 
                           n11252, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_172_port, ZN => 
                           n10961);
   U12558 : AOI22_X1 port map( A1 => n8606, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_44_port, B1 => 
                           n8603, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_140_port, ZN => 
                           n10960);
   U12559 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_396_port, B1 => 
                           n11246, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_300_port, ZN => 
                           n10959);
   U12560 : AOI22_X1 port map( A1 => n8598, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_268_port, B1 => 
                           n11253, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_12_port, ZN => 
                           n10958);
   U12561 : NAND4_X1 port map( A1 => n10961, A2 => n10960, A3 => n10959, A4 => 
                           n10958, ZN => n10962);
   U12562 : OR2_X1 port map( A1 => n10963, A2 => n10962, ZN => 
                           DRAMRF_DATA_OUT(12));
   U12563 : AOI22_X1 port map( A1 => n8585, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_461_port, B1 => 
                           n8593, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_109_port, ZN => 
                           n10967);
   U12564 : AOI22_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_493_port, B1 => 
                           n8587, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_333_port, ZN => 
                           n10966);
   U12565 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_205_port, B1 => 
                           n8591, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_77_port, ZN => 
                           n10965);
   U12566 : AOI22_X1 port map( A1 => n11239, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_365_port, B1 => 
                           n8589, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_237_port, ZN => 
                           n10964);
   U12567 : NAND4_X1 port map( A1 => n10967, A2 => n10966, A3 => n10965, A4 => 
                           n10964, ZN => n10973);
   U12568 : AOI22_X1 port map( A1 => n8608, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_429_port, B1 => 
                           n8604, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_141_port, ZN => 
                           n10971);
   U12569 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_397_port, B1 => 
                           n11246, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_301_port, ZN => 
                           n10970);
   U12570 : AOI22_X1 port map( A1 => n8599, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_13_port, B1 => 
                           n8605, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_45_port, ZN => 
                           n10969);
   U12571 : AOI22_X1 port map( A1 => n8598, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_269_port, B1 => 
                           n11252, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_173_port, ZN => 
                           n10968);
   U12572 : NAND4_X1 port map( A1 => n10971, A2 => n10970, A3 => n10969, A4 => 
                           n10968, ZN => n10972);
   U12573 : OR2_X1 port map( A1 => n10973, A2 => n10972, ZN => 
                           DRAMRF_DATA_OUT(13));
   U12574 : AOI22_X1 port map( A1 => n8589, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_238_port, B1 => 
                           n8593, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_110_port, ZN => 
                           n10977);
   U12575 : AOI22_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_494_port, B1 => 
                           n11240, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_334_port, ZN => 
                           n10976);
   U12576 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_462_port, B1 => 
                           n11236, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_78_port, ZN => 
                           n10975);
   U12577 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_366_port, B1 => 
                           n8584, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_206_port, ZN => 
                           n10974);
   U12578 : NAND4_X1 port map( A1 => n10977, A2 => n10976, A3 => n10975, A4 => 
                           n10974, ZN => n10983);
   U12579 : AOI22_X1 port map( A1 => n8600, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_14_port, B1 => 
                           n8601, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_174_port, ZN => 
                           n10981);
   U12580 : AOI22_X1 port map( A1 => n8595, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_302_port, B1 => 
                           n11249, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_270_port, ZN => 
                           n10980);
   U12581 : AOI22_X1 port map( A1 => n11251, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_46_port, B1 => 
                           n8604, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_142_port, ZN => 
                           n10979);
   U12582 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_398_port, B1 => 
                           n8608, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_430_port, ZN => 
                           n10978);
   U12583 : NAND4_X1 port map( A1 => n10981, A2 => n10980, A3 => n10979, A4 => 
                           n10978, ZN => n10982);
   U12584 : OR2_X1 port map( A1 => n10983, A2 => n10982, ZN => 
                           DRAMRF_DATA_OUT(14));
   U12585 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_207_port, B1 => 
                           n11237, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_463_port, ZN => 
                           n10987);
   U12586 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_367_port, B1 => 
                           n8591, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_79_port, ZN => 
                           n10986);
   U12587 : AOI22_X1 port map( A1 => n11235, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_495_port, B1 => 
                           n8590, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_239_port, ZN => 
                           n10985);
   U12588 : AOI22_X1 port map( A1 => n11240, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_335_port, B1 => 
                           n11234, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_111_port, ZN => 
                           n10984);
   U12589 : NAND4_X1 port map( A1 => n10987, A2 => n10986, A3 => n10985, A4 => 
                           n10984, ZN => n10993);
   U12590 : AOI22_X1 port map( A1 => n11249, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_271_port, B1 => 
                           n11251, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_47_port, ZN => 
                           n10991);
   U12591 : AOI22_X1 port map( A1 => n8596, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_303_port, B1 => 
                           n11248, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_143_port, ZN => 
                           n10990);
   U12592 : AOI22_X1 port map( A1 => n8599, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_15_port, B1 => 
                           n8607, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_431_port, ZN => 
                           n10989);
   U12593 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_399_port, B1 => 
                           n8601, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_175_port, ZN => 
                           n10988);
   U12594 : NAND4_X1 port map( A1 => n10991, A2 => n10990, A3 => n10989, A4 => 
                           n10988, ZN => n10992);
   U12595 : OR2_X1 port map( A1 => n10993, A2 => n10992, ZN => 
                           DRAMRF_DATA_OUT(15));
   U12596 : AOI22_X1 port map( A1 => n8585, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_464_port, B1 => 
                           n8587, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_336_port, ZN => 
                           n10997);
   U12597 : AOI22_X1 port map( A1 => n8584, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_208_port, B1 => 
                           n8589, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_240_port, ZN => 
                           n10996);
   U12598 : AOI22_X1 port map( A1 => n11239, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_368_port, B1 => 
                           n8592, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_112_port, ZN => 
                           n10995);
   U12599 : AOI22_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_496_port, B1 => 
                           n11236, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_80_port, ZN => 
                           n10994);
   U12600 : NAND4_X1 port map( A1 => n10997, A2 => n10996, A3 => n10995, A4 => 
                           n10994, ZN => n11003);
   U12601 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_400_port, B1 => 
                           n8597, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_272_port, ZN => 
                           n11001);
   U12602 : AOI22_X1 port map( A1 => n8606, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_48_port, B1 => 
                           n8603, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_144_port, ZN => 
                           n11000);
   U12603 : AOI22_X1 port map( A1 => n11246, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_304_port, B1 => 
                           n8599, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_16_port, ZN => 
                           n10999);
   U12604 : AOI22_X1 port map( A1 => n8607, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_432_port, B1 => 
                           n8602, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_176_port, ZN => 
                           n10998);
   U12605 : NAND4_X1 port map( A1 => n11001, A2 => n11000, A3 => n10999, A4 => 
                           n10998, ZN => n11002);
   U12606 : OR2_X1 port map( A1 => n11003, A2 => n11002, ZN => 
                           DRAMRF_DATA_OUT(16));
   U12607 : AOI22_X1 port map( A1 => n8586, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_465_port, B1 => 
                           n8588, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_337_port, ZN => 
                           n11007);
   U12608 : AOI22_X1 port map( A1 => n8584, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_209_port, B1 => 
                           n11238, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_241_port, ZN => 
                           n11006);
   U12609 : AOI22_X1 port map( A1 => n11235, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_497_port, B1 => 
                           n11239, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_369_port, ZN => 
                           n11005);
   U12610 : AOI22_X1 port map( A1 => n8591, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_81_port, B1 => 
                           n11234, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_113_port, ZN => 
                           n11004);
   U12611 : NAND4_X1 port map( A1 => n11007, A2 => n11006, A3 => n11005, A4 => 
                           n11004, ZN => n11013);
   U12612 : AOI22_X1 port map( A1 => n11253, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_17_port, B1 => 
                           n11248, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_145_port, ZN => 
                           n11011);
   U12613 : AOI22_X1 port map( A1 => n8596, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_305_port, B1 => 
                           n11252, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_177_port, ZN => 
                           n11010);
   U12614 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_401_port, B1 => 
                           n11250, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_433_port, ZN => 
                           n11009);
   U12615 : AOI22_X1 port map( A1 => n11249, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_273_port, B1 => 
                           n8605, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_49_port, ZN => 
                           n11008);
   U12616 : NAND4_X1 port map( A1 => n11011, A2 => n11010, A3 => n11009, A4 => 
                           n11008, ZN => n11012);
   U12617 : OR2_X1 port map( A1 => n11013, A2 => n11012, ZN => 
                           DRAMRF_DATA_OUT(17));
   U12618 : AOI22_X1 port map( A1 => n8586, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_466_port, B1 => 
                           n8591, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_82_port, ZN => 
                           n11017);
   U12619 : AOI22_X1 port map( A1 => n11239, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_370_port, B1 => 
                           n8584, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_210_port, ZN => 
                           n11016);
   U12620 : AOI22_X1 port map( A1 => n8589, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_242_port, B1 => 
                           n8593, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_114_port, ZN => 
                           n11015);
   U12621 : AOI22_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_498_port, B1 => 
                           n8588, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_338_port, ZN => 
                           n11014);
   U12622 : NAND4_X1 port map( A1 => n11017, A2 => n11016, A3 => n11015, A4 => 
                           n11014, ZN => n11023);
   U12623 : AOI22_X1 port map( A1 => n8599, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_18_port, B1 => 
                           n8607, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_434_port, ZN => 
                           n11021);
   U12624 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_402_port, B1 => 
                           n8597, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_274_port, ZN => 
                           n11020);
   U12625 : AOI22_X1 port map( A1 => n8605, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_50_port, B1 => 
                           n8602, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_178_port, ZN => 
                           n11019);
   U12626 : AOI22_X1 port map( A1 => n8595, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_306_port, B1 => 
                           n8604, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_146_port, ZN => 
                           n11018);
   U12627 : NAND4_X1 port map( A1 => n11021, A2 => n11020, A3 => n11019, A4 => 
                           n11018, ZN => n11022);
   U12628 : OR2_X1 port map( A1 => n11023, A2 => n11022, ZN => 
                           DRAMRF_DATA_OUT(18));
   U12629 : AOI22_X1 port map( A1 => n11235, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_499_port, B1 => 
                           n11241, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_211_port, ZN => 
                           n11027);
   U12630 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_371_port, B1 => 
                           n8589, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_243_port, ZN => 
                           n11026);
   U12631 : AOI22_X1 port map( A1 => n8588, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_339_port, B1 => 
                           n11234, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_115_port, ZN => 
                           n11025);
   U12632 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_467_port, B1 => 
                           n11236, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_83_port, ZN => 
                           n11024);
   U12633 : NAND4_X1 port map( A1 => n11027, A2 => n11026, A3 => n11025, A4 => 
                           n11024, ZN => n11033);
   U12634 : AOI22_X1 port map( A1 => n8597, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_275_port, B1 => 
                           n8608, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_435_port, ZN => 
                           n11031);
   U12635 : AOI22_X1 port map( A1 => n8596, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_307_port, B1 => 
                           n11248, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_147_port, ZN => 
                           n11030);
   U12636 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_403_port, B1 => 
                           n8606, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_51_port, ZN => 
                           n11029);
   U12637 : AOI22_X1 port map( A1 => n8600, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_19_port, B1 => 
                           n8601, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_179_port, ZN => 
                           n11028);
   U12638 : NAND4_X1 port map( A1 => n11031, A2 => n11030, A3 => n11029, A4 => 
                           n11028, ZN => n11032);
   U12639 : OR2_X1 port map( A1 => n11033, A2 => n11032, ZN => 
                           DRAMRF_DATA_OUT(19));
   U12640 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_449_port, B1 => 
                           n8591, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_65_port, ZN => 
                           n11037);
   U12641 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_353_port, B1 => 
                           n8592, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_97_port, ZN => 
                           n11036);
   U12642 : AOI22_X1 port map( A1 => n8587, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_321_port, B1 => 
                           n8590, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_225_port, ZN => 
                           n11035);
   U12643 : AOI22_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_481_port, B1 => 
                           n11241, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_193_port, ZN => 
                           n11034);
   U12644 : NAND4_X1 port map( A1 => n11037, A2 => n11036, A3 => n11035, A4 => 
                           n11034, ZN => n11043);
   U12645 : AOI22_X1 port map( A1 => n8600, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_1_port, B1 => 
                           n8606, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_33_port, ZN => 
                           n11041);
   U12646 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_385_port, B1 => 
                           n8608, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_417_port, ZN => 
                           n11040);
   U12647 : AOI22_X1 port map( A1 => n8598, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_257_port, B1 => 
                           n8603, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_129_port, ZN => 
                           n11039);
   U12648 : AOI22_X1 port map( A1 => n11246, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_289_port, B1 => 
                           n8602, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_161_port, ZN => 
                           n11038);
   U12649 : NAND4_X1 port map( A1 => n11041, A2 => n11040, A3 => n11039, A4 => 
                           n11038, ZN => n11042);
   U12650 : OR2_X1 port map( A1 => n11043, A2 => n11042, ZN => 
                           DRAMRF_DATA_OUT(1));
   U12651 : AOI22_X1 port map( A1 => n11239, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_372_port, B1 => 
                           n8590, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_244_port, ZN => 
                           n11047);
   U12652 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_212_port, B1 => 
                           n11237, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_468_port, ZN => 
                           n11046);
   U12653 : AOI22_X1 port map( A1 => n11236, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_84_port, B1 => 
                           n8592, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_116_port, ZN => 
                           n11045);
   U12654 : AOI22_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_500_port, B1 => 
                           n11240, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_340_port, ZN => 
                           n11044);
   U12655 : NAND4_X1 port map( A1 => n11047, A2 => n11046, A3 => n11045, A4 => 
                           n11044, ZN => n11053);
   U12656 : AOI22_X1 port map( A1 => n11246, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_308_port, B1 => 
                           n11251, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_52_port, ZN => 
                           n11051);
   U12657 : AOI22_X1 port map( A1 => n11253, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_20_port, B1 => 
                           n11250, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_436_port, ZN => 
                           n11050);
   U12658 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_404_port, B1 => 
                           n11252, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_180_port, ZN => 
                           n11049);
   U12659 : AOI22_X1 port map( A1 => n8597, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_276_port, B1 => 
                           n8603, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_148_port, ZN => 
                           n11048);
   U12660 : NAND4_X1 port map( A1 => n11051, A2 => n11050, A3 => n11049, A4 => 
                           n11048, ZN => n11052);
   U12661 : OR2_X1 port map( A1 => n11053, A2 => n11052, ZN => 
                           DRAMRF_DATA_OUT(20));
   U12662 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_213_port, B1 => 
                           n11236, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_85_port, ZN => 
                           n11057);
   U12663 : AOI22_X1 port map( A1 => n11239, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_373_port, B1 => 
                           n8593, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_117_port, ZN => 
                           n11056);
   U12664 : AOI22_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_501_port, B1 => 
                           n8585, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_469_port, ZN => 
                           n11055);
   U12665 : AOI22_X1 port map( A1 => n8588, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_341_port, B1 => 
                           n11238, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_245_port, ZN => 
                           n11054);
   U12666 : NAND4_X1 port map( A1 => n11057, A2 => n11056, A3 => n11055, A4 => 
                           n11054, ZN => n11063);
   U12667 : AOI22_X1 port map( A1 => n8608, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_437_port, B1 => 
                           n8604, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_149_port, ZN => 
                           n11061);
   U12668 : AOI22_X1 port map( A1 => n8595, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_309_port, B1 => 
                           n8599, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_21_port, ZN => 
                           n11060);
   U12669 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_405_port, B1 => 
                           n11251, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_53_port, ZN => 
                           n11059);
   U12670 : AOI22_X1 port map( A1 => n11249, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_277_port, B1 => 
                           n11252, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_181_port, ZN => 
                           n11058);
   U12671 : NAND4_X1 port map( A1 => n11061, A2 => n11060, A3 => n11059, A4 => 
                           n11058, ZN => n11062);
   U12672 : OR2_X1 port map( A1 => n11063, A2 => n11062, ZN => 
                           DRAMRF_DATA_OUT(21));
   U12673 : AOI22_X1 port map( A1 => n8584, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_214_port, B1 => 
                           n8593, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_118_port, ZN => 
                           n11067);
   U12674 : AOI22_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_502_port, B1 => 
                           n11240, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_342_port, ZN => 
                           n11066);
   U12675 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_374_port, B1 => 
                           n11238, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_246_port, ZN => 
                           n11065);
   U12676 : AOI22_X1 port map( A1 => n8585, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_470_port, B1 => 
                           n8591, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_86_port, ZN => 
                           n11064);
   U12677 : NAND4_X1 port map( A1 => n11067, A2 => n11066, A3 => n11065, A4 => 
                           n11064, ZN => n11073);
   U12678 : AOI22_X1 port map( A1 => n8597, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_278_port, B1 => 
                           n11250, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_438_port, ZN => 
                           n11071);
   U12679 : AOI22_X1 port map( A1 => n8595, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_310_port, B1 => 
                           n8604, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_150_port, ZN => 
                           n11070);
   U12680 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_406_port, B1 => 
                           n8600, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_22_port, ZN => 
                           n11069);
   U12681 : AOI22_X1 port map( A1 => n8606, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_54_port, B1 => 
                           n8601, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_182_port, ZN => 
                           n11068);
   U12682 : NAND4_X1 port map( A1 => n11071, A2 => n11070, A3 => n11069, A4 => 
                           n11068, ZN => n11072);
   U12683 : OR2_X1 port map( A1 => n11073, A2 => n11072, ZN => 
                           DRAMRF_DATA_OUT(22));
   U12684 : AOI22_X1 port map( A1 => n8584, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_215_port, B1 => 
                           n11236, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_87_port, ZN => 
                           n11077);
   U12685 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_375_port, B1 => 
                           n8585, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_471_port, ZN => 
                           n11076);
   U12686 : AOI22_X1 port map( A1 => n8590, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_247_port, B1 => 
                           n11234, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_119_port, ZN => 
                           n11075);
   U12687 : AOI22_X1 port map( A1 => n11235, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_503_port, B1 => 
                           n8587, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_343_port, ZN => 
                           n11074);
   U12688 : NAND4_X1 port map( A1 => n11077, A2 => n11076, A3 => n11075, A4 => 
                           n11074, ZN => n11083);
   U12689 : AOI22_X1 port map( A1 => n8596, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_311_port, B1 => 
                           n11248, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_151_port, ZN => 
                           n11081);
   U12690 : AOI22_X1 port map( A1 => n8598, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_279_port, B1 => 
                           n8607, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_439_port, ZN => 
                           n11080);
   U12691 : AOI22_X1 port map( A1 => n11253, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_23_port, B1 => 
                           n8605, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_55_port, ZN => 
                           n11079);
   U12692 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_407_port, B1 => 
                           n8601, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_183_port, ZN => 
                           n11078);
   U12693 : NAND4_X1 port map( A1 => n11081, A2 => n11080, A3 => n11079, A4 => 
                           n11078, ZN => n11082);
   U12694 : OR2_X1 port map( A1 => n11083, A2 => n11082, ZN => 
                           DRAMRF_DATA_OUT(23));
   U12695 : AOI22_X1 port map( A1 => n11239, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_376_port, B1 => 
                           n8591, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_88_port, ZN => 
                           n11087);
   U12696 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_216_port, B1 => 
                           n8586, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_472_port, ZN => 
                           n11086);
   U12697 : AOI22_X1 port map( A1 => n11240, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_344_port, B1 => 
                           n8592, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_120_port, ZN => 
                           n11085);
   U12698 : AOI22_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_504_port, B1 => 
                           n8589, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_248_port, ZN => 
                           n11084);
   U12699 : NAND4_X1 port map( A1 => n11087, A2 => n11086, A3 => n11085, A4 => 
                           n11084, ZN => n11093);
   U12700 : AOI22_X1 port map( A1 => n11246, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_312_port, B1 => 
                           n8598, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_280_port, ZN => 
                           n11091);
   U12701 : AOI22_X1 port map( A1 => n8602, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_184_port, B1 => 
                           n8603, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_152_port, ZN => 
                           n11090);
   U12702 : AOI22_X1 port map( A1 => n8599, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_24_port, B1 => 
                           n8606, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_56_port, ZN => 
                           n11089);
   U12703 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_408_port, B1 => 
                           n8608, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_440_port, ZN => 
                           n11088);
   U12704 : NAND4_X1 port map( A1 => n11091, A2 => n11090, A3 => n11089, A4 => 
                           n11088, ZN => n11092);
   U12705 : OR2_X1 port map( A1 => n11093, A2 => n11092, ZN => 
                           DRAMRF_DATA_OUT(24));
   U12706 : AOI22_X1 port map( A1 => n8591, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_89_port, B1 => 
                           n11234, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_121_port, ZN => 
                           n11097);
   U12707 : AOI22_X1 port map( A1 => n11235, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_505_port, B1 => 
                           n8583, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_377_port, ZN => 
                           n11096);
   U12708 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_217_port, B1 => 
                           n8588, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_345_port, ZN => 
                           n11095);
   U12709 : AOI22_X1 port map( A1 => n8586, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_473_port, B1 => 
                           n8590, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_249_port, ZN => 
                           n11094);
   U12710 : NAND4_X1 port map( A1 => n11097, A2 => n11096, A3 => n11095, A4 => 
                           n11094, ZN => n11103);
   U12711 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_409_port, B1 => 
                           n11253, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_25_port, ZN => 
                           n11101);
   U12712 : AOI22_X1 port map( A1 => n8596, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_313_port, B1 => 
                           n8602, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_185_port, ZN => 
                           n11100);
   U12713 : AOI22_X1 port map( A1 => n8598, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_281_port, B1 => 
                           n8605, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_57_port, ZN => 
                           n11099);
   U12714 : AOI22_X1 port map( A1 => n11250, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_441_port, B1 => 
                           n11248, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_153_port, ZN => 
                           n11098);
   U12715 : NAND4_X1 port map( A1 => n11101, A2 => n11100, A3 => n11099, A4 => 
                           n11098, ZN => n11102);
   U12716 : OR2_X1 port map( A1 => n11103, A2 => n11102, ZN => 
                           DRAMRF_DATA_OUT(25));
   U12717 : AOI22_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_506_port, B1 => 
                           n8587, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_346_port, ZN => 
                           n11107);
   U12718 : AOI22_X1 port map( A1 => n11239, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_378_port, B1 => 
                           n8593, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_122_port, ZN => 
                           n11106);
   U12719 : AOI22_X1 port map( A1 => n8584, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_218_port, B1 => 
                           n8589, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_250_port, ZN => 
                           n11105);
   U12720 : AOI22_X1 port map( A1 => n8585, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_474_port, B1 => 
                           n11236, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_90_port, ZN => 
                           n11104);
   U12721 : NAND4_X1 port map( A1 => n11107, A2 => n11106, A3 => n11105, A4 => 
                           n11104, ZN => n11113);
   U12722 : AOI22_X1 port map( A1 => n8595, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_314_port, B1 => 
                           n11251, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_58_port, ZN => 
                           n11111);
   U12723 : AOI22_X1 port map( A1 => n11250, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_442_port, B1 => 
                           n11252, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_186_port, ZN => 
                           n11110);
   U12724 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_410_port, B1 => 
                           n11249, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_282_port, ZN => 
                           n11109);
   U12725 : AOI22_X1 port map( A1 => n8600, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_26_port, B1 => 
                           n8604, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_154_port, ZN => 
                           n11108);
   U12726 : NAND4_X1 port map( A1 => n11111, A2 => n11110, A3 => n11109, A4 => 
                           n11108, ZN => n11112);
   U12727 : OR2_X1 port map( A1 => n11113, A2 => n11112, ZN => 
                           DRAMRF_DATA_OUT(26));
   U12728 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_379_port, B1 => 
                           n11240, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_347_port, ZN => 
                           n11117);
   U12729 : AOI22_X1 port map( A1 => n11235, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_507_port, B1 => 
                           n11234, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_123_port, ZN => 
                           n11116);
   U12730 : AOI22_X1 port map( A1 => n8584, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_219_port, B1 => 
                           n11237, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_475_port, ZN => 
                           n11115);
   U12731 : AOI22_X1 port map( A1 => n11238, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_251_port, B1 => 
                           n8591, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_91_port, ZN => 
                           n11114);
   U12732 : NAND4_X1 port map( A1 => n11117, A2 => n11116, A3 => n11115, A4 => 
                           n11114, ZN => n11123);
   U12733 : AOI22_X1 port map( A1 => n11251, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_59_port, B1 => 
                           n11248, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_155_port, ZN => 
                           n11121);
   U12734 : AOI22_X1 port map( A1 => n8596, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_315_port, B1 => 
                           n8598, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_283_port, ZN => 
                           n11120);
   U12735 : AOI22_X1 port map( A1 => n8607, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_443_port, B1 => 
                           n8602, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_187_port, ZN => 
                           n11119);
   U12736 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_411_port, B1 => 
                           n8600, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_27_port, ZN => 
                           n11118);
   U12737 : NAND4_X1 port map( A1 => n11121, A2 => n11120, A3 => n11119, A4 => 
                           n11118, ZN => n11122);
   U12738 : OR2_X1 port map( A1 => n11123, A2 => n11122, ZN => 
                           DRAMRF_DATA_OUT(27));
   U12739 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_220_port, B1 => 
                           n8587, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_348_port, ZN => 
                           n11127);
   U12740 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_380_port, B1 => 
                           n8592, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_124_port, ZN => 
                           n11126);
   U12741 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_476_port, B1 => 
                           n11236, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_92_port, ZN => 
                           n11125);
   U12742 : AOI22_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_508_port, B1 => 
                           n11238, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_252_port, ZN => 
                           n11124);
   U12743 : NAND4_X1 port map( A1 => n11127, A2 => n11126, A3 => n11125, A4 => 
                           n11124, ZN => n11133);
   U12744 : AOI22_X1 port map( A1 => n11251, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_60_port, B1 => 
                           n8601, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_188_port, ZN => 
                           n11131);
   U12745 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_412_port, B1 => 
                           n8595, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_316_port, ZN => 
                           n11130);
   U12746 : AOI22_X1 port map( A1 => n8607, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_444_port, B1 => 
                           n8603, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_156_port, ZN => 
                           n11129);
   U12747 : AOI22_X1 port map( A1 => n11249, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_284_port, B1 => 
                           n8599, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_28_port, ZN => 
                           n11128);
   U12748 : NAND4_X1 port map( A1 => n11131, A2 => n11130, A3 => n11129, A4 => 
                           n11128, ZN => n11132);
   U12749 : OR2_X1 port map( A1 => n11133, A2 => n11132, ZN => 
                           DRAMRF_DATA_OUT(28));
   U12750 : AOI22_X1 port map( A1 => n8585, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_477_port, B1 => 
                           n8591, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_93_port, ZN => 
                           n11137);
   U12751 : AOI22_X1 port map( A1 => n11239, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_381_port, B1 => 
                           n8592, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_125_port, ZN => 
                           n11136);
   U12752 : AOI22_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_509_port, B1 => 
                           n8589, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_253_port, ZN => 
                           n11135);
   U12753 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_221_port, B1 => 
                           n8588, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_349_port, ZN => 
                           n11134);
   U12754 : NAND4_X1 port map( A1 => n11137, A2 => n11136, A3 => n11135, A4 => 
                           n11134, ZN => n11143);
   U12755 : AOI22_X1 port map( A1 => n11246, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_317_port, B1 => 
                           n8597, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_285_port, ZN => 
                           n11141);
   U12756 : AOI22_X1 port map( A1 => n8599, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_29_port, B1 => 
                           n8603, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_157_port, ZN => 
                           n11140);
   U12757 : AOI22_X1 port map( A1 => n8605, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_61_port, B1 => 
                           n8607, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_445_port, ZN => 
                           n11139);
   U12758 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_413_port, B1 => 
                           n8602, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_189_port, ZN => 
                           n11138);
   U12759 : NAND4_X1 port map( A1 => n11141, A2 => n11140, A3 => n11139, A4 => 
                           n11138, ZN => n11142);
   U12760 : OR2_X1 port map( A1 => n11143, A2 => n11142, ZN => 
                           DRAMRF_DATA_OUT(29));
   U12761 : AOI22_X1 port map( A1 => n11240, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_322_port, B1 => 
                           n8593, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_98_port, ZN => 
                           n11147);
   U12762 : AOI22_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_482_port, B1 => 
                           n11236, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_66_port, ZN => 
                           n11146);
   U12763 : AOI22_X1 port map( A1 => n11239, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_354_port, B1 => 
                           n8590, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_226_port, ZN => 
                           n11145);
   U12764 : AOI22_X1 port map( A1 => n8584, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_194_port, B1 => 
                           n8586, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_450_port, ZN => 
                           n11144);
   U12765 : NAND4_X1 port map( A1 => n11147, A2 => n11146, A3 => n11145, A4 => 
                           n11144, ZN => n11153);
   U12766 : AOI22_X1 port map( A1 => n11253, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_2_port, B1 => 
                           n8605, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_34_port, ZN => 
                           n11151);
   U12767 : AOI22_X1 port map( A1 => n8608, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_418_port, B1 => 
                           n8604, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_130_port, ZN => 
                           n11150);
   U12768 : AOI22_X1 port map( A1 => n11246, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_290_port, B1 => 
                           n8598, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_258_port, ZN => 
                           n11149);
   U12769 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_386_port, B1 => 
                           n11252, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_162_port, ZN => 
                           n11148);
   U12770 : NAND4_X1 port map( A1 => n11151, A2 => n11150, A3 => n11149, A4 => 
                           n11148, ZN => n11152);
   U12771 : OR2_X1 port map( A1 => n11153, A2 => n11152, ZN => 
                           DRAMRF_DATA_OUT(2));
   U12772 : AOI22_X1 port map( A1 => n8587, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_350_port, B1 => 
                           n8591, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_94_port, ZN => 
                           n11157);
   U12773 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_382_port, B1 => 
                           n8585, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_478_port, ZN => 
                           n11156);
   U12774 : AOI22_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_510_port, B1 => 
                           n8593, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_126_port, ZN => 
                           n11155);
   U12775 : AOI22_X1 port map( A1 => n8584, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_222_port, B1 => 
                           n8590, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_254_port, ZN => 
                           n11154);
   U12776 : NAND4_X1 port map( A1 => n11157, A2 => n11156, A3 => n11155, A4 => 
                           n11154, ZN => n11163);
   U12777 : AOI22_X1 port map( A1 => n8599, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_30_port, B1 => 
                           n11252, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_190_port, ZN => 
                           n11161);
   U12778 : AOI22_X1 port map( A1 => n11249, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_286_port, B1 => 
                           n8604, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_158_port, ZN => 
                           n11160);
   U12779 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_414_port, B1 => 
                           n11250, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_446_port, ZN => 
                           n11159);
   U12780 : AOI22_X1 port map( A1 => n8595, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_318_port, B1 => 
                           n8606, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_62_port, ZN => 
                           n11158);
   U12781 : NAND4_X1 port map( A1 => n11161, A2 => n11160, A3 => n11159, A4 => 
                           n11158, ZN => n11162);
   U12782 : OR2_X1 port map( A1 => n11163, A2 => n11162, ZN => 
                           DRAMRF_DATA_OUT(30));
   U12783 : AOI22_X1 port map( A1 => n8586, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_479_port, B1 => 
                           n11236, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_95_port, ZN => 
                           n11167);
   U12784 : AOI22_X1 port map( A1 => n11235, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_511_port, B1 => 
                           n11234, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_127_port, ZN => 
                           n11166);
   U12785 : AOI22_X1 port map( A1 => n8587, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_351_port, B1 => 
                           n11238, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_255_port, ZN => 
                           n11165);
   U12786 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_383_port, B1 => 
                           n8584, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_223_port, ZN => 
                           n11164);
   U12787 : NAND4_X1 port map( A1 => n11167, A2 => n11166, A3 => n11165, A4 => 
                           n11164, ZN => n11173);
   U12788 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_415_port, B1 => 
                           n11248, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_159_port, ZN => 
                           n11171);
   U12789 : AOI22_X1 port map( A1 => n8595, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_319_port, B1 => 
                           n8606, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_63_port, ZN => 
                           n11170);
   U12790 : AOI22_X1 port map( A1 => n8600, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_31_port, B1 => 
                           n8601, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_191_port, ZN => 
                           n11169);
   U12791 : AOI22_X1 port map( A1 => n8597, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_287_port, B1 => 
                           n8607, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_447_port, ZN => 
                           n11168);
   U12792 : NAND4_X1 port map( A1 => n11171, A2 => n11170, A3 => n11169, A4 => 
                           n11168, ZN => n11172);
   U12793 : OR2_X1 port map( A1 => n11173, A2 => n11172, ZN => 
                           DRAMRF_DATA_OUT(31));
   U12794 : AOI22_X1 port map( A1 => n11239, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_355_port, B1 => 
                           n11238, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_227_port, ZN => 
                           n11177);
   U12795 : AOI22_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_483_port, B1 => 
                           n8592, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_99_port, ZN => 
                           n11176);
   U12796 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_195_port, B1 => 
                           n8591, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_67_port, ZN => 
                           n11175);
   U12797 : AOI22_X1 port map( A1 => n8586, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_451_port, B1 => 
                           n8588, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_323_port, ZN => 
                           n11174);
   U12798 : NAND4_X1 port map( A1 => n11177, A2 => n11176, A3 => n11175, A4 => 
                           n11174, ZN => n11183);
   U12799 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_387_port, B1 => 
                           n8596, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_291_port, ZN => 
                           n11181);
   U12800 : AOI22_X1 port map( A1 => n8598, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_259_port, B1 => 
                           n8603, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_131_port, ZN => 
                           n11180);
   U12801 : AOI22_X1 port map( A1 => n8605, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_35_port, B1 => 
                           n8601, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_163_port, ZN => 
                           n11179);
   U12802 : AOI22_X1 port map( A1 => n8600, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_3_port, B1 => 
                           n8608, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_419_port, ZN => 
                           n11178);
   U12803 : NAND4_X1 port map( A1 => n11181, A2 => n11180, A3 => n11179, A4 => 
                           n11178, ZN => n11182);
   U12804 : OR2_X1 port map( A1 => n11183, A2 => n11182, ZN => 
                           DRAMRF_DATA_OUT(3));
   U12805 : AOI22_X1 port map( A1 => n8588, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_324_port, B1 => 
                           n11234, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_100_port, ZN => 
                           n11187);
   U12806 : AOI22_X1 port map( A1 => n11235, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_484_port, B1 => 
                           n8583, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_356_port, ZN => 
                           n11186);
   U12807 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_452_port, B1 => 
                           n8589, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_228_port, ZN => 
                           n11185);
   U12808 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_196_port, B1 => 
                           n11236, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_68_port, ZN => 
                           n11184);
   U12809 : NAND4_X1 port map( A1 => n11187, A2 => n11186, A3 => n11185, A4 => 
                           n11184, ZN => n11193);
   U12810 : AOI22_X1 port map( A1 => n8597, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_260_port, B1 => 
                           n11248, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_132_port, ZN => 
                           n11191);
   U12811 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_388_port, B1 => 
                           n8602, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_164_port, ZN => 
                           n11190);
   U12812 : AOI22_X1 port map( A1 => n11253, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_4_port, B1 => 
                           n8608, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_420_port, ZN => 
                           n11189);
   U12813 : AOI22_X1 port map( A1 => n8596, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_292_port, B1 => 
                           n11251, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_36_port, ZN => 
                           n11188);
   U12814 : NAND4_X1 port map( A1 => n11191, A2 => n11190, A3 => n11189, A4 => 
                           n11188, ZN => n11192);
   U12815 : OR2_X1 port map( A1 => n11193, A2 => n11192, ZN => 
                           DRAMRF_DATA_OUT(4));
   U12816 : AOI22_X1 port map( A1 => n11239, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_357_port, B1 => 
                           n8591, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_69_port, ZN => 
                           n11197);
   U12817 : AOI22_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_485_port, B1 => 
                           n8584, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_197_port, ZN => 
                           n11196);
   U12818 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_453_port, B1 => 
                           n11240, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_325_port, ZN => 
                           n11195);
   U12819 : AOI22_X1 port map( A1 => n8590, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_229_port, B1 => 
                           n8593, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_101_port, ZN => 
                           n11194);
   U12820 : NAND4_X1 port map( A1 => n11197, A2 => n11196, A3 => n11195, A4 => 
                           n11194, ZN => n11203);
   U12821 : AOI22_X1 port map( A1 => n11246, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_293_port, B1 => 
                           n11251, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_37_port, ZN => 
                           n11201);
   U12822 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_389_port, B1 => 
                           n11252, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_165_port, ZN => 
                           n11200);
   U12823 : AOI22_X1 port map( A1 => n11249, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_261_port, B1 => 
                           n8600, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_5_port, ZN => 
                           n11199);
   U12824 : AOI22_X1 port map( A1 => n11250, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_421_port, B1 => 
                           n8604, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_133_port, ZN => 
                           n11198);
   U12825 : NAND4_X1 port map( A1 => n11201, A2 => n11200, A3 => n11199, A4 => 
                           n11198, ZN => n11202);
   U12826 : OR2_X1 port map( A1 => n11203, A2 => n11202, ZN => 
                           DRAMRF_DATA_OUT(5));
   U12827 : AOI22_X1 port map( A1 => n11235, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_486_port, B1 => 
                           n8590, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_230_port, ZN => 
                           n11207);
   U12828 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_358_port, B1 => 
                           n8586, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_454_port, ZN => 
                           n11206);
   U12829 : AOI22_X1 port map( A1 => n11236, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_70_port, B1 => 
                           n11234, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_102_port, ZN => 
                           n11205);
   U12830 : AOI22_X1 port map( A1 => n8584, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_198_port, B1 => 
                           n11240, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_326_port, ZN => 
                           n11204);
   U12831 : NAND4_X1 port map( A1 => n11207, A2 => n11206, A3 => n11205, A4 => 
                           n11204, ZN => n11213);
   U12832 : AOI22_X1 port map( A1 => n8606, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_38_port, B1 => 
                           n8602, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_166_port, ZN => 
                           n11211);
   U12833 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_390_port, B1 => 
                           n11253, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_6_port, ZN => 
                           n11210);
   U12834 : AOI22_X1 port map( A1 => n8597, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_262_port, B1 => 
                           n11250, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_422_port, ZN => 
                           n11209);
   U12835 : AOI22_X1 port map( A1 => n8596, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_294_port, B1 => 
                           n11248, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_134_port, ZN => 
                           n11208);
   U12836 : NAND4_X1 port map( A1 => n11211, A2 => n11210, A3 => n11209, A4 => 
                           n11208, ZN => n11212);
   U12837 : OR2_X1 port map( A1 => n11213, A2 => n11212, ZN => 
                           DRAMRF_DATA_OUT(6));
   U12838 : AOI22_X1 port map( A1 => n11240, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_327_port, B1 => 
                           n11236, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_71_port, ZN => 
                           n11217);
   U12839 : AOI22_X1 port map( A1 => n8589, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_231_port, B1 => 
                           n8592, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_103_port, ZN => 
                           n11216);
   U12840 : AOI22_X1 port map( A1 => n8584, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_199_port, B1 => 
                           n11237, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_455_port, ZN => 
                           n11215);
   U12841 : AOI22_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_487_port, B1 => 
                           n11239, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_359_port, ZN => 
                           n11214);
   U12842 : NAND4_X1 port map( A1 => n11217, A2 => n11216, A3 => n11215, A4 => 
                           n11214, ZN => n11223);
   U12843 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_391_port, B1 => 
                           n8605, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_39_port, ZN => 
                           n11221);
   U12844 : AOI22_X1 port map( A1 => n8598, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_263_port, B1 => 
                           n11250, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_423_port, ZN => 
                           n11220);
   U12845 : AOI22_X1 port map( A1 => n11253, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_7_port, B1 => 
                           n8603, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_135_port, ZN => 
                           n11219);
   U12846 : AOI22_X1 port map( A1 => n8595, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_295_port, B1 => 
                           n8601, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_167_port, ZN => 
                           n11218);
   U12847 : NAND4_X1 port map( A1 => n11221, A2 => n11220, A3 => n11219, A4 => 
                           n11218, ZN => n11222);
   U12848 : OR2_X1 port map( A1 => n11223, A2 => n11222, ZN => 
                           DRAMRF_DATA_OUT(7));
   U12849 : AOI22_X1 port map( A1 => n8583, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_360_port, B1 => 
                           n11241, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_200_port, ZN => 
                           n11227);
   U12850 : AOI22_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_488_port, B1 => 
                           n8587, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_328_port, ZN => 
                           n11226);
   U12851 : AOI22_X1 port map( A1 => n8590, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_232_port, B1 => 
                           n8591, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_72_port, ZN => 
                           n11225);
   U12852 : AOI22_X1 port map( A1 => n8585, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_456_port, B1 => 
                           n8592, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_104_port, ZN => 
                           n11224);
   U12853 : NAND4_X1 port map( A1 => n11227, A2 => n11226, A3 => n11225, A4 => 
                           n11224, ZN => n11233);
   U12854 : AOI22_X1 port map( A1 => n8599, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_8_port, B1 => 
                           n8603, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_136_port, ZN => 
                           n11231);
   U12855 : AOI22_X1 port map( A1 => n8596, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_296_port, B1 => 
                           n8606, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_40_port, ZN => 
                           n11230);
   U12856 : AOI22_X1 port map( A1 => n8594, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_392_port, B1 => 
                           n8607, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_424_port, ZN => 
                           n11229);
   U12857 : AOI22_X1 port map( A1 => n8598, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_264_port, B1 => 
                           n8602, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_168_port, ZN => 
                           n11228);
   U12858 : NAND4_X1 port map( A1 => n11231, A2 => n11230, A3 => n11229, A4 => 
                           n11228, ZN => n11232);
   U12859 : OR2_X1 port map( A1 => n11233, A2 => n11232, ZN => 
                           DRAMRF_DATA_OUT(8));
   U12860 : AOI22_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_489_port, B1 => 
                           n8593, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_105_port, ZN => 
                           n11245);
   U12861 : AOI22_X1 port map( A1 => n8586, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_457_port, B1 => 
                           n11236, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_73_port, ZN => 
                           n11244);
   U12862 : AOI22_X1 port map( A1 => n11239, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_361_port, B1 => 
                           n8589, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_233_port, ZN => 
                           n11243);
   U12863 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_201_port, B1 => 
                           n8588, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_329_port, ZN => 
                           n11242);
   U12864 : NAND4_X1 port map( A1 => n11245, A2 => n11244, A3 => n11243, A4 => 
                           n11242, ZN => n11259);
   U12865 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_393_port, B1 => 
                           n8595, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_297_port, ZN => 
                           n11257);
   U12866 : AOI22_X1 port map( A1 => n11249, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_265_port, B1 => 
                           n8604, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_137_port, ZN => 
                           n11256);
   U12867 : AOI22_X1 port map( A1 => n11251, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_41_port, B1 => 
                           n8608, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_425_port, ZN => 
                           n11255);
   U12868 : AOI22_X1 port map( A1 => n8600, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_9_port, B1 => 
                           n11252, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_169_port, ZN => 
                           n11254);
   U12869 : NAND4_X1 port map( A1 => n11257, A2 => n11256, A3 => n11255, A4 => 
                           n11254, ZN => n11258);
   U12870 : OR2_X1 port map( A1 => n11259, A2 => n11258, ZN => 
                           DRAMRF_DATA_OUT(9));
   U12871 : NOR2_X1 port map( A1 => n495, A2 => n393, ZN => DRAM_ADDRESS_0_port
                           );
   U12872 : AOI21_X1 port map( B1 => n392, B2 => n393, A => n496, ZN => 
                           DRAM_ADDRESS_1_port);
   U12873 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(8), B1 =>
                           DataPath_i_REG_ME_DATA_DATAMEM_8_port, B2 => n11305,
                           ZN => n11327);
   U12874 : OAI21_X1 port map( B1 => DATA_SIZE_0_port, B2 => DATA_SIZE_1_port, 
                           A => i_DATAMEM_RM, ZN => n11300);
   U12875 : NOR4_X1 port map( A1 => n8388, A2 => n11270, A3 => n11347, A4 => 
                           n496, ZN => n11285);
   U12876 : INV_X1 port map( A => n11285, ZN => n11310);
   U12877 : NAND2_X1 port map( A1 => n495, A2 => n11331, ZN => n11260);
   U12878 : MUX2_X1 port map( A => DRAM_DATA_IN(24), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_24_port, S => n11305,
                           Z => n11365);
   U12879 : AOI22_X1 port map( A1 => n11304, A2 => n11365, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_0_port, B2 => n11305,
                           ZN => n11264);
   U12880 : NAND2_X1 port map( A1 => n11373, A2 => n8376, ZN => n11261);
   U12881 : NAND3_X1 port map( A1 => i_DATAMEM_RM, A2 => n496, A3 => n11373, ZN
                           => n11262);
   U12882 : INV_X1 port map( A => n11370, ZN => n11295);
   U12883 : OAI21_X1 port map( B1 => n495, B2 => n11262, A => n11295, ZN => 
                           n11306);
   U12884 : MUX2_X1 port map( A => DRAM_DATA_IN(16), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_16_port, S => n11305,
                           Z => n11302);
   U12885 : AOI22_X1 port map( A1 => DRAM_DATA_IN(0), A2 => n11307, B1 => 
                           n11306, B2 => n11302, ZN => n11263);
   U12886 : OAI211_X1 port map( C1 => n11327, C2 => n11310, A => n11264, B => 
                           n11263, ZN => DRAM_DATA_OUT_0_port);
   U12887 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(15), B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_15_port, B2 => 
                           n11305, ZN => n11296);
   U12888 : AOI22_X1 port map( A1 => DRAM_DATA_IN(7), A2 => n11307, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_7_port, B2 => n11305,
                           ZN => n11266);
   U12889 : MUX2_X1 port map( A => DRAM_DATA_IN(31), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_31_port, S => n11305,
                           Z => n11294);
   U12890 : MUX2_X1 port map( A => DRAM_DATA_IN(23), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_23_port, S => n11305,
                           Z => n11324);
   U12891 : AOI22_X1 port map( A1 => n11304, A2 => n11294, B1 => n11324, B2 => 
                           n11306, ZN => n11265);
   U12892 : OAI211_X1 port map( C1 => n11296, C2 => n11310, A => n11266, B => 
                           n11265, ZN => DRAM_DATA_OUT_7_port);
   U12893 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(10), B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_10_port, B2 => 
                           n11305, ZN => n11269);
   U12894 : AOI22_X1 port map( A1 => DRAM_DATA_IN(2), A2 => n11307, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_2_port, B2 => n11305,
                           ZN => n11268);
   U12895 : MUX2_X1 port map( A => DRAM_DATA_IN(26), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_26_port, S => n11305,
                           Z => n11333);
   U12896 : MUX2_X1 port map( A => DRAM_DATA_IN(18), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_18_port, S => n11305,
                           Z => n11313);
   U12897 : AOI22_X1 port map( A1 => n11304, A2 => n11333, B1 => n11306, B2 => 
                           n11313, ZN => n11267);
   U12898 : OAI211_X1 port map( C1 => n11269, C2 => n11310, A => n11268, B => 
                           n11267, ZN => DRAM_DATA_OUT_2_port);
   U12899 : NOR2_X1 port map( A1 => n11331, A2 => n11269, ZN => n11334);
   U12900 : AOI21_X1 port map( B1 => n11370, B2 => n11333, A => n11334, ZN => 
                           n11271);
   U12901 : NAND3_X1 port map( A1 => n11373, A2 => n8382, A3 => 
                           DRAM_DATA_OUT_7_port, ZN => n11325);
   U12902 : AOI21_X1 port map( B1 => n11355, B2 => DRAM_DATA_OUT_2_port, A => 
                           n11329, ZN => n11336);
   U12903 : OAI21_X1 port map( B1 => n11373, B2 => n11271, A => n11336, ZN => 
                           DRAM_DATA_OUT_10_port);
   U12904 : INV_X1 port map( A => n11306, ZN => n11288);
   U12905 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(19), B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_19_port, B2 => 
                           n11305, ZN => n11316);
   U12906 : MUX2_X1 port map( A => DRAM_DATA_IN(27), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_27_port, S => n11305,
                           Z => n11337);
   U12907 : AOI22_X1 port map( A1 => n11304, A2 => n11337, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_3_port, B2 => n11305,
                           ZN => n11273);
   U12908 : MUX2_X1 port map( A => DRAM_DATA_IN(11), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_11_port, S => n11305,
                           Z => n11274);
   U12909 : AOI22_X1 port map( A1 => n11285, A2 => n11274, B1 => n11307, B2 => 
                           DRAM_DATA_IN(3), ZN => n11272);
   U12910 : OAI211_X1 port map( C1 => n11288, C2 => n11316, A => n11273, B => 
                           n11272, ZN => DRAM_DATA_OUT_3_port);
   U12911 : NAND2_X1 port map( A1 => n11347, A2 => n11274, ZN => n11339);
   U12912 : INV_X1 port map( A => n11339, ZN => n11275);
   U12913 : AOI21_X1 port map( B1 => n11370, B2 => n11337, A => n11275, ZN => 
                           n11277);
   U12914 : NAND2_X1 port map( A1 => n11355, A2 => DRAM_DATA_OUT_3_port, ZN => 
                           n11276);
   U12915 : INV_X1 port map( A => n11329, ZN => n11291);
   U12916 : OAI211_X1 port map( C1 => n11373, C2 => n11277, A => n11276, B => 
                           n11291, ZN => DRAM_DATA_OUT_11_port);
   U12917 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(12), B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_12_port, B2 => 
                           n11305, ZN => n11280);
   U12918 : MUX2_X1 port map( A => DRAM_DATA_IN(28), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_28_port, S => n11305,
                           Z => n11340);
   U12919 : AOI22_X1 port map( A1 => n11304, A2 => n11340, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_4_port, B2 => n11305,
                           ZN => n11279);
   U12920 : MUX2_X1 port map( A => DRAM_DATA_IN(20), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_20_port, S => n11305,
                           Z => n11317);
   U12921 : AOI22_X1 port map( A1 => DRAM_DATA_IN(4), A2 => n11307, B1 => 
                           n11306, B2 => n11317, ZN => n11278);
   U12922 : OAI211_X1 port map( C1 => n11280, C2 => n11310, A => n11279, B => 
                           n11278, ZN => DRAM_DATA_OUT_4_port);
   U12923 : NOR2_X1 port map( A1 => n11331, A2 => n11280, ZN => n11341);
   U12924 : AOI21_X1 port map( B1 => n11370, B2 => n11340, A => n11341, ZN => 
                           n11281);
   U12925 : AOI21_X1 port map( B1 => n11355, B2 => DRAM_DATA_OUT_4_port, A => 
                           n11329, ZN => n11345);
   U12926 : OAI21_X1 port map( B1 => n11373, B2 => n11281, A => n11345, ZN => 
                           DRAM_DATA_OUT_12_port);
   U12927 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(21), B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_21_port, B2 => 
                           n11305, ZN => n11320);
   U12928 : MUX2_X1 port map( A => DRAM_DATA_IN(13), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_13_port, S => n11305,
                           Z => n11346);
   U12929 : AOI22_X1 port map( A1 => n11285, A2 => n11346, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_5_port, B2 => n11305,
                           ZN => n11283);
   U12930 : MUX2_X1 port map( A => DRAM_DATA_IN(29), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_29_port, S => n11305,
                           Z => n11349);
   U12931 : AOI22_X1 port map( A1 => n11304, A2 => n11349, B1 => n11307, B2 => 
                           DRAM_DATA_IN(5), ZN => n11282);
   U12932 : OAI211_X1 port map( C1 => n11288, C2 => n11320, A => n11283, B => 
                           n11282, ZN => DRAM_DATA_OUT_5_port);
   U12933 : AOI22_X1 port map( A1 => n11370, A2 => n11349, B1 => n11347, B2 => 
                           n11346, ZN => n11284);
   U12934 : AOI21_X1 port map( B1 => n11355, B2 => DRAM_DATA_OUT_5_port, A => 
                           n11329, ZN => n11351);
   U12935 : OAI21_X1 port map( B1 => n11373, B2 => n11284, A => n11351, ZN => 
                           DRAM_DATA_OUT_13_port);
   U12936 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(22), B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_22_port, B2 => 
                           n11305, ZN => n11322);
   U12937 : MUX2_X1 port map( A => DRAM_DATA_IN(14), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_14_port, S => n11305,
                           Z => n11289);
   U12938 : AOI22_X1 port map( A1 => n11285, A2 => n11289, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_6_port, B2 => n11305,
                           ZN => n11287);
   U12939 : MUX2_X1 port map( A => DRAM_DATA_IN(30), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_30_port, S => n11305,
                           Z => n11353);
   U12940 : AOI22_X1 port map( A1 => n11304, A2 => n11353, B1 => n11307, B2 => 
                           DRAM_DATA_IN(6), ZN => n11286);
   U12941 : OAI211_X1 port map( C1 => n11288, C2 => n11322, A => n11287, B => 
                           n11286, ZN => DRAM_DATA_OUT_6_port);
   U12942 : NAND2_X1 port map( A1 => n11347, A2 => n11289, ZN => n11359);
   U12943 : INV_X1 port map( A => n11359, ZN => n11290);
   U12944 : AOI21_X1 port map( B1 => n11370, B2 => n11353, A => n11290, ZN => 
                           n11293);
   U12945 : NAND2_X1 port map( A1 => n11355, A2 => DRAM_DATA_OUT_6_port, ZN => 
                           n11292);
   U12946 : OAI211_X1 port map( C1 => n11373, C2 => n11293, A => n11292, B => 
                           n11291, ZN => DRAM_DATA_OUT_14_port);
   U12947 : INV_X1 port map( A => n11294, ZN => n11363);
   U12948 : OAI22_X1 port map( A1 => n11331, A2 => n11296, B1 => n11363, B2 => 
                           n11295, ZN => n11298);
   U12949 : INV_X1 port map( A => n11298, ZN => n11297);
   U12950 : OAI211_X1 port map( C1 => n8382, C2 => n11305, A => n11373, B => 
                           DRAM_DATA_OUT_7_port, ZN => n11361);
   U12951 : OAI21_X1 port map( B1 => n11373, B2 => n11297, A => n11361, ZN => 
                           DRAM_DATA_OUT_15_port);
   U12952 : NOR2_X1 port map( A1 => n392, A2 => DATA_SIZE_1_port, ZN => n11299)
                           ;
   U12953 : OAI211_X1 port map( C1 => n8382, C2 => n11305, A => n11299, B => 
                           n11298, ZN => n11360);
   U12954 : NOR2_X1 port map( A1 => n11305, A2 => n11360, ZN => n11348);
   U12955 : NAND3_X1 port map( A1 => n11305, A2 => DATA_SIZE_0_port, A3 => n393
                           , ZN => n11358);
   U12956 : NOR2_X1 port map( A1 => n11355, A2 => n11342, ZN => n11301);
   U12957 : NAND2_X1 port map( A1 => n11301, A2 => n11300, ZN => n11362);
   U12958 : INV_X1 port map( A => n11301, ZN => n11323);
   U12959 : AOI22_X1 port map( A1 => n11354, A2 => n11302, B1 => 
                           DRAM_DATA_OUT_0_port, B2 => n11323, ZN => n11303);
   U12960 : NAND2_X1 port map( A1 => n11357, A2 => n11303, ZN => 
                           DRAM_DATA_OUT_16_port);
   U12961 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(9), B1 =>
                           DataPath_i_REG_ME_DATA_DATAMEM_9_port, B2 => n11305,
                           ZN => n11330);
   U12962 : MUX2_X1 port map( A => DRAM_DATA_IN(25), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_25_port, S => n11305,
                           Z => n11369);
   U12963 : AOI22_X1 port map( A1 => n11304, A2 => n11369, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_1_port, B2 => n11305,
                           ZN => n11309);
   U12964 : MUX2_X1 port map( A => DRAM_DATA_IN(17), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_17_port, S => n11305,
                           Z => n11311);
   U12965 : AOI22_X1 port map( A1 => DRAM_DATA_IN(1), A2 => n11307, B1 => 
                           n11306, B2 => n11311, ZN => n11308);
   U12966 : OAI211_X1 port map( C1 => n11330, C2 => n11310, A => n11309, B => 
                           n11308, ZN => DRAM_DATA_OUT_1_port);
   U12967 : AOI22_X1 port map( A1 => n11354, A2 => n11311, B1 => 
                           DRAM_DATA_OUT_1_port, B2 => n11323, ZN => n11312);
   U12968 : NAND2_X1 port map( A1 => n11357, A2 => n11312, ZN => 
                           DRAM_DATA_OUT_17_port);
   U12969 : AOI22_X1 port map( A1 => n11354, A2 => n11313, B1 => 
                           DRAM_DATA_OUT_2_port, B2 => n11323, ZN => n11314);
   U12970 : NAND2_X1 port map( A1 => n11357, A2 => n11314, ZN => 
                           DRAM_DATA_OUT_18_port);
   U12971 : NAND2_X1 port map( A1 => n11323, A2 => DRAM_DATA_OUT_3_port, ZN => 
                           n11315);
   U12972 : OAI211_X1 port map( C1 => n11316, C2 => n11362, A => n11357, B => 
                           n11315, ZN => DRAM_DATA_OUT_19_port);
   U12973 : AOI22_X1 port map( A1 => n11354, A2 => n11317, B1 => 
                           DRAM_DATA_OUT_4_port, B2 => n11323, ZN => n11318);
   U12974 : NAND2_X1 port map( A1 => n11357, A2 => n11318, ZN => 
                           DRAM_DATA_OUT_20_port);
   U12975 : NAND2_X1 port map( A1 => DRAM_DATA_OUT_5_port, A2 => n11323, ZN => 
                           n11319);
   U12976 : OAI211_X1 port map( C1 => n11320, C2 => n11362, A => n11357, B => 
                           n11319, ZN => DRAM_DATA_OUT_21_port);
   U12977 : NAND2_X1 port map( A1 => n11323, A2 => DRAM_DATA_OUT_6_port, ZN => 
                           n11321);
   U12978 : OAI211_X1 port map( C1 => n11322, C2 => n11362, A => n11357, B => 
                           n11321, ZN => DRAM_DATA_OUT_22_port);
   U12979 : AOI22_X1 port map( A1 => n11354, A2 => n11324, B1 => 
                           DRAM_DATA_OUT_7_port, B2 => n11323, ZN => n11326);
   U12980 : INV_X1 port map( A => n11348, ZN => n11343);
   U12981 : NAND3_X1 port map( A1 => n11326, A2 => n11325, A3 => n11343, ZN => 
                           DRAM_DATA_OUT_23_port);
   U12982 : AOI21_X1 port map( B1 => n11355, B2 => DRAM_DATA_OUT_0_port, A => 
                           n11329, ZN => n11366);
   U12983 : NOR2_X1 port map( A1 => n11331, A2 => n11327, ZN => n11364);
   U12984 : AOI22_X1 port map( A1 => n11342, A2 => n11364, B1 => n11354, B2 => 
                           n11365, ZN => n11328);
   U12985 : NAND3_X1 port map( A1 => n11366, A2 => n11328, A3 => n11343, ZN => 
                           DRAM_DATA_OUT_24_port);
   U12986 : AOI21_X1 port map( B1 => n11355, B2 => DRAM_DATA_OUT_1_port, A => 
                           n11329, ZN => n11371);
   U12987 : NOR2_X1 port map( A1 => n11331, A2 => n11330, ZN => n11368);
   U12988 : AOI22_X1 port map( A1 => n11342, A2 => n11368, B1 => n11354, B2 => 
                           n11369, ZN => n11332);
   U12989 : NAND3_X1 port map( A1 => n11371, A2 => n11332, A3 => n11343, ZN => 
                           DRAM_DATA_OUT_25_port);
   U12990 : AOI22_X1 port map( A1 => n11342, A2 => n11334, B1 => n11354, B2 => 
                           n11333, ZN => n11335);
   U12991 : NAND3_X1 port map( A1 => n11336, A2 => n11335, A3 => n11343, ZN => 
                           DRAM_DATA_OUT_26_port);
   U12992 : AOI22_X1 port map( A1 => n11355, A2 => DRAM_DATA_OUT_3_port, B1 => 
                           n11354, B2 => n11337, ZN => n11338);
   U12993 : OAI211_X1 port map( C1 => n11339, C2 => n11358, A => n11357, B => 
                           n11338, ZN => DRAM_DATA_OUT_27_port);
   U12994 : AOI22_X1 port map( A1 => n11342, A2 => n11341, B1 => n11354, B2 => 
                           n11340, ZN => n11344);
   U12995 : NAND3_X1 port map( A1 => n11345, A2 => n11344, A3 => n11343, ZN => 
                           DRAM_DATA_OUT_28_port);
   U12996 : NAND2_X1 port map( A1 => n11347, A2 => n11346, ZN => n11352);
   U12997 : AOI21_X1 port map( B1 => n11354, B2 => n11349, A => n11348, ZN => 
                           n11350);
   U12998 : OAI211_X1 port map( C1 => n11358, C2 => n11352, A => n11351, B => 
                           n11350, ZN => DRAM_DATA_OUT_29_port);
   U12999 : AOI22_X1 port map( A1 => n11355, A2 => DRAM_DATA_OUT_6_port, B1 => 
                           n11354, B2 => n11353, ZN => n11356);
   U13000 : OAI211_X1 port map( C1 => n11359, C2 => n11358, A => n11357, B => 
                           n11356, ZN => DRAM_DATA_OUT_30_port);
   U13001 : OAI211_X1 port map( C1 => n11363, C2 => n11362, A => n11361, B => 
                           n11360, ZN => DRAM_DATA_OUT_31_port);
   U13002 : AOI21_X1 port map( B1 => n11370, B2 => n11365, A => n11364, ZN => 
                           n11367);
   U13003 : OAI21_X1 port map( B1 => n11373, B2 => n11367, A => n11366, ZN => 
                           DRAM_DATA_OUT_8_port);
   U13004 : AOI21_X1 port map( B1 => n11370, B2 => n11369, A => n11368, ZN => 
                           n11372);
   U13005 : OAI21_X1 port map( B1 => n11373, B2 => n11372, A => n11371, ZN => 
                           DRAM_DATA_OUT_9_port);
   U13006 : NAND2_X1 port map( A1 => DataPath_RF_POP_ADDRGEN_curr_state_0_port,
                           A2 => n851, ZN => n11374);
   U13007 : OAI21_X1 port map( B1 => n11376, B2 => n852, A => n12057, ZN => 
                           n11417);
   U13008 : OR2_X1 port map( A1 => RST, A2 => n11417, ZN => 
                           DataPath_RF_POP_ADDRGEN_N46);
   U13009 : OAI22_X1 port map( A1 => n11376, A2 => n853, B1 => n852, B2 => 
                           n12047, ZN => n5830);
   U13010 : OAI22_X1 port map( A1 => n11376, A2 => n854, B1 => n853, B2 => 
                           n12047, ZN => n5794);
   U13011 : OAI22_X1 port map( A1 => n11376, A2 => n855, B1 => n854, B2 => 
                           n12047, ZN => n5758);
   U13012 : OAI22_X1 port map( A1 => n11376, A2 => n856, B1 => n855, B2 => 
                           n12047, ZN => n5722);
   U13013 : OAI22_X1 port map( A1 => n11376, A2 => n857, B1 => n856, B2 => 
                           n12047, ZN => n5686);
   U13014 : OAI22_X1 port map( A1 => n11376, A2 => n858, B1 => n857, B2 => 
                           n12047, ZN => n5650);
   U13015 : OAI22_X1 port map( A1 => n11376, A2 => n859, B1 => n858, B2 => 
                           n12047, ZN => n5614);
   U13016 : OAI22_X1 port map( A1 => n11376, A2 => n860, B1 => n859, B2 => 
                           n12047, ZN => n6146);
   U13017 : OAI22_X1 port map( A1 => n11376, A2 => n861, B1 => n860, B2 => 
                           n12047, ZN => n6126);
   U13018 : OAI22_X1 port map( A1 => n11376, A2 => n862, B1 => n861, B2 => 
                           n12047, ZN => n6089);
   U13019 : OAI22_X1 port map( A1 => n11376, A2 => n863, B1 => n862, B2 => 
                           n12047, ZN => n6052);
   U13020 : OAI22_X1 port map( A1 => n11376, A2 => n864, B1 => n863, B2 => 
                           n12047, ZN => n6015);
   U13021 : OAI22_X1 port map( A1 => n11376, A2 => n865, B1 => n864, B2 => 
                           n12047, ZN => n5978);
   U13022 : OAI22_X1 port map( A1 => n11376, A2 => n866, B1 => n865, B2 => 
                           n12047, ZN => n5941);
   U13023 : AOI22_X1 port map( A1 => DataPath_RF_POP_ADDRGEN_curr_addr_15_port,
                           A2 => n12057, B1 => n11377, B2 => n8401, ZN => 
                           n12059);
   U13024 : NOR2_X1 port map( A1 => RST, A2 => n12059, ZN => 
                           DataPath_RF_POP_ADDRGEN_N61);
   U13025 : NOR2_X1 port map( A1 => RST, A2 => n12045, ZN => n11393);
   U13026 : OAI21_X1 port map( B1 => n10855, B2 => n8437, A => n11393, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N46);
   U13027 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, B1 => 
                           n11391, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, ZN => 
                           n11378);
   U13028 : NOR2_X1 port map( A1 => RST, A2 => n11378, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N47);
   U13029 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, B1 => 
                           n11391, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, ZN => 
                           n11379);
   U13030 : NOR2_X1 port map( A1 => RST, A2 => n11379, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N48);
   U13031 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, B1 => 
                           n11391, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, ZN => 
                           n11380);
   U13032 : NOR2_X1 port map( A1 => RST, A2 => n11380, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N49);
   U13033 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, B1 => 
                           n11391, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, ZN => 
                           n11381);
   U13034 : NOR2_X1 port map( A1 => RST, A2 => n11381, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N50);
   U13035 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, B1 => 
                           n11391, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, ZN => 
                           n11382);
   U13036 : NOR2_X1 port map( A1 => RST, A2 => n11382, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N51);
   U13037 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, B1 => 
                           n11391, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, ZN => 
                           n11383);
   U13038 : NOR2_X1 port map( A1 => RST, A2 => n11383, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N52);
   U13039 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, B1 => 
                           n11391, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, ZN => 
                           n11384);
   U13040 : NOR2_X1 port map( A1 => RST, A2 => n11384, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N53);
   U13041 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, B1 => 
                           n11391, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, ZN => 
                           n11385);
   U13042 : NOR2_X1 port map( A1 => RST, A2 => n11385, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N54);
   U13043 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, B1 => 
                           n11391, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, ZN => 
                           n11386);
   U13044 : NOR2_X1 port map( A1 => RST, A2 => n11386, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N55);
   U13045 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, B1 => 
                           n11391, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, ZN => 
                           n11387);
   U13046 : NOR2_X1 port map( A1 => RST, A2 => n11387, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N56);
   U13047 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, B1 => 
                           n11391, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, ZN => 
                           n11388);
   U13048 : NOR2_X1 port map( A1 => RST, A2 => n11388, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N57);
   U13049 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, B1 => 
                           n11391, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, ZN => 
                           n11389);
   U13050 : NOR2_X1 port map( A1 => RST, A2 => n11389, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N58);
   U13051 : AOI22_X1 port map( A1 => n10855, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, B2 => 
                           n11391, ZN => n11390);
   U13052 : NOR2_X1 port map( A1 => RST, A2 => n11390, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N59);
   U13053 : AOI22_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_addr_14_port
                           , A2 => n11391, B1 => n10855, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, ZN => 
                           n11392);
   U13054 : NOR2_X1 port map( A1 => RST, A2 => n11392, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N60);
   U13055 : INV_X1 port map( A => n11393, ZN => n12046);
   U13056 : NOR2_X1 port map( A1 => n11394, A2 => n12046, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N61);
   U13057 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_10_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N14);
   U13058 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_12_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N16);
   U13059 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_14_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N18);
   U13060 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_15_port, A2 => 
                           n8689, ZN => DataPath_RF_RDPORT0_OUTLATCH_N19);
   U13061 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_16_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N20);
   U13062 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_17_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N21);
   U13063 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_18_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N22);
   U13064 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_19_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N23);
   U13065 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_21_port, A2 => 
                           n8688, ZN => DataPath_RF_RDPORT0_OUTLATCH_N25);
   U13066 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_23_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N27);
   U13067 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_24_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N28);
   U13068 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_25_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N29);
   U13069 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_26_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N30);
   U13070 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_27_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N31);
   U13071 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_28_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N32);
   U13072 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_29_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N33);
   U13073 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_30_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N34);
   U13074 : AND2_X1 port map( A1 => DataPath_RF_internal_out1_1_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT0_OUTLATCH_N5);
   U13075 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_10_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N14);
   U13076 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_12_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N16);
   U13077 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_14_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N18);
   U13078 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_15_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N19);
   U13079 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_16_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N20);
   U13080 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_17_port, A2 => 
                           n8695, ZN => DataPath_RF_RDPORT1_OUTLATCH_N21);
   U13081 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_18_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N22);
   U13082 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_19_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N23);
   U13083 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_22_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N26);
   U13084 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_23_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N27);
   U13085 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_24_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N28);
   U13086 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_25_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N29);
   U13087 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_26_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N30);
   U13088 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_27_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N31);
   U13089 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_28_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N32);
   U13090 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_29_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N33);
   U13091 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_30_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N34);
   U13092 : AND2_X1 port map( A1 => DataPath_RF_internal_out2_2_port, A2 => 
                           n8694, ZN => DataPath_RF_RDPORT1_OUTLATCH_N6);
   U13093 : NAND2_X1 port map( A1 => n11889, A2 => n11413, ZN => n11824);
   U13094 : NAND2_X1 port map( A1 => n11889, A2 => n11414, ZN => n11823);
   U13095 : OAI22_X1 port map( A1 => n577, A2 => n11824, B1 => n8441, B2 => 
                           n11823, ZN => n11396);
   U13096 : MUX2_X1 port map( A => DRAMRF_DATA_IN(16), B => 
                           DataPath_WRF_CUhw_curr_data_16_port, S => n10868, Z 
                           => n11754);
   U13097 : NAND2_X1 port map( A1 => n8692, A2 => n11754, ZN => n3341);
   U13098 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2288_port, B1 => n12159,
                           B2 => n8669, ZN => n6142);
   U13099 : MUX2_X1 port map( A => DRAMRF_DATA_IN(17), B => 
                           DataPath_WRF_CUhw_curr_data_17_port, S => n10868, Z 
                           => n11633);
   U13100 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2289_port, B1 => n12160,
                           B2 => n8669, ZN => n6141);
   U13101 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(18), B1
                           => DataPath_WRF_CUhw_curr_data_18_port, B2 => n10868
                           , ZN => n11755);
   U13102 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2290_port, B1 => n12161,
                           B2 => n8669, ZN => n6140);
   U13103 : MUX2_X1 port map( A => DRAMRF_DATA_IN(19), B => 
                           DataPath_WRF_CUhw_curr_data_19_port, S => n10868, Z 
                           => n11756);
   U13104 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2291_port, B1 => n12162,
                           B2 => n8669, ZN => n6139);
   U13105 : MUX2_X1 port map( A => DRAMRF_DATA_IN(20), B => 
                           DataPath_WRF_CUhw_curr_data_20_port, S => n10868, Z 
                           => n11757);
   U13106 : AOI22_X1 port map( A1 => n8679, A2 => 
                           DataPath_i_REG_LDSTR_OUT_20_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_20_port, B2 => n8411, ZN 
                           => n11936);
   U13107 : AOI22_X1 port map( A1 => n12193, A2 => 
                           DataPath_RF_bus_reg_dataout_2292_port, B1 => n12163,
                           B2 => n8669, ZN => n6138);
   U13108 : MUX2_X1 port map( A => DRAMRF_DATA_IN(21), B => 
                           DataPath_WRF_CUhw_curr_data_21_port, S => n10868, Z 
                           => n11758);
   U13109 : AOI22_X1 port map( A1 => n8679, A2 => 
                           DataPath_i_REG_LDSTR_OUT_21_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_21_port, B2 => n8411, ZN 
                           => n11937);
   U13110 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2293_port, B1 => n12164,
                           B2 => n8669, ZN => n6137);
   U13111 : MUX2_X1 port map( A => DRAMRF_DATA_IN(22), B => 
                           DataPath_WRF_CUhw_curr_data_22_port, S => n10868, Z 
                           => n11759);
   U13112 : AOI22_X1 port map( A1 => n8679, A2 => 
                           DataPath_i_REG_LDSTR_OUT_22_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_22_port, B2 => n8411, ZN 
                           => n11938);
   U13113 : AOI22_X1 port map( A1 => n12193, A2 => 
                           DataPath_RF_bus_reg_dataout_2294_port, B1 => n12165,
                           B2 => n8669, ZN => n6136);
   U13114 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(23), B1
                           => DataPath_WRF_CUhw_curr_data_23_port, B2 => n10868
                           , ZN => n11968);
   U13115 : AOI22_X1 port map( A1 => n8679, A2 => 
                           DataPath_i_REG_LDSTR_OUT_23_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_23_port, B2 => n8411, ZN 
                           => n11939);
   U13116 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2295_port, B1 => n12166,
                           B2 => n8669, ZN => n6135);
   U13117 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(24), B1
                           => DataPath_WRF_CUhw_curr_data_24_port, B2 => n10868
                           , ZN => n11969);
   U13118 : AOI22_X1 port map( A1 => n8679, A2 => 
                           DataPath_i_REG_LDSTR_OUT_24_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_24_port, B2 => n8411, ZN 
                           => n11940);
   U13119 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2296_port, B1 => n12167,
                           B2 => n8669, ZN => n6134);
   U13120 : MUX2_X1 port map( A => DRAMRF_DATA_IN(25), B => 
                           DataPath_WRF_CUhw_curr_data_25_port, S => n10868, Z 
                           => n11760);
   U13121 : AOI22_X1 port map( A1 => n8679, A2 => 
                           DataPath_i_REG_LDSTR_OUT_25_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_25_port, B2 => n8411, ZN 
                           => n11941);
   U13122 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2297_port, B1 => n12168,
                           B2 => n8669, ZN => n6133);
   U13123 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(26), B1
                           => DataPath_WRF_CUhw_curr_data_26_port, B2 => n10868
                           , ZN => n11970);
   U13124 : AOI22_X1 port map( A1 => n8679, A2 => 
                           DataPath_i_REG_LDSTR_OUT_26_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_26_port, B2 => n8411, ZN 
                           => n11942);
   U13125 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2298_port, B1 => n12169,
                           B2 => n8669, ZN => n6132);
   U13126 : MUX2_X1 port map( A => DRAMRF_DATA_IN(27), B => 
                           DataPath_WRF_CUhw_curr_data_27_port, S => n10868, Z 
                           => n11761);
   U13127 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2299_port, B1 => n12170,
                           B2 => n8669, ZN => n6131);
   U13128 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(28), B1
                           => DataPath_WRF_CUhw_curr_data_28_port, B2 => n10868
                           , ZN => n11971);
   U13129 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_28_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_28_port, B2 => n8411, ZN 
                           => n11944);
   U13130 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2300_port, B1 => n12171,
                           B2 => n8669, ZN => n6130);
   U13131 : MUX2_X1 port map( A => DRAMRF_DATA_IN(29), B => 
                           DataPath_WRF_CUhw_curr_data_29_port, S => n10868, Z 
                           => n11762);
   U13132 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_29_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_29_port, B2 => n8411, ZN 
                           => n11945);
   U13133 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2301_port, B1 => n12172,
                           B2 => n8669, ZN => n6129);
   U13134 : MUX2_X1 port map( A => DRAMRF_DATA_IN(30), B => 
                           DataPath_WRF_CUhw_curr_data_30_port, S => n10868, Z 
                           => n11763);
   U13135 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_30_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_30_port, B2 => n8411, ZN 
                           => n11946);
   U13136 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2302_port, B1 => n12173,
                           B2 => n8669, ZN => n6128);
   U13137 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_31_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_31_port, B2 => n8411, ZN 
                           => n11949);
   U13138 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(31), B1
                           => DataPath_WRF_CUhw_curr_data_31_port, B2 => n10868
                           , ZN => n11764);
   U13139 : OR2_X1 port map( A1 => RST, A2 => n11764, ZN => n3324);
   U13140 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2303_port, B1 => n12175,
                           B2 => n8669, ZN => n6127);
   U13141 : NAND2_X1 port map( A1 => n11893, A2 => n11413, ZN => n11829);
   U13142 : NAND2_X1 port map( A1 => n11893, A2 => n11414, ZN => n11828);
   U13143 : OAI22_X1 port map( A1 => n577, A2 => n11829, B1 => n8441, B2 => 
                           n11828, ZN => n11397);
   U13144 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(0), B1 
                           => DataPath_WRF_CUhw_curr_data_0_port, B2 => n10868,
                           ZN => n11956);
   U13145 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_0_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_0_port, B2 => n8680, ZN =>
                           n11916);
   U13146 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2240_port, B1 => n12177,
                           B2 => n11398, ZN => n6123);
   U13147 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(1), B1 
                           => DataPath_WRF_CUhw_curr_data_1_port, B2 => n10868,
                           ZN => n11957);
   U13148 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_1_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_1_port, B2 => n8411, ZN =>
                           n11917);
   U13149 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2241_port, B1 => n12178,
                           B2 => n11398, ZN => n6122);
   U13150 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(2), B1 
                           => DataPath_WRF_CUhw_curr_data_2_port, B2 => n10868,
                           ZN => n11958);
   U13151 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_2_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_2_port, B2 => n8680, ZN =>
                           n11918);
   U13152 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2242_port, B1 => n12179,
                           B2 => n11398, ZN => n6121);
   U13153 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(3), B1 
                           => DataPath_WRF_CUhw_curr_data_3_port, B2 => n10868,
                           ZN => n11959);
   U13154 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_3_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_3_port, B2 => n8680, ZN =>
                           n11919);
   U13155 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2243_port, B1 => n12180,
                           B2 => n11398, ZN => n6120);
   U13156 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(4), B1 
                           => DataPath_WRF_CUhw_curr_data_4_port, B2 => n10868,
                           ZN => n11960);
   U13157 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_4_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_4_port, B2 => n8411, ZN =>
                           n11920);
   U13158 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2244_port, B1 => n12181,
                           B2 => n11398, ZN => n6119);
   U13159 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(5), B1 
                           => DataPath_WRF_CUhw_curr_data_5_port, B2 => n10868,
                           ZN => n11961);
   U13160 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_5_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_5_port, B2 => n8411, ZN =>
                           n11921);
   U13161 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2245_port, B1 => n12182,
                           B2 => n11398, ZN => n6118);
   U13162 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(6), B1 
                           => DataPath_WRF_CUhw_curr_data_6_port, B2 => n10868,
                           ZN => n11962);
   U13163 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_6_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_6_port, B2 => n8411, ZN =>
                           n11922);
   U13164 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2246_port, B1 => n12183,
                           B2 => n11398, ZN => n6117);
   U13165 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(7), B1 
                           => DataPath_WRF_CUhw_curr_data_7_port, B2 => n10868,
                           ZN => n11750);
   U13166 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2247_port, B1 => n12184,
                           B2 => n11398, ZN => n6116);
   U13167 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(8), B1 
                           => DataPath_WRF_CUhw_curr_data_8_port, B2 => n10868,
                           ZN => n11963);
   U13168 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_8_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_8_port, B2 => n8680, ZN =>
                           n11924);
   U13169 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2248_port, B1 => n12185,
                           B2 => n11398, ZN => n6115);
   U13170 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(9), B1 
                           => DataPath_WRF_CUhw_curr_data_9_port, B2 => n10868,
                           ZN => n11964);
   U13171 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_9_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_9_port, B2 => n8411, ZN =>
                           n11925);
   U13172 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2249_port, B1 => n12186,
                           B2 => n11398, ZN => n6114);
   U13173 : MUX2_X1 port map( A => DRAMRF_DATA_IN(10), B => 
                           DataPath_WRF_CUhw_curr_data_10_port, S => n10868, Z 
                           => n11751);
   U13174 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2250_port, B1 => n12187,
                           B2 => n11398, ZN => n6113);
   U13175 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(11), B1
                           => DataPath_WRF_CUhw_curr_data_11_port, B2 => n10868
                           , ZN => n11965);
   U13176 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_11_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_11_port, B2 => n8411, ZN 
                           => n11927);
   U13177 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2251_port, B1 => n12188,
                           B2 => n11398, ZN => n6112);
   U13178 : MUX2_X1 port map( A => DRAMRF_DATA_IN(12), B => 
                           DataPath_WRF_CUhw_curr_data_12_port, S => n10868, Z 
                           => n11752);
   U13179 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2252_port, B1 => n12189,
                           B2 => n11398, ZN => n6111);
   U13180 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(13), B1
                           => DataPath_WRF_CUhw_curr_data_13_port, B2 => n10868
                           , ZN => n11966);
   U13181 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_13_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_13_port, B2 => n8411, ZN 
                           => n11929);
   U13182 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2253_port, B1 => n12190,
                           B2 => n11398, ZN => n6110);
   U13183 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => DRAMRF_DATA_IN(14), B1
                           => DataPath_WRF_CUhw_curr_data_14_port, B2 => n10868
                           , ZN => n11967);
   U13184 : AOI22_X1 port map( A1 => n8301, A2 => 
                           DataPath_i_REG_LDSTR_OUT_14_port, B1 => 
                           DataPath_i_REG_MEM_ALUOUT_14_port, B2 => n8411, ZN 
                           => n11930);
   U13185 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2254_port, B1 => n12191,
                           B2 => n11398, ZN => n6109);
   U13186 : MUX2_X1 port map( A => DRAMRF_DATA_IN(15), B => 
                           DataPath_WRF_CUhw_curr_data_15_port, S => n10868, Z 
                           => n11631);
   U13187 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2255_port, B1 => n12192,
                           B2 => n11398, ZN => n6108);
   U13188 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2256_port, B1 => n12159,
                           B2 => n11398, ZN => n6107);
   U13189 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2257_port, B1 => n12160,
                           B2 => n11398, ZN => n6106);
   U13190 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2258_port, B1 => n12161,
                           B2 => n11398, ZN => n6105);
   U13191 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2259_port, B1 => n12162,
                           B2 => n11398, ZN => n6104);
   U13192 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2260_port, B1 => n12163,
                           B2 => n11398, ZN => n6103);
   U13193 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2261_port, B1 => n12164,
                           B2 => n11398, ZN => n6102);
   U13194 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2262_port, B1 => n12165,
                           B2 => n11398, ZN => n6101);
   U13195 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2263_port, B1 => n12166,
                           B2 => n11398, ZN => n6100);
   U13196 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2264_port, B1 => n12167,
                           B2 => n11398, ZN => n6099);
   U13197 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2265_port, B1 => n12168,
                           B2 => n11398, ZN => n6098);
   U13198 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2266_port, B1 => n12169,
                           B2 => n11398, ZN => n6097);
   U13199 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2267_port, B1 => n12170,
                           B2 => n11398, ZN => n6096);
   U13200 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2268_port, B1 => n12171,
                           B2 => n11398, ZN => n6095);
   U13201 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2269_port, B1 => n12172,
                           B2 => n11398, ZN => n6094);
   U13202 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2270_port, B1 => n12173,
                           B2 => n11398, ZN => n6093);
   U13203 : AOI22_X1 port map( A1 => n8506, A2 => 
                           DataPath_RF_bus_reg_dataout_2271_port, B1 => n12175,
                           B2 => n11398, ZN => n6090);
   U13204 : NAND2_X1 port map( A1 => n11897, A2 => n11414, ZN => n11552);
   U13205 : NAND2_X1 port map( A1 => n11897, A2 => n11413, ZN => n11833);
   U13206 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2208_port, B1 => n12177,
                           B2 => n11401, ZN => n6086);
   U13207 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2209_port, B1 => n12178,
                           B2 => n11401, ZN => n6085);
   U13208 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2210_port, B1 => n12179,
                           B2 => n11401, ZN => n6084);
   U13209 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2211_port, B1 => n12180,
                           B2 => n11401, ZN => n6083);
   U13210 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2212_port, B1 => n12181,
                           B2 => n11401, ZN => n6082);
   U13211 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2213_port, B1 => n12182,
                           B2 => n11401, ZN => n6081);
   U13212 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2214_port, B1 => n12183,
                           B2 => n11401, ZN => n6080);
   U13213 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2215_port, B1 => n12184,
                           B2 => n11401, ZN => n6079);
   U13214 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2216_port, B1 => n12185,
                           B2 => n11401, ZN => n6078);
   U13215 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2217_port, B1 => n12186,
                           B2 => n11401, ZN => n6077);
   U13216 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2218_port, B1 => n12187,
                           B2 => n11401, ZN => n6076);
   U13217 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2219_port, B1 => n12188,
                           B2 => n11401, ZN => n6075);
   U13218 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2220_port, B1 => n12189,
                           B2 => n11401, ZN => n6074);
   U13219 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2221_port, B1 => n12190,
                           B2 => n11401, ZN => n6073);
   U13220 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2222_port, B1 => n12191,
                           B2 => n11401, ZN => n6072);
   U13221 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2223_port, B1 => n12192,
                           B2 => n11401, ZN => n6071);
   U13222 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2224_port, B1 => n12159,
                           B2 => n11401, ZN => n6070);
   U13223 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2225_port, B1 => n12160,
                           B2 => n11401, ZN => n6069);
   U13224 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2226_port, B1 => n12161,
                           B2 => n11401, ZN => n6068);
   U13225 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2227_port, B1 => n12162,
                           B2 => n11401, ZN => n6067);
   U13226 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2228_port, B1 => n12163,
                           B2 => n11401, ZN => n6066);
   U13227 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2229_port, B1 => n12164,
                           B2 => n11401, ZN => n6065);
   U13228 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2230_port, B1 => n12165,
                           B2 => n11401, ZN => n6064);
   U13229 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2231_port, B1 => n12166,
                           B2 => n11401, ZN => n6063);
   U13230 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2232_port, B1 => n12167,
                           B2 => n11401, ZN => n6062);
   U13231 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2233_port, B1 => n12168,
                           B2 => n11401, ZN => n6061);
   U13232 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2234_port, B1 => n12169,
                           B2 => n11401, ZN => n6060);
   U13233 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2235_port, B1 => n12170,
                           B2 => n11401, ZN => n6059);
   U13234 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2236_port, B1 => n12171,
                           B2 => n11401, ZN => n6058);
   U13235 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2237_port, B1 => n12172,
                           B2 => n11401, ZN => n6057);
   U13236 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2238_port, B1 => n12173,
                           B2 => n11401, ZN => n6056);
   U13237 : AOI22_X1 port map( A1 => n11402, A2 => 
                           DataPath_RF_bus_reg_dataout_2239_port, B1 => n12175,
                           B2 => n11401, ZN => n6053);
   U13238 : NAND2_X1 port map( A1 => n11901, A2 => n11413, ZN => n11839);
   U13239 : NAND2_X1 port map( A1 => n11901, A2 => n11414, ZN => n11838);
   U13240 : OAI22_X1 port map( A1 => n577, A2 => n11839, B1 => n8441, B2 => 
                           n11838, ZN => n11403);
   U13241 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2176_port, B1 => n12177,
                           B2 => n11404, ZN => n6049);
   U13242 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2177_port, B1 => n12178,
                           B2 => n11404, ZN => n6048);
   U13243 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2178_port, B1 => n12179,
                           B2 => n11404, ZN => n6047);
   U13244 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2179_port, B1 => n12180,
                           B2 => n11404, ZN => n6046);
   U13245 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2180_port, B1 => n12181,
                           B2 => n11404, ZN => n6045);
   U13246 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2181_port, B1 => n12182,
                           B2 => n11404, ZN => n6044);
   U13247 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2182_port, B1 => n12183,
                           B2 => n11404, ZN => n6043);
   U13248 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2183_port, B1 => n12184,
                           B2 => n11404, ZN => n6042);
   U13249 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2184_port, B1 => n12185,
                           B2 => n11404, ZN => n6041);
   U13250 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2185_port, B1 => n12186,
                           B2 => n11404, ZN => n6040);
   U13251 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2186_port, B1 => n12187,
                           B2 => n11404, ZN => n6039);
   U13252 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2187_port, B1 => n12188,
                           B2 => n11404, ZN => n6038);
   U13253 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2188_port, B1 => n12189,
                           B2 => n11404, ZN => n6037);
   U13254 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2189_port, B1 => n12190,
                           B2 => n11404, ZN => n6036);
   U13255 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2190_port, B1 => n12191,
                           B2 => n11404, ZN => n6035);
   U13256 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2191_port, B1 => n12192,
                           B2 => n11404, ZN => n6034);
   U13257 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2192_port, B1 => n12159,
                           B2 => n11404, ZN => n6033);
   U13258 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2193_port, B1 => n12160,
                           B2 => n11404, ZN => n6032);
   U13259 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2194_port, B1 => n12161,
                           B2 => n11404, ZN => n6031);
   U13260 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2195_port, B1 => n12162,
                           B2 => n11404, ZN => n6030);
   U13261 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2196_port, B1 => n12163,
                           B2 => n11404, ZN => n6029);
   U13262 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2197_port, B1 => n12164,
                           B2 => n11404, ZN => n6028);
   U13263 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2198_port, B1 => n12165,
                           B2 => n11404, ZN => n6027);
   U13264 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2199_port, B1 => n12166,
                           B2 => n11404, ZN => n6026);
   U13265 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2200_port, B1 => n12167,
                           B2 => n11404, ZN => n6025);
   U13266 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2201_port, B1 => n12168,
                           B2 => n11404, ZN => n6024);
   U13267 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2202_port, B1 => n12169,
                           B2 => n11404, ZN => n6023);
   U13268 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2203_port, B1 => n12170,
                           B2 => n11404, ZN => n6022);
   U13269 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2204_port, B1 => n12171,
                           B2 => n11404, ZN => n6021);
   U13270 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2205_port, B1 => n12172,
                           B2 => n11404, ZN => n6020);
   U13271 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2206_port, B1 => n12173,
                           B2 => n11404, ZN => n6019);
   U13272 : AOI22_X1 port map( A1 => n8507, A2 => 
                           DataPath_RF_bus_reg_dataout_2207_port, B1 => n12175,
                           B2 => n11404, ZN => n6016);
   U13273 : NAND2_X1 port map( A1 => n11905, A2 => n11414, ZN => n11589);
   U13274 : NAND2_X1 port map( A1 => n11905, A2 => n11413, ZN => n11842);
   U13275 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2144_port, B1 => n12177,
                           B2 => n11407, ZN => n6012);
   U13276 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2145_port, B1 => n12178,
                           B2 => n11407, ZN => n6011);
   U13277 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2146_port, B1 => n12179,
                           B2 => n11407, ZN => n6010);
   U13278 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2147_port, B1 => n12180,
                           B2 => n11407, ZN => n6009);
   U13279 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2148_port, B1 => n12181,
                           B2 => n11407, ZN => n6008);
   U13280 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2149_port, B1 => n12182,
                           B2 => n11407, ZN => n6007);
   U13281 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2150_port, B1 => n12183,
                           B2 => n11407, ZN => n6006);
   U13282 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2151_port, B1 => n12184,
                           B2 => n11407, ZN => n6005);
   U13283 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2152_port, B1 => n12185,
                           B2 => n11407, ZN => n6004);
   U13284 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2153_port, B1 => n12186,
                           B2 => n11407, ZN => n6003);
   U13285 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2154_port, B1 => n12187,
                           B2 => n11407, ZN => n6002);
   U13286 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2155_port, B1 => n12188,
                           B2 => n11407, ZN => n6001);
   U13287 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2156_port, B1 => n12189,
                           B2 => n11407, ZN => n6000);
   U13288 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2157_port, B1 => n12190,
                           B2 => n11407, ZN => n5999);
   U13289 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2158_port, B1 => n12191,
                           B2 => n11407, ZN => n5998);
   U13290 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2159_port, B1 => n12192,
                           B2 => n11407, ZN => n5997);
   U13291 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2160_port, B1 => n12159,
                           B2 => n11407, ZN => n5996);
   U13292 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2161_port, B1 => n12160,
                           B2 => n11407, ZN => n5995);
   U13293 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2162_port, B1 => n12161,
                           B2 => n11407, ZN => n5994);
   U13294 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2163_port, B1 => n12162,
                           B2 => n11407, ZN => n5993);
   U13295 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2164_port, B1 => n12163,
                           B2 => n11407, ZN => n5992);
   U13296 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2165_port, B1 => n12164,
                           B2 => n11407, ZN => n5991);
   U13297 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2166_port, B1 => n12165,
                           B2 => n11407, ZN => n5990);
   U13298 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2167_port, B1 => n12166,
                           B2 => n11407, ZN => n5989);
   U13299 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2168_port, B1 => n12167,
                           B2 => n11407, ZN => n5988);
   U13300 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2169_port, B1 => n12168,
                           B2 => n11407, ZN => n5987);
   U13301 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2170_port, B1 => n12169,
                           B2 => n11407, ZN => n5986);
   U13302 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2171_port, B1 => n12170,
                           B2 => n11407, ZN => n5985);
   U13303 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2172_port, B1 => n12171,
                           B2 => n11407, ZN => n5984);
   U13304 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2173_port, B1 => n12172,
                           B2 => n11407, ZN => n5983);
   U13305 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2174_port, B1 => n12173,
                           B2 => n11407, ZN => n5982);
   U13306 : AOI22_X1 port map( A1 => n11408, A2 => 
                           DataPath_RF_bus_reg_dataout_2175_port, B1 => n12175,
                           B2 => n11407, ZN => n5979);
   U13307 : NAND2_X1 port map( A1 => n11909, A2 => n11413, ZN => n11848);
   U13308 : NAND2_X1 port map( A1 => n11909, A2 => n11414, ZN => n11847);
   U13309 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2112_port, B1 => n12177,
                           B2 => n11409, ZN => n5975);
   U13310 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2113_port, B1 => n12178,
                           B2 => n11409, ZN => n5974);
   U13311 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2114_port, B1 => n12179,
                           B2 => n11409, ZN => n5973);
   U13312 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2115_port, B1 => n12180,
                           B2 => n11409, ZN => n5972);
   U13313 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2116_port, B1 => n12181,
                           B2 => n11409, ZN => n5971);
   U13314 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2117_port, B1 => n12182,
                           B2 => n11409, ZN => n5970);
   U13315 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2118_port, B1 => n12183,
                           B2 => n11409, ZN => n5969);
   U13316 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2119_port, B1 => n12184,
                           B2 => n11409, ZN => n5968);
   U13317 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2120_port, B1 => n12185,
                           B2 => n11409, ZN => n5967);
   U13318 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2121_port, B1 => n12186,
                           B2 => n11409, ZN => n5966);
   U13319 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2122_port, B1 => n12187,
                           B2 => n11409, ZN => n5965);
   U13320 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2123_port, B1 => n12188,
                           B2 => n11409, ZN => n5964);
   U13321 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2124_port, B1 => n12189,
                           B2 => n11409, ZN => n5963);
   U13322 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2125_port, B1 => n12190,
                           B2 => n11409, ZN => n5962);
   U13323 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2126_port, B1 => n12191,
                           B2 => n11409, ZN => n5961);
   U13324 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2127_port, B1 => n12192,
                           B2 => n11409, ZN => n5960);
   U13325 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2128_port, B1 => n12159,
                           B2 => n11409, ZN => n5959);
   U13326 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2129_port, B1 => n12160,
                           B2 => n11409, ZN => n5958);
   U13327 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2130_port, B1 => n12161,
                           B2 => n11409, ZN => n5957);
   U13328 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2131_port, B1 => n12162,
                           B2 => n11409, ZN => n5956);
   U13329 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2132_port, B1 => n12163,
                           B2 => n11409, ZN => n5955);
   U13330 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2133_port, B1 => n12164,
                           B2 => n11409, ZN => n5954);
   U13331 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2134_port, B1 => n12165,
                           B2 => n11409, ZN => n5953);
   U13332 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2135_port, B1 => n12166,
                           B2 => n11409, ZN => n5952);
   U13333 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2136_port, B1 => n12167,
                           B2 => n11409, ZN => n5951);
   U13334 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2137_port, B1 => n12168,
                           B2 => n11409, ZN => n5950);
   U13335 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2138_port, B1 => n12169,
                           B2 => n11409, ZN => n5949);
   U13336 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2139_port, B1 => n12170,
                           B2 => n11409, ZN => n5948);
   U13337 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2140_port, B1 => n12171,
                           B2 => n11409, ZN => n5947);
   U13338 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2141_port, B1 => n12172,
                           B2 => n11409, ZN => n5946);
   U13339 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2142_port, B1 => n12173,
                           B2 => n11409, ZN => n5945);
   U13340 : AOI22_X1 port map( A1 => n8508, A2 => 
                           DataPath_RF_bus_reg_dataout_2143_port, B1 => n12175,
                           B2 => n11409, ZN => n5942);
   U13341 : NAND2_X1 port map( A1 => n11914, A2 => n11413, ZN => n11852);
   U13342 : NAND2_X1 port map( A1 => n11914, A2 => n11414, ZN => n11851);
   U13343 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2080_port, B1 => n12177,
                           B2 => n11411, ZN => n5938);
   U13344 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2081_port, B1 => n12178,
                           B2 => n11411, ZN => n5937);
   U13345 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2082_port, B1 => n12179,
                           B2 => n11411, ZN => n5936);
   U13346 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2083_port, B1 => n12180,
                           B2 => n11411, ZN => n5935);
   U13347 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2084_port, B1 => n12181,
                           B2 => n11411, ZN => n5934);
   U13348 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2085_port, B1 => n12182,
                           B2 => n11411, ZN => n5933);
   U13349 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2086_port, B1 => n12183,
                           B2 => n11411, ZN => n5932);
   U13350 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2087_port, B1 => n12184,
                           B2 => n11411, ZN => n5931);
   U13351 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2088_port, B1 => n12185,
                           B2 => n11411, ZN => n5930);
   U13352 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2089_port, B1 => n12186,
                           B2 => n11411, ZN => n5929);
   U13353 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2090_port, B1 => n12187,
                           B2 => n11411, ZN => n5928);
   U13354 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2091_port, B1 => n12188,
                           B2 => n11411, ZN => n5927);
   U13355 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2092_port, B1 => n12189,
                           B2 => n11411, ZN => n5926);
   U13356 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2093_port, B1 => n12190,
                           B2 => n11411, ZN => n5925);
   U13357 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2094_port, B1 => n12191,
                           B2 => n11411, ZN => n5924);
   U13358 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2095_port, B1 => n12192,
                           B2 => n11411, ZN => n5923);
   U13359 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2096_port, B1 => n12159,
                           B2 => n11411, ZN => n5922);
   U13360 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2097_port, B1 => n12160,
                           B2 => n11411, ZN => n5921);
   U13361 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2098_port, B1 => n12161,
                           B2 => n11411, ZN => n5920);
   U13362 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2099_port, B1 => n12162,
                           B2 => n11411, ZN => n5919);
   U13363 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2100_port, B1 => n12163,
                           B2 => n11411, ZN => n5918);
   U13364 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2101_port, B1 => n12164,
                           B2 => n11411, ZN => n5917);
   U13365 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2102_port, B1 => n12165,
                           B2 => n11411, ZN => n5916);
   U13366 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2103_port, B1 => n12166,
                           B2 => n11411, ZN => n5915);
   U13367 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2104_port, B1 => n12167,
                           B2 => n11411, ZN => n5914);
   U13368 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2105_port, B1 => n12168,
                           B2 => n11411, ZN => n5913);
   U13369 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2106_port, B1 => n12169,
                           B2 => n11411, ZN => n5912);
   U13370 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2107_port, B1 => n12170,
                           B2 => n11411, ZN => n5911);
   U13371 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2108_port, B1 => n12171,
                           B2 => n11411, ZN => n5910);
   U13372 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2109_port, B1 => n12172,
                           B2 => n11411, ZN => n5909);
   U13373 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2110_port, B1 => n12173,
                           B2 => n11411, ZN => n5908);
   U13374 : AOI22_X1 port map( A1 => n8509, A2 => 
                           DataPath_RF_bus_reg_dataout_2111_port, B1 => n12175,
                           B2 => n11411, ZN => n5905);
   U13375 : NAND2_X1 port map( A1 => n11455, A2 => n11413, ZN => n11856);
   U13376 : NAND2_X1 port map( A1 => n11455, A2 => n11414, ZN => n11855);
   U13377 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2048_port, B1 => n12177,
                           B2 => n11415, ZN => n5900);
   U13378 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2049_port, B1 => n12178,
                           B2 => n11415, ZN => n5899);
   U13379 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2050_port, B1 => n12179,
                           B2 => n11415, ZN => n5898);
   U13380 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2051_port, B1 => n12180,
                           B2 => n11415, ZN => n5897);
   U13381 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2052_port, B1 => n12181,
                           B2 => n11415, ZN => n5896);
   U13382 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2053_port, B1 => n12182,
                           B2 => n11415, ZN => n5895);
   U13383 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2054_port, B1 => n12183,
                           B2 => n11415, ZN => n5894);
   U13384 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2055_port, B1 => n12184,
                           B2 => n11415, ZN => n5893);
   U13385 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2056_port, B1 => n12185,
                           B2 => n11415, ZN => n5892);
   U13386 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2057_port, B1 => n12186,
                           B2 => n11415, ZN => n5891);
   U13387 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2058_port, B1 => n12187,
                           B2 => n11415, ZN => n5890);
   U13388 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2059_port, B1 => n12188,
                           B2 => n11415, ZN => n5889);
   U13389 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2060_port, B1 => n12189,
                           B2 => n11415, ZN => n5888);
   U13390 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2061_port, B1 => n12190,
                           B2 => n11415, ZN => n5887);
   U13391 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2062_port, B1 => n12191,
                           B2 => n11415, ZN => n5886);
   U13392 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2063_port, B1 => n12192,
                           B2 => n11415, ZN => n5885);
   U13393 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2064_port, B1 => n12159,
                           B2 => n11415, ZN => n5884);
   U13394 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2065_port, B1 => n12160,
                           B2 => n11415, ZN => n5883);
   U13395 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2066_port, B1 => n12161,
                           B2 => n11415, ZN => n5882);
   U13396 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2067_port, B1 => n12162,
                           B2 => n11415, ZN => n5881);
   U13397 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2068_port, B1 => n12163,
                           B2 => n11415, ZN => n5880);
   U13398 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2069_port, B1 => n12164,
                           B2 => n11415, ZN => n5879);
   U13399 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2070_port, B1 => n12165,
                           B2 => n11415, ZN => n5878);
   U13400 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2071_port, B1 => n12166,
                           B2 => n11415, ZN => n5877);
   U13401 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2072_port, B1 => n12167,
                           B2 => n11415, ZN => n5876);
   U13402 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2073_port, B1 => n12168,
                           B2 => n11415, ZN => n5875);
   U13403 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2074_port, B1 => n12169,
                           B2 => n11415, ZN => n5874);
   U13404 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2075_port, B1 => n12170,
                           B2 => n11415, ZN => n5873);
   U13405 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2076_port, B1 => n12171,
                           B2 => n11415, ZN => n5872);
   U13406 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2077_port, B1 => n12172,
                           B2 => n11415, ZN => n5871);
   U13407 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2078_port, B1 => n12173,
                           B2 => n11415, ZN => n5870);
   U13408 : AOI22_X1 port map( A1 => n8510, A2 => 
                           DataPath_RF_bus_reg_dataout_2079_port, B1 => n12175,
                           B2 => n11415, ZN => n5867);
   U13409 : NAND2_X1 port map( A1 => n11889, A2 => n11456, ZN => n12094);
   U13410 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2016_port, A2 
                           => n8609, B1 => n11420, B2 => n11432, ZN => n5864);
   U13411 : AOI22_X1 port map( A1 => n11420, A2 => n11433, B1 => n11419, B2 => 
                           DataPath_RF_bus_reg_dataout_2017_port, ZN => n5863);
   U13412 : AOI22_X1 port map( A1 => n11420, A2 => n11434, B1 => n11419, B2 => 
                           DataPath_RF_bus_reg_dataout_2018_port, ZN => n5862);
   U13413 : AOI22_X1 port map( A1 => n11420, A2 => n11435, B1 => n8609, B2 => 
                           DataPath_RF_bus_reg_dataout_2019_port, ZN => n5861);
   U13414 : AOI22_X1 port map( A1 => n11420, A2 => n11436, B1 => n8609, B2 => 
                           DataPath_RF_bus_reg_dataout_2020_port, ZN => n5860);
   U13415 : AOI22_X1 port map( A1 => n11420, A2 => n11437, B1 => n8609, B2 => 
                           DataPath_RF_bus_reg_dataout_2021_port, ZN => n5859);
   U13416 : AOI22_X1 port map( A1 => n11420, A2 => n11438, B1 => n8609, B2 => 
                           DataPath_RF_bus_reg_dataout_2022_port, ZN => n5858);
   U13417 : AOI22_X1 port map( A1 => n11420, A2 => n11439, B1 => n8609, B2 => 
                           DataPath_RF_bus_reg_dataout_2023_port, ZN => n5857);
   U13418 : AOI22_X1 port map( A1 => n11420, A2 => n11440, B1 => n8609, B2 => 
                           DataPath_RF_bus_reg_dataout_2024_port, ZN => n5856);
   U13419 : AOI22_X1 port map( A1 => n11420, A2 => n11441, B1 => n11419, B2 => 
                           DataPath_RF_bus_reg_dataout_2025_port, ZN => n5855);
   U13420 : NAND2_X1 port map( A1 => n8692, A2 => n11751, ZN => n3347);
   U13421 : OAI22_X1 port map( A1 => n11419, A2 => n11488, B1 => 
                           DataPath_RF_bus_reg_dataout_2026_port, B2 => n11418,
                           ZN => n5854);
   U13422 : AOI22_X1 port map( A1 => n11420, A2 => n11442, B1 => n11419, B2 => 
                           DataPath_RF_bus_reg_dataout_2027_port, ZN => n5853);
   U13423 : NAND2_X1 port map( A1 => n8692, A2 => n11752, ZN => n3345);
   U13424 : OAI22_X1 port map( A1 => n8609, A2 => n11490, B1 => 
                           DataPath_RF_bus_reg_dataout_2028_port, B2 => n11418,
                           ZN => n5852);
   U13425 : AOI22_X1 port map( A1 => n11420, A2 => n11443, B1 => n8609, B2 => 
                           DataPath_RF_bus_reg_dataout_2029_port, ZN => n5851);
   U13426 : AOI22_X1 port map( A1 => n11420, A2 => n11444, B1 => n8609, B2 => 
                           DataPath_RF_bus_reg_dataout_2030_port, ZN => n5850);
   U13427 : NAND2_X1 port map( A1 => n8692, A2 => n11631, ZN => n3342);
   U13428 : OAI22_X1 port map( A1 => n8609, A2 => n7807, B1 => 
                           DataPath_RF_bus_reg_dataout_2031_port, B2 => n11418,
                           ZN => n5849);
   U13429 : OAI22_X1 port map( A1 => n8609, A2 => n11494, B1 => 
                           DataPath_RF_bus_reg_dataout_2032_port, B2 => n11418,
                           ZN => n5848);
   U13430 : NAND2_X1 port map( A1 => n8692, A2 => n11633, ZN => n3340);
   U13431 : OAI22_X1 port map( A1 => n11419, A2 => n11495, B1 => 
                           DataPath_RF_bus_reg_dataout_2033_port, B2 => n11418,
                           ZN => n5847);
   U13432 : AOI22_X1 port map( A1 => n11420, A2 => n11445, B1 => n8609, B2 => 
                           DataPath_RF_bus_reg_dataout_2034_port, ZN => n5846);
   U13433 : NAND2_X1 port map( A1 => n8692, A2 => n11756, ZN => n3338);
   U13434 : OAI22_X1 port map( A1 => n11419, A2 => n11497, B1 => 
                           DataPath_RF_bus_reg_dataout_2035_port, B2 => n11418,
                           ZN => n5845);
   U13435 : NAND2_X1 port map( A1 => n8693, A2 => n11757, ZN => n3337);
   U13436 : OAI22_X1 port map( A1 => n8609, A2 => n11498, B1 => 
                           DataPath_RF_bus_reg_dataout_2036_port, B2 => n11418,
                           ZN => n5844);
   U13437 : NAND2_X1 port map( A1 => n8692, A2 => n11758, ZN => n3336);
   U13438 : OAI22_X1 port map( A1 => n8609, A2 => n11499, B1 => 
                           DataPath_RF_bus_reg_dataout_2037_port, B2 => n11418,
                           ZN => n5843);
   U13439 : NAND2_X1 port map( A1 => n8692, A2 => n11759, ZN => n3335);
   U13440 : OAI22_X1 port map( A1 => n8609, A2 => n11500, B1 => 
                           DataPath_RF_bus_reg_dataout_2038_port, B2 => n11418,
                           ZN => n5842);
   U13441 : AOI22_X1 port map( A1 => n11420, A2 => n11446, B1 => n8609, B2 => 
                           DataPath_RF_bus_reg_dataout_2039_port, ZN => n5841);
   U13442 : AOI22_X1 port map( A1 => n11420, A2 => n11447, B1 => n8609, B2 => 
                           DataPath_RF_bus_reg_dataout_2040_port, ZN => n5840);
   U13443 : NAND2_X1 port map( A1 => n8693, A2 => n11760, ZN => n3332);
   U13444 : OAI22_X1 port map( A1 => n11419, A2 => n11503, B1 => 
                           DataPath_RF_bus_reg_dataout_2041_port, B2 => n11418,
                           ZN => n5839);
   U13445 : AOI22_X1 port map( A1 => n11420, A2 => n11448, B1 => n11419, B2 => 
                           DataPath_RF_bus_reg_dataout_2042_port, ZN => n5838);
   U13446 : NAND2_X1 port map( A1 => n8693, A2 => n11761, ZN => n3330);
   U13447 : OAI22_X1 port map( A1 => n8609, A2 => n11505, B1 => 
                           DataPath_RF_bus_reg_dataout_2043_port, B2 => n11418,
                           ZN => n5837);
   U13448 : AOI22_X1 port map( A1 => n11420, A2 => n11421, B1 => n11419, B2 => 
                           DataPath_RF_bus_reg_dataout_2044_port, ZN => n5836);
   U13449 : NAND2_X1 port map( A1 => n8692, A2 => n11762, ZN => n3328);
   U13450 : OAI22_X1 port map( A1 => n8609, A2 => n11507, B1 => 
                           DataPath_RF_bus_reg_dataout_2045_port, B2 => n11418,
                           ZN => n5835);
   U13451 : NAND2_X1 port map( A1 => n8693, A2 => n11763, ZN => n3327);
   U13452 : OAI22_X1 port map( A1 => n8609, A2 => n11508, B1 => 
                           DataPath_RF_bus_reg_dataout_2046_port, B2 => n11418,
                           ZN => n5834);
   U13453 : AOI22_X1 port map( A1 => n11420, A2 => n11450, B1 => n11419, B2 => 
                           DataPath_RF_bus_reg_dataout_2047_port, ZN => n5831);
   U13454 : OAI22_X1 port map( A1 => n11478, A2 => n8610, B1 => 
                           DataPath_RF_bus_reg_dataout_1984_port, B2 => n8511, 
                           ZN => n5828);
   U13455 : OAI22_X1 port map( A1 => n8610, A2 => n11479, B1 => 
                           DataPath_RF_bus_reg_dataout_1985_port, B2 => n11422,
                           ZN => n5827);
   U13456 : OAI22_X1 port map( A1 => n8610, A2 => n11480, B1 => 
                           DataPath_RF_bus_reg_dataout_1986_port, B2 => n11422,
                           ZN => n5826);
   U13457 : OAI22_X1 port map( A1 => n8610, A2 => n11481, B1 => 
                           DataPath_RF_bus_reg_dataout_1987_port, B2 => n8511, 
                           ZN => n5825);
   U13458 : OAI22_X1 port map( A1 => n11423, A2 => n11482, B1 => 
                           DataPath_RF_bus_reg_dataout_1988_port, B2 => n8511, 
                           ZN => n5824);
   U13459 : OAI22_X1 port map( A1 => n11423, A2 => n11483, B1 => 
                           DataPath_RF_bus_reg_dataout_1989_port, B2 => n11422,
                           ZN => n5823);
   U13460 : OAI22_X1 port map( A1 => n8610, A2 => n11484, B1 => 
                           DataPath_RF_bus_reg_dataout_1990_port, B2 => n11422,
                           ZN => n5822);
   U13461 : OAI22_X1 port map( A1 => n8610, A2 => n11485, B1 => 
                           DataPath_RF_bus_reg_dataout_1991_port, B2 => n8511, 
                           ZN => n5821);
   U13462 : OAI22_X1 port map( A1 => n8610, A2 => n11486, B1 => 
                           DataPath_RF_bus_reg_dataout_1992_port, B2 => n8511, 
                           ZN => n5820);
   U13463 : OAI22_X1 port map( A1 => n11423, A2 => n11487, B1 => 
                           DataPath_RF_bus_reg_dataout_1993_port, B2 => n11422,
                           ZN => n5819);
   U13464 : AOI22_X1 port map( A1 => n11488, A2 => n8511, B1 => n8610, B2 => 
                           DataPath_RF_bus_reg_dataout_1994_port, ZN => n5818);
   U13465 : OAI22_X1 port map( A1 => n8610, A2 => n11489, B1 => 
                           DataPath_RF_bus_reg_dataout_1995_port, B2 => n11422,
                           ZN => n5817);
   U13466 : AOI22_X1 port map( A1 => n11490, A2 => n11422, B1 => n11423, B2 => 
                           DataPath_RF_bus_reg_dataout_1996_port, ZN => n5816);
   U13467 : OAI22_X1 port map( A1 => n8610, A2 => n11491, B1 => 
                           DataPath_RF_bus_reg_dataout_1997_port, B2 => n8511, 
                           ZN => n5815);
   U13468 : OAI22_X1 port map( A1 => n8610, A2 => n11492, B1 => 
                           DataPath_RF_bus_reg_dataout_1998_port, B2 => n8511, 
                           ZN => n5814);
   U13469 : OAI22_X1 port map( A1 => n7807, A2 => n8610, B1 => 
                           DataPath_RF_bus_reg_dataout_1999_port, B2 => n11422,
                           ZN => n5813);
   U13470 : OAI22_X1 port map( A1 => n11494, A2 => n8610, B1 => 
                           DataPath_RF_bus_reg_dataout_2000_port, B2 => n8511, 
                           ZN => n5812);
   U13471 : OAI22_X1 port map( A1 => n11423, A2 => n11495, B1 => 
                           DataPath_RF_bus_reg_dataout_2001_port, B2 => n8511, 
                           ZN => n5811);
   U13472 : OAI22_X1 port map( A1 => n11423, A2 => n11496, B1 => 
                           DataPath_RF_bus_reg_dataout_2002_port, B2 => n8511, 
                           ZN => n5810);
   U13473 : OAI22_X1 port map( A1 => n8610, A2 => n11497, B1 => 
                           DataPath_RF_bus_reg_dataout_2003_port, B2 => n11422,
                           ZN => n5809);
   U13474 : OAI22_X1 port map( A1 => n11498, A2 => n11423, B1 => 
                           DataPath_RF_bus_reg_dataout_2004_port, B2 => n8511, 
                           ZN => n5808);
   U13475 : OAI22_X1 port map( A1 => n8610, A2 => n11499, B1 => 
                           DataPath_RF_bus_reg_dataout_2005_port, B2 => n8511, 
                           ZN => n5807);
   U13476 : OAI22_X1 port map( A1 => n11500, A2 => n11423, B1 => 
                           DataPath_RF_bus_reg_dataout_2006_port, B2 => n8511, 
                           ZN => n5806);
   U13477 : OAI22_X1 port map( A1 => n8610, A2 => n11501, B1 => 
                           DataPath_RF_bus_reg_dataout_2007_port, B2 => n11422,
                           ZN => n5805);
   U13478 : OAI22_X1 port map( A1 => n11423, A2 => n11502, B1 => 
                           DataPath_RF_bus_reg_dataout_2008_port, B2 => n11422,
                           ZN => n5804);
   U13479 : AOI22_X1 port map( A1 => n11503, A2 => n11422, B1 => n8610, B2 => 
                           DataPath_RF_bus_reg_dataout_2009_port, ZN => n5803);
   U13480 : OAI22_X1 port map( A1 => n8610, A2 => n11504, B1 => 
                           DataPath_RF_bus_reg_dataout_2010_port, B2 => n8511, 
                           ZN => n5802);
   U13481 : OAI22_X1 port map( A1 => n8610, A2 => n11505, B1 => 
                           DataPath_RF_bus_reg_dataout_2011_port, B2 => n8511, 
                           ZN => n5801);
   U13482 : OAI22_X1 port map( A1 => n8610, A2 => n11506, B1 => 
                           DataPath_RF_bus_reg_dataout_2012_port, B2 => n8511, 
                           ZN => n5800);
   U13483 : OAI22_X1 port map( A1 => n11423, A2 => n11507, B1 => 
                           DataPath_RF_bus_reg_dataout_2013_port, B2 => n11422,
                           ZN => n5799);
   U13484 : OAI22_X1 port map( A1 => n11423, A2 => n11508, B1 => 
                           DataPath_RF_bus_reg_dataout_2014_port, B2 => n8511, 
                           ZN => n5798);
   U13485 : OAI22_X1 port map( A1 => n8610, A2 => n11510, B1 => 
                           DataPath_RF_bus_reg_dataout_2015_port, B2 => n8511, 
                           ZN => n5795);
   U13486 : NAND2_X1 port map( A1 => n11456, A2 => n11897, ZN => n12112);
   U13487 : AOI22_X1 port map( A1 => n11478, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1952_port, ZN => n5792);
   U13488 : AOI22_X1 port map( A1 => n11479, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1953_port, ZN => n5791);
   U13489 : AOI22_X1 port map( A1 => n11480, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1954_port, ZN => n5790);
   U13490 : AOI22_X1 port map( A1 => n11481, A2 => n7801, B1 => n11425, B2 => 
                           DataPath_RF_bus_reg_dataout_1955_port, ZN => n5789);
   U13491 : AOI22_X1 port map( A1 => n11482, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1956_port, ZN => n5788);
   U13492 : AOI22_X1 port map( A1 => n11483, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1957_port, ZN => n5787);
   U13493 : AOI22_X1 port map( A1 => n11484, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1958_port, ZN => n5786);
   U13494 : AOI22_X1 port map( A1 => n11485, A2 => n7801, B1 => n11425, B2 => 
                           DataPath_RF_bus_reg_dataout_1959_port, ZN => n5785);
   U13495 : AOI22_X1 port map( A1 => n11486, A2 => n7801, B1 => n11425, B2 => 
                           DataPath_RF_bus_reg_dataout_1960_port, ZN => n5784);
   U13496 : AOI22_X1 port map( A1 => n11487, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1961_port, ZN => n5783);
   U13497 : OAI22_X1 port map( A1 => n11488, A2 => n8611, B1 => 
                           DataPath_RF_bus_reg_dataout_1962_port, B2 => n7801, 
                           ZN => n5782);
   U13498 : AOI22_X1 port map( A1 => n11489, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1963_port, ZN => n5781);
   U13499 : OAI22_X1 port map( A1 => n11490, A2 => n8611, B1 => 
                           DataPath_RF_bus_reg_dataout_1964_port, B2 => n7801, 
                           ZN => n5780);
   U13500 : AOI22_X1 port map( A1 => n11491, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1965_port, ZN => n5779);
   U13501 : AOI22_X1 port map( A1 => n11492, A2 => n7801, B1 => n11425, B2 => 
                           DataPath_RF_bus_reg_dataout_1966_port, ZN => n5778);
   U13502 : AOI22_X1 port map( A1 => n7807, A2 => n7801, B1 => n11425, B2 => 
                           DataPath_RF_bus_reg_dataout_1967_port, ZN => n5777);
   U13503 : AOI22_X1 port map( A1 => n11494, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1968_port, ZN => n5776);
   U13504 : INV_X1 port map( A => n11425, ZN => n11424);
   U13505 : AOI22_X1 port map( A1 => n8611, A2 => 
                           DataPath_RF_bus_reg_dataout_1969_port, B1 => n11495,
                           B2 => n11424, ZN => n5775);
   U13506 : AOI22_X1 port map( A1 => n11496, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1970_port, ZN => n5774);
   U13507 : AOI22_X1 port map( A1 => n8611, A2 => 
                           DataPath_RF_bus_reg_dataout_1971_port, B1 => n11497,
                           B2 => n11424, ZN => n5773);
   U13508 : AOI22_X1 port map( A1 => n11498, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1972_port, ZN => n5772);
   U13509 : AOI22_X1 port map( A1 => n8611, A2 => 
                           DataPath_RF_bus_reg_dataout_1973_port, B1 => n11499,
                           B2 => n11424, ZN => n5771);
   U13510 : AOI22_X1 port map( A1 => n11500, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1974_port, ZN => n5770);
   U13511 : AOI22_X1 port map( A1 => n11501, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1975_port, ZN => n5769);
   U13512 : AOI22_X1 port map( A1 => n11502, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1976_port, ZN => n5768);
   U13513 : OAI22_X1 port map( A1 => n11503, A2 => n11425, B1 => 
                           DataPath_RF_bus_reg_dataout_1977_port, B2 => n7801, 
                           ZN => n5767);
   U13514 : AOI22_X1 port map( A1 => n11504, A2 => n7801, B1 => n11425, B2 => 
                           DataPath_RF_bus_reg_dataout_1978_port, ZN => n5766);
   U13515 : AOI22_X1 port map( A1 => n11425, A2 => 
                           DataPath_RF_bus_reg_dataout_1979_port, B1 => n11505,
                           B2 => n11424, ZN => n5765);
   U13516 : AOI22_X1 port map( A1 => n11506, A2 => n7801, B1 => n11425, B2 => 
                           DataPath_RF_bus_reg_dataout_1980_port, ZN => n5764);
   U13517 : AOI22_X1 port map( A1 => n11425, A2 => 
                           DataPath_RF_bus_reg_dataout_1981_port, B1 => n11507,
                           B2 => n11424, ZN => n5763);
   U13518 : AOI22_X1 port map( A1 => n8611, A2 => 
                           DataPath_RF_bus_reg_dataout_1982_port, B1 => n11508,
                           B2 => n11424, ZN => n5762);
   U13519 : AOI22_X1 port map( A1 => n11510, A2 => n7801, B1 => n8611, B2 => 
                           DataPath_RF_bus_reg_dataout_1983_port, ZN => n5759);
   U13520 : NAND2_X1 port map( A1 => n11456, A2 => n11901, ZN => n12115);
   U13521 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1920_port, B1 => n11478,
                           B2 => n11428, ZN => n5756);
   U13522 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1921_port, B1 => n11479,
                           B2 => n11428, ZN => n5755);
   U13523 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1922_port, B1 => n11480,
                           B2 => n11428, ZN => n5754);
   U13524 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1923_port, B1 => n11481,
                           B2 => n11428, ZN => n5753);
   U13525 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1924_port, B1 => n11482,
                           B2 => n11428, ZN => n5752);
   U13526 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1925_port, B1 => n11483,
                           B2 => n11428, ZN => n5751);
   U13527 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1926_port, B1 => n11484,
                           B2 => n11428, ZN => n5750);
   U13528 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1927_port, B1 => n11485,
                           B2 => n11428, ZN => n5749);
   U13529 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1928_port, B1 => n11486,
                           B2 => n11428, ZN => n5748);
   U13530 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1929_port, B1 => n11487,
                           B2 => n11428, ZN => n5747);
   U13531 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1930_port, B1 => n11488,
                           B2 => n11428, ZN => n5746);
   U13532 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1931_port, B1 => n11489,
                           B2 => n11428, ZN => n5745);
   U13533 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1932_port, B1 => n11490,
                           B2 => n11428, ZN => n5744);
   U13534 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1933_port, B1 => n11491,
                           B2 => n11428, ZN => n5743);
   U13535 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1934_port, B1 => n11492,
                           B2 => n11428, ZN => n5742);
   U13536 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1935_port, B1 => n7807, 
                           B2 => n11428, ZN => n5741);
   U13537 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1936_port, B1 => n11494,
                           B2 => n11428, ZN => n5740);
   U13538 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1937_port, B1 => n11495,
                           B2 => n11428, ZN => n5739);
   U13539 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1938_port, B1 => n11496,
                           B2 => n11428, ZN => n5738);
   U13540 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1939_port, B1 => n11497,
                           B2 => n11428, ZN => n5737);
   U13541 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1940_port, B1 => n11498,
                           B2 => n11428, ZN => n5736);
   U13542 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1941_port, B1 => n11499,
                           B2 => n11428, ZN => n5735);
   U13543 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1942_port, B1 => n11500,
                           B2 => n11428, ZN => n5734);
   U13544 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1943_port, B1 => n11501,
                           B2 => n11428, ZN => n5733);
   U13545 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1944_port, B1 => n11502,
                           B2 => n11428, ZN => n5732);
   U13546 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1945_port, B1 => n11503,
                           B2 => n11428, ZN => n5731);
   U13547 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1946_port, B1 => n11504,
                           B2 => n11428, ZN => n5730);
   U13548 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1947_port, B1 => n11505,
                           B2 => n11428, ZN => n5729);
   U13549 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1948_port, B1 => n11506,
                           B2 => n11428, ZN => n5728);
   U13550 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1949_port, B1 => n11507,
                           B2 => n11428, ZN => n5727);
   U13551 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1950_port, B1 => n11508,
                           B2 => n11428, ZN => n5726);
   U13552 : AOI22_X1 port map( A1 => n8612, A2 => 
                           DataPath_RF_bus_reg_dataout_1951_port, B1 => n11510,
                           B2 => n11428, ZN => n5723);
   U13553 : NAND2_X1 port map( A1 => n11456, A2 => n11905, ZN => n12118);
   U13554 : OAI22_X1 port map( A1 => n11478, A2 => n11431, B1 => 
                           DataPath_RF_bus_reg_dataout_1888_port, B2 => n11430,
                           ZN => n5720);
   U13555 : OAI22_X1 port map( A1 => n11479, A2 => n8613, B1 => 
                           DataPath_RF_bus_reg_dataout_1889_port, B2 => n11430,
                           ZN => n5719);
   U13556 : OAI22_X1 port map( A1 => n11480, A2 => n8613, B1 => 
                           DataPath_RF_bus_reg_dataout_1890_port, B2 => n8512, 
                           ZN => n5718);
   U13557 : OAI22_X1 port map( A1 => n11481, A2 => n8613, B1 => 
                           DataPath_RF_bus_reg_dataout_1891_port, B2 => n8512, 
                           ZN => n5717);
   U13558 : AOI22_X1 port map( A1 => n11482, A2 => n11430, B1 => n11431, B2 => 
                           DataPath_RF_bus_reg_dataout_1892_port, ZN => n5716);
   U13559 : OAI22_X1 port map( A1 => n11483, A2 => n11431, B1 => 
                           DataPath_RF_bus_reg_dataout_1893_port, B2 => n11430,
                           ZN => n5715);
   U13560 : AOI22_X1 port map( A1 => n11484, A2 => n8512, B1 => n8613, B2 => 
                           DataPath_RF_bus_reg_dataout_1894_port, ZN => n5714);
   U13561 : OAI22_X1 port map( A1 => n11485, A2 => n8613, B1 => 
                           DataPath_RF_bus_reg_dataout_1895_port, B2 => n11430,
                           ZN => n5713);
   U13562 : AOI22_X1 port map( A1 => n11486, A2 => n8512, B1 => n8613, B2 => 
                           DataPath_RF_bus_reg_dataout_1896_port, ZN => n5712);
   U13563 : OAI22_X1 port map( A1 => n11487, A2 => n8613, B1 => 
                           DataPath_RF_bus_reg_dataout_1897_port, B2 => n8512, 
                           ZN => n5711);
   U13564 : AOI22_X1 port map( A1 => n11488, A2 => n11430, B1 => n8613, B2 => 
                           DataPath_RF_bus_reg_dataout_1898_port, ZN => n5710);
   U13565 : OAI22_X1 port map( A1 => n11489, A2 => n8613, B1 => 
                           DataPath_RF_bus_reg_dataout_1899_port, B2 => n8512, 
                           ZN => n5709);
   U13566 : AOI22_X1 port map( A1 => n11490, A2 => n11430, B1 => n11431, B2 => 
                           DataPath_RF_bus_reg_dataout_1900_port, ZN => n5708);
   U13567 : AOI22_X1 port map( A1 => n11491, A2 => n8512, B1 => n8613, B2 => 
                           DataPath_RF_bus_reg_dataout_1901_port, ZN => n5707);
   U13568 : OAI22_X1 port map( A1 => n11492, A2 => n11431, B1 => 
                           DataPath_RF_bus_reg_dataout_1902_port, B2 => n11430,
                           ZN => n5706);
   U13569 : OAI22_X1 port map( A1 => n7807, A2 => n11431, B1 => 
                           DataPath_RF_bus_reg_dataout_1903_port, B2 => n8512, 
                           ZN => n5705);
   U13570 : AOI22_X1 port map( A1 => n11494, A2 => n8512, B1 => n8613, B2 => 
                           DataPath_RF_bus_reg_dataout_1904_port, ZN => n5704);
   U13571 : OAI22_X1 port map( A1 => n8613, A2 => n11495, B1 => 
                           DataPath_RF_bus_reg_dataout_1905_port, B2 => n8512, 
                           ZN => n5703);
   U13572 : OAI22_X1 port map( A1 => n11496, A2 => n8613, B1 => 
                           DataPath_RF_bus_reg_dataout_1906_port, B2 => n8512, 
                           ZN => n5702);
   U13573 : OAI22_X1 port map( A1 => n8613, A2 => n11497, B1 => 
                           DataPath_RF_bus_reg_dataout_1907_port, B2 => n8512, 
                           ZN => n5701);
   U13574 : OAI22_X1 port map( A1 => n11498, A2 => n8613, B1 => 
                           DataPath_RF_bus_reg_dataout_1908_port, B2 => n8512, 
                           ZN => n5700);
   U13575 : OAI22_X1 port map( A1 => n8613, A2 => n11499, B1 => 
                           DataPath_RF_bus_reg_dataout_1909_port, B2 => n8512, 
                           ZN => n5699);
   U13576 : OAI22_X1 port map( A1 => n11500, A2 => n8613, B1 => 
                           DataPath_RF_bus_reg_dataout_1910_port, B2 => n8512, 
                           ZN => n5698);
   U13577 : OAI22_X1 port map( A1 => n11501, A2 => n11431, B1 => 
                           DataPath_RF_bus_reg_dataout_1911_port, B2 => n11430,
                           ZN => n5697);
   U13578 : OAI22_X1 port map( A1 => n11502, A2 => n8613, B1 => 
                           DataPath_RF_bus_reg_dataout_1912_port, B2 => n11430,
                           ZN => n5696);
   U13579 : AOI22_X1 port map( A1 => n11503, A2 => n11430, B1 => n11431, B2 => 
                           DataPath_RF_bus_reg_dataout_1913_port, ZN => n5695);
   U13580 : OAI22_X1 port map( A1 => n11504, A2 => n8613, B1 => 
                           DataPath_RF_bus_reg_dataout_1914_port, B2 => n8512, 
                           ZN => n5694);
   U13581 : OAI22_X1 port map( A1 => n11431, A2 => n11505, B1 => 
                           DataPath_RF_bus_reg_dataout_1915_port, B2 => n8512, 
                           ZN => n5693);
   U13582 : OAI22_X1 port map( A1 => n11506, A2 => n8613, B1 => 
                           DataPath_RF_bus_reg_dataout_1916_port, B2 => n11430,
                           ZN => n5692);
   U13583 : OAI22_X1 port map( A1 => n11431, A2 => n11507, B1 => 
                           DataPath_RF_bus_reg_dataout_1917_port, B2 => n11430,
                           ZN => n5691);
   U13584 : OAI22_X1 port map( A1 => n8613, A2 => n11508, B1 => 
                           DataPath_RF_bus_reg_dataout_1918_port, B2 => n8512, 
                           ZN => n5690);
   U13585 : OAI22_X1 port map( A1 => n11510, A2 => n11431, B1 => 
                           DataPath_RF_bus_reg_dataout_1919_port, B2 => n8512, 
                           ZN => n5687);
   U13586 : NAND2_X1 port map( A1 => n11456, A2 => n11909, ZN => n12121);
   U13587 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1856_port, A2 
                           => n8614, B1 => n11451, B2 => n11432, ZN => n5684);
   U13588 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1857_port, A2 
                           => n8614, B1 => n11451, B2 => n11433, ZN => n5683);
   U13589 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1858_port, A2 
                           => n8614, B1 => n11451, B2 => n11434, ZN => n5682);
   U13590 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1859_port, A2 
                           => n8614, B1 => n11451, B2 => n11435, ZN => n5681);
   U13591 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1860_port, A2 
                           => n11452, B1 => n11451, B2 => n11436, ZN => n5680);
   U13592 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1861_port, A2 
                           => n8614, B1 => n11451, B2 => n11437, ZN => n5679);
   U13593 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1862_port, A2 
                           => n11452, B1 => n11451, B2 => n11438, ZN => n5678);
   U13594 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1863_port, A2 
                           => n8614, B1 => n11451, B2 => n11439, ZN => n5677);
   U13595 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1864_port, A2 
                           => n8614, B1 => n11451, B2 => n11440, ZN => n5676);
   U13596 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1865_port, A2 
                           => n8614, B1 => n11451, B2 => n11441, ZN => n5675);
   U13597 : OAI22_X1 port map( A1 => n11488, A2 => n8614, B1 => 
                           DataPath_RF_bus_reg_dataout_1866_port, B2 => n11449,
                           ZN => n5674);
   U13598 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1867_port, A2 
                           => n11452, B1 => n11451, B2 => n11442, ZN => n5673);
   U13599 : OAI22_X1 port map( A1 => n11490, A2 => n11452, B1 => 
                           DataPath_RF_bus_reg_dataout_1868_port, B2 => n11449,
                           ZN => n5672);
   U13600 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1869_port, A2 
                           => n11452, B1 => n11451, B2 => n11443, ZN => n5671);
   U13601 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1870_port, A2 
                           => n8614, B1 => n11451, B2 => n11444, ZN => n5670);
   U13602 : OAI22_X1 port map( A1 => n7807, A2 => n11452, B1 => 
                           DataPath_RF_bus_reg_dataout_1871_port, B2 => n11449,
                           ZN => n5669);
   U13603 : AOI22_X1 port map( A1 => n11494, A2 => n11449, B1 => n8614, B2 => 
                           DataPath_RF_bus_reg_dataout_1872_port, ZN => n5668);
   U13604 : OAI22_X1 port map( A1 => n8614, A2 => n11495, B1 => 
                           DataPath_RF_bus_reg_dataout_1873_port, B2 => n11449,
                           ZN => n5667);
   U13605 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1874_port, A2 
                           => n11452, B1 => n11451, B2 => n11445, ZN => n5666);
   U13606 : OAI22_X1 port map( A1 => n11452, A2 => n11497, B1 => 
                           DataPath_RF_bus_reg_dataout_1875_port, B2 => n11449,
                           ZN => n5665);
   U13607 : AOI22_X1 port map( A1 => n11498, A2 => n11449, B1 => n8614, B2 => 
                           DataPath_RF_bus_reg_dataout_1876_port, ZN => n5664);
   U13608 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1877_port, A2 
                           => n8614, B1 => n11499, B2 => n11449, ZN => n5663);
   U13609 : AOI22_X1 port map( A1 => n11500, A2 => n11449, B1 => n8614, B2 => 
                           DataPath_RF_bus_reg_dataout_1878_port, ZN => n5662);
   U13610 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1879_port, A2 
                           => n8614, B1 => n11451, B2 => n11446, ZN => n5661);
   U13611 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1880_port, A2 
                           => n8614, B1 => n11451, B2 => n11447, ZN => n5660);
   U13612 : AOI22_X1 port map( A1 => n11503, A2 => n11449, B1 => n11452, B2 => 
                           DataPath_RF_bus_reg_dataout_1881_port, ZN => n5659);
   U13613 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1882_port, A2 
                           => n8614, B1 => n11451, B2 => n11448, ZN => n5658);
   U13614 : OAI22_X1 port map( A1 => n8614, A2 => n11505, B1 => 
                           DataPath_RF_bus_reg_dataout_1883_port, B2 => n11449,
                           ZN => n5657);
   U13615 : AOI22_X1 port map( A1 => n11506, A2 => n11449, B1 => n11452, B2 => 
                           DataPath_RF_bus_reg_dataout_1884_port, ZN => n5656);
   U13616 : OAI22_X1 port map( A1 => n11452, A2 => n11507, B1 => 
                           DataPath_RF_bus_reg_dataout_1885_port, B2 => n11449,
                           ZN => n5655);
   U13617 : OAI22_X1 port map( A1 => n8614, A2 => n11508, B1 => 
                           DataPath_RF_bus_reg_dataout_1886_port, B2 => n11449,
                           ZN => n5654);
   U13618 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1887_port, A2 
                           => n8614, B1 => n11451, B2 => n11450, ZN => n5651);
   U13619 : NAND2_X1 port map( A1 => n11456, A2 => n11914, ZN => n12155);
   U13620 : OAI22_X1 port map( A1 => n11478, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1824_port, B2 => n8513, 
                           ZN => n5648);
   U13621 : OAI22_X1 port map( A1 => n11479, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1825_port, B2 => n11453,
                           ZN => n5647);
   U13622 : OAI22_X1 port map( A1 => n11480, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1826_port, B2 => n11453,
                           ZN => n5646);
   U13623 : OAI22_X1 port map( A1 => n11481, A2 => n11454, B1 => 
                           DataPath_RF_bus_reg_dataout_1827_port, B2 => n8513, 
                           ZN => n5645);
   U13624 : OAI22_X1 port map( A1 => n11482, A2 => n11454, B1 => 
                           DataPath_RF_bus_reg_dataout_1828_port, B2 => n8513, 
                           ZN => n5644);
   U13625 : OAI22_X1 port map( A1 => n11483, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1829_port, B2 => n11453,
                           ZN => n5643);
   U13626 : OAI22_X1 port map( A1 => n11484, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1830_port, B2 => n11453,
                           ZN => n5642);
   U13627 : OAI22_X1 port map( A1 => n11485, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1831_port, B2 => n8513, 
                           ZN => n5641);
   U13628 : OAI22_X1 port map( A1 => n11486, A2 => n11454, B1 => 
                           DataPath_RF_bus_reg_dataout_1832_port, B2 => n8513, 
                           ZN => n5640);
   U13629 : OAI22_X1 port map( A1 => n11487, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1833_port, B2 => n11453,
                           ZN => n5639);
   U13630 : AOI22_X1 port map( A1 => n11488, A2 => n11453, B1 => n11454, B2 => 
                           DataPath_RF_bus_reg_dataout_1834_port, ZN => n5638);
   U13631 : OAI22_X1 port map( A1 => n11489, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1835_port, B2 => n11453,
                           ZN => n5637);
   U13632 : AOI22_X1 port map( A1 => n11490, A2 => n8513, B1 => n8615, B2 => 
                           DataPath_RF_bus_reg_dataout_1836_port, ZN => n5636);
   U13633 : OAI22_X1 port map( A1 => n11491, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1837_port, B2 => n8513, 
                           ZN => n5635);
   U13634 : OAI22_X1 port map( A1 => n11492, A2 => n11454, B1 => 
                           DataPath_RF_bus_reg_dataout_1838_port, B2 => n8513, 
                           ZN => n5634);
   U13635 : OAI22_X1 port map( A1 => n7807, A2 => n11454, B1 => 
                           DataPath_RF_bus_reg_dataout_1839_port, B2 => n11453,
                           ZN => n5633);
   U13636 : OAI22_X1 port map( A1 => n11494, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1840_port, B2 => n8513, 
                           ZN => n5632);
   U13637 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1841_port, A2 
                           => n8615, B1 => n11495, B2 => n8513, ZN => n5631);
   U13638 : AOI22_X1 port map( A1 => n11496, A2 => n8513, B1 => n8615, B2 => 
                           DataPath_RF_bus_reg_dataout_1842_port, ZN => n5630);
   U13639 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1843_port, A2 
                           => n11454, B1 => n11497, B2 => n8513, ZN => n5629);
   U13640 : OAI22_X1 port map( A1 => n11498, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1844_port, B2 => n8513, 
                           ZN => n5628);
   U13641 : OAI22_X1 port map( A1 => n11454, A2 => n11499, B1 => 
                           DataPath_RF_bus_reg_dataout_1845_port, B2 => n8513, 
                           ZN => n5627);
   U13642 : OAI22_X1 port map( A1 => n11500, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1846_port, B2 => n11453,
                           ZN => n5626);
   U13643 : OAI22_X1 port map( A1 => n11501, A2 => n11454, B1 => 
                           DataPath_RF_bus_reg_dataout_1847_port, B2 => n11453,
                           ZN => n5625);
   U13644 : OAI22_X1 port map( A1 => n11502, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1848_port, B2 => n8513, 
                           ZN => n5624);
   U13645 : AOI22_X1 port map( A1 => n11503, A2 => n11453, B1 => n11454, B2 => 
                           DataPath_RF_bus_reg_dataout_1849_port, ZN => n5623);
   U13646 : OAI22_X1 port map( A1 => n11504, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1850_port, B2 => n8513, 
                           ZN => n5622);
   U13647 : OAI22_X1 port map( A1 => n8615, A2 => n11505, B1 => 
                           DataPath_RF_bus_reg_dataout_1851_port, B2 => n11453,
                           ZN => n5621);
   U13648 : OAI22_X1 port map( A1 => n11506, A2 => n8615, B1 => 
                           DataPath_RF_bus_reg_dataout_1852_port, B2 => n11453,
                           ZN => n5620);
   U13649 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1853_port, A2 
                           => n8615, B1 => n11507, B2 => n8513, ZN => n5619);
   U13650 : OAI22_X1 port map( A1 => n8615, A2 => n11508, B1 => 
                           DataPath_RF_bus_reg_dataout_1854_port, B2 => n8513, 
                           ZN => n5618);
   U13651 : OAI22_X1 port map( A1 => n11510, A2 => n11454, B1 => 
                           DataPath_RF_bus_reg_dataout_1855_port, B2 => n8513, 
                           ZN => n5615);
   U13652 : NAND2_X1 port map( A1 => n11456, A2 => n11455, ZN => n12158);
   U13653 : OAI22_X1 port map( A1 => n11478, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1792_port, B2 => n11458,
                           ZN => n5609);
   U13654 : OAI22_X1 port map( A1 => n11479, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1793_port, B2 => n11458,
                           ZN => n5608);
   U13655 : OAI22_X1 port map( A1 => n11480, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1794_port, B2 => n8514, 
                           ZN => n5607);
   U13656 : OAI22_X1 port map( A1 => n11481, A2 => n11457, B1 => 
                           DataPath_RF_bus_reg_dataout_1795_port, B2 => n8514, 
                           ZN => n5606);
   U13657 : OAI22_X1 port map( A1 => n11482, A2 => n11457, B1 => 
                           DataPath_RF_bus_reg_dataout_1796_port, B2 => n11458,
                           ZN => n5605);
   U13658 : OAI22_X1 port map( A1 => n11483, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1797_port, B2 => n11458,
                           ZN => n5604);
   U13659 : OAI22_X1 port map( A1 => n11484, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1798_port, B2 => n8514, 
                           ZN => n5603);
   U13660 : OAI22_X1 port map( A1 => n11485, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1799_port, B2 => n8514, 
                           ZN => n5602);
   U13661 : OAI22_X1 port map( A1 => n11486, A2 => n11457, B1 => 
                           DataPath_RF_bus_reg_dataout_1800_port, B2 => n11458,
                           ZN => n5601);
   U13662 : OAI22_X1 port map( A1 => n11487, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1801_port, B2 => n11458,
                           ZN => n5600);
   U13663 : AOI22_X1 port map( A1 => n11488, A2 => n11458, B1 => n8616, B2 => 
                           DataPath_RF_bus_reg_dataout_1802_port, ZN => n5599);
   U13664 : OAI22_X1 port map( A1 => n11489, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1803_port, B2 => n8514, 
                           ZN => n5598);
   U13665 : AOI22_X1 port map( A1 => n11490, A2 => n8514, B1 => n11457, B2 => 
                           DataPath_RF_bus_reg_dataout_1804_port, ZN => n5597);
   U13666 : OAI22_X1 port map( A1 => n11491, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1805_port, B2 => n8514, 
                           ZN => n5596);
   U13667 : OAI22_X1 port map( A1 => n11492, A2 => n11457, B1 => 
                           DataPath_RF_bus_reg_dataout_1806_port, B2 => n11458,
                           ZN => n5595);
   U13668 : OAI22_X1 port map( A1 => n7807, A2 => n11457, B1 => 
                           DataPath_RF_bus_reg_dataout_1807_port, B2 => n8514, 
                           ZN => n5594);
   U13669 : OAI22_X1 port map( A1 => n11494, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1808_port, B2 => n8514, 
                           ZN => n5593);
   U13670 : OAI22_X1 port map( A1 => n8616, A2 => n11495, B1 => 
                           DataPath_RF_bus_reg_dataout_1809_port, B2 => n8514, 
                           ZN => n5592);
   U13671 : OAI22_X1 port map( A1 => n11496, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1810_port, B2 => n11458,
                           ZN => n5591);
   U13672 : OAI22_X1 port map( A1 => n8616, A2 => n11497, B1 => 
                           DataPath_RF_bus_reg_dataout_1811_port, B2 => n8514, 
                           ZN => n5590);
   U13673 : OAI22_X1 port map( A1 => n11498, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1812_port, B2 => n8514, 
                           ZN => n5589);
   U13674 : OAI22_X1 port map( A1 => n8616, A2 => n11499, B1 => 
                           DataPath_RF_bus_reg_dataout_1813_port, B2 => n8514, 
                           ZN => n5588);
   U13675 : OAI22_X1 port map( A1 => n11500, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1814_port, B2 => n8514, 
                           ZN => n5587);
   U13676 : OAI22_X1 port map( A1 => n11501, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1815_port, B2 => n11458,
                           ZN => n5586);
   U13677 : OAI22_X1 port map( A1 => n11502, A2 => n11457, B1 => 
                           DataPath_RF_bus_reg_dataout_1816_port, B2 => n8514, 
                           ZN => n5585);
   U13678 : AOI22_X1 port map( A1 => n11503, A2 => n8514, B1 => n8616, B2 => 
                           DataPath_RF_bus_reg_dataout_1817_port, ZN => n5584);
   U13679 : OAI22_X1 port map( A1 => n11504, A2 => n8616, B1 => 
                           DataPath_RF_bus_reg_dataout_1818_port, B2 => n8514, 
                           ZN => n5583);
   U13680 : OAI22_X1 port map( A1 => n11457, A2 => n11505, B1 => 
                           DataPath_RF_bus_reg_dataout_1819_port, B2 => n11458,
                           ZN => n5582);
   U13681 : OAI22_X1 port map( A1 => n11506, A2 => n11457, B1 => 
                           DataPath_RF_bus_reg_dataout_1820_port, B2 => n11458,
                           ZN => n5581);
   U13682 : OAI22_X1 port map( A1 => n11457, A2 => n11507, B1 => 
                           DataPath_RF_bus_reg_dataout_1821_port, B2 => n8514, 
                           ZN => n5580);
   U13683 : OAI22_X1 port map( A1 => n8616, A2 => n11508, B1 => 
                           DataPath_RF_bus_reg_dataout_1822_port, B2 => n8514, 
                           ZN => n5579);
   U13684 : AOI22_X1 port map( A1 => n11510, A2 => n11458, B1 => n11457, B2 => 
                           DataPath_RF_bus_reg_dataout_1823_port, ZN => n5576);
   U13685 : OAI22_X1 port map( A1 => n577, A2 => n11823, B1 => n11824, B2 => 
                           n11596, ZN => n11459);
   U13686 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1760_port, B1 => n11478,
                           B2 => n11460, ZN => n5574);
   U13687 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1761_port, B1 => n11479,
                           B2 => n11460, ZN => n5573);
   U13688 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1762_port, B1 => n11480,
                           B2 => n11460, ZN => n5572);
   U13689 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1763_port, B1 => n11481,
                           B2 => n11460, ZN => n5571);
   U13690 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1764_port, B1 => n11482,
                           B2 => n11460, ZN => n5570);
   U13691 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1765_port, B1 => n11483,
                           B2 => n11460, ZN => n5569);
   U13692 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1766_port, B1 => n11484,
                           B2 => n11460, ZN => n5568);
   U13693 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1767_port, B1 => n11485,
                           B2 => n11460, ZN => n5567);
   U13694 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1768_port, B1 => n11486,
                           B2 => n11460, ZN => n5566);
   U13695 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1769_port, B1 => n11487,
                           B2 => n11460, ZN => n5565);
   U13696 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1770_port, B1 => n11488,
                           B2 => n11460, ZN => n5564);
   U13697 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1771_port, B1 => n11489,
                           B2 => n11460, ZN => n5563);
   U13698 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1772_port, B1 => n11490,
                           B2 => n11460, ZN => n5562);
   U13699 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1773_port, B1 => n11491,
                           B2 => n11460, ZN => n5561);
   U13700 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1774_port, B1 => n11492,
                           B2 => n11460, ZN => n5560);
   U13701 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1775_port, B1 => n7807, 
                           B2 => n11460, ZN => n5559);
   U13702 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1776_port, B1 => n11494,
                           B2 => n11460, ZN => n5558);
   U13703 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1777_port, B1 => n11495,
                           B2 => n11460, ZN => n5557);
   U13704 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1778_port, B1 => n11496,
                           B2 => n11460, ZN => n5556);
   U13705 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1779_port, B1 => n11497,
                           B2 => n11460, ZN => n5555);
   U13706 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1780_port, B1 => n11498,
                           B2 => n11460, ZN => n5554);
   U13707 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1781_port, B1 => n11499,
                           B2 => n11460, ZN => n5553);
   U13708 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1782_port, B1 => n11500,
                           B2 => n11460, ZN => n5552);
   U13709 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1783_port, B1 => n11501,
                           B2 => n11460, ZN => n5551);
   U13710 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1784_port, B1 => n11502,
                           B2 => n11460, ZN => n5550);
   U13711 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1785_port, B1 => n11503,
                           B2 => n11460, ZN => n5549);
   U13712 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1786_port, B1 => n11504,
                           B2 => n11460, ZN => n5548);
   U13713 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1787_port, B1 => n11505,
                           B2 => n11460, ZN => n5547);
   U13714 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1788_port, B1 => n11506,
                           B2 => n11460, ZN => n5546);
   U13715 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1789_port, B1 => n11507,
                           B2 => n11460, ZN => n5545);
   U13716 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1790_port, B1 => n11508,
                           B2 => n11460, ZN => n5544);
   U13717 : AOI22_X1 port map( A1 => n8515, A2 => 
                           DataPath_RF_bus_reg_dataout_1791_port, B1 => n11510,
                           B2 => n11460, ZN => n5541);
   U13718 : OAI22_X1 port map( A1 => n577, A2 => n11828, B1 => n11829, B2 => 
                           n11596, ZN => n11462);
   U13719 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1728_port, B1 => n11478,
                           B2 => n11463, ZN => n5539);
   U13720 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1729_port, B1 => n11479,
                           B2 => n11463, ZN => n5538);
   U13721 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1730_port, B1 => n11480,
                           B2 => n11463, ZN => n5537);
   U13722 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1731_port, B1 => n11481,
                           B2 => n11463, ZN => n5536);
   U13723 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1732_port, B1 => n11482,
                           B2 => n11463, ZN => n5535);
   U13724 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1733_port, B1 => n11483,
                           B2 => n11463, ZN => n5534);
   U13725 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1734_port, B1 => n11484,
                           B2 => n11463, ZN => n5533);
   U13726 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1735_port, B1 => n11485,
                           B2 => n11463, ZN => n5532);
   U13727 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1736_port, B1 => n11486,
                           B2 => n11463, ZN => n5531);
   U13728 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1737_port, B1 => n11487,
                           B2 => n11463, ZN => n5530);
   U13729 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1738_port, B1 => n11488,
                           B2 => n11463, ZN => n5529);
   U13730 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1739_port, B1 => n11489,
                           B2 => n11463, ZN => n5528);
   U13731 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1740_port, B1 => n11490,
                           B2 => n11463, ZN => n5527);
   U13732 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1741_port, B1 => n11491,
                           B2 => n11463, ZN => n5526);
   U13733 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1742_port, B1 => n11492,
                           B2 => n11463, ZN => n5525);
   U13734 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1743_port, B1 => n7807, 
                           B2 => n11463, ZN => n5524);
   U13735 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1744_port, B1 => n11494,
                           B2 => n11463, ZN => n5523);
   U13736 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1745_port, B1 => n11495,
                           B2 => n11463, ZN => n5522);
   U13737 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1746_port, B1 => n11496,
                           B2 => n11463, ZN => n5521);
   U13738 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1747_port, B1 => n11497,
                           B2 => n11463, ZN => n5520);
   U13739 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1748_port, B1 => n11498,
                           B2 => n11463, ZN => n5519);
   U13740 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1749_port, B1 => n11499,
                           B2 => n11463, ZN => n5518);
   U13741 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1750_port, B1 => n11500,
                           B2 => n11463, ZN => n5517);
   U13742 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1751_port, B1 => n11501,
                           B2 => n11463, ZN => n5516);
   U13743 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1752_port, B1 => n11502,
                           B2 => n11463, ZN => n5515);
   U13744 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1753_port, B1 => n11503,
                           B2 => n11463, ZN => n5514);
   U13745 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1754_port, B1 => n11504,
                           B2 => n11463, ZN => n5513);
   U13746 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1755_port, B1 => n11505,
                           B2 => n11463, ZN => n5512);
   U13747 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1756_port, B1 => n11506,
                           B2 => n11463, ZN => n5511);
   U13748 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1757_port, B1 => n11507,
                           B2 => n11463, ZN => n5510);
   U13749 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1758_port, B1 => n11508,
                           B2 => n11463, ZN => n5509);
   U13750 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_1759_port, B1 => n11510,
                           B2 => n11463, ZN => n5506);
   U13751 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1696_port, B1 => n11478,
                           B2 => n11466, ZN => n5504);
   U13752 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1697_port, B1 => n11479,
                           B2 => n11466, ZN => n5503);
   U13753 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1698_port, B1 => n11480,
                           B2 => n11466, ZN => n5502);
   U13754 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1699_port, B1 => n11481,
                           B2 => n11466, ZN => n5501);
   U13755 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1700_port, B1 => n11482,
                           B2 => n11466, ZN => n5500);
   U13756 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1701_port, B1 => n11483,
                           B2 => n11466, ZN => n5499);
   U13757 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1702_port, B1 => n11484,
                           B2 => n11466, ZN => n5498);
   U13758 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1703_port, B1 => n11485,
                           B2 => n11466, ZN => n5497);
   U13759 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1704_port, B1 => n11486,
                           B2 => n11466, ZN => n5496);
   U13760 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1705_port, B1 => n11487,
                           B2 => n11466, ZN => n5495);
   U13761 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1706_port, B1 => n11488,
                           B2 => n11466, ZN => n5494);
   U13762 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1707_port, B1 => n11489,
                           B2 => n11466, ZN => n5493);
   U13763 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1708_port, B1 => n11490,
                           B2 => n11466, ZN => n5492);
   U13764 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1709_port, B1 => n11491,
                           B2 => n11466, ZN => n5491);
   U13765 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1710_port, B1 => n11492,
                           B2 => n11466, ZN => n5490);
   U13766 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1711_port, B1 => n7807, 
                           B2 => n11466, ZN => n5489);
   U13767 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1712_port, B1 => n11494,
                           B2 => n11466, ZN => n5488);
   U13768 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1713_port, B1 => n11495,
                           B2 => n11466, ZN => n5487);
   U13769 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1714_port, B1 => n11496,
                           B2 => n11466, ZN => n5486);
   U13770 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1715_port, B1 => n11497,
                           B2 => n11466, ZN => n5485);
   U13771 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1716_port, B1 => n11498,
                           B2 => n11466, ZN => n5484);
   U13772 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1717_port, B1 => n11499,
                           B2 => n11466, ZN => n5483);
   U13773 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1718_port, B1 => n11500,
                           B2 => n11466, ZN => n5482);
   U13774 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1719_port, B1 => n11501,
                           B2 => n11466, ZN => n5481);
   U13775 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1720_port, B1 => n11502,
                           B2 => n11466, ZN => n5480);
   U13776 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1721_port, B1 => n11503,
                           B2 => n11466, ZN => n5479);
   U13777 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1722_port, B1 => n11504,
                           B2 => n11466, ZN => n5478);
   U13778 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1723_port, B1 => n11505,
                           B2 => n11466, ZN => n5477);
   U13779 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1724_port, B1 => n11506,
                           B2 => n11466, ZN => n5476);
   U13780 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1725_port, B1 => n11507,
                           B2 => n11466, ZN => n5475);
   U13781 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1726_port, B1 => n11508,
                           B2 => n11466, ZN => n5474);
   U13782 : AOI22_X1 port map( A1 => n11467, A2 => 
                           DataPath_RF_bus_reg_dataout_1727_port, B1 => n11510,
                           B2 => n11466, ZN => n5471);
   U13783 : OAI22_X1 port map( A1 => n577, A2 => n11838, B1 => n11839, B2 => 
                           n11596, ZN => n11468);
   U13784 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1664_port, B1 => n11478,
                           B2 => n11469, ZN => n5469);
   U13785 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1665_port, B1 => n11479,
                           B2 => n11469, ZN => n5468);
   U13786 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1666_port, B1 => n11480,
                           B2 => n11469, ZN => n5467);
   U13787 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1667_port, B1 => n11481,
                           B2 => n11469, ZN => n5466);
   U13788 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1668_port, B1 => n11482,
                           B2 => n11469, ZN => n5465);
   U13789 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1669_port, B1 => n11483,
                           B2 => n11469, ZN => n5464);
   U13790 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1670_port, B1 => n11484,
                           B2 => n11469, ZN => n5463);
   U13791 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1671_port, B1 => n11485,
                           B2 => n11469, ZN => n5462);
   U13792 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1672_port, B1 => n11486,
                           B2 => n11469, ZN => n5461);
   U13793 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1673_port, B1 => n11487,
                           B2 => n11469, ZN => n5460);
   U13794 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1674_port, B1 => n11488,
                           B2 => n11469, ZN => n5459);
   U13795 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1675_port, B1 => n11489,
                           B2 => n11469, ZN => n5458);
   U13796 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1676_port, B1 => n11490,
                           B2 => n11469, ZN => n5457);
   U13797 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1677_port, B1 => n11491,
                           B2 => n11469, ZN => n5456);
   U13798 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1678_port, B1 => n11492,
                           B2 => n11469, ZN => n5455);
   U13799 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1679_port, B1 => n7807, 
                           B2 => n11469, ZN => n5454);
   U13800 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1680_port, B1 => n11494,
                           B2 => n11469, ZN => n5453);
   U13801 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1681_port, B1 => n11495,
                           B2 => n11469, ZN => n5452);
   U13802 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1682_port, B1 => n11496,
                           B2 => n11469, ZN => n5451);
   U13803 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1683_port, B1 => n11497,
                           B2 => n11469, ZN => n5450);
   U13804 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1684_port, B1 => n11498,
                           B2 => n11469, ZN => n5449);
   U13805 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1685_port, B1 => n11499,
                           B2 => n11469, ZN => n5448);
   U13806 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1686_port, B1 => n11500,
                           B2 => n11469, ZN => n5447);
   U13807 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1687_port, B1 => n11501,
                           B2 => n11469, ZN => n5446);
   U13808 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1688_port, B1 => n11502,
                           B2 => n11469, ZN => n5445);
   U13809 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1689_port, B1 => n11503,
                           B2 => n11469, ZN => n5444);
   U13810 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1690_port, B1 => n11504,
                           B2 => n11469, ZN => n5443);
   U13811 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1691_port, B1 => n11505,
                           B2 => n11469, ZN => n5442);
   U13812 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1692_port, B1 => n11506,
                           B2 => n11469, ZN => n5441);
   U13813 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1693_port, B1 => n11507,
                           B2 => n11469, ZN => n5440);
   U13814 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1694_port, B1 => n11508,
                           B2 => n11469, ZN => n5439);
   U13815 : AOI22_X1 port map( A1 => n8517, A2 => 
                           DataPath_RF_bus_reg_dataout_1695_port, B1 => n11510,
                           B2 => n11469, ZN => n5436);
   U13816 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1632_port, B1 => n11478,
                           B2 => n11472, ZN => n5434);
   U13817 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1633_port, B1 => n11479,
                           B2 => n11472, ZN => n5433);
   U13818 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1634_port, B1 => n11480,
                           B2 => n11472, ZN => n5432);
   U13819 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1635_port, B1 => n11481,
                           B2 => n11472, ZN => n5431);
   U13820 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1636_port, B1 => n11482,
                           B2 => n11472, ZN => n5430);
   U13821 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1637_port, B1 => n11483,
                           B2 => n11472, ZN => n5429);
   U13822 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1638_port, B1 => n11484,
                           B2 => n11472, ZN => n5428);
   U13823 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1639_port, B1 => n11485,
                           B2 => n11472, ZN => n5427);
   U13824 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1640_port, B1 => n11486,
                           B2 => n11472, ZN => n5426);
   U13825 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1641_port, B1 => n11487,
                           B2 => n11472, ZN => n5425);
   U13826 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1642_port, B1 => n11488,
                           B2 => n11472, ZN => n5424);
   U13827 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1643_port, B1 => n11489,
                           B2 => n11472, ZN => n5423);
   U13828 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1644_port, B1 => n11490,
                           B2 => n11472, ZN => n5422);
   U13829 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1645_port, B1 => n11491,
                           B2 => n11472, ZN => n5421);
   U13830 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1646_port, B1 => n11492,
                           B2 => n11472, ZN => n5420);
   U13831 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1647_port, B1 => n7807, 
                           B2 => n11472, ZN => n5419);
   U13832 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1648_port, B1 => n11494,
                           B2 => n11472, ZN => n5418);
   U13833 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1649_port, B1 => n11495,
                           B2 => n11472, ZN => n5417);
   U13834 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1650_port, B1 => n11496,
                           B2 => n11472, ZN => n5416);
   U13835 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1651_port, B1 => n11497,
                           B2 => n11472, ZN => n5415);
   U13836 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1652_port, B1 => n11498,
                           B2 => n11472, ZN => n5414);
   U13837 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1653_port, B1 => n11499,
                           B2 => n11472, ZN => n5413);
   U13838 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1654_port, B1 => n11500,
                           B2 => n11472, ZN => n5412);
   U13839 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1655_port, B1 => n11501,
                           B2 => n11472, ZN => n5411);
   U13840 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1656_port, B1 => n11502,
                           B2 => n11472, ZN => n5410);
   U13841 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1657_port, B1 => n11503,
                           B2 => n11472, ZN => n5409);
   U13842 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1658_port, B1 => n11504,
                           B2 => n11472, ZN => n5408);
   U13843 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1659_port, B1 => n11505,
                           B2 => n11472, ZN => n5407);
   U13844 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1660_port, B1 => n11506,
                           B2 => n11472, ZN => n5406);
   U13845 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1661_port, B1 => n11507,
                           B2 => n11472, ZN => n5405);
   U13846 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1662_port, B1 => n11508,
                           B2 => n11472, ZN => n5404);
   U13847 : AOI22_X1 port map( A1 => n11473, A2 => 
                           DataPath_RF_bus_reg_dataout_1663_port, B1 => n11510,
                           B2 => n11472, ZN => n5401);
   U13848 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1600_port, B1 => n11478,
                           B2 => n11474, ZN => n5399);
   U13849 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1601_port, B1 => n11479,
                           B2 => n11474, ZN => n5398);
   U13850 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1602_port, B1 => n11480,
                           B2 => n11474, ZN => n5397);
   U13851 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1603_port, B1 => n11481,
                           B2 => n11474, ZN => n5396);
   U13852 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1604_port, B1 => n11482,
                           B2 => n11474, ZN => n5395);
   U13853 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1605_port, B1 => n11483,
                           B2 => n11474, ZN => n5394);
   U13854 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1606_port, B1 => n11484,
                           B2 => n11474, ZN => n5393);
   U13855 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1607_port, B1 => n11485,
                           B2 => n11474, ZN => n5392);
   U13856 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1608_port, B1 => n11486,
                           B2 => n11474, ZN => n5391);
   U13857 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1609_port, B1 => n11487,
                           B2 => n11474, ZN => n5390);
   U13858 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1610_port, B1 => n11488,
                           B2 => n11474, ZN => n5389);
   U13859 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1611_port, B1 => n11489,
                           B2 => n11474, ZN => n5388);
   U13860 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1612_port, B1 => n11490,
                           B2 => n11474, ZN => n5387);
   U13861 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1613_port, B1 => n11491,
                           B2 => n11474, ZN => n5386);
   U13862 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1614_port, B1 => n11492,
                           B2 => n11474, ZN => n5385);
   U13863 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1615_port, B1 => n7807, 
                           B2 => n11474, ZN => n5384);
   U13864 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1616_port, B1 => n11494,
                           B2 => n11474, ZN => n5383);
   U13865 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1617_port, B1 => n11495,
                           B2 => n11474, ZN => n5382);
   U13866 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1618_port, B1 => n11496,
                           B2 => n11474, ZN => n5381);
   U13867 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1619_port, B1 => n11497,
                           B2 => n11474, ZN => n5380);
   U13868 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1620_port, B1 => n11498,
                           B2 => n11474, ZN => n5379);
   U13869 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1621_port, B1 => n11499,
                           B2 => n11474, ZN => n5378);
   U13870 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1622_port, B1 => n11500,
                           B2 => n11474, ZN => n5377);
   U13871 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1623_port, B1 => n11501,
                           B2 => n11474, ZN => n5376);
   U13872 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1624_port, B1 => n11502,
                           B2 => n11474, ZN => n5375);
   U13873 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1625_port, B1 => n11503,
                           B2 => n11474, ZN => n5374);
   U13874 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1626_port, B1 => n11504,
                           B2 => n11474, ZN => n5373);
   U13875 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1627_port, B1 => n11505,
                           B2 => n11474, ZN => n5372);
   U13876 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1628_port, B1 => n11506,
                           B2 => n11474, ZN => n5371);
   U13877 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1629_port, B1 => n11507,
                           B2 => n11474, ZN => n5370);
   U13878 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1630_port, B1 => n11508,
                           B2 => n11474, ZN => n5369);
   U13879 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_1631_port, B1 => n11510,
                           B2 => n11474, ZN => n5366);
   U13880 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1568_port, B1 => n11478,
                           B2 => n11476, ZN => n5364);
   U13881 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1569_port, B1 => n11479,
                           B2 => n11476, ZN => n5363);
   U13882 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1570_port, B1 => n11480,
                           B2 => n11476, ZN => n5362);
   U13883 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1571_port, B1 => n11481,
                           B2 => n11476, ZN => n5361);
   U13884 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1572_port, B1 => n11482,
                           B2 => n11476, ZN => n5360);
   U13885 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1573_port, B1 => n11483,
                           B2 => n11476, ZN => n5359);
   U13886 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1574_port, B1 => n11484,
                           B2 => n11476, ZN => n5358);
   U13887 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1575_port, B1 => n11485,
                           B2 => n11476, ZN => n5357);
   U13888 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1576_port, B1 => n11486,
                           B2 => n11476, ZN => n5356);
   U13889 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1577_port, B1 => n11487,
                           B2 => n11476, ZN => n5355);
   U13890 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1578_port, B1 => n11488,
                           B2 => n11476, ZN => n5354);
   U13891 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1579_port, B1 => n11489,
                           B2 => n11476, ZN => n5353);
   U13892 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1580_port, B1 => n11490,
                           B2 => n11476, ZN => n5352);
   U13893 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1581_port, B1 => n11491,
                           B2 => n11476, ZN => n5351);
   U13894 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1582_port, B1 => n11492,
                           B2 => n11476, ZN => n5350);
   U13895 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1583_port, B1 => n7807, 
                           B2 => n11476, ZN => n5349);
   U13896 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1584_port, B1 => n11494,
                           B2 => n11476, ZN => n5348);
   U13897 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1585_port, B1 => n11495,
                           B2 => n11476, ZN => n5347);
   U13898 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1586_port, B1 => n11496,
                           B2 => n11476, ZN => n5346);
   U13899 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1587_port, B1 => n11497,
                           B2 => n11476, ZN => n5345);
   U13900 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1588_port, B1 => n11498,
                           B2 => n11476, ZN => n5344);
   U13901 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1589_port, B1 => n11499,
                           B2 => n11476, ZN => n5343);
   U13902 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1590_port, B1 => n11500,
                           B2 => n11476, ZN => n5342);
   U13903 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1591_port, B1 => n11501,
                           B2 => n11476, ZN => n5341);
   U13904 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1592_port, B1 => n11502,
                           B2 => n11476, ZN => n5340);
   U13905 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1593_port, B1 => n11503,
                           B2 => n11476, ZN => n5339);
   U13906 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1594_port, B1 => n11504,
                           B2 => n11476, ZN => n5338);
   U13907 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1595_port, B1 => n11505,
                           B2 => n11476, ZN => n5337);
   U13908 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1596_port, B1 => n11506,
                           B2 => n11476, ZN => n5336);
   U13909 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1597_port, B1 => n11507,
                           B2 => n11476, ZN => n5335);
   U13910 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1598_port, B1 => n11508,
                           B2 => n11476, ZN => n5334);
   U13911 : AOI22_X1 port map( A1 => n8519, A2 => 
                           DataPath_RF_bus_reg_dataout_1599_port, B1 => n11510,
                           B2 => n11476, ZN => n5331);
   U13912 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1536_port, B1 => n11478,
                           B2 => n11509, ZN => n5327);
   U13913 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1537_port, B1 => n11479,
                           B2 => n11509, ZN => n5325);
   U13914 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1538_port, B1 => n11480,
                           B2 => n11509, ZN => n5323);
   U13915 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1539_port, B1 => n11481,
                           B2 => n11509, ZN => n5321);
   U13916 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1540_port, B1 => n11482,
                           B2 => n11509, ZN => n5319);
   U13917 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1541_port, B1 => n11483,
                           B2 => n11509, ZN => n5317);
   U13918 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1542_port, B1 => n11484,
                           B2 => n11509, ZN => n5315);
   U13919 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1543_port, B1 => n11485,
                           B2 => n11509, ZN => n5313);
   U13920 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1544_port, B1 => n11486,
                           B2 => n11509, ZN => n5311);
   U13921 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1545_port, B1 => n11487,
                           B2 => n11509, ZN => n5309);
   U13922 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1546_port, B1 => n11488,
                           B2 => n11509, ZN => n5307);
   U13923 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1547_port, B1 => n11489,
                           B2 => n11509, ZN => n5305);
   U13924 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1548_port, B1 => n11490,
                           B2 => n11509, ZN => n5303);
   U13925 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1549_port, B1 => n11491,
                           B2 => n11509, ZN => n5301);
   U13926 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1550_port, B1 => n11492,
                           B2 => n11509, ZN => n5299);
   U13927 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1551_port, B1 => n7807, 
                           B2 => n11509, ZN => n5297);
   U13928 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1552_port, B1 => n11494,
                           B2 => n11509, ZN => n5295);
   U13929 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1553_port, B1 => n11495,
                           B2 => n11509, ZN => n5293);
   U13930 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1554_port, B1 => n11496,
                           B2 => n11509, ZN => n5291);
   U13931 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1555_port, B1 => n11497,
                           B2 => n11509, ZN => n5289);
   U13932 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1556_port, B1 => n11498,
                           B2 => n11509, ZN => n5287);
   U13933 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1557_port, B1 => n11499,
                           B2 => n11509, ZN => n5285);
   U13934 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1558_port, B1 => n11500,
                           B2 => n11509, ZN => n5283);
   U13935 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1559_port, B1 => n11501,
                           B2 => n11509, ZN => n5281);
   U13936 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1560_port, B1 => n11502,
                           B2 => n11509, ZN => n5279);
   U13937 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1561_port, B1 => n11503,
                           B2 => n11509, ZN => n5277);
   U13938 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1562_port, B1 => n11504,
                           B2 => n11509, ZN => n5275);
   U13939 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1563_port, B1 => n11505,
                           B2 => n11509, ZN => n5273);
   U13940 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1564_port, B1 => n11506,
                           B2 => n11509, ZN => n5271);
   U13941 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1565_port, B1 => n11507,
                           B2 => n11509, ZN => n5269);
   U13942 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1566_port, B1 => n11508,
                           B2 => n11509, ZN => n5267);
   U13943 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_1567_port, B1 => n11510,
                           B2 => n11509, ZN => n5263);
   U13944 : AOI22_X1 port map( A1 => n11597, A2 => n11512, B1 => n11513, B2 => 
                           DataPath_RF_bus_reg_dataout_1504_port, ZN => n5261);
   U13945 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1505_port, A2 
                           => n11513, B1 => n11598, B2 => n11512, ZN => n5260);
   U13946 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1506_port, A2 
                           => n8617, B1 => n11599, B2 => n8521, ZN => n5259);
   U13947 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1507_port, A2 
                           => n8617, B1 => n11600, B2 => n8521, ZN => n5258);
   U13948 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1508_port, A2 
                           => n8617, B1 => n11601, B2 => n11512, ZN => n5257);
   U13949 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1509_port, A2 
                           => n11513, B1 => n11602, B2 => n11512, ZN => n5256);
   U13950 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1510_port, A2 
                           => n8617, B1 => n11603, B2 => n8521, ZN => n5255);
   U13951 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1511_port, A2 
                           => n8617, B1 => n11604, B2 => n8521, ZN => n5254);
   U13952 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1512_port, A2 
                           => n8617, B1 => n11605, B2 => n11512, ZN => n5253);
   U13953 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1513_port, A2 
                           => n11513, B1 => n11606, B2 => n11512, ZN => n5252);
   U13954 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1514_port, A2 
                           => n11513, B1 => n11607, B2 => n8521, ZN => n5251);
   U13955 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1515_port, A2 
                           => n8617, B1 => n11608, B2 => n8521, ZN => n5250);
   U13956 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1516_port, A2 
                           => n8617, B1 => n11609, B2 => n11512, ZN => n5249);
   U13957 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1517_port, A2 
                           => n8617, B1 => n11610, B2 => n11512, ZN => n5248);
   U13958 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1518_port, A2 
                           => n8617, B1 => n11611, B2 => n8521, ZN => n5247);
   U13959 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1519_port, A2 
                           => n8617, B1 => n11612, B2 => n8521, ZN => n5246);
   U13960 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1520_port, A2 
                           => n8617, B1 => n11613, B2 => n11512, ZN => n5245);
   U13961 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1521_port, A2 
                           => n8617, B1 => n11614, B2 => n8521, ZN => n5244);
   U13962 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1522_port, A2 
                           => n11513, B1 => n11615, B2 => n8521, ZN => n5243);
   U13963 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1523_port, A2 
                           => n8617, B1 => n11616, B2 => n8521, ZN => n5242);
   U13964 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1524_port, A2 
                           => n11513, B1 => n11617, B2 => n11512, ZN => n5241);
   U13965 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1525_port, A2 
                           => n8617, B1 => n11618, B2 => n8521, ZN => n5240);
   U13966 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1526_port, A2 
                           => n8617, B1 => n11619, B2 => n8521, ZN => n5239);
   U13967 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1527_port, A2 
                           => n11513, B1 => n11620, B2 => n8521, ZN => n5238);
   U13968 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1528_port, A2 
                           => n11513, B1 => n11621, B2 => n11512, ZN => n5237);
   U13969 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1529_port, A2 
                           => n11513, B1 => n11622, B2 => n11512, ZN => n5236);
   U13970 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1530_port, A2 
                           => n8617, B1 => n11623, B2 => n8521, ZN => n5235);
   U13971 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1531_port, A2 
                           => n8617, B1 => n11624, B2 => n8521, ZN => n5234);
   U13972 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1532_port, A2 
                           => n8617, B1 => n11625, B2 => n8521, ZN => n5233);
   U13973 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1533_port, A2 
                           => n11513, B1 => n11626, B2 => n11512, ZN => n5232);
   U13974 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1534_port, A2 
                           => n8617, B1 => n11627, B2 => n8521, ZN => n5231);
   U13975 : OAI22_X1 port map( A1 => n8617, A2 => n11629, B1 => 
                           DataPath_RF_bus_reg_dataout_1535_port, B2 => n11512,
                           ZN => n5228);
   U13976 : AOI22_X1 port map( A1 => n11597, A2 => n8522, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1472_port, ZN => n5226);
   U13977 : AOI22_X1 port map( A1 => n11598, A2 => n11514, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1473_port, ZN => n5225);
   U13978 : AOI22_X1 port map( A1 => n11599, A2 => n11514, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1474_port, ZN => n5224);
   U13979 : AOI22_X1 port map( A1 => n11600, A2 => n8522, B1 => n11515, B2 => 
                           DataPath_RF_bus_reg_dataout_1475_port, ZN => n5223);
   U13980 : AOI22_X1 port map( A1 => n11601, A2 => n8522, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1476_port, ZN => n5222);
   U13981 : AOI22_X1 port map( A1 => n11602, A2 => n11514, B1 => n11515, B2 => 
                           DataPath_RF_bus_reg_dataout_1477_port, ZN => n5221);
   U13982 : AOI22_X1 port map( A1 => n11603, A2 => n11514, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1478_port, ZN => n5220);
   U13983 : AOI22_X1 port map( A1 => n11604, A2 => n8522, B1 => n11515, B2 => 
                           DataPath_RF_bus_reg_dataout_1479_port, ZN => n5219);
   U13984 : AOI22_X1 port map( A1 => n11605, A2 => n8522, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1480_port, ZN => n5218);
   U13985 : AOI22_X1 port map( A1 => n11606, A2 => n11514, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1481_port, ZN => n5217);
   U13986 : AOI22_X1 port map( A1 => n11607, A2 => n11514, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1482_port, ZN => n5216);
   U13987 : AOI22_X1 port map( A1 => n11608, A2 => n8522, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1483_port, ZN => n5215);
   U13988 : AOI22_X1 port map( A1 => n11609, A2 => n8522, B1 => n11515, B2 => 
                           DataPath_RF_bus_reg_dataout_1484_port, ZN => n5214);
   U13989 : AOI22_X1 port map( A1 => n11610, A2 => n11514, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1485_port, ZN => n5213);
   U13990 : AOI22_X1 port map( A1 => n11611, A2 => n11514, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1486_port, ZN => n5212);
   U13991 : AOI22_X1 port map( A1 => n11612, A2 => n8522, B1 => n11515, B2 => 
                           DataPath_RF_bus_reg_dataout_1487_port, ZN => n5211);
   U13992 : AOI22_X1 port map( A1 => n11613, A2 => n8522, B1 => n11515, B2 => 
                           DataPath_RF_bus_reg_dataout_1488_port, ZN => n5210);
   U13993 : AOI22_X1 port map( A1 => n11614, A2 => n11514, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1489_port, ZN => n5209);
   U13994 : AOI22_X1 port map( A1 => n11615, A2 => n11514, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1490_port, ZN => n5208);
   U13995 : AOI22_X1 port map( A1 => n11616, A2 => n8522, B1 => n11515, B2 => 
                           DataPath_RF_bus_reg_dataout_1491_port, ZN => n5207);
   U13996 : AOI22_X1 port map( A1 => n11617, A2 => n8522, B1 => n11515, B2 => 
                           DataPath_RF_bus_reg_dataout_1492_port, ZN => n5206);
   U13997 : AOI22_X1 port map( A1 => n11618, A2 => n11514, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1493_port, ZN => n5205);
   U13998 : AOI22_X1 port map( A1 => n11619, A2 => n11514, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1494_port, ZN => n5204);
   U13999 : AOI22_X1 port map( A1 => n11620, A2 => n8522, B1 => n11515, B2 => 
                           DataPath_RF_bus_reg_dataout_1495_port, ZN => n5203);
   U14000 : AOI22_X1 port map( A1 => n11621, A2 => n8522, B1 => n11515, B2 => 
                           DataPath_RF_bus_reg_dataout_1496_port, ZN => n5202);
   U14001 : AOI22_X1 port map( A1 => n11622, A2 => n11514, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1497_port, ZN => n5201);
   U14002 : AOI22_X1 port map( A1 => n11623, A2 => n8522, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1498_port, ZN => n5200);
   U14003 : AOI22_X1 port map( A1 => n11624, A2 => n8522, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1499_port, ZN => n5199);
   U14004 : AOI22_X1 port map( A1 => n11625, A2 => n8522, B1 => n11515, B2 => 
                           DataPath_RF_bus_reg_dataout_1500_port, ZN => n5198);
   U14005 : AOI22_X1 port map( A1 => n11626, A2 => n8522, B1 => n11515, B2 => 
                           DataPath_RF_bus_reg_dataout_1501_port, ZN => n5197);
   U14006 : AOI22_X1 port map( A1 => n11627, A2 => n8522, B1 => n8618, B2 => 
                           DataPath_RF_bus_reg_dataout_1502_port, ZN => n5196);
   U14007 : OAI22_X1 port map( A1 => n11629, A2 => n8618, B1 => 
                           DataPath_RF_bus_reg_dataout_1503_port, B2 => n8522, 
                           ZN => n5193);
   U14008 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1440_port, A2 
                           => n8619, B1 => n11529, B2 => n11553, ZN => n5191);
   U14009 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1441_port, A2 
                           => n11531, B1 => n11529, B2 => n11554, ZN => n5190);
   U14010 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1442_port, A2 
                           => n8619, B1 => n11529, B2 => n11540, ZN => n5189);
   U14011 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1443_port, A2 
                           => n11531, B1 => n11529, B2 => n11555, ZN => n5188);
   U14012 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1444_port, A2 
                           => n8619, B1 => n11529, B2 => n11556, ZN => n5187);
   U14013 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1445_port, A2 
                           => n8619, B1 => n11529, B2 => n11557, ZN => n5186);
   U14014 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1446_port, A2 
                           => n11531, B1 => n11529, B2 => n11558, ZN => n5185);
   U14015 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1447_port, A2 
                           => n11531, B1 => n11529, B2 => n11559, ZN => n5184);
   U14016 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1448_port, A2 
                           => n11531, B1 => n11529, B2 => n11560, ZN => n5183);
   U14017 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1449_port, A2 
                           => n8619, B1 => n11529, B2 => n11561, ZN => n5182);
   U14018 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1450_port, A2 
                           => n8619, B1 => n11529, B2 => n11562, ZN => n5181);
   U14019 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1451_port, A2 
                           => n11531, B1 => n11529, B2 => n11563, ZN => n5180);
   U14020 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1452_port, A2 
                           => n11531, B1 => n11529, B2 => n11564, ZN => n5179);
   U14021 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1453_port, A2 
                           => n8619, B1 => n11529, B2 => n11565, ZN => n5178);
   U14022 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1454_port, A2 
                           => n8619, B1 => n11529, B2 => n11566, ZN => n5177);
   U14023 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1455_port, A2 
                           => n8619, B1 => n11529, B2 => n11567, ZN => n5176);
   U14024 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1456_port, A2 
                           => n11531, B1 => n11529, B2 => n11568, ZN => n5175);
   U14025 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1457_port, A2 
                           => n11531, B1 => n11529, B2 => n11569, ZN => n5174);
   U14026 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1458_port, A2 
                           => n8619, B1 => n11529, B2 => n11570, ZN => n5173);
   U14027 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1459_port, A2 
                           => n8619, B1 => n11529, B2 => n11571, ZN => n5172);
   U14028 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1460_port, A2 
                           => n8619, B1 => n11529, B2 => n11572, ZN => n5171);
   U14029 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1461_port, A2 
                           => n8619, B1 => n11529, B2 => n11573, ZN => n5170);
   U14030 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1462_port, A2 
                           => n8619, B1 => n11529, B2 => n11574, ZN => n5169);
   U14031 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1463_port, A2 
                           => n8619, B1 => n11529, B2 => n11575, ZN => n5168);
   U14032 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1464_port, A2 
                           => n11531, B1 => n11529, B2 => n11576, ZN => n5167);
   U14033 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1465_port, A2 
                           => n8619, B1 => n11529, B2 => n11577, ZN => n5166);
   U14034 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1466_port, A2 
                           => n8619, B1 => n11529, B2 => n11578, ZN => n5165);
   U14035 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1467_port, A2 
                           => n8619, B1 => n11529, B2 => n11579, ZN => n5164);
   U14036 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1468_port, A2 
                           => n11531, B1 => n11529, B2 => n11580, ZN => n5163);
   U14037 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1469_port, A2 
                           => n8619, B1 => n11529, B2 => n11581, ZN => n5162);
   U14038 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1470_port, A2 
                           => n8619, B1 => n11529, B2 => n11582, ZN => n5161);
   U14039 : OAI22_X1 port map( A1 => n11629, A2 => n8619, B1 => 
                           DataPath_RF_bus_reg_dataout_1471_port, B2 => n11530,
                           ZN => n5158);
   U14040 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1408_port, A2 
                           => n8620, B1 => n11532, B2 => n11553, ZN => n5156);
   U14041 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1409_port, A2 
                           => n11533, B1 => n11532, B2 => n11554, ZN => n5155);
   U14042 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1410_port, A2 
                           => n8620, B1 => n11532, B2 => n11540, ZN => n5154);
   U14043 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1411_port, A2 
                           => n8620, B1 => n11532, B2 => n11555, ZN => n5153);
   U14044 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1412_port, A2 
                           => n8620, B1 => n11532, B2 => n11556, ZN => n5152);
   U14045 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1413_port, A2 
                           => n8620, B1 => n11532, B2 => n11557, ZN => n5151);
   U14046 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1414_port, A2 
                           => n11533, B1 => n11532, B2 => n11558, ZN => n5150);
   U14047 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1415_port, A2 
                           => n8620, B1 => n11532, B2 => n11559, ZN => n5149);
   U14048 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1416_port, A2 
                           => n11533, B1 => n11532, B2 => n11560, ZN => n5148);
   U14049 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1417_port, A2 
                           => n8620, B1 => n11532, B2 => n11561, ZN => n5147);
   U14050 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1418_port, A2 
                           => n11533, B1 => n11532, B2 => n11562, ZN => n5146);
   U14051 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1419_port, A2 
                           => n8620, B1 => n11532, B2 => n11563, ZN => n5145);
   U14052 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1420_port, A2 
                           => n8620, B1 => n11532, B2 => n11564, ZN => n5144);
   U14053 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1421_port, A2 
                           => n8620, B1 => n11532, B2 => n11565, ZN => n5143);
   U14054 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1422_port, A2 
                           => n8620, B1 => n11532, B2 => n11566, ZN => n5142);
   U14055 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1423_port, A2 
                           => n11533, B1 => n11532, B2 => n11567, ZN => n5141);
   U14056 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1424_port, A2 
                           => n8620, B1 => n11532, B2 => n11568, ZN => n5140);
   U14057 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1425_port, A2 
                           => n11533, B1 => n11532, B2 => n11569, ZN => n5139);
   U14058 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1426_port, A2 
                           => n8620, B1 => n11532, B2 => n11570, ZN => n5138);
   U14059 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1427_port, A2 
                           => n11533, B1 => n11532, B2 => n11571, ZN => n5137);
   U14060 : AOI22_X1 port map( A1 => n11617, A2 => n11534, B1 => n8620, B2 => 
                           DataPath_RF_bus_reg_dataout_1428_port, ZN => n5136);
   U14061 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1429_port, A2 
                           => n8620, B1 => n11532, B2 => n11573, ZN => n5135);
   U14062 : AOI22_X1 port map( A1 => n11619, A2 => n11534, B1 => n8620, B2 => 
                           DataPath_RF_bus_reg_dataout_1430_port, ZN => n5134);
   U14063 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1431_port, A2 
                           => n8620, B1 => n11532, B2 => n11575, ZN => n5133);
   U14064 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1432_port, A2 
                           => n8620, B1 => n11532, B2 => n11576, ZN => n5132);
   U14065 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1433_port, A2 
                           => n8620, B1 => n11532, B2 => n11577, ZN => n5131);
   U14066 : AOI22_X1 port map( A1 => n11623, A2 => n11534, B1 => n8620, B2 => 
                           DataPath_RF_bus_reg_dataout_1434_port, ZN => n5130);
   U14067 : AOI22_X1 port map( A1 => n11624, A2 => n11534, B1 => n11533, B2 => 
                           DataPath_RF_bus_reg_dataout_1435_port, ZN => n5129);
   U14068 : AOI22_X1 port map( A1 => n11625, A2 => n11534, B1 => n8620, B2 => 
                           DataPath_RF_bus_reg_dataout_1436_port, ZN => n5128);
   U14069 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1437_port, A2 
                           => n11533, B1 => n11532, B2 => n11581, ZN => n5127);
   U14070 : AOI22_X1 port map( A1 => n11627, A2 => n11534, B1 => n11533, B2 => 
                           DataPath_RF_bus_reg_dataout_1438_port, ZN => n5126);
   U14071 : AOI22_X1 port map( A1 => n11629, A2 => n11534, B1 => n11533, B2 => 
                           DataPath_RF_bus_reg_dataout_1439_port, ZN => n5123);
   U14072 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1376_port, A2 
                           => n8621, B1 => n11535, B2 => n11553, ZN => n5121);
   U14073 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1377_port, A2 
                           => n8621, B1 => n11535, B2 => n11554, ZN => n5120);
   U14074 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1378_port, A2 
                           => n8621, B1 => n11535, B2 => n11540, ZN => n5119);
   U14075 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1379_port, A2 
                           => n11536, B1 => n11535, B2 => n11555, ZN => n5118);
   U14076 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1380_port, A2 
                           => n8621, B1 => n11535, B2 => n11556, ZN => n5117);
   U14077 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1381_port, A2 
                           => n8621, B1 => n11535, B2 => n11557, ZN => n5116);
   U14078 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1382_port, A2 
                           => n8621, B1 => n11535, B2 => n11558, ZN => n5115);
   U14079 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1383_port, A2 
                           => n11536, B1 => n11535, B2 => n11559, ZN => n5114);
   U14080 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1384_port, A2 
                           => n8621, B1 => n11535, B2 => n11560, ZN => n5113);
   U14081 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1385_port, A2 
                           => n8621, B1 => n11535, B2 => n11561, ZN => n5112);
   U14082 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1386_port, A2 
                           => n8621, B1 => n11535, B2 => n11562, ZN => n5111);
   U14083 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1387_port, A2 
                           => n8621, B1 => n11535, B2 => n11563, ZN => n5110);
   U14084 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1388_port, A2 
                           => n11536, B1 => n11535, B2 => n11564, ZN => n5109);
   U14085 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1389_port, A2 
                           => n11536, B1 => n11535, B2 => n11565, ZN => n5108);
   U14086 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1390_port, A2 
                           => n8621, B1 => n11535, B2 => n11566, ZN => n5107);
   U14087 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1391_port, A2 
                           => n8621, B1 => n11535, B2 => n11567, ZN => n5106);
   U14088 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1392_port, A2 
                           => n11536, B1 => n11535, B2 => n11568, ZN => n5105);
   U14089 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1393_port, A2 
                           => n11536, B1 => n11535, B2 => n11569, ZN => n5104);
   U14090 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1394_port, A2 
                           => n8621, B1 => n11535, B2 => n11570, ZN => n5103);
   U14091 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1395_port, A2 
                           => n8621, B1 => n11535, B2 => n11571, ZN => n5102);
   U14092 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1396_port, A2 
                           => n8621, B1 => n11535, B2 => n11572, ZN => n5101);
   U14093 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1397_port, A2 
                           => n11536, B1 => n11535, B2 => n11573, ZN => n5100);
   U14094 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1398_port, A2 
                           => n8621, B1 => n11535, B2 => n11574, ZN => n5099);
   U14095 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1399_port, A2 
                           => n8621, B1 => n11535, B2 => n11575, ZN => n5098);
   U14096 : AOI22_X1 port map( A1 => n11621, A2 => n11537, B1 => n11536, B2 => 
                           DataPath_RF_bus_reg_dataout_1400_port, ZN => n5097);
   U14097 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1401_port, A2 
                           => n8621, B1 => n11535, B2 => n11577, ZN => n5096);
   U14098 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1402_port, A2 
                           => n11536, B1 => n11535, B2 => n11578, ZN => n5095);
   U14099 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1403_port, A2 
                           => n11536, B1 => n11535, B2 => n11579, ZN => n5094);
   U14100 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1404_port, A2 
                           => n8621, B1 => n11535, B2 => n11580, ZN => n5093);
   U14101 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1405_port, A2 
                           => n8621, B1 => n11535, B2 => n11581, ZN => n5092);
   U14102 : AOI22_X1 port map( A1 => n11627, A2 => n11537, B1 => n11536, B2 => 
                           DataPath_RF_bus_reg_dataout_1406_port, ZN => n5091);
   U14103 : AOI22_X1 port map( A1 => n11629, A2 => n11537, B1 => n8621, B2 => 
                           DataPath_RF_bus_reg_dataout_1407_port, ZN => n5088);
   U14104 : OAI22_X1 port map( A1 => n11597, A2 => n11538, B1 => 
                           DataPath_RF_bus_reg_dataout_1344_port, B2 => n8523, 
                           ZN => n5086);
   U14105 : OAI22_X1 port map( A1 => n11598, A2 => n11538, B1 => 
                           DataPath_RF_bus_reg_dataout_1345_port, B2 => n11539,
                           ZN => n5085);
   U14106 : OAI22_X1 port map( A1 => n11599, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1346_port, B2 => n11539,
                           ZN => n5084);
   U14107 : OAI22_X1 port map( A1 => n11600, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1347_port, B2 => n8523, 
                           ZN => n5083);
   U14108 : OAI22_X1 port map( A1 => n11601, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1348_port, B2 => n8523, 
                           ZN => n5082);
   U14109 : OAI22_X1 port map( A1 => n11602, A2 => n11538, B1 => 
                           DataPath_RF_bus_reg_dataout_1349_port, B2 => n11539,
                           ZN => n5081);
   U14110 : OAI22_X1 port map( A1 => n11603, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1350_port, B2 => n11539,
                           ZN => n5080);
   U14111 : OAI22_X1 port map( A1 => n11604, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1351_port, B2 => n8523, 
                           ZN => n5079);
   U14112 : OAI22_X1 port map( A1 => n11605, A2 => n11538, B1 => 
                           DataPath_RF_bus_reg_dataout_1352_port, B2 => n8523, 
                           ZN => n5078);
   U14113 : OAI22_X1 port map( A1 => n11606, A2 => n11538, B1 => 
                           DataPath_RF_bus_reg_dataout_1353_port, B2 => n11539,
                           ZN => n5077);
   U14114 : OAI22_X1 port map( A1 => n11607, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1354_port, B2 => n11539,
                           ZN => n5076);
   U14115 : OAI22_X1 port map( A1 => n11608, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1355_port, B2 => n8523, 
                           ZN => n5075);
   U14116 : OAI22_X1 port map( A1 => n11609, A2 => n11538, B1 => 
                           DataPath_RF_bus_reg_dataout_1356_port, B2 => n8523, 
                           ZN => n5074);
   U14117 : OAI22_X1 port map( A1 => n11610, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1357_port, B2 => n11539,
                           ZN => n5073);
   U14118 : OAI22_X1 port map( A1 => n11611, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1358_port, B2 => n11539,
                           ZN => n5072);
   U14119 : OAI22_X1 port map( A1 => n11612, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1359_port, B2 => n8523, 
                           ZN => n5071);
   U14120 : OAI22_X1 port map( A1 => n11613, A2 => n11538, B1 => 
                           DataPath_RF_bus_reg_dataout_1360_port, B2 => n8523, 
                           ZN => n5070);
   U14121 : OAI22_X1 port map( A1 => n11614, A2 => n11538, B1 => 
                           DataPath_RF_bus_reg_dataout_1361_port, B2 => n11539,
                           ZN => n5069);
   U14122 : OAI22_X1 port map( A1 => n11615, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1362_port, B2 => n11539,
                           ZN => n5068);
   U14123 : OAI22_X1 port map( A1 => n11616, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1363_port, B2 => n8523, 
                           ZN => n5067);
   U14124 : OAI22_X1 port map( A1 => n11617, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1364_port, B2 => n8523, 
                           ZN => n5066);
   U14125 : OAI22_X1 port map( A1 => n11618, A2 => n11538, B1 => 
                           DataPath_RF_bus_reg_dataout_1365_port, B2 => n11539,
                           ZN => n5065);
   U14126 : OAI22_X1 port map( A1 => n11619, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1366_port, B2 => n11539,
                           ZN => n5064);
   U14127 : OAI22_X1 port map( A1 => n11620, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1367_port, B2 => n8523, 
                           ZN => n5063);
   U14128 : OAI22_X1 port map( A1 => n11621, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1368_port, B2 => n8523, 
                           ZN => n5062);
   U14129 : OAI22_X1 port map( A1 => n11622, A2 => n11538, B1 => 
                           DataPath_RF_bus_reg_dataout_1369_port, B2 => n11539,
                           ZN => n5061);
   U14130 : OAI22_X1 port map( A1 => n11623, A2 => n11538, B1 => 
                           DataPath_RF_bus_reg_dataout_1370_port, B2 => n8523, 
                           ZN => n5060);
   U14131 : OAI22_X1 port map( A1 => n11624, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1371_port, B2 => n8523, 
                           ZN => n5059);
   U14132 : OAI22_X1 port map( A1 => n11625, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1372_port, B2 => n8523, 
                           ZN => n5058);
   U14133 : OAI22_X1 port map( A1 => n11626, A2 => n8622, B1 => 
                           DataPath_RF_bus_reg_dataout_1373_port, B2 => n8523, 
                           ZN => n5057);
   U14134 : OAI22_X1 port map( A1 => n11627, A2 => n11538, B1 => 
                           DataPath_RF_bus_reg_dataout_1374_port, B2 => n8523, 
                           ZN => n5056);
   U14135 : AOI22_X1 port map( A1 => n11629, A2 => n11539, B1 => n8622, B2 => 
                           DataPath_RF_bus_reg_dataout_1375_port, ZN => n5053);
   U14136 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1312_port, A2 
                           => n11543, B1 => n11541, B2 => n11553, ZN => n5051);
   U14137 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1313_port, A2 
                           => n8623, B1 => n11541, B2 => n11554, ZN => n5050);
   U14138 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1314_port, A2 
                           => n8623, B1 => n11541, B2 => n11540, ZN => n5049);
   U14139 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1315_port, A2 
                           => n8623, B1 => n11541, B2 => n11555, ZN => n5048);
   U14140 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1316_port, A2 
                           => n11543, B1 => n11541, B2 => n11556, ZN => n5047);
   U14141 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1317_port, A2 
                           => n8623, B1 => n11541, B2 => n11557, ZN => n5046);
   U14142 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1318_port, A2 
                           => n8623, B1 => n11541, B2 => n11558, ZN => n5045);
   U14143 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1319_port, A2 
                           => n11543, B1 => n11541, B2 => n11559, ZN => n5044);
   U14144 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1320_port, A2 
                           => n11543, B1 => n11541, B2 => n11560, ZN => n5043);
   U14145 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1321_port, A2 
                           => n11543, B1 => n11541, B2 => n11561, ZN => n5042);
   U14146 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1322_port, A2 
                           => n8623, B1 => n11541, B2 => n11562, ZN => n5041);
   U14147 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1323_port, A2 
                           => n11543, B1 => n11541, B2 => n11563, ZN => n5040);
   U14148 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1324_port, A2 
                           => n8623, B1 => n11541, B2 => n11564, ZN => n5039);
   U14149 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1325_port, A2 
                           => n11543, B1 => n11541, B2 => n11565, ZN => n5038);
   U14150 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1326_port, A2 
                           => n8623, B1 => n11541, B2 => n11566, ZN => n5037);
   U14151 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1327_port, A2 
                           => n11543, B1 => n11541, B2 => n11567, ZN => n5036);
   U14152 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1328_port, A2 
                           => n11543, B1 => n11541, B2 => n11568, ZN => n5035);
   U14153 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1329_port, A2 
                           => n8623, B1 => n11541, B2 => n11569, ZN => n5034);
   U14154 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1330_port, A2 
                           => n8623, B1 => n11541, B2 => n11570, ZN => n5033);
   U14155 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1331_port, A2 
                           => n8623, B1 => n11541, B2 => n11571, ZN => n5032);
   U14156 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1332_port, A2 
                           => n11543, B1 => n11541, B2 => n11572, ZN => n5031);
   U14157 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1333_port, A2 
                           => n8623, B1 => n11541, B2 => n11573, ZN => n5030);
   U14158 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1334_port, A2 
                           => n8623, B1 => n11541, B2 => n11574, ZN => n5029);
   U14159 : AOI22_X1 port map( A1 => n11620, A2 => n11542, B1 => n8623, B2 => 
                           DataPath_RF_bus_reg_dataout_1335_port, ZN => n5028);
   U14160 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1336_port, A2 
                           => n8623, B1 => n11541, B2 => n11576, ZN => n5027);
   U14161 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1337_port, A2 
                           => n11543, B1 => n11541, B2 => n11577, ZN => n5026);
   U14162 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1338_port, A2 
                           => n8623, B1 => n11541, B2 => n11578, ZN => n5025);
   U14163 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1339_port, A2 
                           => n8623, B1 => n11541, B2 => n11579, ZN => n5024);
   U14164 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1340_port, A2 
                           => n8623, B1 => n11541, B2 => n11580, ZN => n5023);
   U14165 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1341_port, A2 
                           => n8623, B1 => n11541, B2 => n11581, ZN => n5022);
   U14166 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1342_port, A2 
                           => n8623, B1 => n11541, B2 => n11582, ZN => n5021);
   U14167 : OAI22_X1 port map( A1 => n11629, A2 => n8623, B1 => 
                           DataPath_RF_bus_reg_dataout_1343_port, B2 => n11542,
                           ZN => n5018);
   U14168 : OAI22_X1 port map( A1 => n11597, A2 => n11544, B1 => 
                           DataPath_RF_bus_reg_dataout_1280_port, B2 => n8524, 
                           ZN => n5016);
   U14169 : OAI22_X1 port map( A1 => n11598, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1281_port, B2 => n11545,
                           ZN => n5015);
   U14170 : OAI22_X1 port map( A1 => n11599, A2 => n11544, B1 => 
                           DataPath_RF_bus_reg_dataout_1282_port, B2 => n11545,
                           ZN => n5014);
   U14171 : OAI22_X1 port map( A1 => n11600, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1283_port, B2 => n8524, 
                           ZN => n5013);
   U14172 : OAI22_X1 port map( A1 => n11601, A2 => n11544, B1 => 
                           DataPath_RF_bus_reg_dataout_1284_port, B2 => n8524, 
                           ZN => n5012);
   U14173 : OAI22_X1 port map( A1 => n11602, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1285_port, B2 => n11545,
                           ZN => n5011);
   U14174 : OAI22_X1 port map( A1 => n11603, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1286_port, B2 => n11545,
                           ZN => n5010);
   U14175 : OAI22_X1 port map( A1 => n11604, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1287_port, B2 => n8524, 
                           ZN => n5009);
   U14176 : OAI22_X1 port map( A1 => n11605, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1288_port, B2 => n8524, 
                           ZN => n5008);
   U14177 : OAI22_X1 port map( A1 => n11606, A2 => n11544, B1 => 
                           DataPath_RF_bus_reg_dataout_1289_port, B2 => n11545,
                           ZN => n5007);
   U14178 : OAI22_X1 port map( A1 => n11607, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1290_port, B2 => n11545,
                           ZN => n5006);
   U14179 : OAI22_X1 port map( A1 => n11608, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1291_port, B2 => n8524, 
                           ZN => n5005);
   U14180 : AOI22_X1 port map( A1 => n11609, A2 => n8524, B1 => n8624, B2 => 
                           DataPath_RF_bus_reg_dataout_1292_port, ZN => n5004);
   U14181 : OAI22_X1 port map( A1 => n11610, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1293_port, B2 => n8524, 
                           ZN => n5003);
   U14182 : OAI22_X1 port map( A1 => n11611, A2 => n11544, B1 => 
                           DataPath_RF_bus_reg_dataout_1294_port, B2 => n11545,
                           ZN => n5002);
   U14183 : OAI22_X1 port map( A1 => n11612, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1295_port, B2 => n11545,
                           ZN => n5001);
   U14184 : OAI22_X1 port map( A1 => n11613, A2 => n11544, B1 => 
                           DataPath_RF_bus_reg_dataout_1296_port, B2 => n8524, 
                           ZN => n5000);
   U14185 : OAI22_X1 port map( A1 => n11614, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1297_port, B2 => n8524, 
                           ZN => n4999);
   U14186 : OAI22_X1 port map( A1 => n11615, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1298_port, B2 => n11545,
                           ZN => n4998);
   U14187 : OAI22_X1 port map( A1 => n11616, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1299_port, B2 => n11545,
                           ZN => n4997);
   U14188 : OAI22_X1 port map( A1 => n11617, A2 => n11544, B1 => 
                           DataPath_RF_bus_reg_dataout_1300_port, B2 => n8524, 
                           ZN => n4996);
   U14189 : AOI22_X1 port map( A1 => n11618, A2 => n11545, B1 => n8624, B2 => 
                           DataPath_RF_bus_reg_dataout_1301_port, ZN => n4995);
   U14190 : OAI22_X1 port map( A1 => n11619, A2 => n11544, B1 => 
                           DataPath_RF_bus_reg_dataout_1302_port, B2 => n8524, 
                           ZN => n4994);
   U14191 : OAI22_X1 port map( A1 => n11620, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1303_port, B2 => n11545,
                           ZN => n4993);
   U14192 : OAI22_X1 port map( A1 => n11621, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1304_port, B2 => n8524, 
                           ZN => n4992);
   U14193 : OAI22_X1 port map( A1 => n11622, A2 => n11544, B1 => 
                           DataPath_RF_bus_reg_dataout_1305_port, B2 => n8524, 
                           ZN => n4991);
   U14194 : OAI22_X1 port map( A1 => n11623, A2 => n11544, B1 => 
                           DataPath_RF_bus_reg_dataout_1306_port, B2 => n8524, 
                           ZN => n4990);
   U14195 : OAI22_X1 port map( A1 => n11624, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1307_port, B2 => n8524, 
                           ZN => n4989);
   U14196 : OAI22_X1 port map( A1 => n11625, A2 => n8624, B1 => 
                           DataPath_RF_bus_reg_dataout_1308_port, B2 => n8524, 
                           ZN => n4988);
   U14197 : OAI22_X1 port map( A1 => n11626, A2 => n11544, B1 => 
                           DataPath_RF_bus_reg_dataout_1309_port, B2 => n8524, 
                           ZN => n4987);
   U14198 : OAI22_X1 port map( A1 => n11627, A2 => n11544, B1 => 
                           DataPath_RF_bus_reg_dataout_1310_port, B2 => n8524, 
                           ZN => n4986);
   U14199 : AOI22_X1 port map( A1 => n11629, A2 => n11545, B1 => n8624, B2 => 
                           DataPath_RF_bus_reg_dataout_1311_port, ZN => n4983);
   U14200 : OAI22_X1 port map( A1 => n8442, A2 => n11824, B1 => n11596, B2 => 
                           n11823, ZN => n11546);
   U14201 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1248_port, B1 => n11597,
                           B2 => n11547, ZN => n4981);
   U14202 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1249_port, B1 => n11598,
                           B2 => n11547, ZN => n4980);
   U14203 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1250_port, B1 => n11599,
                           B2 => n11547, ZN => n4979);
   U14204 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1251_port, B1 => n11600,
                           B2 => n11547, ZN => n4978);
   U14205 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1252_port, B1 => n11601,
                           B2 => n11547, ZN => n4977);
   U14206 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1253_port, B1 => n11602,
                           B2 => n11547, ZN => n4976);
   U14207 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1254_port, B1 => n11603,
                           B2 => n11547, ZN => n4975);
   U14208 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1255_port, B1 => n11604,
                           B2 => n11547, ZN => n4974);
   U14209 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1256_port, B1 => n11605,
                           B2 => n11547, ZN => n4973);
   U14210 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1257_port, B1 => n11606,
                           B2 => n11547, ZN => n4972);
   U14211 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1258_port, B1 => n11607,
                           B2 => n11547, ZN => n4971);
   U14212 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1259_port, B1 => n11608,
                           B2 => n11547, ZN => n4970);
   U14213 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1260_port, B1 => n11609,
                           B2 => n11547, ZN => n4969);
   U14214 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1261_port, B1 => n11610,
                           B2 => n11547, ZN => n4968);
   U14215 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1262_port, B1 => n11611,
                           B2 => n11547, ZN => n4967);
   U14216 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1263_port, B1 => n11612,
                           B2 => n11547, ZN => n4966);
   U14217 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1264_port, B1 => n11613,
                           B2 => n11547, ZN => n4965);
   U14218 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1265_port, B1 => n11614,
                           B2 => n11547, ZN => n4964);
   U14219 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1266_port, B1 => n11615,
                           B2 => n11547, ZN => n4963);
   U14220 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1267_port, B1 => n11616,
                           B2 => n11547, ZN => n4962);
   U14221 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1268_port, B1 => n11617,
                           B2 => n11547, ZN => n4961);
   U14222 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1269_port, B1 => n11618,
                           B2 => n11547, ZN => n4960);
   U14223 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1270_port, B1 => n11619,
                           B2 => n11547, ZN => n4959);
   U14224 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1271_port, B1 => n11620,
                           B2 => n11547, ZN => n4958);
   U14225 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1272_port, B1 => n11621,
                           B2 => n11547, ZN => n4957);
   U14226 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1273_port, B1 => n11622,
                           B2 => n11547, ZN => n4956);
   U14227 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1274_port, B1 => n11623,
                           B2 => n11547, ZN => n4955);
   U14228 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1275_port, B1 => n11624,
                           B2 => n11547, ZN => n4954);
   U14229 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1276_port, B1 => n11625,
                           B2 => n11547, ZN => n4953);
   U14230 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1277_port, B1 => n11626,
                           B2 => n11547, ZN => n4952);
   U14231 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1278_port, B1 => n11627,
                           B2 => n11547, ZN => n4951);
   U14232 : AOI22_X1 port map( A1 => n8525, A2 => 
                           DataPath_RF_bus_reg_dataout_1279_port, B1 => n11629,
                           B2 => n11547, ZN => n4948);
   U14233 : OAI22_X1 port map( A1 => n8442, A2 => n11829, B1 => n11596, B2 => 
                           n11828, ZN => n11549);
   U14234 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1216_port, B1 => n11597,
                           B2 => n11550, ZN => n4946);
   U14235 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1217_port, B1 => n11598,
                           B2 => n11550, ZN => n4945);
   U14236 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1218_port, B1 => n11599,
                           B2 => n11550, ZN => n4944);
   U14237 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1219_port, B1 => n11600,
                           B2 => n11550, ZN => n4943);
   U14238 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1220_port, B1 => n11601,
                           B2 => n11550, ZN => n4942);
   U14239 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1221_port, B1 => n11602,
                           B2 => n11550, ZN => n4941);
   U14240 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1222_port, B1 => n11603,
                           B2 => n11550, ZN => n4940);
   U14241 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1223_port, B1 => n11604,
                           B2 => n11550, ZN => n4939);
   U14242 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1224_port, B1 => n11605,
                           B2 => n11550, ZN => n4938);
   U14243 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1225_port, B1 => n11606,
                           B2 => n11550, ZN => n4937);
   U14244 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1226_port, B1 => n11607,
                           B2 => n11550, ZN => n4936);
   U14245 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1227_port, B1 => n11608,
                           B2 => n11550, ZN => n4935);
   U14246 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1228_port, B1 => n11609,
                           B2 => n11550, ZN => n4934);
   U14247 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1229_port, B1 => n11610,
                           B2 => n11550, ZN => n4933);
   U14248 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1230_port, B1 => n11611,
                           B2 => n11550, ZN => n4932);
   U14249 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1231_port, B1 => n11612,
                           B2 => n11550, ZN => n4931);
   U14250 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1232_port, B1 => n11613,
                           B2 => n11550, ZN => n4930);
   U14251 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1233_port, B1 => n11614,
                           B2 => n11550, ZN => n4929);
   U14252 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1234_port, B1 => n11615,
                           B2 => n11550, ZN => n4928);
   U14253 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1235_port, B1 => n11616,
                           B2 => n11550, ZN => n4927);
   U14254 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1236_port, B1 => n11617,
                           B2 => n11550, ZN => n4926);
   U14255 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1237_port, B1 => n11618,
                           B2 => n11550, ZN => n4925);
   U14256 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1238_port, B1 => n11619,
                           B2 => n11550, ZN => n4924);
   U14257 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1239_port, B1 => n11620,
                           B2 => n11550, ZN => n4923);
   U14258 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1240_port, B1 => n11621,
                           B2 => n11550, ZN => n4922);
   U14259 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1241_port, B1 => n11622,
                           B2 => n11550, ZN => n4921);
   U14260 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1242_port, B1 => n11623,
                           B2 => n11550, ZN => n4920);
   U14261 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1243_port, B1 => n11624,
                           B2 => n11550, ZN => n4919);
   U14262 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1244_port, B1 => n11625,
                           B2 => n11550, ZN => n4918);
   U14263 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1245_port, B1 => n11626,
                           B2 => n11550, ZN => n4917);
   U14264 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1246_port, B1 => n11627,
                           B2 => n11550, ZN => n4916);
   U14265 : AOI22_X1 port map( A1 => n8526, A2 => 
                           DataPath_RF_bus_reg_dataout_1247_port, B1 => n11629,
                           B2 => n11550, ZN => n4913);
   U14266 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1184_port, A2 
                           => n11585, B1 => n11583, B2 => n11553, ZN => n4911);
   U14267 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1185_port, A2 
                           => n8625, B1 => n11583, B2 => n11554, ZN => n4910);
   U14268 : AOI22_X1 port map( A1 => n11599, A2 => n11584, B1 => n8625, B2 => 
                           DataPath_RF_bus_reg_dataout_1186_port, ZN => n4909);
   U14269 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1187_port, A2 
                           => n8625, B1 => n11583, B2 => n11555, ZN => n4908);
   U14270 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1188_port, A2 
                           => n8625, B1 => n11583, B2 => n11556, ZN => n4907);
   U14271 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1189_port, A2 
                           => n11585, B1 => n11583, B2 => n11557, ZN => n4906);
   U14272 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1190_port, A2 
                           => n8625, B1 => n11583, B2 => n11558, ZN => n4905);
   U14273 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1191_port, A2 
                           => n8625, B1 => n11583, B2 => n11559, ZN => n4904);
   U14274 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1192_port, A2 
                           => n8625, B1 => n11583, B2 => n11560, ZN => n4903);
   U14275 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1193_port, A2 
                           => n11585, B1 => n11583, B2 => n11561, ZN => n4902);
   U14276 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1194_port, A2 
                           => n11585, B1 => n11583, B2 => n11562, ZN => n4901);
   U14277 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1195_port, A2 
                           => n8625, B1 => n11583, B2 => n11563, ZN => n4900);
   U14278 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1196_port, A2 
                           => n11585, B1 => n11583, B2 => n11564, ZN => n4899);
   U14279 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1197_port, A2 
                           => n8625, B1 => n11583, B2 => n11565, ZN => n4898);
   U14280 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1198_port, A2 
                           => n11585, B1 => n11583, B2 => n11566, ZN => n4897);
   U14281 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1199_port, A2 
                           => n8625, B1 => n11583, B2 => n11567, ZN => n4896);
   U14282 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1200_port, A2 
                           => n8625, B1 => n11583, B2 => n11568, ZN => n4895);
   U14283 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1201_port, A2 
                           => n8625, B1 => n11583, B2 => n11569, ZN => n4894);
   U14284 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1202_port, A2 
                           => n11585, B1 => n11583, B2 => n11570, ZN => n4893);
   U14285 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1203_port, A2 
                           => n11585, B1 => n11583, B2 => n11571, ZN => n4892);
   U14286 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1204_port, A2 
                           => n8625, B1 => n11583, B2 => n11572, ZN => n4891);
   U14287 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1205_port, A2 
                           => n8625, B1 => n11583, B2 => n11573, ZN => n4890);
   U14288 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1206_port, A2 
                           => n8625, B1 => n11583, B2 => n11574, ZN => n4889);
   U14289 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1207_port, A2 
                           => n11585, B1 => n11583, B2 => n11575, ZN => n4888);
   U14290 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1208_port, A2 
                           => n8625, B1 => n11583, B2 => n11576, ZN => n4887);
   U14291 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1209_port, A2 
                           => n8625, B1 => n11583, B2 => n11577, ZN => n4886);
   U14292 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1210_port, A2 
                           => n8625, B1 => n11583, B2 => n11578, ZN => n4885);
   U14293 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1211_port, A2 
                           => n11585, B1 => n11583, B2 => n11579, ZN => n4884);
   U14294 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1212_port, A2 
                           => n8625, B1 => n11583, B2 => n11580, ZN => n4883);
   U14295 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1213_port, A2 
                           => n8625, B1 => n11583, B2 => n11581, ZN => n4882);
   U14296 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1214_port, A2 
                           => n8625, B1 => n11583, B2 => n11582, ZN => n4881);
   U14297 : OAI22_X1 port map( A1 => n11629, A2 => n11585, B1 => 
                           DataPath_RF_bus_reg_dataout_1215_port, B2 => n11584,
                           ZN => n4878);
   U14298 : OAI22_X1 port map( A1 => n8442, A2 => n11839, B1 => n11596, B2 => 
                           n11838, ZN => n11586);
   U14299 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1152_port, B1 => n11597,
                           B2 => n11587, ZN => n4876);
   U14300 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1153_port, B1 => n11598,
                           B2 => n11587, ZN => n4875);
   U14301 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1154_port, B1 => n11599,
                           B2 => n11587, ZN => n4874);
   U14302 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1155_port, B1 => n11600,
                           B2 => n11587, ZN => n4873);
   U14303 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1156_port, B1 => n11601,
                           B2 => n11587, ZN => n4872);
   U14304 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1157_port, B1 => n11602,
                           B2 => n11587, ZN => n4871);
   U14305 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1158_port, B1 => n11603,
                           B2 => n11587, ZN => n4870);
   U14306 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1159_port, B1 => n11604,
                           B2 => n11587, ZN => n4869);
   U14307 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1160_port, B1 => n11605,
                           B2 => n11587, ZN => n4868);
   U14308 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1161_port, B1 => n11606,
                           B2 => n11587, ZN => n4867);
   U14309 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1162_port, B1 => n11607,
                           B2 => n11587, ZN => n4866);
   U14310 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1163_port, B1 => n11608,
                           B2 => n11587, ZN => n4865);
   U14311 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1164_port, B1 => n11609,
                           B2 => n11587, ZN => n4864);
   U14312 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1165_port, B1 => n11610,
                           B2 => n11587, ZN => n4863);
   U14313 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1166_port, B1 => n11611,
                           B2 => n11587, ZN => n4862);
   U14314 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1167_port, B1 => n11612,
                           B2 => n11587, ZN => n4861);
   U14315 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1168_port, B1 => n11613,
                           B2 => n11587, ZN => n4860);
   U14316 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1169_port, B1 => n11614,
                           B2 => n11587, ZN => n4859);
   U14317 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1170_port, B1 => n11615,
                           B2 => n11587, ZN => n4858);
   U14318 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1171_port, B1 => n11616,
                           B2 => n11587, ZN => n4857);
   U14319 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1172_port, B1 => n11617,
                           B2 => n11587, ZN => n4856);
   U14320 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1173_port, B1 => n11618,
                           B2 => n11587, ZN => n4855);
   U14321 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1174_port, B1 => n11619,
                           B2 => n11587, ZN => n4854);
   U14322 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1175_port, B1 => n11620,
                           B2 => n11587, ZN => n4853);
   U14323 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1176_port, B1 => n11621,
                           B2 => n11587, ZN => n4852);
   U14324 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1177_port, B1 => n11622,
                           B2 => n11587, ZN => n4851);
   U14325 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1178_port, B1 => n11623,
                           B2 => n11587, ZN => n4850);
   U14326 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1179_port, B1 => n11624,
                           B2 => n11587, ZN => n4849);
   U14327 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1180_port, B1 => n11625,
                           B2 => n11587, ZN => n4848);
   U14328 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1181_port, B1 => n11626,
                           B2 => n11587, ZN => n4847);
   U14329 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1182_port, B1 => n11627,
                           B2 => n11587, ZN => n4846);
   U14330 : AOI22_X1 port map( A1 => n8527, A2 => 
                           DataPath_RF_bus_reg_dataout_1183_port, B1 => n11629,
                           B2 => n11587, ZN => n4843);
   U14331 : AOI22_X1 port map( A1 => n11597, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1120_port, ZN => n4841);
   U14332 : AOI22_X1 port map( A1 => n11598, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1121_port, ZN => n4840);
   U14333 : AOI22_X1 port map( A1 => n11599, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1122_port, ZN => n4839);
   U14334 : AOI22_X1 port map( A1 => n11600, A2 => n11590, B1 => n11591, B2 => 
                           DataPath_RF_bus_reg_dataout_1123_port, ZN => n4838);
   U14335 : AOI22_X1 port map( A1 => n11601, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1124_port, ZN => n4837);
   U14336 : AOI22_X1 port map( A1 => n11602, A2 => n11590, B1 => n11591, B2 => 
                           DataPath_RF_bus_reg_dataout_1125_port, ZN => n4836);
   U14337 : AOI22_X1 port map( A1 => n11603, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1126_port, ZN => n4835);
   U14338 : AOI22_X1 port map( A1 => n11604, A2 => n11590, B1 => n11591, B2 => 
                           DataPath_RF_bus_reg_dataout_1127_port, ZN => n4834);
   U14339 : AOI22_X1 port map( A1 => n11605, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1128_port, ZN => n4833);
   U14340 : AOI22_X1 port map( A1 => n11606, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1129_port, ZN => n4832);
   U14341 : AOI22_X1 port map( A1 => n11607, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1130_port, ZN => n4831);
   U14342 : AOI22_X1 port map( A1 => n11608, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1131_port, ZN => n4830);
   U14343 : AOI22_X1 port map( A1 => n11609, A2 => n11590, B1 => n11591, B2 => 
                           DataPath_RF_bus_reg_dataout_1132_port, ZN => n4829);
   U14344 : AOI22_X1 port map( A1 => n11610, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1133_port, ZN => n4828);
   U14345 : AOI22_X1 port map( A1 => n11611, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1134_port, ZN => n4827);
   U14346 : AOI22_X1 port map( A1 => n11612, A2 => n11590, B1 => n11591, B2 => 
                           DataPath_RF_bus_reg_dataout_1135_port, ZN => n4826);
   U14347 : AOI22_X1 port map( A1 => n11613, A2 => n11590, B1 => n11591, B2 => 
                           DataPath_RF_bus_reg_dataout_1136_port, ZN => n4825);
   U14348 : AOI22_X1 port map( A1 => n11614, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1137_port, ZN => n4824);
   U14349 : AOI22_X1 port map( A1 => n11615, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1138_port, ZN => n4823);
   U14350 : AOI22_X1 port map( A1 => n11616, A2 => n11590, B1 => n11591, B2 => 
                           DataPath_RF_bus_reg_dataout_1139_port, ZN => n4822);
   U14351 : AOI22_X1 port map( A1 => n11617, A2 => n11590, B1 => n11591, B2 => 
                           DataPath_RF_bus_reg_dataout_1140_port, ZN => n4821);
   U14352 : AOI22_X1 port map( A1 => n11618, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1141_port, ZN => n4820);
   U14353 : AOI22_X1 port map( A1 => n11619, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1142_port, ZN => n4819);
   U14354 : AOI22_X1 port map( A1 => n11620, A2 => n11590, B1 => n11591, B2 => 
                           DataPath_RF_bus_reg_dataout_1143_port, ZN => n4818);
   U14355 : AOI22_X1 port map( A1 => n11621, A2 => n11590, B1 => n11591, B2 => 
                           DataPath_RF_bus_reg_dataout_1144_port, ZN => n4817);
   U14356 : AOI22_X1 port map( A1 => n11622, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1145_port, ZN => n4816);
   U14357 : AOI22_X1 port map( A1 => n11623, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1146_port, ZN => n4815);
   U14358 : AOI22_X1 port map( A1 => n11624, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1147_port, ZN => n4814);
   U14359 : AOI22_X1 port map( A1 => n11625, A2 => n11590, B1 => n11591, B2 => 
                           DataPath_RF_bus_reg_dataout_1148_port, ZN => n4813);
   U14360 : AOI22_X1 port map( A1 => n11626, A2 => n11590, B1 => n11591, B2 => 
                           DataPath_RF_bus_reg_dataout_1149_port, ZN => n4812);
   U14361 : AOI22_X1 port map( A1 => n11627, A2 => n11590, B1 => n8626, B2 => 
                           DataPath_RF_bus_reg_dataout_1150_port, ZN => n4811);
   U14362 : OAI22_X1 port map( A1 => n11629, A2 => n8626, B1 => 
                           DataPath_RF_bus_reg_dataout_1151_port, B2 => n11590,
                           ZN => n4808);
   U14363 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1088_port, B1 => n11597,
                           B2 => n11592, ZN => n4806);
   U14364 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1089_port, B1 => n11598,
                           B2 => n11592, ZN => n4805);
   U14365 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1090_port, B1 => n11599,
                           B2 => n11592, ZN => n4804);
   U14366 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1091_port, B1 => n11600,
                           B2 => n11592, ZN => n4803);
   U14367 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1092_port, B1 => n11601,
                           B2 => n11592, ZN => n4802);
   U14368 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1093_port, B1 => n11602,
                           B2 => n11592, ZN => n4801);
   U14369 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1094_port, B1 => n11603,
                           B2 => n11592, ZN => n4800);
   U14370 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1095_port, B1 => n11604,
                           B2 => n11592, ZN => n4799);
   U14371 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1096_port, B1 => n11605,
                           B2 => n11592, ZN => n4798);
   U14372 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1097_port, B1 => n11606,
                           B2 => n11592, ZN => n4797);
   U14373 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1098_port, B1 => n11607,
                           B2 => n11592, ZN => n4796);
   U14374 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1099_port, B1 => n11608,
                           B2 => n11592, ZN => n4795);
   U14375 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1100_port, B1 => n11609,
                           B2 => n11592, ZN => n4794);
   U14376 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1101_port, B1 => n11610,
                           B2 => n11592, ZN => n4793);
   U14377 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1102_port, B1 => n11611,
                           B2 => n11592, ZN => n4792);
   U14378 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1103_port, B1 => n11612,
                           B2 => n11592, ZN => n4791);
   U14379 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1104_port, B1 => n11613,
                           B2 => n11592, ZN => n4790);
   U14380 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1105_port, B1 => n11614,
                           B2 => n11592, ZN => n4789);
   U14381 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1106_port, B1 => n11615,
                           B2 => n11592, ZN => n4788);
   U14382 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1107_port, B1 => n11616,
                           B2 => n11592, ZN => n4787);
   U14383 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1108_port, B1 => n11617,
                           B2 => n11592, ZN => n4786);
   U14384 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1109_port, B1 => n11618,
                           B2 => n11592, ZN => n4785);
   U14385 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1110_port, B1 => n11619,
                           B2 => n11592, ZN => n4784);
   U14386 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1111_port, B1 => n11620,
                           B2 => n11592, ZN => n4783);
   U14387 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1112_port, B1 => n11621,
                           B2 => n11592, ZN => n4782);
   U14388 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1113_port, B1 => n11622,
                           B2 => n11592, ZN => n4781);
   U14389 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1114_port, B1 => n11623,
                           B2 => n11592, ZN => n4780);
   U14390 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1115_port, B1 => n11624,
                           B2 => n11592, ZN => n4779);
   U14391 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1116_port, B1 => n11625,
                           B2 => n11592, ZN => n4778);
   U14392 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1117_port, B1 => n11626,
                           B2 => n11592, ZN => n4777);
   U14393 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1118_port, B1 => n11627,
                           B2 => n11592, ZN => n4776);
   U14394 : AOI22_X1 port map( A1 => n8528, A2 => 
                           DataPath_RF_bus_reg_dataout_1119_port, B1 => n11629,
                           B2 => n11592, ZN => n4773);
   U14395 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1056_port, B1 => n11597,
                           B2 => n11594, ZN => n4771);
   U14396 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1057_port, B1 => n11598,
                           B2 => n11594, ZN => n4770);
   U14397 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1058_port, B1 => n11599,
                           B2 => n11594, ZN => n4769);
   U14398 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1059_port, B1 => n11600,
                           B2 => n11594, ZN => n4768);
   U14399 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1060_port, B1 => n11601,
                           B2 => n11594, ZN => n4767);
   U14400 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1061_port, B1 => n11602,
                           B2 => n11594, ZN => n4766);
   U14401 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1062_port, B1 => n11603,
                           B2 => n11594, ZN => n4765);
   U14402 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1063_port, B1 => n11604,
                           B2 => n11594, ZN => n4764);
   U14403 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1064_port, B1 => n11605,
                           B2 => n11594, ZN => n4763);
   U14404 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1065_port, B1 => n11606,
                           B2 => n11594, ZN => n4762);
   U14405 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1066_port, B1 => n11607,
                           B2 => n11594, ZN => n4761);
   U14406 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1067_port, B1 => n11608,
                           B2 => n11594, ZN => n4760);
   U14407 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1068_port, B1 => n11609,
                           B2 => n11594, ZN => n4759);
   U14408 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1069_port, B1 => n11610,
                           B2 => n11594, ZN => n4758);
   U14409 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1070_port, B1 => n11611,
                           B2 => n11594, ZN => n4757);
   U14410 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1071_port, B1 => n11612,
                           B2 => n11594, ZN => n4756);
   U14411 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1072_port, B1 => n11613,
                           B2 => n11594, ZN => n4755);
   U14412 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1073_port, B1 => n11614,
                           B2 => n11594, ZN => n4754);
   U14413 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1074_port, B1 => n11615,
                           B2 => n11594, ZN => n4753);
   U14414 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1075_port, B1 => n11616,
                           B2 => n11594, ZN => n4752);
   U14415 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1076_port, B1 => n11617,
                           B2 => n11594, ZN => n4751);
   U14416 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1077_port, B1 => n11618,
                           B2 => n11594, ZN => n4750);
   U14417 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1078_port, B1 => n11619,
                           B2 => n11594, ZN => n4749);
   U14418 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1079_port, B1 => n11620,
                           B2 => n11594, ZN => n4748);
   U14419 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1080_port, B1 => n11621,
                           B2 => n11594, ZN => n4747);
   U14420 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1081_port, B1 => n11622,
                           B2 => n11594, ZN => n4746);
   U14421 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1082_port, B1 => n11623,
                           B2 => n11594, ZN => n4745);
   U14422 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1083_port, B1 => n11624,
                           B2 => n11594, ZN => n4744);
   U14423 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1084_port, B1 => n11625,
                           B2 => n11594, ZN => n4743);
   U14424 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1085_port, B1 => n11626,
                           B2 => n11594, ZN => n4742);
   U14425 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1086_port, B1 => n11627,
                           B2 => n11594, ZN => n4741);
   U14426 : AOI22_X1 port map( A1 => n8529, A2 => 
                           DataPath_RF_bus_reg_dataout_1087_port, B1 => n11629,
                           B2 => n11594, ZN => n4738);
   U14427 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1024_port, B1 => n11597,
                           B2 => n11628, ZN => n4734);
   U14428 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1025_port, B1 => n11598,
                           B2 => n11628, ZN => n4732);
   U14429 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1026_port, B1 => n11599,
                           B2 => n11628, ZN => n4730);
   U14430 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1027_port, B1 => n11600,
                           B2 => n11628, ZN => n4728);
   U14431 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1028_port, B1 => n11601,
                           B2 => n11628, ZN => n4726);
   U14432 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1029_port, B1 => n11602,
                           B2 => n11628, ZN => n4724);
   U14433 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1030_port, B1 => n11603,
                           B2 => n11628, ZN => n4722);
   U14434 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1031_port, B1 => n11604,
                           B2 => n11628, ZN => n4720);
   U14435 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1032_port, B1 => n11605,
                           B2 => n11628, ZN => n4718);
   U14436 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1033_port, B1 => n11606,
                           B2 => n11628, ZN => n4716);
   U14437 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1034_port, B1 => n11607,
                           B2 => n11628, ZN => n4714);
   U14438 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1035_port, B1 => n11608,
                           B2 => n11628, ZN => n4712);
   U14439 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1036_port, B1 => n11609,
                           B2 => n11628, ZN => n4710);
   U14440 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1037_port, B1 => n11610,
                           B2 => n11628, ZN => n4708);
   U14441 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1038_port, B1 => n11611,
                           B2 => n11628, ZN => n4706);
   U14442 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1039_port, B1 => n11612,
                           B2 => n11628, ZN => n4704);
   U14443 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1040_port, B1 => n11613,
                           B2 => n11628, ZN => n4702);
   U14444 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1041_port, B1 => n11614,
                           B2 => n11628, ZN => n4700);
   U14445 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1042_port, B1 => n11615,
                           B2 => n11628, ZN => n4698);
   U14446 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1043_port, B1 => n11616,
                           B2 => n11628, ZN => n4696);
   U14447 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1044_port, B1 => n11617,
                           B2 => n11628, ZN => n4694);
   U14448 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1045_port, B1 => n11618,
                           B2 => n11628, ZN => n4692);
   U14449 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1046_port, B1 => n11619,
                           B2 => n11628, ZN => n4690);
   U14450 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1047_port, B1 => n11620,
                           B2 => n11628, ZN => n4688);
   U14451 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1048_port, B1 => n11621,
                           B2 => n11628, ZN => n4686);
   U14452 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1049_port, B1 => n11622,
                           B2 => n11628, ZN => n4684);
   U14453 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1050_port, B1 => n11623,
                           B2 => n11628, ZN => n4682);
   U14454 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1051_port, B1 => n11624,
                           B2 => n11628, ZN => n4680);
   U14455 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1052_port, B1 => n11625,
                           B2 => n11628, ZN => n4678);
   U14456 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1053_port, B1 => n11626,
                           B2 => n11628, ZN => n4676);
   U14457 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1054_port, B1 => n11627,
                           B2 => n11628, ZN => n4674);
   U14458 : AOI22_X1 port map( A1 => n8530, A2 => 
                           DataPath_RF_bus_reg_dataout_1055_port, B1 => n11629,
                           B2 => n11628, ZN => n4670);
   U14459 : AOI22_X1 port map( A1 => n11716, A2 => n11634, B1 => n8627, B2 => 
                           DataPath_RF_bus_reg_dataout_992_port, ZN => n4668);
   U14460 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_993_port, A2 
                           => n8627, B1 => n11717, B2 => n8533, ZN => n4667);
   U14461 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_994_port, A2 
                           => n8627, B1 => n11718, B2 => n11634, ZN => n4666);
   U14462 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_995_port, A2 
                           => n11635, B1 => n11719, B2 => n11634, ZN => n4665);
   U14463 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_996_port, A2 
                           => n8627, B1 => n11720, B2 => n8533, ZN => n4664);
   U14464 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_997_port, A2 
                           => n8627, B1 => n11721, B2 => n8533, ZN => n4663);
   U14465 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_998_port, A2 
                           => n8627, B1 => n11722, B2 => n11634, ZN => n4662);
   U14466 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_999_port, A2 
                           => n11635, B1 => n11723, B2 => n11634, ZN => n4661);
   U14467 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1000_port, A2 
                           => n11635, B1 => n11724, B2 => n8533, ZN => n4660);
   U14468 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1001_port, A2 
                           => n8627, B1 => n11725, B2 => n8533, ZN => n4659);
   U14469 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1002_port, A2 
                           => n8627, B1 => n11726, B2 => n11634, ZN => n4658);
   U14470 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1003_port, A2 
                           => n8627, B1 => n11727, B2 => n11634, ZN => n4657);
   U14471 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1004_port, A2 
                           => n11635, B1 => n11728, B2 => n8533, ZN => n4656);
   U14472 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1005_port, A2 
                           => n8627, B1 => n11729, B2 => n8533, ZN => n4655);
   U14473 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1006_port, A2 
                           => n8627, B1 => n11730, B2 => n11634, ZN => n4654);
   U14474 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1007_port, A2 
                           => n8627, B1 => n11731, B2 => n11634, ZN => n4653);
   U14475 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1008_port, A2 
                           => n11635, B1 => n11732, B2 => n8533, ZN => n4652);
   U14476 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1009_port, A2 
                           => n11635, B1 => n11733, B2 => n8533, ZN => n4651);
   U14477 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1010_port, A2 
                           => n8627, B1 => n11734, B2 => n11634, ZN => n4650);
   U14478 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1011_port, A2 
                           => n8627, B1 => n11735, B2 => n11634, ZN => n4649);
   U14479 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1012_port, A2 
                           => n8627, B1 => n11736, B2 => n8533, ZN => n4648);
   U14480 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1013_port, A2 
                           => n11635, B1 => n11737, B2 => n8533, ZN => n4647);
   U14481 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1014_port, A2 
                           => n8627, B1 => n11738, B2 => n11634, ZN => n4646);
   U14482 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1015_port, A2 
                           => n8627, B1 => n11739, B2 => n11634, ZN => n4645);
   U14483 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1016_port, A2 
                           => n11635, B1 => n11740, B2 => n8533, ZN => n4644);
   U14484 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1017_port, A2 
                           => n11635, B1 => n11741, B2 => n8533, ZN => n4643);
   U14485 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1018_port, A2 
                           => n8627, B1 => n11742, B2 => n11634, ZN => n4642);
   U14486 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1019_port, A2 
                           => n8627, B1 => n11743, B2 => n8533, ZN => n4641);
   U14487 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1020_port, A2 
                           => n11635, B1 => n11744, B2 => n8533, ZN => n4640);
   U14488 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1021_port, A2 
                           => n11635, B1 => n11745, B2 => n8533, ZN => n4639);
   U14489 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1022_port, A2 
                           => n8627, B1 => n11746, B2 => n8533, ZN => n4638);
   U14490 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1023_port, A2 
                           => n8627, B1 => n11748, B2 => n8533, ZN => n4635);
   U14491 : OAI22_X1 port map( A1 => n11716, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_960_port, B2 => n11636, 
                           ZN => n4633);
   U14492 : OAI22_X1 port map( A1 => n11717, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_961_port, B2 => n11636, 
                           ZN => n4632);
   U14493 : OAI22_X1 port map( A1 => n11718, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_962_port, B2 => n8534, 
                           ZN => n4631);
   U14494 : OAI22_X1 port map( A1 => n11719, A2 => n11637, B1 => 
                           DataPath_RF_bus_reg_dataout_963_port, B2 => n8534, 
                           ZN => n4630);
   U14495 : OAI22_X1 port map( A1 => n11720, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_964_port, B2 => n11636, 
                           ZN => n4629);
   U14496 : OAI22_X1 port map( A1 => n11721, A2 => n11637, B1 => 
                           DataPath_RF_bus_reg_dataout_965_port, B2 => n11636, 
                           ZN => n4628);
   U14497 : OAI22_X1 port map( A1 => n11722, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_966_port, B2 => n8534, 
                           ZN => n4627);
   U14498 : OAI22_X1 port map( A1 => n11723, A2 => n11637, B1 => 
                           DataPath_RF_bus_reg_dataout_967_port, B2 => n8534, 
                           ZN => n4626);
   U14499 : OAI22_X1 port map( A1 => n11724, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_968_port, B2 => n11636, 
                           ZN => n4625);
   U14500 : OAI22_X1 port map( A1 => n11725, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_969_port, B2 => n11636, 
                           ZN => n4624);
   U14501 : OAI22_X1 port map( A1 => n11726, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_970_port, B2 => n8534, 
                           ZN => n4623);
   U14502 : OAI22_X1 port map( A1 => n11727, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_971_port, B2 => n8534, 
                           ZN => n4622);
   U14503 : OAI22_X1 port map( A1 => n11728, A2 => n11637, B1 => 
                           DataPath_RF_bus_reg_dataout_972_port, B2 => n11636, 
                           ZN => n4621);
   U14504 : OAI22_X1 port map( A1 => n11729, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_973_port, B2 => n11636, 
                           ZN => n4620);
   U14505 : OAI22_X1 port map( A1 => n11730, A2 => n11637, B1 => 
                           DataPath_RF_bus_reg_dataout_974_port, B2 => n8534, 
                           ZN => n4619);
   U14506 : OAI22_X1 port map( A1 => n11731, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_975_port, B2 => n8534, 
                           ZN => n4618);
   U14507 : OAI22_X1 port map( A1 => n11732, A2 => n11637, B1 => 
                           DataPath_RF_bus_reg_dataout_976_port, B2 => n11636, 
                           ZN => n4617);
   U14508 : OAI22_X1 port map( A1 => n11733, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_977_port, B2 => n11636, 
                           ZN => n4616);
   U14509 : OAI22_X1 port map( A1 => n11734, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_978_port, B2 => n8534, 
                           ZN => n4615);
   U14510 : OAI22_X1 port map( A1 => n11735, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_979_port, B2 => n8534, 
                           ZN => n4614);
   U14511 : OAI22_X1 port map( A1 => n11736, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_980_port, B2 => n11636, 
                           ZN => n4613);
   U14512 : OAI22_X1 port map( A1 => n11737, A2 => n11637, B1 => 
                           DataPath_RF_bus_reg_dataout_981_port, B2 => n11636, 
                           ZN => n4612);
   U14513 : OAI22_X1 port map( A1 => n11738, A2 => n11637, B1 => 
                           DataPath_RF_bus_reg_dataout_982_port, B2 => n8534, 
                           ZN => n4611);
   U14514 : OAI22_X1 port map( A1 => n11739, A2 => n11637, B1 => 
                           DataPath_RF_bus_reg_dataout_983_port, B2 => n8534, 
                           ZN => n4610);
   U14515 : OAI22_X1 port map( A1 => n11740, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_984_port, B2 => n11636, 
                           ZN => n4609);
   U14516 : OAI22_X1 port map( A1 => n11741, A2 => n11637, B1 => 
                           DataPath_RF_bus_reg_dataout_985_port, B2 => n8534, 
                           ZN => n4608);
   U14517 : OAI22_X1 port map( A1 => n11742, A2 => n11637, B1 => 
                           DataPath_RF_bus_reg_dataout_986_port, B2 => n8534, 
                           ZN => n4607);
   U14518 : OAI22_X1 port map( A1 => n11743, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_987_port, B2 => n8534, 
                           ZN => n4606);
   U14519 : OAI22_X1 port map( A1 => n11744, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_988_port, B2 => n8534, 
                           ZN => n4605);
   U14520 : OAI22_X1 port map( A1 => n11745, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_989_port, B2 => n8534, 
                           ZN => n4604);
   U14521 : OAI22_X1 port map( A1 => n11746, A2 => n8628, B1 => 
                           DataPath_RF_bus_reg_dataout_990_port, B2 => n8534, 
                           ZN => n4603);
   U14522 : OAI22_X1 port map( A1 => n11748, A2 => n11637, B1 => 
                           DataPath_RF_bus_reg_dataout_991_port, B2 => n8534, 
                           ZN => n4600);
   U14523 : OAI22_X1 port map( A1 => n11716, A2 => n8629, B1 => 
                           DataPath_RF_bus_reg_dataout_928_port, B2 => n11638, 
                           ZN => n4598);
   U14524 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_929_port, A2 
                           => n8629, B1 => n11652, B2 => n11665, ZN => n4597);
   U14525 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_930_port, A2 
                           => n8629, B1 => n11652, B2 => n11666, ZN => n4596);
   U14526 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_931_port, A2 
                           => n8629, B1 => n11652, B2 => n11667, ZN => n4595);
   U14527 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_932_port, A2 
                           => n11653, B1 => n11652, B2 => n11668, ZN => n4594);
   U14528 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_933_port, A2 
                           => n8629, B1 => n11652, B2 => n11669, ZN => n4593);
   U14529 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_934_port, A2 
                           => n11653, B1 => n11652, B2 => n11670, ZN => n4592);
   U14530 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_935_port, A2 
                           => n8629, B1 => n11652, B2 => n11671, ZN => n4591);
   U14531 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_936_port, A2 
                           => n11653, B1 => n11652, B2 => n11672, ZN => n4590);
   U14532 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_937_port, A2 
                           => n11653, B1 => n11652, B2 => n11673, ZN => n4589);
   U14533 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_938_port, A2 
                           => n8629, B1 => n11652, B2 => n11674, ZN => n4588);
   U14534 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_939_port, A2 
                           => n8629, B1 => n11652, B2 => n11675, ZN => n4587);
   U14535 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_940_port, A2 
                           => n8629, B1 => n11652, B2 => n11676, ZN => n4586);
   U14536 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_941_port, A2 
                           => n8629, B1 => n11652, B2 => n11677, ZN => n4585);
   U14537 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_942_port, A2 
                           => n8629, B1 => n11652, B2 => n11678, ZN => n4584);
   U14538 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_943_port, A2 
                           => n8629, B1 => n11652, B2 => n11679, ZN => n4583);
   U14539 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_944_port, A2 
                           => n8629, B1 => n11652, B2 => n11680, ZN => n4582);
   U14540 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_945_port, A2 
                           => n11653, B1 => n11652, B2 => n11681, ZN => n4581);
   U14541 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_946_port, A2 
                           => n11653, B1 => n11652, B2 => n11682, ZN => n4580);
   U14542 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_947_port, A2 
                           => n8629, B1 => n11652, B2 => n11683, ZN => n4579);
   U14543 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_948_port, A2 
                           => n8629, B1 => n11652, B2 => n11684, ZN => n4578);
   U14544 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_949_port, A2 
                           => n8629, B1 => n11652, B2 => n11685, ZN => n4577);
   U14545 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_950_port, A2 
                           => n11653, B1 => n11652, B2 => n11686, ZN => n4576);
   U14546 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_951_port, A2 
                           => n8629, B1 => n11652, B2 => n11687, ZN => n4575);
   U14547 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_952_port, A2 
                           => n11653, B1 => n11652, B2 => n11688, ZN => n4574);
   U14548 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_953_port, A2 
                           => n8629, B1 => n11652, B2 => n11689, ZN => n4573);
   U14549 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_954_port, A2 
                           => n11653, B1 => n11652, B2 => n11690, ZN => n4572);
   U14550 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_955_port, A2 
                           => n11653, B1 => n11652, B2 => n11691, ZN => n4571);
   U14551 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_956_port, A2 
                           => n8629, B1 => n11652, B2 => n11657, ZN => n4570);
   U14552 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_957_port, A2 
                           => n8629, B1 => n11652, B2 => n11658, ZN => n4569);
   U14553 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_958_port, A2 
                           => n8629, B1 => n11652, B2 => n11693, ZN => n4568);
   U14554 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_959_port, A2 
                           => n11653, B1 => n11652, B2 => n11694, ZN => n4565);
   U14555 : OAI22_X1 port map( A1 => n11716, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_896_port, B2 => n11654, 
                           ZN => n4563);
   U14556 : OAI22_X1 port map( A1 => n11717, A2 => n11655, B1 => 
                           DataPath_RF_bus_reg_dataout_897_port, B2 => n11654, 
                           ZN => n4562);
   U14557 : OAI22_X1 port map( A1 => n11718, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_898_port, B2 => n8535, 
                           ZN => n4561);
   U14558 : OAI22_X1 port map( A1 => n11719, A2 => n11655, B1 => 
                           DataPath_RF_bus_reg_dataout_899_port, B2 => n8535, 
                           ZN => n4560);
   U14559 : OAI22_X1 port map( A1 => n11720, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_900_port, B2 => n11654, 
                           ZN => n4559);
   U14560 : OAI22_X1 port map( A1 => n11721, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_901_port, B2 => n11654, 
                           ZN => n4558);
   U14561 : OAI22_X1 port map( A1 => n11722, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_902_port, B2 => n8535, 
                           ZN => n4557);
   U14562 : OAI22_X1 port map( A1 => n11723, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_903_port, B2 => n8535, 
                           ZN => n4556);
   U14563 : OAI22_X1 port map( A1 => n11724, A2 => n11655, B1 => 
                           DataPath_RF_bus_reg_dataout_904_port, B2 => n11654, 
                           ZN => n4555);
   U14564 : AOI22_X1 port map( A1 => n11725, A2 => n11654, B1 => n8630, B2 => 
                           DataPath_RF_bus_reg_dataout_905_port, ZN => n4554);
   U14565 : OAI22_X1 port map( A1 => n11726, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_906_port, B2 => n11654, 
                           ZN => n4553);
   U14566 : OAI22_X1 port map( A1 => n11727, A2 => n11655, B1 => 
                           DataPath_RF_bus_reg_dataout_907_port, B2 => n8535, 
                           ZN => n4552);
   U14567 : OAI22_X1 port map( A1 => n11728, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_908_port, B2 => n8535, 
                           ZN => n4551);
   U14568 : OAI22_X1 port map( A1 => n11729, A2 => n11655, B1 => 
                           DataPath_RF_bus_reg_dataout_909_port, B2 => n11654, 
                           ZN => n4550);
   U14569 : OAI22_X1 port map( A1 => n11730, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_910_port, B2 => n11654, 
                           ZN => n4549);
   U14570 : OAI22_X1 port map( A1 => n11731, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_911_port, B2 => n8535, 
                           ZN => n4548);
   U14571 : AOI22_X1 port map( A1 => n11732, A2 => n8535, B1 => n8630, B2 => 
                           DataPath_RF_bus_reg_dataout_912_port, ZN => n4547);
   U14572 : OAI22_X1 port map( A1 => n11733, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_913_port, B2 => n8535, 
                           ZN => n4546);
   U14573 : OAI22_X1 port map( A1 => n11734, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_914_port, B2 => n11654, 
                           ZN => n4545);
   U14574 : AOI22_X1 port map( A1 => n11735, A2 => n8535, B1 => n11655, B2 => 
                           DataPath_RF_bus_reg_dataout_915_port, ZN => n4544);
   U14575 : OAI22_X1 port map( A1 => n11736, A2 => n11655, B1 => 
                           DataPath_RF_bus_reg_dataout_916_port, B2 => n11654, 
                           ZN => n4543);
   U14576 : OAI22_X1 port map( A1 => n11737, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_917_port, B2 => n8535, 
                           ZN => n4542);
   U14577 : OAI22_X1 port map( A1 => n11738, A2 => n11655, B1 => 
                           DataPath_RF_bus_reg_dataout_918_port, B2 => n8535, 
                           ZN => n4541);
   U14578 : OAI22_X1 port map( A1 => n11739, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_919_port, B2 => n11654, 
                           ZN => n4540);
   U14579 : OAI22_X1 port map( A1 => n11740, A2 => n11655, B1 => 
                           DataPath_RF_bus_reg_dataout_920_port, B2 => n8535, 
                           ZN => n4539);
   U14580 : OAI22_X1 port map( A1 => n11741, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_921_port, B2 => n8535, 
                           ZN => n4538);
   U14581 : AOI22_X1 port map( A1 => n11742, A2 => n11654, B1 => n11655, B2 => 
                           DataPath_RF_bus_reg_dataout_922_port, ZN => n4537);
   U14582 : OAI22_X1 port map( A1 => n11743, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_923_port, B2 => n8535, 
                           ZN => n4536);
   U14583 : OAI22_X1 port map( A1 => n11744, A2 => n11655, B1 => 
                           DataPath_RF_bus_reg_dataout_924_port, B2 => n8535, 
                           ZN => n4535);
   U14584 : OAI22_X1 port map( A1 => n11745, A2 => n11655, B1 => 
                           DataPath_RF_bus_reg_dataout_925_port, B2 => n8535, 
                           ZN => n4534);
   U14585 : OAI22_X1 port map( A1 => n11746, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_926_port, B2 => n8535, 
                           ZN => n4533);
   U14586 : OAI22_X1 port map( A1 => n11748, A2 => n8630, B1 => 
                           DataPath_RF_bus_reg_dataout_927_port, B2 => n8535, 
                           ZN => n4530);
   U14587 : OAI22_X1 port map( A1 => n11716, A2 => n8631, B1 => 
                           DataPath_RF_bus_reg_dataout_864_port, B2 => n11656, 
                           ZN => n4528);
   U14588 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_865_port, A2 
                           => n8631, B1 => n11659, B2 => n11665, ZN => n4527);
   U14589 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_866_port, A2 
                           => n8631, B1 => n11659, B2 => n11666, ZN => n4526);
   U14590 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_867_port, A2 
                           => n11660, B1 => n11659, B2 => n11667, ZN => n4525);
   U14591 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_868_port, A2 
                           => n8631, B1 => n11659, B2 => n11668, ZN => n4524);
   U14592 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_869_port, A2 
                           => n8631, B1 => n11659, B2 => n11669, ZN => n4523);
   U14593 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_870_port, A2 
                           => n8631, B1 => n11659, B2 => n11670, ZN => n4522);
   U14594 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_871_port, A2 
                           => n11660, B1 => n11659, B2 => n11671, ZN => n4521);
   U14595 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_872_port, A2 
                           => n8631, B1 => n11659, B2 => n11672, ZN => n4520);
   U14596 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_873_port, A2 
                           => n8631, B1 => n11659, B2 => n11673, ZN => n4519);
   U14597 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_874_port, A2 
                           => n8631, B1 => n11659, B2 => n11674, ZN => n4518);
   U14598 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_875_port, A2 
                           => n11660, B1 => n11659, B2 => n11675, ZN => n4517);
   U14599 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_876_port, A2 
                           => n11660, B1 => n11659, B2 => n11676, ZN => n4516);
   U14600 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_877_port, A2 
                           => n8631, B1 => n11659, B2 => n11677, ZN => n4515);
   U14601 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_878_port, A2 
                           => n8631, B1 => n11659, B2 => n11678, ZN => n4514);
   U14602 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_879_port, A2 
                           => n8631, B1 => n11659, B2 => n11679, ZN => n4513);
   U14603 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_880_port, A2 
                           => n11660, B1 => n11659, B2 => n11680, ZN => n4512);
   U14604 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_881_port, A2 
                           => n8631, B1 => n11659, B2 => n11681, ZN => n4511);
   U14605 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_882_port, A2 
                           => n8631, B1 => n11659, B2 => n11682, ZN => n4510);
   U14606 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_883_port, A2 
                           => n11660, B1 => n11659, B2 => n11683, ZN => n4509);
   U14607 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_884_port, A2 
                           => n11660, B1 => n11659, B2 => n11684, ZN => n4508);
   U14608 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_885_port, A2 
                           => n8631, B1 => n11659, B2 => n11685, ZN => n4507);
   U14609 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_886_port, A2 
                           => n8631, B1 => n11659, B2 => n11686, ZN => n4506);
   U14610 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_887_port, A2 
                           => n8631, B1 => n11659, B2 => n11687, ZN => n4505);
   U14611 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_888_port, A2 
                           => n8631, B1 => n11659, B2 => n11688, ZN => n4504);
   U14612 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_889_port, A2 
                           => n8631, B1 => n11659, B2 => n11689, ZN => n4503);
   U14613 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_890_port, A2 
                           => n8631, B1 => n11659, B2 => n11690, ZN => n4502);
   U14614 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_891_port, A2 
                           => n11660, B1 => n11659, B2 => n11691, ZN => n4501);
   U14615 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_892_port, A2 
                           => n11660, B1 => n11659, B2 => n11657, ZN => n4500);
   U14616 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_893_port, A2 
                           => n8631, B1 => n11659, B2 => n11658, ZN => n4499);
   U14617 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_894_port, A2 
                           => n8631, B1 => n11659, B2 => n11693, ZN => n4498);
   U14618 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_895_port, A2 
                           => n11660, B1 => n11659, B2 => n11694, ZN => n4495);
   U14619 : OAI22_X1 port map( A1 => n11716, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_832_port, B2 => n11662, 
                           ZN => n4493);
   U14620 : OAI22_X1 port map( A1 => n11717, A2 => n11661, B1 => 
                           DataPath_RF_bus_reg_dataout_833_port, B2 => n11662, 
                           ZN => n4492);
   U14621 : OAI22_X1 port map( A1 => n11718, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_834_port, B2 => n8536, 
                           ZN => n4491);
   U14622 : OAI22_X1 port map( A1 => n11719, A2 => n11661, B1 => 
                           DataPath_RF_bus_reg_dataout_835_port, B2 => n8536, 
                           ZN => n4490);
   U14623 : OAI22_X1 port map( A1 => n11720, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_836_port, B2 => n11662, 
                           ZN => n4489);
   U14624 : OAI22_X1 port map( A1 => n11721, A2 => n11661, B1 => 
                           DataPath_RF_bus_reg_dataout_837_port, B2 => n11662, 
                           ZN => n4488);
   U14625 : OAI22_X1 port map( A1 => n11722, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_838_port, B2 => n8536, 
                           ZN => n4487);
   U14626 : OAI22_X1 port map( A1 => n11723, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_839_port, B2 => n8536, 
                           ZN => n4486);
   U14627 : OAI22_X1 port map( A1 => n11724, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_840_port, B2 => n11662, 
                           ZN => n4485);
   U14628 : OAI22_X1 port map( A1 => n11725, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_841_port, B2 => n11662, 
                           ZN => n4484);
   U14629 : OAI22_X1 port map( A1 => n11726, A2 => n11661, B1 => 
                           DataPath_RF_bus_reg_dataout_842_port, B2 => n8536, 
                           ZN => n4483);
   U14630 : OAI22_X1 port map( A1 => n11727, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_843_port, B2 => n8536, 
                           ZN => n4482);
   U14631 : OAI22_X1 port map( A1 => n11728, A2 => n11661, B1 => 
                           DataPath_RF_bus_reg_dataout_844_port, B2 => n11662, 
                           ZN => n4481);
   U14632 : OAI22_X1 port map( A1 => n11729, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_845_port, B2 => n11662, 
                           ZN => n4480);
   U14633 : OAI22_X1 port map( A1 => n11730, A2 => n11661, B1 => 
                           DataPath_RF_bus_reg_dataout_846_port, B2 => n8536, 
                           ZN => n4479);
   U14634 : OAI22_X1 port map( A1 => n11731, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_847_port, B2 => n8536, 
                           ZN => n4478);
   U14635 : OAI22_X1 port map( A1 => n11732, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_848_port, B2 => n11662, 
                           ZN => n4477);
   U14636 : OAI22_X1 port map( A1 => n11733, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_849_port, B2 => n11662, 
                           ZN => n4476);
   U14637 : OAI22_X1 port map( A1 => n11734, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_850_port, B2 => n8536, 
                           ZN => n4475);
   U14638 : OAI22_X1 port map( A1 => n11735, A2 => n11661, B1 => 
                           DataPath_RF_bus_reg_dataout_851_port, B2 => n8536, 
                           ZN => n4474);
   U14639 : OAI22_X1 port map( A1 => n11736, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_852_port, B2 => n11662, 
                           ZN => n4473);
   U14640 : OAI22_X1 port map( A1 => n11737, A2 => n11661, B1 => 
                           DataPath_RF_bus_reg_dataout_853_port, B2 => n11662, 
                           ZN => n4472);
   U14641 : OAI22_X1 port map( A1 => n11738, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_854_port, B2 => n8536, 
                           ZN => n4471);
   U14642 : OAI22_X1 port map( A1 => n11739, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_855_port, B2 => n8536, 
                           ZN => n4470);
   U14643 : OAI22_X1 port map( A1 => n11740, A2 => n11661, B1 => 
                           DataPath_RF_bus_reg_dataout_856_port, B2 => n11662, 
                           ZN => n4469);
   U14644 : OAI22_X1 port map( A1 => n11741, A2 => n11661, B1 => 
                           DataPath_RF_bus_reg_dataout_857_port, B2 => n8536, 
                           ZN => n4468);
   U14645 : OAI22_X1 port map( A1 => n11742, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_858_port, B2 => n8536, 
                           ZN => n4467);
   U14646 : OAI22_X1 port map( A1 => n11743, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_859_port, B2 => n8536, 
                           ZN => n4466);
   U14647 : AOI22_X1 port map( A1 => n11744, A2 => n8536, B1 => n11661, B2 => 
                           DataPath_RF_bus_reg_dataout_860_port, ZN => n4465);
   U14648 : OAI22_X1 port map( A1 => n11745, A2 => n11661, B1 => 
                           DataPath_RF_bus_reg_dataout_861_port, B2 => n8536, 
                           ZN => n4464);
   U14649 : OAI22_X1 port map( A1 => n11746, A2 => n8632, B1 => 
                           DataPath_RF_bus_reg_dataout_862_port, B2 => n8536, 
                           ZN => n4463);
   U14650 : AOI22_X1 port map( A1 => n11748, A2 => n11662, B1 => n8632, B2 => 
                           DataPath_RF_bus_reg_dataout_863_port, ZN => n4460);
   U14651 : AOI22_X1 port map( A1 => n11716, A2 => n11664, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_800_port, ZN => n4458);
   U14652 : AOI22_X1 port map( A1 => n11717, A2 => n8537, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_801_port, ZN => n4457);
   U14653 : AOI22_X1 port map( A1 => n11718, A2 => n8537, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_802_port, ZN => n4456);
   U14654 : AOI22_X1 port map( A1 => n11719, A2 => n11664, B1 => n11663, B2 => 
                           DataPath_RF_bus_reg_dataout_803_port, ZN => n4455);
   U14655 : AOI22_X1 port map( A1 => n11720, A2 => n11664, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_804_port, ZN => n4454);
   U14656 : AOI22_X1 port map( A1 => n11721, A2 => n8537, B1 => n11663, B2 => 
                           DataPath_RF_bus_reg_dataout_805_port, ZN => n4453);
   U14657 : AOI22_X1 port map( A1 => n11722, A2 => n8537, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_806_port, ZN => n4452);
   U14658 : AOI22_X1 port map( A1 => n11723, A2 => n11664, B1 => n11663, B2 => 
                           DataPath_RF_bus_reg_dataout_807_port, ZN => n4451);
   U14659 : AOI22_X1 port map( A1 => n11724, A2 => n11664, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_808_port, ZN => n4450);
   U14660 : AOI22_X1 port map( A1 => n11725, A2 => n8537, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_809_port, ZN => n4449);
   U14661 : AOI22_X1 port map( A1 => n11726, A2 => n8537, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_810_port, ZN => n4448);
   U14662 : AOI22_X1 port map( A1 => n11727, A2 => n11664, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_811_port, ZN => n4447);
   U14663 : AOI22_X1 port map( A1 => n11728, A2 => n11664, B1 => n11663, B2 => 
                           DataPath_RF_bus_reg_dataout_812_port, ZN => n4446);
   U14664 : AOI22_X1 port map( A1 => n11729, A2 => n8537, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_813_port, ZN => n4445);
   U14665 : AOI22_X1 port map( A1 => n11730, A2 => n8537, B1 => n11663, B2 => 
                           DataPath_RF_bus_reg_dataout_814_port, ZN => n4444);
   U14666 : AOI22_X1 port map( A1 => n11731, A2 => n11664, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_815_port, ZN => n4443);
   U14667 : AOI22_X1 port map( A1 => n11732, A2 => n11664, B1 => n11663, B2 => 
                           DataPath_RF_bus_reg_dataout_816_port, ZN => n4442);
   U14668 : AOI22_X1 port map( A1 => n11733, A2 => n8537, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_817_port, ZN => n4441);
   U14669 : AOI22_X1 port map( A1 => n11734, A2 => n8537, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_818_port, ZN => n4440);
   U14670 : AOI22_X1 port map( A1 => n11735, A2 => n11664, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_819_port, ZN => n4439);
   U14671 : AOI22_X1 port map( A1 => n11736, A2 => n11664, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_820_port, ZN => n4438);
   U14672 : AOI22_X1 port map( A1 => n11737, A2 => n8537, B1 => n11663, B2 => 
                           DataPath_RF_bus_reg_dataout_821_port, ZN => n4437);
   U14673 : AOI22_X1 port map( A1 => n11738, A2 => n8537, B1 => n11663, B2 => 
                           DataPath_RF_bus_reg_dataout_822_port, ZN => n4436);
   U14674 : AOI22_X1 port map( A1 => n11739, A2 => n11664, B1 => n11663, B2 => 
                           DataPath_RF_bus_reg_dataout_823_port, ZN => n4435);
   U14675 : AOI22_X1 port map( A1 => n11740, A2 => n11664, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_824_port, ZN => n4434);
   U14676 : AOI22_X1 port map( A1 => n11741, A2 => n8537, B1 => n11663, B2 => 
                           DataPath_RF_bus_reg_dataout_825_port, ZN => n4433);
   U14677 : AOI22_X1 port map( A1 => n11742, A2 => n8537, B1 => n11663, B2 => 
                           DataPath_RF_bus_reg_dataout_826_port, ZN => n4432);
   U14678 : AOI22_X1 port map( A1 => n11743, A2 => n8537, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_827_port, ZN => n4431);
   U14679 : AOI22_X1 port map( A1 => n11744, A2 => n8537, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_828_port, ZN => n4430);
   U14680 : AOI22_X1 port map( A1 => n11745, A2 => n8537, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_829_port, ZN => n4429);
   U14681 : AOI22_X1 port map( A1 => n11746, A2 => n8537, B1 => n8633, B2 => 
                           DataPath_RF_bus_reg_dataout_830_port, ZN => n4428);
   U14682 : AOI22_X1 port map( A1 => n11748, A2 => n8537, B1 => n11663, B2 => 
                           DataPath_RF_bus_reg_dataout_831_port, ZN => n4425);
   U14683 : OAI22_X1 port map( A1 => n11716, A2 => n8634, B1 => 
                           DataPath_RF_bus_reg_dataout_768_port, B2 => n11692, 
                           ZN => n4423);
   U14684 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_769_port, A2 
                           => n11696, B1 => n11695, B2 => n11665, ZN => n4422);
   U14685 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_770_port, A2 
                           => n8634, B1 => n11695, B2 => n11666, ZN => n4421);
   U14686 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_771_port, A2 
                           => n8634, B1 => n11695, B2 => n11667, ZN => n4420);
   U14687 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_772_port, A2 
                           => n8634, B1 => n11695, B2 => n11668, ZN => n4419);
   U14688 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_773_port, A2 
                           => n11696, B1 => n11695, B2 => n11669, ZN => n4418);
   U14689 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_774_port, A2 
                           => n8634, B1 => n11695, B2 => n11670, ZN => n4417);
   U14690 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_775_port, A2 
                           => n8634, B1 => n11695, B2 => n11671, ZN => n4416);
   U14691 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_776_port, A2 
                           => n8634, B1 => n11695, B2 => n11672, ZN => n4415);
   U14692 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_777_port, A2 
                           => n11696, B1 => n11695, B2 => n11673, ZN => n4414);
   U14693 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_778_port, A2 
                           => n8634, B1 => n11695, B2 => n11674, ZN => n4413);
   U14694 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_779_port, A2 
                           => n8634, B1 => n11695, B2 => n11675, ZN => n4412);
   U14695 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_780_port, A2 
                           => n11696, B1 => n11695, B2 => n11676, ZN => n4411);
   U14696 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_781_port, A2 
                           => n8634, B1 => n11695, B2 => n11677, ZN => n4410);
   U14697 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_782_port, A2 
                           => n8634, B1 => n11695, B2 => n11678, ZN => n4409);
   U14698 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_783_port, A2 
                           => n8634, B1 => n11695, B2 => n11679, ZN => n4408);
   U14699 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_784_port, A2 
                           => n11696, B1 => n11695, B2 => n11680, ZN => n4407);
   U14700 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_785_port, A2 
                           => n8634, B1 => n11695, B2 => n11681, ZN => n4406);
   U14701 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_786_port, A2 
                           => n8634, B1 => n11695, B2 => n11682, ZN => n4405);
   U14702 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_787_port, A2 
                           => n8634, B1 => n11695, B2 => n11683, ZN => n4404);
   U14703 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_788_port, A2 
                           => n11696, B1 => n11695, B2 => n11684, ZN => n4403);
   U14704 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_789_port, A2 
                           => n11696, B1 => n11695, B2 => n11685, ZN => n4402);
   U14705 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_790_port, A2 
                           => n8634, B1 => n11695, B2 => n11686, ZN => n4401);
   U14706 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_791_port, A2 
                           => n8634, B1 => n11695, B2 => n11687, ZN => n4400);
   U14707 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_792_port, A2 
                           => n8634, B1 => n11695, B2 => n11688, ZN => n4399);
   U14708 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_793_port, A2 
                           => n11696, B1 => n11695, B2 => n11689, ZN => n4398);
   U14709 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_794_port, A2 
                           => n8634, B1 => n11695, B2 => n11690, ZN => n4397);
   U14710 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_795_port, A2 
                           => n8634, B1 => n11695, B2 => n11691, ZN => n4396);
   U14711 : AOI22_X1 port map( A1 => n11744, A2 => n11692, B1 => n8634, B2 => 
                           DataPath_RF_bus_reg_dataout_796_port, ZN => n4395);
   U14712 : AOI22_X1 port map( A1 => n11745, A2 => n11692, B1 => n8634, B2 => 
                           DataPath_RF_bus_reg_dataout_797_port, ZN => n4394);
   U14713 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_798_port, A2 
                           => n11696, B1 => n11695, B2 => n11693, ZN => n4393);
   U14714 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_799_port, A2 
                           => n11696, B1 => n11695, B2 => n11694, ZN => n4390);
   U14715 : OAI22_X1 port map( A1 => n8442, A2 => n11823, B1 => n8299, B2 => 
                           n11824, ZN => n11697);
   U14716 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_736_port, B1 => n11716, 
                           B2 => n11698, ZN => n4388);
   U14717 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_737_port, B1 => n11717, 
                           B2 => n11698, ZN => n4387);
   U14718 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_738_port, B1 => n11718, 
                           B2 => n11698, ZN => n4386);
   U14719 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_739_port, B1 => n11719, 
                           B2 => n11698, ZN => n4385);
   U14720 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_740_port, B1 => n11720, 
                           B2 => n11698, ZN => n4384);
   U14721 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_741_port, B1 => n11721, 
                           B2 => n11698, ZN => n4383);
   U14722 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_742_port, B1 => n11722, 
                           B2 => n11698, ZN => n4382);
   U14723 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_743_port, B1 => n11723, 
                           B2 => n11698, ZN => n4381);
   U14724 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_744_port, B1 => n11724, 
                           B2 => n11698, ZN => n4380);
   U14725 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_745_port, B1 => n11725, 
                           B2 => n11698, ZN => n4379);
   U14726 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_746_port, B1 => n11726, 
                           B2 => n11698, ZN => n4378);
   U14727 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_747_port, B1 => n11727, 
                           B2 => n11698, ZN => n4377);
   U14728 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_748_port, B1 => n11728, 
                           B2 => n11698, ZN => n4376);
   U14729 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_749_port, B1 => n11729, 
                           B2 => n11698, ZN => n4375);
   U14730 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_750_port, B1 => n11730, 
                           B2 => n11698, ZN => n4374);
   U14731 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_751_port, B1 => n11731, 
                           B2 => n11698, ZN => n4373);
   U14732 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_752_port, B1 => n11732, 
                           B2 => n11698, ZN => n4372);
   U14733 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_753_port, B1 => n11733, 
                           B2 => n11698, ZN => n4371);
   U14734 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_754_port, B1 => n11734, 
                           B2 => n11698, ZN => n4370);
   U14735 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_755_port, B1 => n11735, 
                           B2 => n11698, ZN => n4369);
   U14736 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_756_port, B1 => n11736, 
                           B2 => n11698, ZN => n4368);
   U14737 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_757_port, B1 => n11737, 
                           B2 => n11698, ZN => n4367);
   U14738 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_758_port, B1 => n11738, 
                           B2 => n11698, ZN => n4366);
   U14739 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_759_port, B1 => n11739, 
                           B2 => n11698, ZN => n4365);
   U14740 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_760_port, B1 => n11740, 
                           B2 => n11698, ZN => n4364);
   U14741 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_761_port, B1 => n11741, 
                           B2 => n11698, ZN => n4363);
   U14742 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_762_port, B1 => n11742, 
                           B2 => n11698, ZN => n4362);
   U14743 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_763_port, B1 => n11743, 
                           B2 => n11698, ZN => n4361);
   U14744 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_764_port, B1 => n11744, 
                           B2 => n11698, ZN => n4360);
   U14745 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_765_port, B1 => n11745, 
                           B2 => n11698, ZN => n4359);
   U14746 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_766_port, B1 => n11746, 
                           B2 => n11698, ZN => n4358);
   U14747 : AOI22_X1 port map( A1 => n8538, A2 => 
                           DataPath_RF_bus_reg_dataout_767_port, B1 => n11748, 
                           B2 => n11698, ZN => n4355);
   U14748 : OAI22_X1 port map( A1 => n8442, A2 => n11828, B1 => n8299, B2 => 
                           n11829, ZN => n11700);
   U14749 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_704_port, B1 => n11716, 
                           B2 => n11701, ZN => n4353);
   U14750 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_705_port, B1 => n11717, 
                           B2 => n11701, ZN => n4352);
   U14751 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_706_port, B1 => n11718, 
                           B2 => n11701, ZN => n4351);
   U14752 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_707_port, B1 => n11719, 
                           B2 => n11701, ZN => n4350);
   U14753 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_708_port, B1 => n11720, 
                           B2 => n11701, ZN => n4349);
   U14754 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_709_port, B1 => n11721, 
                           B2 => n11701, ZN => n4348);
   U14755 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_710_port, B1 => n11722, 
                           B2 => n11701, ZN => n4347);
   U14756 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_711_port, B1 => n11723, 
                           B2 => n11701, ZN => n4346);
   U14757 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_712_port, B1 => n11724, 
                           B2 => n11701, ZN => n4345);
   U14758 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_713_port, B1 => n11725, 
                           B2 => n11701, ZN => n4344);
   U14759 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_714_port, B1 => n11726, 
                           B2 => n11701, ZN => n4343);
   U14760 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_715_port, B1 => n11727, 
                           B2 => n11701, ZN => n4342);
   U14761 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_716_port, B1 => n11728, 
                           B2 => n11701, ZN => n4341);
   U14762 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_717_port, B1 => n11729, 
                           B2 => n11701, ZN => n4340);
   U14763 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_718_port, B1 => n11730, 
                           B2 => n11701, ZN => n4339);
   U14764 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_719_port, B1 => n11731, 
                           B2 => n11701, ZN => n4338);
   U14765 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_720_port, B1 => n11732, 
                           B2 => n11701, ZN => n4337);
   U14766 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_721_port, B1 => n11733, 
                           B2 => n11701, ZN => n4336);
   U14767 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_722_port, B1 => n11734, 
                           B2 => n11701, ZN => n4335);
   U14768 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_723_port, B1 => n11735, 
                           B2 => n11701, ZN => n4334);
   U14769 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_724_port, B1 => n11736, 
                           B2 => n11701, ZN => n4333);
   U14770 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_725_port, B1 => n11737, 
                           B2 => n11701, ZN => n4332);
   U14771 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_726_port, B1 => n11738, 
                           B2 => n11701, ZN => n4331);
   U14772 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_727_port, B1 => n11739, 
                           B2 => n11701, ZN => n4330);
   U14773 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_728_port, B1 => n11740, 
                           B2 => n11701, ZN => n4329);
   U14774 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_729_port, B1 => n11741, 
                           B2 => n11701, ZN => n4328);
   U14775 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_730_port, B1 => n11742, 
                           B2 => n11701, ZN => n4327);
   U14776 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_731_port, B1 => n11743, 
                           B2 => n11701, ZN => n4326);
   U14777 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_732_port, B1 => n11744, 
                           B2 => n11701, ZN => n4325);
   U14778 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_733_port, B1 => n11745, 
                           B2 => n11701, ZN => n4324);
   U14779 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_734_port, B1 => n11746, 
                           B2 => n11701, ZN => n4323);
   U14780 : AOI22_X1 port map( A1 => n8539, A2 => 
                           DataPath_RF_bus_reg_dataout_735_port, B1 => n11748, 
                           B2 => n11701, ZN => n4320);
   U14781 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_672_port, B1 => n11716, 
                           B2 => n11704, ZN => n4318);
   U14782 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_673_port, B1 => n11717, 
                           B2 => n11704, ZN => n4317);
   U14783 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_674_port, B1 => n11718, 
                           B2 => n11704, ZN => n4316);
   U14784 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_675_port, B1 => n11719, 
                           B2 => n11704, ZN => n4315);
   U14785 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_676_port, B1 => n11720, 
                           B2 => n11704, ZN => n4314);
   U14786 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_677_port, B1 => n11721, 
                           B2 => n11704, ZN => n4313);
   U14787 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_678_port, B1 => n11722, 
                           B2 => n11704, ZN => n4312);
   U14788 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_679_port, B1 => n11723, 
                           B2 => n11704, ZN => n4311);
   U14789 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_680_port, B1 => n11724, 
                           B2 => n11704, ZN => n4310);
   U14790 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_681_port, B1 => n11725, 
                           B2 => n11704, ZN => n4309);
   U14791 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_682_port, B1 => n11726, 
                           B2 => n11704, ZN => n4308);
   U14792 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_683_port, B1 => n11727, 
                           B2 => n11704, ZN => n4307);
   U14793 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_684_port, B1 => n11728, 
                           B2 => n11704, ZN => n4306);
   U14794 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_685_port, B1 => n11729, 
                           B2 => n11704, ZN => n4305);
   U14795 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_686_port, B1 => n11730, 
                           B2 => n11704, ZN => n4304);
   U14796 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_687_port, B1 => n11731, 
                           B2 => n11704, ZN => n4303);
   U14797 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_688_port, B1 => n11732, 
                           B2 => n11704, ZN => n4302);
   U14798 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_689_port, B1 => n11733, 
                           B2 => n11704, ZN => n4301);
   U14799 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_690_port, B1 => n11734, 
                           B2 => n11704, ZN => n4300);
   U14800 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_691_port, B1 => n11735, 
                           B2 => n11704, ZN => n4299);
   U14801 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_692_port, B1 => n11736, 
                           B2 => n11704, ZN => n4298);
   U14802 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_693_port, B1 => n11737, 
                           B2 => n11704, ZN => n4297);
   U14803 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_694_port, B1 => n11738, 
                           B2 => n11704, ZN => n4296);
   U14804 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_695_port, B1 => n11739, 
                           B2 => n11704, ZN => n4295);
   U14805 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_696_port, B1 => n11740, 
                           B2 => n11704, ZN => n4294);
   U14806 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_697_port, B1 => n11741, 
                           B2 => n11704, ZN => n4293);
   U14807 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_698_port, B1 => n11742, 
                           B2 => n11704, ZN => n4292);
   U14808 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_699_port, B1 => n11743, 
                           B2 => n11704, ZN => n4291);
   U14809 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_700_port, B1 => n11744, 
                           B2 => n11704, ZN => n4290);
   U14810 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_701_port, B1 => n11745, 
                           B2 => n11704, ZN => n4289);
   U14811 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_702_port, B1 => n11746, 
                           B2 => n11704, ZN => n4288);
   U14812 : AOI22_X1 port map( A1 => n11705, A2 => 
                           DataPath_RF_bus_reg_dataout_703_port, B1 => n11748, 
                           B2 => n11704, ZN => n4285);
   U14813 : OAI22_X1 port map( A1 => n8442, A2 => n11838, B1 => n8299, B2 => 
                           n11839, ZN => n11706);
   U14814 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_640_port, B1 => n11716, 
                           B2 => n11707, ZN => n4283);
   U14815 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_641_port, B1 => n11717, 
                           B2 => n11707, ZN => n4282);
   U14816 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_642_port, B1 => n11718, 
                           B2 => n11707, ZN => n4281);
   U14817 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_643_port, B1 => n11719, 
                           B2 => n11707, ZN => n4280);
   U14818 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_644_port, B1 => n11720, 
                           B2 => n11707, ZN => n4279);
   U14819 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_645_port, B1 => n11721, 
                           B2 => n11707, ZN => n4278);
   U14820 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_646_port, B1 => n11722, 
                           B2 => n11707, ZN => n4277);
   U14821 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_647_port, B1 => n11723, 
                           B2 => n11707, ZN => n4276);
   U14822 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_648_port, B1 => n11724, 
                           B2 => n11707, ZN => n4275);
   U14823 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_649_port, B1 => n11725, 
                           B2 => n11707, ZN => n4274);
   U14824 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_650_port, B1 => n11726, 
                           B2 => n11707, ZN => n4273);
   U14825 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_651_port, B1 => n11727, 
                           B2 => n11707, ZN => n4272);
   U14826 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_652_port, B1 => n11728, 
                           B2 => n11707, ZN => n4271);
   U14827 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_653_port, B1 => n11729, 
                           B2 => n11707, ZN => n4270);
   U14828 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_654_port, B1 => n11730, 
                           B2 => n11707, ZN => n4269);
   U14829 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_655_port, B1 => n11731, 
                           B2 => n11707, ZN => n4268);
   U14830 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_656_port, B1 => n11732, 
                           B2 => n11707, ZN => n4267);
   U14831 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_657_port, B1 => n11733, 
                           B2 => n11707, ZN => n4266);
   U14832 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_658_port, B1 => n11734, 
                           B2 => n11707, ZN => n4265);
   U14833 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_659_port, B1 => n11735, 
                           B2 => n11707, ZN => n4264);
   U14834 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_660_port, B1 => n11736, 
                           B2 => n11707, ZN => n4263);
   U14835 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_661_port, B1 => n11737, 
                           B2 => n11707, ZN => n4262);
   U14836 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_662_port, B1 => n11738, 
                           B2 => n11707, ZN => n4261);
   U14837 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_663_port, B1 => n11739, 
                           B2 => n11707, ZN => n4260);
   U14838 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_664_port, B1 => n11740, 
                           B2 => n11707, ZN => n4259);
   U14839 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_665_port, B1 => n11741, 
                           B2 => n11707, ZN => n4258);
   U14840 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_666_port, B1 => n11742, 
                           B2 => n11707, ZN => n4257);
   U14841 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_667_port, B1 => n11743, 
                           B2 => n11707, ZN => n4256);
   U14842 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_668_port, B1 => n11744, 
                           B2 => n11707, ZN => n4255);
   U14843 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_669_port, B1 => n11745, 
                           B2 => n11707, ZN => n4254);
   U14844 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_670_port, B1 => n11746, 
                           B2 => n11707, ZN => n4253);
   U14845 : AOI22_X1 port map( A1 => n8540, A2 => 
                           DataPath_RF_bus_reg_dataout_671_port, B1 => n11748, 
                           B2 => n11707, ZN => n4250);
   U14846 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_608_port, B1 => n11716, 
                           B2 => n11710, ZN => n4248);
   U14847 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_609_port, B1 => n11717, 
                           B2 => n11710, ZN => n4247);
   U14848 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_610_port, B1 => n11718, 
                           B2 => n11710, ZN => n4246);
   U14849 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_611_port, B1 => n11719, 
                           B2 => n11710, ZN => n4245);
   U14850 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_612_port, B1 => n11720, 
                           B2 => n11710, ZN => n4244);
   U14851 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_613_port, B1 => n11721, 
                           B2 => n11710, ZN => n4243);
   U14852 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_614_port, B1 => n11722, 
                           B2 => n11710, ZN => n4242);
   U14853 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_615_port, B1 => n11723, 
                           B2 => n11710, ZN => n4241);
   U14854 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_616_port, B1 => n11724, 
                           B2 => n11710, ZN => n4240);
   U14855 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_617_port, B1 => n11725, 
                           B2 => n11710, ZN => n4239);
   U14856 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_618_port, B1 => n11726, 
                           B2 => n11710, ZN => n4238);
   U14857 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_619_port, B1 => n11727, 
                           B2 => n11710, ZN => n4237);
   U14858 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_620_port, B1 => n11728, 
                           B2 => n11710, ZN => n4236);
   U14859 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_621_port, B1 => n11729, 
                           B2 => n11710, ZN => n4235);
   U14860 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_622_port, B1 => n11730, 
                           B2 => n11710, ZN => n4234);
   U14861 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_623_port, B1 => n11731, 
                           B2 => n11710, ZN => n4233);
   U14862 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_624_port, B1 => n11732, 
                           B2 => n11710, ZN => n4232);
   U14863 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_625_port, B1 => n11733, 
                           B2 => n11710, ZN => n4231);
   U14864 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_626_port, B1 => n11734, 
                           B2 => n11710, ZN => n4230);
   U14865 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_627_port, B1 => n11735, 
                           B2 => n11710, ZN => n4229);
   U14866 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_628_port, B1 => n11736, 
                           B2 => n11710, ZN => n4228);
   U14867 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_629_port, B1 => n11737, 
                           B2 => n11710, ZN => n4227);
   U14868 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_630_port, B1 => n11738, 
                           B2 => n11710, ZN => n4226);
   U14869 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_631_port, B1 => n11739, 
                           B2 => n11710, ZN => n4225);
   U14870 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_632_port, B1 => n11740, 
                           B2 => n11710, ZN => n4224);
   U14871 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_633_port, B1 => n11741, 
                           B2 => n11710, ZN => n4223);
   U14872 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_634_port, B1 => n11742, 
                           B2 => n11710, ZN => n4222);
   U14873 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_635_port, B1 => n11743, 
                           B2 => n11710, ZN => n4221);
   U14874 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_636_port, B1 => n11744, 
                           B2 => n11710, ZN => n4220);
   U14875 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_637_port, B1 => n11745, 
                           B2 => n11710, ZN => n4219);
   U14876 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_638_port, B1 => n11746, 
                           B2 => n11710, ZN => n4218);
   U14877 : AOI22_X1 port map( A1 => n11711, A2 => 
                           DataPath_RF_bus_reg_dataout_639_port, B1 => n11748, 
                           B2 => n11710, ZN => n4215);
   U14878 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_576_port, B1 => n11716, 
                           B2 => n11712, ZN => n4213);
   U14879 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_577_port, B1 => n11717, 
                           B2 => n11712, ZN => n4212);
   U14880 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_578_port, B1 => n11718, 
                           B2 => n11712, ZN => n4211);
   U14881 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_579_port, B1 => n11719, 
                           B2 => n11712, ZN => n4210);
   U14882 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_580_port, B1 => n11720, 
                           B2 => n11712, ZN => n4209);
   U14883 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_581_port, B1 => n11721, 
                           B2 => n11712, ZN => n4208);
   U14884 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_582_port, B1 => n11722, 
                           B2 => n11712, ZN => n4207);
   U14885 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_583_port, B1 => n11723, 
                           B2 => n11712, ZN => n4206);
   U14886 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_584_port, B1 => n11724, 
                           B2 => n11712, ZN => n4205);
   U14887 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_585_port, B1 => n11725, 
                           B2 => n11712, ZN => n4204);
   U14888 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_586_port, B1 => n11726, 
                           B2 => n11712, ZN => n4203);
   U14889 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_587_port, B1 => n11727, 
                           B2 => n11712, ZN => n4202);
   U14890 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_588_port, B1 => n11728, 
                           B2 => n11712, ZN => n4201);
   U14891 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_589_port, B1 => n11729, 
                           B2 => n11712, ZN => n4200);
   U14892 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_590_port, B1 => n11730, 
                           B2 => n11712, ZN => n4199);
   U14893 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_591_port, B1 => n11731, 
                           B2 => n11712, ZN => n4198);
   U14894 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_592_port, B1 => n11732, 
                           B2 => n11712, ZN => n4197);
   U14895 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_593_port, B1 => n11733, 
                           B2 => n11712, ZN => n4196);
   U14896 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_594_port, B1 => n11734, 
                           B2 => n11712, ZN => n4195);
   U14897 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_595_port, B1 => n11735, 
                           B2 => n11712, ZN => n4194);
   U14898 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_596_port, B1 => n11736, 
                           B2 => n11712, ZN => n4193);
   U14899 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_597_port, B1 => n11737, 
                           B2 => n11712, ZN => n4192);
   U14900 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_598_port, B1 => n11738, 
                           B2 => n11712, ZN => n4191);
   U14901 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_599_port, B1 => n11739, 
                           B2 => n11712, ZN => n4190);
   U14902 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_600_port, B1 => n11740, 
                           B2 => n11712, ZN => n4189);
   U14903 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_601_port, B1 => n11741, 
                           B2 => n11712, ZN => n4188);
   U14904 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_602_port, B1 => n11742, 
                           B2 => n11712, ZN => n4187);
   U14905 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_603_port, B1 => n11743, 
                           B2 => n11712, ZN => n4186);
   U14906 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_604_port, B1 => n11744, 
                           B2 => n11712, ZN => n4185);
   U14907 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_605_port, B1 => n11745, 
                           B2 => n11712, ZN => n4184);
   U14908 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_606_port, B1 => n11746, 
                           B2 => n11712, ZN => n4183);
   U14909 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_bus_reg_dataout_607_port, B1 => n11748, 
                           B2 => n11712, ZN => n4180);
   U14910 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_544_port, B1 => n11716, 
                           B2 => n11714, ZN => n4178);
   U14911 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_545_port, B1 => n11717, 
                           B2 => n11714, ZN => n4177);
   U14912 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_546_port, B1 => n11718, 
                           B2 => n11714, ZN => n4176);
   U14913 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_547_port, B1 => n11719, 
                           B2 => n11714, ZN => n4175);
   U14914 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_548_port, B1 => n11720, 
                           B2 => n11714, ZN => n4174);
   U14915 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_549_port, B1 => n11721, 
                           B2 => n11714, ZN => n4173);
   U14916 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_550_port, B1 => n11722, 
                           B2 => n11714, ZN => n4172);
   U14917 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_551_port, B1 => n11723, 
                           B2 => n11714, ZN => n4171);
   U14918 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_552_port, B1 => n11724, 
                           B2 => n11714, ZN => n4170);
   U14919 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_553_port, B1 => n11725, 
                           B2 => n11714, ZN => n4169);
   U14920 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_554_port, B1 => n11726, 
                           B2 => n11714, ZN => n4168);
   U14921 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_555_port, B1 => n11727, 
                           B2 => n11714, ZN => n4167);
   U14922 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_556_port, B1 => n11728, 
                           B2 => n11714, ZN => n4166);
   U14923 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_557_port, B1 => n11729, 
                           B2 => n11714, ZN => n4165);
   U14924 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_558_port, B1 => n11730, 
                           B2 => n11714, ZN => n4164);
   U14925 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_559_port, B1 => n11731, 
                           B2 => n11714, ZN => n4163);
   U14926 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_560_port, B1 => n11732, 
                           B2 => n11714, ZN => n4162);
   U14927 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_561_port, B1 => n11733, 
                           B2 => n11714, ZN => n4161);
   U14928 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_562_port, B1 => n11734, 
                           B2 => n11714, ZN => n4160);
   U14929 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_563_port, B1 => n11735, 
                           B2 => n11714, ZN => n4159);
   U14930 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_564_port, B1 => n11736, 
                           B2 => n11714, ZN => n4158);
   U14931 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_565_port, B1 => n11737, 
                           B2 => n11714, ZN => n4157);
   U14932 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_566_port, B1 => n11738, 
                           B2 => n11714, ZN => n4156);
   U14933 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_567_port, B1 => n11739, 
                           B2 => n11714, ZN => n4155);
   U14934 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_568_port, B1 => n11740, 
                           B2 => n11714, ZN => n4154);
   U14935 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_569_port, B1 => n11741, 
                           B2 => n11714, ZN => n4153);
   U14936 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_570_port, B1 => n11742, 
                           B2 => n11714, ZN => n4152);
   U14937 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_571_port, B1 => n11743, 
                           B2 => n11714, ZN => n4151);
   U14938 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_572_port, B1 => n11744, 
                           B2 => n11714, ZN => n4150);
   U14939 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_573_port, B1 => n11745, 
                           B2 => n11714, ZN => n4149);
   U14940 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_574_port, B1 => n11746, 
                           B2 => n11714, ZN => n4148);
   U14941 : AOI22_X1 port map( A1 => n8542, A2 => 
                           DataPath_RF_bus_reg_dataout_575_port, B1 => n11748, 
                           B2 => n11714, ZN => n4145);
   U14942 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_512_port, B1 => n11716, 
                           B2 => n11747, ZN => n4141);
   U14943 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_513_port, B1 => n11717, 
                           B2 => n11747, ZN => n4139);
   U14944 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_514_port, B1 => n11718, 
                           B2 => n11747, ZN => n4137);
   U14945 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_515_port, B1 => n11719, 
                           B2 => n11747, ZN => n4135);
   U14946 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_516_port, B1 => n11720, 
                           B2 => n11747, ZN => n4133);
   U14947 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_517_port, B1 => n11721, 
                           B2 => n11747, ZN => n4131);
   U14948 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_518_port, B1 => n11722, 
                           B2 => n11747, ZN => n4129);
   U14949 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_519_port, B1 => n11723, 
                           B2 => n11747, ZN => n4127);
   U14950 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_520_port, B1 => n11724, 
                           B2 => n11747, ZN => n4125);
   U14951 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_521_port, B1 => n11725, 
                           B2 => n11747, ZN => n4123);
   U14952 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_522_port, B1 => n11726, 
                           B2 => n11747, ZN => n4121);
   U14953 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_523_port, B1 => n11727, 
                           B2 => n11747, ZN => n4119);
   U14954 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_524_port, B1 => n11728, 
                           B2 => n11747, ZN => n4117);
   U14955 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_525_port, B1 => n11729, 
                           B2 => n11747, ZN => n4115);
   U14956 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_526_port, B1 => n11730, 
                           B2 => n11747, ZN => n4113);
   U14957 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_527_port, B1 => n11731, 
                           B2 => n11747, ZN => n4111);
   U14958 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_528_port, B1 => n11732, 
                           B2 => n11747, ZN => n4109);
   U14959 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_529_port, B1 => n11733, 
                           B2 => n11747, ZN => n4107);
   U14960 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_530_port, B1 => n11734, 
                           B2 => n11747, ZN => n4105);
   U14961 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_531_port, B1 => n11735, 
                           B2 => n11747, ZN => n4103);
   U14962 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_532_port, B1 => n11736, 
                           B2 => n11747, ZN => n4101);
   U14963 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_533_port, B1 => n11737, 
                           B2 => n11747, ZN => n4099);
   U14964 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_534_port, B1 => n11738, 
                           B2 => n11747, ZN => n4097);
   U14965 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_535_port, B1 => n11739, 
                           B2 => n11747, ZN => n4095);
   U14966 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_536_port, B1 => n11740, 
                           B2 => n11747, ZN => n4093);
   U14967 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_537_port, B1 => n11741, 
                           B2 => n11747, ZN => n4091);
   U14968 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_538_port, B1 => n11742, 
                           B2 => n11747, ZN => n4089);
   U14969 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_539_port, B1 => n11743, 
                           B2 => n11747, ZN => n4087);
   U14970 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_540_port, B1 => n11744, 
                           B2 => n11747, ZN => n4085);
   U14971 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_541_port, B1 => n11745, 
                           B2 => n11747, ZN => n4083);
   U14972 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_542_port, B1 => n11746, 
                           B2 => n11747, ZN => n4081);
   U14973 : AOI22_X1 port map( A1 => n8543, A2 => 
                           DataPath_RF_bus_reg_dataout_543_port, B1 => n11748, 
                           B2 => n11747, ZN => n4077);
   U14974 : OAI22_X1 port map( A1 => n11858, A2 => n8635, B1 => 
                           DataPath_RF_bus_reg_dataout_480_port, B2 => n7802, 
                           ZN => n4074);
   U14975 : OAI22_X1 port map( A1 => n8635, A2 => n11859, B1 => 
                           DataPath_RF_bus_reg_dataout_481_port, B2 => n7802, 
                           ZN => n4072);
   U14976 : OAI22_X1 port map( A1 => n8635, A2 => n11860, B1 => 
                           DataPath_RF_bus_reg_dataout_482_port, B2 => n7802, 
                           ZN => n4070);
   U14977 : OAI22_X1 port map( A1 => n8635, A2 => n11861, B1 => 
                           DataPath_RF_bus_reg_dataout_483_port, B2 => n7802, 
                           ZN => n4068);
   U14978 : OAI22_X1 port map( A1 => n11766, A2 => n11862, B1 => 
                           DataPath_RF_bus_reg_dataout_484_port, B2 => n7802, 
                           ZN => n4066);
   U14979 : OAI22_X1 port map( A1 => n11766, A2 => n11863, B1 => 
                           DataPath_RF_bus_reg_dataout_485_port, B2 => n7802, 
                           ZN => n4064);
   U14980 : OAI22_X1 port map( A1 => n11766, A2 => n11864, B1 => 
                           DataPath_RF_bus_reg_dataout_486_port, B2 => n7802, 
                           ZN => n4062);
   U14981 : OR2_X1 port map( A1 => RST, A2 => n11750, ZN => n3350);
   U14982 : OAI22_X1 port map( A1 => n8635, A2 => n11865, B1 => 
                           DataPath_RF_bus_reg_dataout_487_port, B2 => n7802, 
                           ZN => n4060);
   U14983 : OAI22_X1 port map( A1 => n8635, A2 => n11866, B1 => 
                           DataPath_RF_bus_reg_dataout_488_port, B2 => n7802, 
                           ZN => n4058);
   U14984 : OAI22_X1 port map( A1 => n8635, A2 => n11867, B1 => 
                           DataPath_RF_bus_reg_dataout_489_port, B2 => n7802, 
                           ZN => n4056);
   U14985 : OAI22_X1 port map( A1 => n8635, A2 => n11868, B1 => 
                           DataPath_RF_bus_reg_dataout_490_port, B2 => n7802, 
                           ZN => n4054);
   U14986 : OAI22_X1 port map( A1 => n8635, A2 => n11869, B1 => 
                           DataPath_RF_bus_reg_dataout_491_port, B2 => n7802, 
                           ZN => n4052);
   U14987 : OAI22_X1 port map( A1 => n8635, A2 => n11870, B1 => 
                           DataPath_RF_bus_reg_dataout_492_port, B2 => n7802, 
                           ZN => n4050);
   U14988 : OAI22_X1 port map( A1 => n11766, A2 => n11871, B1 => 
                           DataPath_RF_bus_reg_dataout_493_port, B2 => n7802, 
                           ZN => n4048);
   U14989 : OAI22_X1 port map( A1 => n11766, A2 => n11872, B1 => 
                           DataPath_RF_bus_reg_dataout_494_port, B2 => n7802, 
                           ZN => n4046);
   U14990 : OAI22_X1 port map( A1 => n11766, A2 => n7808, B1 => 
                           DataPath_RF_bus_reg_dataout_495_port, B2 => n7802, 
                           ZN => n4044);
   U14991 : OAI22_X1 port map( A1 => n8635, A2 => n11874, B1 => 
                           DataPath_RF_bus_reg_dataout_496_port, B2 => n7802, 
                           ZN => n4042);
   U14992 : OAI22_X1 port map( A1 => n8635, A2 => n11875, B1 => 
                           DataPath_RF_bus_reg_dataout_497_port, B2 => n7802, 
                           ZN => n4040);
   U14993 : OR2_X1 port map( A1 => RST, A2 => n11755, ZN => n3339);
   U14994 : OAI22_X1 port map( A1 => n8635, A2 => n11876, B1 => 
                           DataPath_RF_bus_reg_dataout_498_port, B2 => n7802, 
                           ZN => n4038);
   U14995 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_499_port, A2 
                           => n8635, B1 => n11877, B2 => n7802, ZN => n4036);
   U14996 : OAI22_X1 port map( A1 => n11766, A2 => n11878, B1 => 
                           DataPath_RF_bus_reg_dataout_500_port, B2 => n7802, 
                           ZN => n4034);
   U14997 : OAI22_X1 port map( A1 => n8635, A2 => n11879, B1 => 
                           DataPath_RF_bus_reg_dataout_501_port, B2 => n7802, 
                           ZN => n4032);
   U14998 : OAI22_X1 port map( A1 => n8635, A2 => n11880, B1 => 
                           DataPath_RF_bus_reg_dataout_502_port, B2 => n7802, 
                           ZN => n4030);
   U14999 : OAI22_X1 port map( A1 => n11766, A2 => n11881, B1 => 
                           DataPath_RF_bus_reg_dataout_503_port, B2 => n7802, 
                           ZN => n4028);
   U15000 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_504_port, A2 
                           => n8635, B1 => n11882, B2 => n7802, ZN => n4026);
   U15001 : OAI22_X1 port map( A1 => n8635, A2 => n11883, B1 => 
                           DataPath_RF_bus_reg_dataout_505_port, B2 => n7802, 
                           ZN => n4024);
   U15002 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_506_port, A2 
                           => n11766, B1 => n11884, B2 => n7802, ZN => n4022);
   U15003 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_507_port, A2 
                           => n11766, B1 => n11885, B2 => n7802, ZN => n4020);
   U15004 : OAI22_X1 port map( A1 => n11766, A2 => n11886, B1 => 
                           DataPath_RF_bus_reg_dataout_508_port, B2 => n7802, 
                           ZN => n4018);
   U15005 : OAI22_X1 port map( A1 => n8635, A2 => n11887, B1 => 
                           DataPath_RF_bus_reg_dataout_509_port, B2 => n7802, 
                           ZN => n4016);
   U15006 : OAI22_X1 port map( A1 => n8635, A2 => n11888, B1 => 
                           DataPath_RF_bus_reg_dataout_510_port, B2 => n7802, 
                           ZN => n4014);
   U15007 : OAI22_X1 port map( A1 => n8635, A2 => n12017, B1 => 
                           DataPath_RF_bus_reg_dataout_511_port, B2 => n7802, 
                           ZN => n4010);
   U15008 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_448_port, A2 
                           => n8636, B1 => n11779, B2 => n11783, ZN => n4008);
   U15009 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_449_port, A2 
                           => n8636, B1 => n11779, B2 => n11784, ZN => n4007);
   U15010 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_450_port, A2 
                           => n8636, B1 => n11779, B2 => n11785, ZN => n4006);
   U15011 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_451_port, A2 
                           => n11780, B1 => n11779, B2 => n11767, ZN => n4005);
   U15012 : OAI22_X1 port map( A1 => n11862, A2 => n8636, B1 => 
                           DataPath_RF_bus_reg_dataout_452_port, B2 => n11774, 
                           ZN => n4004);
   U15013 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_453_port, A2 
                           => n11780, B1 => n11779, B2 => n11787, ZN => n4003);
   U15014 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_454_port, A2 
                           => n8636, B1 => n11779, B2 => n11788, ZN => n4002);
   U15015 : OAI22_X1 port map( A1 => n11865, A2 => n8636, B1 => 
                           DataPath_RF_bus_reg_dataout_455_port, B2 => n11774, 
                           ZN => n4001);
   U15016 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_456_port, A2 
                           => n8636, B1 => n11779, B2 => n11789, ZN => n4000);
   U15017 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_457_port, A2 
                           => n8636, B1 => n11779, B2 => n11790, ZN => n3999);
   U15018 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_458_port, A2 
                           => n11780, B1 => n11779, B2 => n11791, ZN => n3998);
   U15019 : OAI22_X1 port map( A1 => n11869, A2 => n8636, B1 => 
                           DataPath_RF_bus_reg_dataout_459_port, B2 => n11774, 
                           ZN => n3997);
   U15020 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_460_port, A2 
                           => n8636, B1 => n11779, B2 => n11793, ZN => n3996);
   U15021 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_461_port, A2 
                           => n8636, B1 => n11779, B2 => n11794, ZN => n3995);
   U15022 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_462_port, A2 
                           => n8636, B1 => n11779, B2 => n11795, ZN => n3994);
   U15023 : OAI22_X1 port map( A1 => n7808, A2 => n11780, B1 => 
                           DataPath_RF_bus_reg_dataout_463_port, B2 => n11774, 
                           ZN => n3993);
   U15024 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_464_port, A2 
                           => n11780, B1 => n11779, B2 => n11771, ZN => n3992);
   U15025 : OAI22_X1 port map( A1 => n11875, A2 => n8636, B1 => 
                           DataPath_RF_bus_reg_dataout_465_port, B2 => n11774, 
                           ZN => n3991);
   U15026 : OAI22_X1 port map( A1 => n11876, A2 => n8636, B1 => 
                           DataPath_RF_bus_reg_dataout_466_port, B2 => n11774, 
                           ZN => n3990);
   U15027 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_467_port, A2 
                           => n11780, B1 => n11779, B2 => n11797, ZN => n3989);
   U15028 : OAI22_X1 port map( A1 => n11878, A2 => n8636, B1 => 
                           DataPath_RF_bus_reg_dataout_468_port, B2 => n11774, 
                           ZN => n3988);
   U15029 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_469_port, A2 
                           => n8636, B1 => n11779, B2 => n11800, ZN => n3987);
   U15030 : OAI22_X1 port map( A1 => n11880, A2 => n11780, B1 => 
                           DataPath_RF_bus_reg_dataout_470_port, B2 => n11774, 
                           ZN => n3986);
   U15031 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_471_port, A2 
                           => n8636, B1 => n11779, B2 => n11803, ZN => n3985);
   U15032 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_472_port, A2 
                           => n8636, B1 => n11779, B2 => n11804, ZN => n3984);
   U15033 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_473_port, A2 
                           => n11780, B1 => n11779, B2 => n11805, ZN => n3983);
   U15034 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_474_port, A2 
                           => n8636, B1 => n11779, B2 => n11806, ZN => n3982);
   U15035 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_475_port, A2 
                           => n11780, B1 => n11779, B2 => n11807, ZN => n3981);
   U15036 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_476_port, A2 
                           => n8636, B1 => n11779, B2 => n11808, ZN => n3980);
   U15037 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_477_port, A2 
                           => n11780, B1 => n11779, B2 => n11809, ZN => n3979);
   U15038 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_478_port, A2 
                           => n8636, B1 => n11779, B2 => n11810, ZN => n3978);
   U15039 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_479_port, A2 
                           => n11780, B1 => n11779, B2 => n11811, ZN => n3975);
   U15040 : OAI22_X1 port map( A1 => n11858, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_416_port, B2 => n7803, 
                           ZN => n3973);
   U15041 : OAI22_X1 port map( A1 => n11859, A2 => n11782, B1 => 
                           DataPath_RF_bus_reg_dataout_417_port, B2 => n7803, 
                           ZN => n3972);
   U15042 : OAI22_X1 port map( A1 => n11860, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_418_port, B2 => n7803, 
                           ZN => n3971);
   U15043 : OAI22_X1 port map( A1 => n11861, A2 => n11782, B1 => 
                           DataPath_RF_bus_reg_dataout_419_port, B2 => n7803, 
                           ZN => n3970);
   U15044 : OAI22_X1 port map( A1 => n11862, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_420_port, B2 => n7803, 
                           ZN => n3969);
   U15045 : OAI22_X1 port map( A1 => n11863, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_421_port, B2 => n7803, 
                           ZN => n3968);
   U15046 : OAI22_X1 port map( A1 => n11864, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_422_port, B2 => n7803, 
                           ZN => n3967);
   U15047 : OAI22_X1 port map( A1 => n11865, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_423_port, B2 => n7803, 
                           ZN => n3966);
   U15048 : OAI22_X1 port map( A1 => n11866, A2 => n11782, B1 => 
                           DataPath_RF_bus_reg_dataout_424_port, B2 => n7803, 
                           ZN => n3965);
   U15049 : OAI22_X1 port map( A1 => n11867, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_425_port, B2 => n7803, 
                           ZN => n3964);
   U15050 : OAI22_X1 port map( A1 => n11868, A2 => n11782, B1 => 
                           DataPath_RF_bus_reg_dataout_426_port, B2 => n7803, 
                           ZN => n3963);
   U15051 : OAI22_X1 port map( A1 => n11869, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_427_port, B2 => n7803, 
                           ZN => n3962);
   U15052 : OAI22_X1 port map( A1 => n11870, A2 => n11782, B1 => 
                           DataPath_RF_bus_reg_dataout_428_port, B2 => n7803, 
                           ZN => n3961);
   U15053 : AOI22_X1 port map( A1 => n11871, A2 => n7803, B1 => n11782, B2 => 
                           DataPath_RF_bus_reg_dataout_429_port, ZN => n3960);
   U15054 : AOI22_X1 port map( A1 => n11872, A2 => n7803, B1 => n8637, B2 => 
                           DataPath_RF_bus_reg_dataout_430_port, ZN => n3959);
   U15055 : OAI22_X1 port map( A1 => n7808, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_431_port, B2 => n7803, 
                           ZN => n3958);
   U15056 : OAI22_X1 port map( A1 => n11874, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_432_port, B2 => n7803, 
                           ZN => n3957);
   U15057 : OAI22_X1 port map( A1 => n11875, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_433_port, B2 => n7803, 
                           ZN => n3956);
   U15058 : AOI22_X1 port map( A1 => n11876, A2 => n7803, B1 => n8637, B2 => 
                           DataPath_RF_bus_reg_dataout_434_port, ZN => n3955);
   U15059 : OAI22_X1 port map( A1 => n11877, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_435_port, B2 => n7803, 
                           ZN => n3954);
   U15060 : OAI22_X1 port map( A1 => n11878, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_436_port, B2 => n7803, 
                           ZN => n3953);
   U15061 : OAI22_X1 port map( A1 => n11879, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_437_port, B2 => n7803, 
                           ZN => n3952);
   U15062 : AOI22_X1 port map( A1 => n11880, A2 => n7803, B1 => n11782, B2 => 
                           DataPath_RF_bus_reg_dataout_438_port, ZN => n3951);
   U15063 : OAI22_X1 port map( A1 => n11881, A2 => n11782, B1 => 
                           DataPath_RF_bus_reg_dataout_439_port, B2 => n7803, 
                           ZN => n3950);
   U15064 : OAI22_X1 port map( A1 => n11882, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_440_port, B2 => n7803, 
                           ZN => n3949);
   U15065 : OAI22_X1 port map( A1 => n11883, A2 => n11782, B1 => 
                           DataPath_RF_bus_reg_dataout_441_port, B2 => n7803, 
                           ZN => n3948);
   U15066 : OAI22_X1 port map( A1 => n11884, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_442_port, B2 => n7803, 
                           ZN => n3947);
   U15067 : OAI22_X1 port map( A1 => n11885, A2 => n11782, B1 => 
                           DataPath_RF_bus_reg_dataout_443_port, B2 => n7803, 
                           ZN => n3946);
   U15068 : OAI22_X1 port map( A1 => n11886, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_444_port, B2 => n7803, 
                           ZN => n3945);
   U15069 : OAI22_X1 port map( A1 => n11887, A2 => n8637, B1 => 
                           DataPath_RF_bus_reg_dataout_445_port, B2 => n7803, 
                           ZN => n3944);
   U15070 : OAI22_X1 port map( A1 => n11888, A2 => n11782, B1 => 
                           DataPath_RF_bus_reg_dataout_446_port, B2 => n7803, 
                           ZN => n3943);
   U15071 : OAI22_X1 port map( A1 => n12017, A2 => n11782, B1 => 
                           DataPath_RF_bus_reg_dataout_447_port, B2 => n7803, 
                           ZN => n3940);
   U15072 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_384_port, A2 
                           => n8638, B1 => n11812, B2 => n11783, ZN => n3938);
   U15073 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_385_port, A2 
                           => n8638, B1 => n11812, B2 => n11784, ZN => n3937);
   U15074 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_386_port, A2 
                           => n8638, B1 => n11812, B2 => n11785, ZN => n3936);
   U15075 : OAI22_X1 port map( A1 => n11861, A2 => n11813, B1 => 
                           DataPath_RF_bus_reg_dataout_387_port, B2 => n11796, 
                           ZN => n3935);
   U15076 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_388_port, A2 
                           => n11813, B1 => n11812, B2 => n11786, ZN => n3934);
   U15077 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_389_port, A2 
                           => n8638, B1 => n11812, B2 => n11787, ZN => n3933);
   U15078 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_390_port, A2 
                           => n8638, B1 => n11812, B2 => n11788, ZN => n3932);
   U15079 : OAI22_X1 port map( A1 => n11865, A2 => n8638, B1 => 
                           DataPath_RF_bus_reg_dataout_391_port, B2 => n11796, 
                           ZN => n3931);
   U15080 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_392_port, A2 
                           => n8638, B1 => n11812, B2 => n11789, ZN => n3930);
   U15081 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_393_port, A2 
                           => n11813, B1 => n11812, B2 => n11790, ZN => n3929);
   U15082 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_394_port, A2 
                           => n11813, B1 => n11812, B2 => n11791, ZN => n3928);
   U15083 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_395_port, A2 
                           => n8638, B1 => n11812, B2 => n11792, ZN => n3927);
   U15084 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_396_port, A2 
                           => n8638, B1 => n11812, B2 => n11793, ZN => n3926);
   U15085 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_397_port, A2 
                           => n8638, B1 => n11812, B2 => n11794, ZN => n3925);
   U15086 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_398_port, A2 
                           => n11813, B1 => n11812, B2 => n11795, ZN => n3924);
   U15087 : OAI22_X1 port map( A1 => n7808, A2 => n8638, B1 => 
                           DataPath_RF_bus_reg_dataout_399_port, B2 => n11796, 
                           ZN => n3923);
   U15088 : OAI22_X1 port map( A1 => n11874, A2 => n8638, B1 => 
                           DataPath_RF_bus_reg_dataout_400_port, B2 => n11796, 
                           ZN => n3922);
   U15089 : OAI22_X1 port map( A1 => n11875, A2 => n11813, B1 => 
                           DataPath_RF_bus_reg_dataout_401_port, B2 => n11796, 
                           ZN => n3921);
   U15090 : OAI22_X1 port map( A1 => n11876, A2 => n8638, B1 => 
                           DataPath_RF_bus_reg_dataout_402_port, B2 => n11796, 
                           ZN => n3920);
   U15091 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_403_port, A2 
                           => n8638, B1 => n11812, B2 => n11797, ZN => n3919);
   U15092 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_404_port, A2 
                           => n8638, B1 => n11812, B2 => n11799, ZN => n3918);
   U15093 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_405_port, A2 
                           => n8638, B1 => n11812, B2 => n11800, ZN => n3917);
   U15094 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_406_port, A2 
                           => n11813, B1 => n11812, B2 => n11802, ZN => n3916);
   U15095 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_407_port, A2 
                           => n11813, B1 => n11812, B2 => n11803, ZN => n3915);
   U15096 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_408_port, A2 
                           => n8638, B1 => n11812, B2 => n11804, ZN => n3914);
   U15097 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_409_port, A2 
                           => n8638, B1 => n11812, B2 => n11805, ZN => n3913);
   U15098 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_410_port, A2 
                           => n11813, B1 => n11812, B2 => n11806, ZN => n3912);
   U15099 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_411_port, A2 
                           => n11813, B1 => n11812, B2 => n11807, ZN => n3911);
   U15100 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_412_port, A2 
                           => n11813, B1 => n11812, B2 => n11808, ZN => n3910);
   U15101 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_413_port, A2 
                           => n8638, B1 => n11812, B2 => n11809, ZN => n3909);
   U15102 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_414_port, A2 
                           => n8638, B1 => n11812, B2 => n11810, ZN => n3908);
   U15103 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_415_port, A2 
                           => n8638, B1 => n11812, B2 => n11811, ZN => n3905);
   U15104 : OAI22_X1 port map( A1 => n11858, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_352_port, B2 => n7805, 
                           ZN => n3903);
   U15105 : OAI22_X1 port map( A1 => n11859, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_353_port, B2 => n7805, 
                           ZN => n3902);
   U15106 : OAI22_X1 port map( A1 => n11860, A2 => n11815, B1 => 
                           DataPath_RF_bus_reg_dataout_354_port, B2 => n7805, 
                           ZN => n3901);
   U15107 : OAI22_X1 port map( A1 => n11861, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_355_port, B2 => n7805, 
                           ZN => n3900);
   U15108 : OAI22_X1 port map( A1 => n11862, A2 => n11815, B1 => 
                           DataPath_RF_bus_reg_dataout_356_port, B2 => n7805, 
                           ZN => n3899);
   U15109 : OAI22_X1 port map( A1 => n11863, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_357_port, B2 => n7805, 
                           ZN => n3898);
   U15110 : OAI22_X1 port map( A1 => n11864, A2 => n11815, B1 => 
                           DataPath_RF_bus_reg_dataout_358_port, B2 => n7805, 
                           ZN => n3897);
   U15111 : OAI22_X1 port map( A1 => n11865, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_359_port, B2 => n7805, 
                           ZN => n3896);
   U15112 : OAI22_X1 port map( A1 => n11866, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_360_port, B2 => n7805, 
                           ZN => n3895);
   U15113 : OAI22_X1 port map( A1 => n11867, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_361_port, B2 => n7805, 
                           ZN => n3894);
   U15114 : OAI22_X1 port map( A1 => n11868, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_362_port, B2 => n7805, 
                           ZN => n3893);
   U15115 : OAI22_X1 port map( A1 => n11869, A2 => n11815, B1 => 
                           DataPath_RF_bus_reg_dataout_363_port, B2 => n7805, 
                           ZN => n3892);
   U15116 : OAI22_X1 port map( A1 => n11870, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_364_port, B2 => n7805, 
                           ZN => n3891);
   U15117 : OAI22_X1 port map( A1 => n11871, A2 => n11815, B1 => 
                           DataPath_RF_bus_reg_dataout_365_port, B2 => n7805, 
                           ZN => n3890);
   U15118 : OAI22_X1 port map( A1 => n11872, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_366_port, B2 => n7805, 
                           ZN => n3889);
   U15119 : OAI22_X1 port map( A1 => n7808, A2 => n11815, B1 => 
                           DataPath_RF_bus_reg_dataout_367_port, B2 => n7805, 
                           ZN => n3888);
   U15120 : OAI22_X1 port map( A1 => n11874, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_368_port, B2 => n7805, 
                           ZN => n3887);
   U15121 : OAI22_X1 port map( A1 => n11875, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_369_port, B2 => n7805, 
                           ZN => n3886);
   U15122 : AOI22_X1 port map( A1 => n11876, A2 => n7805, B1 => n8639, B2 => 
                           DataPath_RF_bus_reg_dataout_370_port, ZN => n3885);
   U15123 : OAI22_X1 port map( A1 => n11877, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_371_port, B2 => n7805, 
                           ZN => n3884);
   U15124 : OAI22_X1 port map( A1 => n11878, A2 => n11815, B1 => 
                           DataPath_RF_bus_reg_dataout_372_port, B2 => n7805, 
                           ZN => n3883);
   U15125 : OAI22_X1 port map( A1 => n11879, A2 => n11815, B1 => 
                           DataPath_RF_bus_reg_dataout_373_port, B2 => n7805, 
                           ZN => n3882);
   U15126 : OAI22_X1 port map( A1 => n11880, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_374_port, B2 => n7805, 
                           ZN => n3881);
   U15127 : OAI22_X1 port map( A1 => n11881, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_375_port, B2 => n7805, 
                           ZN => n3880);
   U15128 : OAI22_X1 port map( A1 => n11882, A2 => n11815, B1 => 
                           DataPath_RF_bus_reg_dataout_376_port, B2 => n7805, 
                           ZN => n3879);
   U15129 : OAI22_X1 port map( A1 => n11883, A2 => n11815, B1 => 
                           DataPath_RF_bus_reg_dataout_377_port, B2 => n7805, 
                           ZN => n3878);
   U15130 : OAI22_X1 port map( A1 => n11884, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_378_port, B2 => n7805, 
                           ZN => n3877);
   U15131 : OAI22_X1 port map( A1 => n11885, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_379_port, B2 => n7805, 
                           ZN => n3876);
   U15132 : OAI22_X1 port map( A1 => n11886, A2 => n11815, B1 => 
                           DataPath_RF_bus_reg_dataout_380_port, B2 => n7805, 
                           ZN => n3875);
   U15133 : OAI22_X1 port map( A1 => n11887, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_381_port, B2 => n7805, 
                           ZN => n3874);
   U15134 : OAI22_X1 port map( A1 => n11888, A2 => n11815, B1 => 
                           DataPath_RF_bus_reg_dataout_382_port, B2 => n7805, 
                           ZN => n3873);
   U15135 : OAI22_X1 port map( A1 => n12017, A2 => n8639, B1 => 
                           DataPath_RF_bus_reg_dataout_383_port, B2 => n7805, 
                           ZN => n3870);
   U15136 : AOI22_X1 port map( A1 => n11818, A2 => 
                           DataPath_RF_bus_reg_dataout_320_port, B1 => n11858, 
                           B2 => n8497, ZN => n3868);
   U15137 : AOI22_X1 port map( A1 => n11818, A2 => 
                           DataPath_RF_bus_reg_dataout_321_port, B1 => n11859, 
                           B2 => n8497, ZN => n3867);
   U15138 : AOI22_X1 port map( A1 => n11818, A2 => 
                           DataPath_RF_bus_reg_dataout_322_port, B1 => n11860, 
                           B2 => n8497, ZN => n3866);
   U15139 : AOI22_X1 port map( A1 => n11818, A2 => 
                           DataPath_RF_bus_reg_dataout_323_port, B1 => n11861, 
                           B2 => n8497, ZN => n3865);
   U15140 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_324_port, B1 => n11862, 
                           B2 => n11817, ZN => n3864);
   U15141 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_325_port, B1 => n11863, 
                           B2 => n11817, ZN => n3863);
   U15142 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_326_port, B1 => n11864, 
                           B2 => n11817, ZN => n3862);
   U15143 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_327_port, B1 => n11865, 
                           B2 => n11817, ZN => n3861);
   U15144 : AOI22_X1 port map( A1 => n11818, A2 => 
                           DataPath_RF_bus_reg_dataout_328_port, B1 => n11866, 
                           B2 => n11817, ZN => n3860);
   U15145 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_329_port, B1 => n11867, 
                           B2 => n11817, ZN => n3859);
   U15146 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_330_port, B1 => n11868, 
                           B2 => n11817, ZN => n3858);
   U15147 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_331_port, B1 => n11869, 
                           B2 => n11817, ZN => n3857);
   U15148 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_332_port, B1 => n11870, 
                           B2 => n8497, ZN => n3856);
   U15149 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_333_port, B1 => n11871, 
                           B2 => n8497, ZN => n3855);
   U15150 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_334_port, B1 => n11872, 
                           B2 => n8497, ZN => n3854);
   U15151 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_335_port, B1 => n7808, 
                           B2 => n8497, ZN => n3853);
   U15152 : AOI22_X1 port map( A1 => n11818, A2 => 
                           DataPath_RF_bus_reg_dataout_336_port, B1 => n11874, 
                           B2 => n8497, ZN => n3852);
   U15153 : AOI22_X1 port map( A1 => n11818, A2 => 
                           DataPath_RF_bus_reg_dataout_337_port, B1 => n11875, 
                           B2 => n8497, ZN => n3851);
   U15154 : AOI22_X1 port map( A1 => n11818, A2 => 
                           DataPath_RF_bus_reg_dataout_338_port, B1 => n11876, 
                           B2 => n8497, ZN => n3850);
   U15155 : AOI22_X1 port map( A1 => n11818, A2 => 
                           DataPath_RF_bus_reg_dataout_339_port, B1 => n11877, 
                           B2 => n8497, ZN => n3849);
   U15156 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_340_port, B1 => n11878, 
                           B2 => n8497, ZN => n3848);
   U15157 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_341_port, B1 => n11879, 
                           B2 => n8497, ZN => n3847);
   U15158 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_342_port, B1 => n11880, 
                           B2 => n8497, ZN => n3846);
   U15159 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_343_port, B1 => n11881, 
                           B2 => n8497, ZN => n3845);
   U15160 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_344_port, B1 => n11882, 
                           B2 => n8497, ZN => n3844);
   U15161 : AOI22_X1 port map( A1 => n11818, A2 => 
                           DataPath_RF_bus_reg_dataout_345_port, B1 => n11883, 
                           B2 => n11817, ZN => n3843);
   U15162 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_346_port, B1 => n11884, 
                           B2 => n8497, ZN => n3842);
   U15163 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_347_port, B1 => n11885, 
                           B2 => n11817, ZN => n3841);
   U15164 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_348_port, B1 => n11886, 
                           B2 => n8497, ZN => n3840);
   U15165 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_349_port, B1 => n11887, 
                           B2 => n8497, ZN => n3839);
   U15166 : AOI22_X1 port map( A1 => n11818, A2 => 
                           DataPath_RF_bus_reg_dataout_350_port, B1 => n11888, 
                           B2 => n11817, ZN => n3838);
   U15167 : AOI22_X1 port map( A1 => n8640, A2 => 
                           DataPath_RF_bus_reg_dataout_351_port, B1 => n12017, 
                           B2 => n8497, ZN => n3835);
   U15168 : AOI22_X1 port map( A1 => n11858, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_288_port, ZN => n3833);
   U15169 : AOI22_X1 port map( A1 => n11859, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_289_port, ZN => n3832);
   U15170 : AOI22_X1 port map( A1 => n11860, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_290_port, ZN => n3831);
   U15171 : AOI22_X1 port map( A1 => n11861, A2 => n7804, B1 => n11819, B2 => 
                           DataPath_RF_bus_reg_dataout_291_port, ZN => n3830);
   U15172 : AOI22_X1 port map( A1 => n11862, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_292_port, ZN => n3829);
   U15173 : AOI22_X1 port map( A1 => n11863, A2 => n7804, B1 => n11819, B2 => 
                           DataPath_RF_bus_reg_dataout_293_port, ZN => n3828);
   U15174 : AOI22_X1 port map( A1 => n11864, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_294_port, ZN => n3827);
   U15175 : AOI22_X1 port map( A1 => n11865, A2 => n7804, B1 => n11819, B2 => 
                           DataPath_RF_bus_reg_dataout_295_port, ZN => n3826);
   U15176 : AOI22_X1 port map( A1 => n11866, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_296_port, ZN => n3825);
   U15177 : AOI22_X1 port map( A1 => n11867, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_297_port, ZN => n3824);
   U15178 : AOI22_X1 port map( A1 => n11868, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_298_port, ZN => n3823);
   U15179 : AOI22_X1 port map( A1 => n11869, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_299_port, ZN => n3822);
   U15180 : AOI22_X1 port map( A1 => n11870, A2 => n7804, B1 => n11819, B2 => 
                           DataPath_RF_bus_reg_dataout_300_port, ZN => n3821);
   U15181 : AOI22_X1 port map( A1 => n11871, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_301_port, ZN => n3820);
   U15182 : AOI22_X1 port map( A1 => n11872, A2 => n7804, B1 => n11819, B2 => 
                           DataPath_RF_bus_reg_dataout_302_port, ZN => n3819);
   U15183 : AOI22_X1 port map( A1 => n7808, A2 => n7804, B1 => n11819, B2 => 
                           DataPath_RF_bus_reg_dataout_303_port, ZN => n3818);
   U15184 : AOI22_X1 port map( A1 => n11874, A2 => n7804, B1 => n11819, B2 => 
                           DataPath_RF_bus_reg_dataout_304_port, ZN => n3817);
   U15185 : AOI22_X1 port map( A1 => n11875, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_305_port, ZN => n3816);
   U15186 : OAI22_X1 port map( A1 => n11876, A2 => n8641, B1 => 
                           DataPath_RF_bus_reg_dataout_306_port, B2 => n7804, 
                           ZN => n3815);
   U15187 : AOI22_X1 port map( A1 => n11877, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_307_port, ZN => n3814);
   U15188 : AOI22_X1 port map( A1 => n11878, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_308_port, ZN => n3813);
   U15189 : AOI22_X1 port map( A1 => n11879, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_309_port, ZN => n3812);
   U15190 : AOI22_X1 port map( A1 => n11880, A2 => n7804, B1 => n11819, B2 => 
                           DataPath_RF_bus_reg_dataout_310_port, ZN => n3811);
   U15191 : AOI22_X1 port map( A1 => n11881, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_311_port, ZN => n3810);
   U15192 : AOI22_X1 port map( A1 => n11882, A2 => n7804, B1 => n11819, B2 => 
                           DataPath_RF_bus_reg_dataout_312_port, ZN => n3809);
   U15193 : AOI22_X1 port map( A1 => n11883, A2 => n7804, B1 => n11819, B2 => 
                           DataPath_RF_bus_reg_dataout_313_port, ZN => n3808);
   U15194 : AOI22_X1 port map( A1 => n11884, A2 => n7804, B1 => n11819, B2 => 
                           DataPath_RF_bus_reg_dataout_314_port, ZN => n3807);
   U15195 : AOI22_X1 port map( A1 => n11885, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_315_port, ZN => n3806);
   U15196 : AOI22_X1 port map( A1 => n11886, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_316_port, ZN => n3805);
   U15197 : AOI22_X1 port map( A1 => n11887, A2 => n7804, B1 => n11819, B2 => 
                           DataPath_RF_bus_reg_dataout_317_port, ZN => n3804);
   U15198 : AOI22_X1 port map( A1 => n11888, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_318_port, ZN => n3803);
   U15199 : AOI22_X1 port map( A1 => n12017, A2 => n7804, B1 => n8641, B2 => 
                           DataPath_RF_bus_reg_dataout_319_port, ZN => n3800);
   U15200 : OAI22_X1 port map( A1 => n11858, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_256_port, B2 => n7806, 
                           ZN => n3798);
   U15201 : OAI22_X1 port map( A1 => n11859, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_257_port, B2 => n7806, 
                           ZN => n3797);
   U15202 : OAI22_X1 port map( A1 => n11860, A2 => n11822, B1 => 
                           DataPath_RF_bus_reg_dataout_258_port, B2 => n7806, 
                           ZN => n3796);
   U15203 : OAI22_X1 port map( A1 => n11861, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_259_port, B2 => n7806, 
                           ZN => n3795);
   U15204 : OAI22_X1 port map( A1 => n11862, A2 => n11822, B1 => 
                           DataPath_RF_bus_reg_dataout_260_port, B2 => n7806, 
                           ZN => n3794);
   U15205 : OAI22_X1 port map( A1 => n11863, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_261_port, B2 => n7806, 
                           ZN => n3793);
   U15206 : OAI22_X1 port map( A1 => n11864, A2 => n11822, B1 => 
                           DataPath_RF_bus_reg_dataout_262_port, B2 => n7806, 
                           ZN => n3792);
   U15207 : OAI22_X1 port map( A1 => n11865, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_263_port, B2 => n7806, 
                           ZN => n3791);
   U15208 : OAI22_X1 port map( A1 => n11866, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_264_port, B2 => n7806, 
                           ZN => n3790);
   U15209 : OAI22_X1 port map( A1 => n11867, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_265_port, B2 => n7806, 
                           ZN => n3789);
   U15210 : OAI22_X1 port map( A1 => n11868, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_266_port, B2 => n7806, 
                           ZN => n3788);
   U15211 : OAI22_X1 port map( A1 => n11869, A2 => n11822, B1 => 
                           DataPath_RF_bus_reg_dataout_267_port, B2 => n7806, 
                           ZN => n3787);
   U15212 : OAI22_X1 port map( A1 => n11870, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_268_port, B2 => n7806, 
                           ZN => n3786);
   U15213 : OAI22_X1 port map( A1 => n11871, A2 => n11822, B1 => 
                           DataPath_RF_bus_reg_dataout_269_port, B2 => n7806, 
                           ZN => n3785);
   U15214 : OAI22_X1 port map( A1 => n11872, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_270_port, B2 => n7806, 
                           ZN => n3784);
   U15215 : OAI22_X1 port map( A1 => n7808, A2 => n11822, B1 => 
                           DataPath_RF_bus_reg_dataout_271_port, B2 => n7806, 
                           ZN => n3783);
   U15216 : OAI22_X1 port map( A1 => n11874, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_272_port, B2 => n7806, 
                           ZN => n3782);
   U15217 : OAI22_X1 port map( A1 => n11875, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_273_port, B2 => n7806, 
                           ZN => n3781);
   U15218 : AOI22_X1 port map( A1 => n11876, A2 => n7806, B1 => n8642, B2 => 
                           DataPath_RF_bus_reg_dataout_274_port, ZN => n3780);
   U15219 : OAI22_X1 port map( A1 => n11877, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_275_port, B2 => n7806, 
                           ZN => n3779);
   U15220 : OAI22_X1 port map( A1 => n11878, A2 => n11822, B1 => 
                           DataPath_RF_bus_reg_dataout_276_port, B2 => n7806, 
                           ZN => n3778);
   U15221 : OAI22_X1 port map( A1 => n11879, A2 => n11822, B1 => 
                           DataPath_RF_bus_reg_dataout_277_port, B2 => n7806, 
                           ZN => n3777);
   U15222 : OAI22_X1 port map( A1 => n11880, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_278_port, B2 => n7806, 
                           ZN => n3776);
   U15223 : OAI22_X1 port map( A1 => n11881, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_279_port, B2 => n7806, 
                           ZN => n3775);
   U15224 : OAI22_X1 port map( A1 => n11882, A2 => n11822, B1 => 
                           DataPath_RF_bus_reg_dataout_280_port, B2 => n7806, 
                           ZN => n3774);
   U15225 : OAI22_X1 port map( A1 => n11883, A2 => n11822, B1 => 
                           DataPath_RF_bus_reg_dataout_281_port, B2 => n7806, 
                           ZN => n3773);
   U15226 : OAI22_X1 port map( A1 => n11884, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_282_port, B2 => n7806, 
                           ZN => n3772);
   U15227 : OAI22_X1 port map( A1 => n11885, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_283_port, B2 => n7806, 
                           ZN => n3771);
   U15228 : OAI22_X1 port map( A1 => n11886, A2 => n11822, B1 => 
                           DataPath_RF_bus_reg_dataout_284_port, B2 => n7806, 
                           ZN => n3770);
   U15229 : OAI22_X1 port map( A1 => n11887, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_285_port, B2 => n7806, 
                           ZN => n3769);
   U15230 : OAI22_X1 port map( A1 => n11888, A2 => n11822, B1 => 
                           DataPath_RF_bus_reg_dataout_286_port, B2 => n7806, 
                           ZN => n3768);
   U15231 : OAI22_X1 port map( A1 => n12017, A2 => n8642, B1 => 
                           DataPath_RF_bus_reg_dataout_287_port, B2 => n7806, 
                           ZN => n3765);
   U15232 : OAI22_X1 port map( A1 => n8441, A2 => n11824, B1 => n8299, B2 => 
                           n11823, ZN => n11825);
   U15233 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_224_port, B1 => n11858, 
                           B2 => n11826, ZN => n3760);
   U15234 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_225_port, B1 => n11859, 
                           B2 => n11826, ZN => n3759);
   U15235 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_226_port, B1 => n11860, 
                           B2 => n11826, ZN => n3758);
   U15236 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_227_port, B1 => n11861, 
                           B2 => n11826, ZN => n3757);
   U15237 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_228_port, B1 => n11862, 
                           B2 => n11826, ZN => n3756);
   U15238 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_229_port, B1 => n11863, 
                           B2 => n11826, ZN => n3755);
   U15239 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_230_port, B1 => n11864, 
                           B2 => n11826, ZN => n3754);
   U15240 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_231_port, B1 => n11865, 
                           B2 => n11826, ZN => n3753);
   U15241 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_232_port, B1 => n11866, 
                           B2 => n11826, ZN => n3752);
   U15242 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_233_port, B1 => n11867, 
                           B2 => n11826, ZN => n3751);
   U15243 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_234_port, B1 => n11868, 
                           B2 => n11826, ZN => n3750);
   U15244 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_235_port, B1 => n11869, 
                           B2 => n11826, ZN => n3749);
   U15245 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_236_port, B1 => n11870, 
                           B2 => n11826, ZN => n3748);
   U15246 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_237_port, B1 => n11871, 
                           B2 => n11826, ZN => n3747);
   U15247 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_238_port, B1 => n11872, 
                           B2 => n11826, ZN => n3746);
   U15248 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_239_port, B1 => n7808, 
                           B2 => n11826, ZN => n3745);
   U15249 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_240_port, B1 => n11874, 
                           B2 => n11826, ZN => n3744);
   U15250 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_241_port, B1 => n11875, 
                           B2 => n11826, ZN => n3743);
   U15251 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_242_port, B1 => n11876, 
                           B2 => n11826, ZN => n3742);
   U15252 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_243_port, B1 => n11877, 
                           B2 => n11826, ZN => n3741);
   U15253 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_244_port, B1 => n11878, 
                           B2 => n11826, ZN => n3740);
   U15254 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_245_port, B1 => n11879, 
                           B2 => n11826, ZN => n3739);
   U15255 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_246_port, B1 => n11880, 
                           B2 => n11826, ZN => n3738);
   U15256 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_247_port, B1 => n11881, 
                           B2 => n11826, ZN => n3737);
   U15257 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_248_port, B1 => n11882, 
                           B2 => n11826, ZN => n3736);
   U15258 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_249_port, B1 => n11883, 
                           B2 => n11826, ZN => n3735);
   U15259 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_250_port, B1 => n11884, 
                           B2 => n11826, ZN => n3734);
   U15260 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_251_port, B1 => n11885, 
                           B2 => n11826, ZN => n3733);
   U15261 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_252_port, B1 => n11886, 
                           B2 => n11826, ZN => n3732);
   U15262 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_253_port, B1 => n11887, 
                           B2 => n11826, ZN => n3731);
   U15263 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_254_port, B1 => n11888, 
                           B2 => n11826, ZN => n3730);
   U15264 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_255_port, B1 => n12017, 
                           B2 => n11826, ZN => n3727);
   U15265 : OAI22_X1 port map( A1 => n8441, A2 => n11829, B1 => n8299, B2 => 
                           n11828, ZN => n11830);
   U15266 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_192_port, B1 => n11858, 
                           B2 => n11831, ZN => n3722);
   U15267 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_193_port, B1 => n11859, 
                           B2 => n11831, ZN => n3721);
   U15268 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_194_port, B1 => n11860, 
                           B2 => n11831, ZN => n3720);
   U15269 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_195_port, B1 => n11861, 
                           B2 => n11831, ZN => n3719);
   U15270 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_196_port, B1 => n11862, 
                           B2 => n11831, ZN => n3718);
   U15271 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_197_port, B1 => n11863, 
                           B2 => n11831, ZN => n3717);
   U15272 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_198_port, B1 => n11864, 
                           B2 => n11831, ZN => n3716);
   U15273 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_199_port, B1 => n11865, 
                           B2 => n11831, ZN => n3715);
   U15274 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_200_port, B1 => n11866, 
                           B2 => n11831, ZN => n3714);
   U15275 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_201_port, B1 => n11867, 
                           B2 => n11831, ZN => n3713);
   U15276 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_202_port, B1 => n11868, 
                           B2 => n11831, ZN => n3712);
   U15277 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_203_port, B1 => n11869, 
                           B2 => n11831, ZN => n3711);
   U15278 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_204_port, B1 => n11870, 
                           B2 => n11831, ZN => n3710);
   U15279 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_205_port, B1 => n11871, 
                           B2 => n11831, ZN => n3709);
   U15280 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_206_port, B1 => n11872, 
                           B2 => n11831, ZN => n3708);
   U15281 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_207_port, B1 => n7808, 
                           B2 => n11831, ZN => n3707);
   U15282 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_208_port, B1 => n11874, 
                           B2 => n11831, ZN => n3706);
   U15283 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_209_port, B1 => n11875, 
                           B2 => n11831, ZN => n3705);
   U15284 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_210_port, B1 => n11876, 
                           B2 => n11831, ZN => n3704);
   U15285 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_211_port, B1 => n11877, 
                           B2 => n11831, ZN => n3703);
   U15286 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_212_port, B1 => n11878, 
                           B2 => n11831, ZN => n3702);
   U15287 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_213_port, B1 => n11879, 
                           B2 => n11831, ZN => n3701);
   U15288 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_214_port, B1 => n11880, 
                           B2 => n11831, ZN => n3700);
   U15289 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_215_port, B1 => n11881, 
                           B2 => n11831, ZN => n3699);
   U15290 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_216_port, B1 => n11882, 
                           B2 => n11831, ZN => n3698);
   U15291 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_217_port, B1 => n11883, 
                           B2 => n11831, ZN => n3697);
   U15292 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_218_port, B1 => n11884, 
                           B2 => n11831, ZN => n3696);
   U15293 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_219_port, B1 => n11885, 
                           B2 => n11831, ZN => n3695);
   U15294 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_220_port, B1 => n11886, 
                           B2 => n11831, ZN => n3694);
   U15295 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_221_port, B1 => n11887, 
                           B2 => n11831, ZN => n3693);
   U15296 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_222_port, B1 => n11888, 
                           B2 => n11831, ZN => n3692);
   U15297 : AOI22_X1 port map( A1 => n8546, A2 => 
                           DataPath_RF_bus_reg_dataout_223_port, B1 => n12017, 
                           B2 => n11831, ZN => n3689);
   U15298 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_160_port, B1 => n11858, 
                           B2 => n11836, ZN => n3684);
   U15299 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_161_port, B1 => n11859, 
                           B2 => n11836, ZN => n3683);
   U15300 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_162_port, B1 => n11860, 
                           B2 => n11836, ZN => n3682);
   U15301 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_163_port, B1 => n11861, 
                           B2 => n11836, ZN => n3681);
   U15302 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_164_port, B1 => n11862, 
                           B2 => n11836, ZN => n3680);
   U15303 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_165_port, B1 => n11863, 
                           B2 => n11836, ZN => n3679);
   U15304 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_166_port, B1 => n11864, 
                           B2 => n11836, ZN => n3678);
   U15305 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_167_port, B1 => n11865, 
                           B2 => n11836, ZN => n3677);
   U15306 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_168_port, B1 => n11866, 
                           B2 => n11836, ZN => n3676);
   U15307 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_169_port, B1 => n11867, 
                           B2 => n11836, ZN => n3675);
   U15308 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_170_port, B1 => n11868, 
                           B2 => n11836, ZN => n3674);
   U15309 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_171_port, B1 => n11869, 
                           B2 => n11836, ZN => n3673);
   U15310 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_172_port, B1 => n11870, 
                           B2 => n11836, ZN => n3672);
   U15311 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_173_port, B1 => n11871, 
                           B2 => n11836, ZN => n3671);
   U15312 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_174_port, B1 => n11872, 
                           B2 => n11836, ZN => n3670);
   U15313 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_175_port, B1 => n7808, 
                           B2 => n11836, ZN => n3669);
   U15314 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_176_port, B1 => n11874, 
                           B2 => n11836, ZN => n3668);
   U15315 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_177_port, B1 => n11875, 
                           B2 => n11836, ZN => n3667);
   U15316 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_178_port, B1 => n11876, 
                           B2 => n11836, ZN => n3666);
   U15317 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_179_port, B1 => n11877, 
                           B2 => n11836, ZN => n3665);
   U15318 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_180_port, B1 => n11878, 
                           B2 => n11836, ZN => n3664);
   U15319 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_181_port, B1 => n11879, 
                           B2 => n11836, ZN => n3663);
   U15320 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_182_port, B1 => n11880, 
                           B2 => n11836, ZN => n3662);
   U15321 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_183_port, B1 => n11881, 
                           B2 => n11836, ZN => n3661);
   U15322 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_184_port, B1 => n11882, 
                           B2 => n11836, ZN => n3660);
   U15323 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_185_port, B1 => n11883, 
                           B2 => n11836, ZN => n3659);
   U15324 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_186_port, B1 => n11884, 
                           B2 => n11836, ZN => n3658);
   U15325 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_187_port, B1 => n11885, 
                           B2 => n11836, ZN => n3657);
   U15326 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_188_port, B1 => n11886, 
                           B2 => n11836, ZN => n3656);
   U15327 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_189_port, B1 => n11887, 
                           B2 => n11836, ZN => n3655);
   U15328 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_190_port, B1 => n11888, 
                           B2 => n11836, ZN => n3654);
   U15329 : AOI22_X1 port map( A1 => n11837, A2 => 
                           DataPath_RF_bus_reg_dataout_191_port, B1 => n12017, 
                           B2 => n11836, ZN => n3651);
   U15330 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_128_port, B1 => n11858, 
                           B2 => n11840, ZN => n3646);
   U15331 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_129_port, B1 => n11859, 
                           B2 => n11840, ZN => n3645);
   U15332 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_130_port, B1 => n11860, 
                           B2 => n11840, ZN => n3644);
   U15333 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_131_port, B1 => n11861, 
                           B2 => n11840, ZN => n3643);
   U15334 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_132_port, B1 => n11862, 
                           B2 => n11840, ZN => n3642);
   U15335 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_133_port, B1 => n11863, 
                           B2 => n11840, ZN => n3641);
   U15336 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_134_port, B1 => n11864, 
                           B2 => n11840, ZN => n3640);
   U15337 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_135_port, B1 => n11865, 
                           B2 => n11840, ZN => n3639);
   U15338 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_136_port, B1 => n11866, 
                           B2 => n11840, ZN => n3638);
   U15339 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_137_port, B1 => n11867, 
                           B2 => n11840, ZN => n3637);
   U15340 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_138_port, B1 => n11868, 
                           B2 => n11840, ZN => n3636);
   U15341 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_139_port, B1 => n11869, 
                           B2 => n11840, ZN => n3635);
   U15342 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_140_port, B1 => n11870, 
                           B2 => n11840, ZN => n3634);
   U15343 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_141_port, B1 => n11871, 
                           B2 => n11840, ZN => n3633);
   U15344 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_142_port, B1 => n11872, 
                           B2 => n11840, ZN => n3632);
   U15345 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_143_port, B1 => n7808, 
                           B2 => n11840, ZN => n3631);
   U15346 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_144_port, B1 => n11874, 
                           B2 => n11840, ZN => n3630);
   U15347 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_145_port, B1 => n11875, 
                           B2 => n11840, ZN => n3629);
   U15348 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_146_port, B1 => n11876, 
                           B2 => n11840, ZN => n3628);
   U15349 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_147_port, B1 => n11877, 
                           B2 => n11840, ZN => n3627);
   U15350 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_148_port, B1 => n11878, 
                           B2 => n11840, ZN => n3626);
   U15351 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_149_port, B1 => n11879, 
                           B2 => n11840, ZN => n3625);
   U15352 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_150_port, B1 => n11880, 
                           B2 => n11840, ZN => n3624);
   U15353 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_151_port, B1 => n11881, 
                           B2 => n11840, ZN => n3623);
   U15354 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_152_port, B1 => n11882, 
                           B2 => n11840, ZN => n3622);
   U15355 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_153_port, B1 => n11883, 
                           B2 => n11840, ZN => n3621);
   U15356 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_154_port, B1 => n11884, 
                           B2 => n11840, ZN => n3620);
   U15357 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_155_port, B1 => n11885, 
                           B2 => n11840, ZN => n3619);
   U15358 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_156_port, B1 => n11886, 
                           B2 => n11840, ZN => n3618);
   U15359 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_157_port, B1 => n11887, 
                           B2 => n11840, ZN => n3617);
   U15360 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_158_port, B1 => n11888, 
                           B2 => n11840, ZN => n3616);
   U15361 : AOI22_X1 port map( A1 => n8547, A2 => 
                           DataPath_RF_bus_reg_dataout_159_port, B1 => n12017, 
                           B2 => n11840, ZN => n3613);
   U15362 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_96_port, B1 => n11858, 
                           B2 => n11845, ZN => n3608);
   U15363 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_97_port, B1 => n11859, 
                           B2 => n11845, ZN => n3607);
   U15364 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_98_port, B1 => n11860, 
                           B2 => n11845, ZN => n3606);
   U15365 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_99_port, B1 => n11861, 
                           B2 => n11845, ZN => n3605);
   U15366 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_100_port, B1 => n11862, 
                           B2 => n11845, ZN => n3604);
   U15367 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_101_port, B1 => n11863, 
                           B2 => n11845, ZN => n3603);
   U15368 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_102_port, B1 => n11864, 
                           B2 => n11845, ZN => n3602);
   U15369 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_103_port, B1 => n11865, 
                           B2 => n11845, ZN => n3601);
   U15370 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_104_port, B1 => n11866, 
                           B2 => n11845, ZN => n3600);
   U15371 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_105_port, B1 => n11867, 
                           B2 => n11845, ZN => n3599);
   U15372 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_106_port, B1 => n11868, 
                           B2 => n11845, ZN => n3598);
   U15373 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_107_port, B1 => n11869, 
                           B2 => n11845, ZN => n3597);
   U15374 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_108_port, B1 => n11870, 
                           B2 => n11845, ZN => n3596);
   U15375 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_109_port, B1 => n11871, 
                           B2 => n11845, ZN => n3595);
   U15376 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_110_port, B1 => n11872, 
                           B2 => n11845, ZN => n3594);
   U15377 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_111_port, B1 => n7808, 
                           B2 => n11845, ZN => n3593);
   U15378 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_112_port, B1 => n11874, 
                           B2 => n11845, ZN => n3592);
   U15379 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_113_port, B1 => n11875, 
                           B2 => n11845, ZN => n3591);
   U15380 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_114_port, B1 => n11876, 
                           B2 => n11845, ZN => n3590);
   U15381 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_115_port, B1 => n11877, 
                           B2 => n11845, ZN => n3589);
   U15382 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_116_port, B1 => n11878, 
                           B2 => n11845, ZN => n3588);
   U15383 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_117_port, B1 => n11879, 
                           B2 => n11845, ZN => n3587);
   U15384 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_118_port, B1 => n11880, 
                           B2 => n11845, ZN => n3586);
   U15385 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_119_port, B1 => n11881, 
                           B2 => n11845, ZN => n3585);
   U15386 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_120_port, B1 => n11882, 
                           B2 => n11845, ZN => n3584);
   U15387 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_121_port, B1 => n11883, 
                           B2 => n11845, ZN => n3583);
   U15388 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_122_port, B1 => n11884, 
                           B2 => n11845, ZN => n3582);
   U15389 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_123_port, B1 => n11885, 
                           B2 => n11845, ZN => n3581);
   U15390 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_124_port, B1 => n11886, 
                           B2 => n11845, ZN => n3580);
   U15391 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_125_port, B1 => n11887, 
                           B2 => n11845, ZN => n3579);
   U15392 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_126_port, B1 => n11888, 
                           B2 => n11845, ZN => n3578);
   U15393 : AOI22_X1 port map( A1 => n11846, A2 => 
                           DataPath_RF_bus_reg_dataout_127_port, B1 => n12017, 
                           B2 => n11845, ZN => n3575);
   U15394 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_64_port, B1 => n11858, 
                           B2 => n11849, ZN => n3570);
   U15395 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_65_port, B1 => n11859, 
                           B2 => n11849, ZN => n3569);
   U15396 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_66_port, B1 => n11860, 
                           B2 => n11849, ZN => n3568);
   U15397 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_67_port, B1 => n11861, 
                           B2 => n11849, ZN => n3567);
   U15398 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_68_port, B1 => n11862, 
                           B2 => n11849, ZN => n3566);
   U15399 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_69_port, B1 => n11863, 
                           B2 => n11849, ZN => n3565);
   U15400 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_70_port, B1 => n11864, 
                           B2 => n11849, ZN => n3564);
   U15401 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_71_port, B1 => n11865, 
                           B2 => n11849, ZN => n3563);
   U15402 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_72_port, B1 => n11866, 
                           B2 => n11849, ZN => n3562);
   U15403 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_73_port, B1 => n11867, 
                           B2 => n11849, ZN => n3561);
   U15404 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_74_port, B1 => n11868, 
                           B2 => n11849, ZN => n3560);
   U15405 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_75_port, B1 => n11869, 
                           B2 => n11849, ZN => n3559);
   U15406 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_76_port, B1 => n11870, 
                           B2 => n11849, ZN => n3558);
   U15407 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_77_port, B1 => n11871, 
                           B2 => n11849, ZN => n3557);
   U15408 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_78_port, B1 => n11872, 
                           B2 => n11849, ZN => n3556);
   U15409 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_79_port, B1 => n7808, B2
                           => n11849, ZN => n3555);
   U15410 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_80_port, B1 => n11874, 
                           B2 => n11849, ZN => n3554);
   U15411 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_81_port, B1 => n11875, 
                           B2 => n11849, ZN => n3553);
   U15412 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_82_port, B1 => n11876, 
                           B2 => n11849, ZN => n3552);
   U15413 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_83_port, B1 => n11877, 
                           B2 => n11849, ZN => n3551);
   U15414 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_84_port, B1 => n11878, 
                           B2 => n11849, ZN => n3550);
   U15415 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_85_port, B1 => n11879, 
                           B2 => n11849, ZN => n3549);
   U15416 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_86_port, B1 => n11880, 
                           B2 => n11849, ZN => n3548);
   U15417 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_87_port, B1 => n11881, 
                           B2 => n11849, ZN => n3547);
   U15418 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_88_port, B1 => n11882, 
                           B2 => n11849, ZN => n3546);
   U15419 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_89_port, B1 => n11883, 
                           B2 => n11849, ZN => n3545);
   U15420 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_90_port, B1 => n11884, 
                           B2 => n11849, ZN => n3544);
   U15421 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_91_port, B1 => n11885, 
                           B2 => n11849, ZN => n3543);
   U15422 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_92_port, B1 => n11886, 
                           B2 => n11849, ZN => n3542);
   U15423 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_93_port, B1 => n11887, 
                           B2 => n11849, ZN => n3541);
   U15424 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_94_port, B1 => n11888, 
                           B2 => n11849, ZN => n3540);
   U15425 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_95_port, B1 => n12017, 
                           B2 => n11849, ZN => n3537);
   U15426 : OAI22_X1 port map( A1 => n8441, A2 => n11852, B1 => n8299, B2 => 
                           n11851, ZN => n11853);
   U15427 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_32_port, B1 => n11858, 
                           B2 => n8644, ZN => n3532);
   U15428 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_33_port, B1 => n11859, 
                           B2 => n8644, ZN => n3531);
   U15429 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_34_port, B1 => n11860, 
                           B2 => n8644, ZN => n3530);
   U15430 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_35_port, B1 => n11861, 
                           B2 => n8644, ZN => n3529);
   U15431 : AOI22_X1 port map( A1 => n11854, A2 => 
                           DataPath_RF_bus_reg_dataout_36_port, B1 => n11862, 
                           B2 => n8644, ZN => n3528);
   U15432 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_37_port, B1 => n11863, 
                           B2 => n8644, ZN => n3527);
   U15433 : AOI22_X1 port map( A1 => n11854, A2 => 
                           DataPath_RF_bus_reg_dataout_38_port, B1 => n11864, 
                           B2 => n8644, ZN => n3526);
   U15434 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_39_port, B1 => n11865, 
                           B2 => n8644, ZN => n3525);
   U15435 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_40_port, B1 => n11866, 
                           B2 => n8644, ZN => n3524);
   U15436 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_41_port, B1 => n11867, 
                           B2 => n8644, ZN => n3523);
   U15437 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_42_port, B1 => n11868, 
                           B2 => n8644, ZN => n3522);
   U15438 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_43_port, B1 => n11869, 
                           B2 => n8644, ZN => n3521);
   U15439 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_44_port, B1 => n11870, 
                           B2 => n8644, ZN => n3520);
   U15440 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_45_port, B1 => n11871, 
                           B2 => n8644, ZN => n3519);
   U15441 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_46_port, B1 => n11872, 
                           B2 => n8644, ZN => n3518);
   U15442 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_47_port, B1 => n7808, B2
                           => n8644, ZN => n3517);
   U15443 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_48_port, B1 => n11874, 
                           B2 => n8644, ZN => n3516);
   U15444 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_49_port, B1 => n11875, 
                           B2 => n8644, ZN => n3515);
   U15445 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_50_port, B1 => n11876, 
                           B2 => n8644, ZN => n3514);
   U15446 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_51_port, B1 => n11877, 
                           B2 => n8644, ZN => n3513);
   U15447 : AOI22_X1 port map( A1 => n11854, A2 => 
                           DataPath_RF_bus_reg_dataout_52_port, B1 => n11878, 
                           B2 => n8644, ZN => n3512);
   U15448 : AOI22_X1 port map( A1 => n11854, A2 => 
                           DataPath_RF_bus_reg_dataout_53_port, B1 => n11879, 
                           B2 => n8644, ZN => n3511);
   U15449 : AOI22_X1 port map( A1 => n11854, A2 => 
                           DataPath_RF_bus_reg_dataout_54_port, B1 => n11880, 
                           B2 => n8644, ZN => n3510);
   U15450 : AOI22_X1 port map( A1 => n11854, A2 => 
                           DataPath_RF_bus_reg_dataout_55_port, B1 => n11881, 
                           B2 => n8644, ZN => n3509);
   U15451 : AOI22_X1 port map( A1 => n11854, A2 => 
                           DataPath_RF_bus_reg_dataout_56_port, B1 => n11882, 
                           B2 => n8644, ZN => n3508);
   U15452 : AOI22_X1 port map( A1 => n11854, A2 => 
                           DataPath_RF_bus_reg_dataout_57_port, B1 => n11883, 
                           B2 => n8644, ZN => n3507);
   U15453 : AOI22_X1 port map( A1 => n11854, A2 => 
                           DataPath_RF_bus_reg_dataout_58_port, B1 => n11884, 
                           B2 => n8644, ZN => n3506);
   U15454 : AOI22_X1 port map( A1 => n11854, A2 => 
                           DataPath_RF_bus_reg_dataout_59_port, B1 => n11885, 
                           B2 => n8644, ZN => n3505);
   U15455 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_60_port, B1 => n11886, 
                           B2 => n8644, ZN => n3504);
   U15456 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_61_port, B1 => n11887, 
                           B2 => n8644, ZN => n3503);
   U15457 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_62_port, B1 => n11888, 
                           B2 => n8644, ZN => n3502);
   U15458 : AOI22_X1 port map( A1 => n8643, A2 => 
                           DataPath_RF_bus_reg_dataout_63_port, B1 => n12017, 
                           B2 => n8644, ZN => n3499);
   U15459 : OAI22_X1 port map( A1 => n8441, A2 => n11856, B1 => n8299, B2 => 
                           n11855, ZN => n11857);
   U15460 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_0_port, B1 => n11858, B2
                           => n8653, ZN => n3492);
   U15461 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_1_port, B1 => n11859, B2
                           => n8653, ZN => n3490);
   U15462 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_2_port, B1 => n11860, B2
                           => n8653, ZN => n3488);
   U15463 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_3_port, B1 => n11861, B2
                           => n8653, ZN => n3486);
   U15464 : AOI22_X1 port map( A1 => n12018, A2 => 
                           DataPath_RF_bus_reg_dataout_4_port, B1 => n11862, B2
                           => n8653, ZN => n3484);
   U15465 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_5_port, B1 => n11863, B2
                           => n8653, ZN => n3482);
   U15466 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_6_port, B1 => n11864, B2
                           => n8653, ZN => n3480);
   U15467 : AOI22_X1 port map( A1 => n12018, A2 => 
                           DataPath_RF_bus_reg_dataout_7_port, B1 => n11865, B2
                           => n8653, ZN => n3478);
   U15468 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_8_port, B1 => n11866, B2
                           => n8653, ZN => n3476);
   U15469 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_9_port, B1 => n11867, B2
                           => n8653, ZN => n3474);
   U15470 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_10_port, B1 => n11868, 
                           B2 => n8653, ZN => n3472);
   U15471 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_11_port, B1 => n11869, 
                           B2 => n8653, ZN => n3470);
   U15472 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_12_port, B1 => n11870, 
                           B2 => n8653, ZN => n3468);
   U15473 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_13_port, B1 => n11871, 
                           B2 => n8653, ZN => n3466);
   U15474 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_14_port, B1 => n11872, 
                           B2 => n8653, ZN => n3464);
   U15475 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_15_port, B1 => n7808, B2
                           => n8653, ZN => n3462);
   U15476 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_16_port, B1 => n11874, 
                           B2 => n8653, ZN => n3460);
   U15477 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_17_port, B1 => n11875, 
                           B2 => n8653, ZN => n3458);
   U15478 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_18_port, B1 => n11876, 
                           B2 => n8653, ZN => n3456);
   U15479 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_19_port, B1 => n11877, 
                           B2 => n8653, ZN => n3454);
   U15480 : AOI22_X1 port map( A1 => n12018, A2 => 
                           DataPath_RF_bus_reg_dataout_20_port, B1 => n11878, 
                           B2 => n8653, ZN => n3452);
   U15481 : AOI22_X1 port map( A1 => n12018, A2 => 
                           DataPath_RF_bus_reg_dataout_21_port, B1 => n11879, 
                           B2 => n8653, ZN => n3450);
   U15482 : AOI22_X1 port map( A1 => n12018, A2 => 
                           DataPath_RF_bus_reg_dataout_22_port, B1 => n11880, 
                           B2 => n8653, ZN => n3448);
   U15483 : AOI22_X1 port map( A1 => n12018, A2 => 
                           DataPath_RF_bus_reg_dataout_23_port, B1 => n11881, 
                           B2 => n8653, ZN => n3446);
   U15484 : AOI22_X1 port map( A1 => n12018, A2 => 
                           DataPath_RF_bus_reg_dataout_24_port, B1 => n11882, 
                           B2 => n8653, ZN => n3444);
   U15485 : AOI22_X1 port map( A1 => n12018, A2 => 
                           DataPath_RF_bus_reg_dataout_25_port, B1 => n11883, 
                           B2 => n8653, ZN => n3442);
   U15486 : AOI22_X1 port map( A1 => n12018, A2 => 
                           DataPath_RF_bus_reg_dataout_26_port, B1 => n11884, 
                           B2 => n8653, ZN => n3440);
   U15487 : AOI22_X1 port map( A1 => n12018, A2 => 
                           DataPath_RF_bus_reg_dataout_27_port, B1 => n11885, 
                           B2 => n8653, ZN => n3438);
   U15488 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_28_port, B1 => n11886, 
                           B2 => n8653, ZN => n3436);
   U15489 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_29_port, B1 => n11887, 
                           B2 => n8653, ZN => n3434);
   U15490 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_30_port, B1 => n11888, 
                           B2 => n8653, ZN => n3432);
   U15491 : NAND2_X1 port map( A1 => n11889, A2 => n11913, ZN => n11890);
   U15492 : OAI22_X1 port map( A1 => n11916, A2 => n11892, B1 => n788, B2 => 
                           n11891, ZN => n6991);
   U15493 : OAI22_X1 port map( A1 => n11917, A2 => n11892, B1 => n789, B2 => 
                           n11891, ZN => n6990);
   U15494 : OAI22_X1 port map( A1 => n11918, A2 => n11892, B1 => n790, B2 => 
                           n11891, ZN => n6989);
   U15495 : OAI22_X1 port map( A1 => n11919, A2 => n11892, B1 => n791, B2 => 
                           n11891, ZN => n6988);
   U15496 : OAI22_X1 port map( A1 => n11920, A2 => n11892, B1 => n792, B2 => 
                           n11891, ZN => n6987);
   U15497 : OAI22_X1 port map( A1 => n11921, A2 => n11892, B1 => n793, B2 => 
                           n11891, ZN => n6986);
   U15498 : OAI22_X1 port map( A1 => n11922, A2 => n11892, B1 => n794, B2 => 
                           n11891, ZN => n6985);
   U15499 : OAI22_X1 port map( A1 => n11923, A2 => n11892, B1 => n795, B2 => 
                           n11891, ZN => n6984);
   U15500 : OAI22_X1 port map( A1 => n11924, A2 => n11892, B1 => n796, B2 => 
                           n11891, ZN => n6983);
   U15501 : OAI22_X1 port map( A1 => n11925, A2 => n11892, B1 => n797, B2 => 
                           n11891, ZN => n6982);
   U15502 : OAI22_X1 port map( A1 => n11926, A2 => n11892, B1 => n798, B2 => 
                           n11891, ZN => n6981);
   U15503 : OAI22_X1 port map( A1 => n11927, A2 => n11892, B1 => n799, B2 => 
                           n11891, ZN => n6980);
   U15504 : OAI22_X1 port map( A1 => n11928, A2 => n8645, B1 => n800, B2 => 
                           n11891, ZN => n6979);
   U15505 : OAI22_X1 port map( A1 => n11929, A2 => n8645, B1 => n801, B2 => 
                           n11891, ZN => n6978);
   U15506 : OAI22_X1 port map( A1 => n11930, A2 => n8645, B1 => n802, B2 => 
                           n11891, ZN => n6977);
   U15507 : OAI22_X1 port map( A1 => n11931, A2 => n8645, B1 => n803, B2 => 
                           n11891, ZN => n6976);
   U15508 : OAI22_X1 port map( A1 => n11932, A2 => n8645, B1 => n804, B2 => 
                           n11891, ZN => n6975);
   U15509 : OAI22_X1 port map( A1 => n11933, A2 => n8645, B1 => n805, B2 => 
                           n11891, ZN => n6974);
   U15510 : OAI22_X1 port map( A1 => n11934, A2 => n8645, B1 => n806, B2 => 
                           n11891, ZN => n6973);
   U15511 : OAI22_X1 port map( A1 => n11935, A2 => n8645, B1 => n807, B2 => 
                           n11891, ZN => n6972);
   U15512 : OAI22_X1 port map( A1 => n11936, A2 => n8645, B1 => n808, B2 => 
                           n11891, ZN => n6971);
   U15513 : OAI22_X1 port map( A1 => n11937, A2 => n8645, B1 => n809, B2 => 
                           n11891, ZN => n6970);
   U15514 : OAI22_X1 port map( A1 => n11938, A2 => n8645, B1 => n810, B2 => 
                           n11891, ZN => n6969);
   U15515 : OAI22_X1 port map( A1 => n11939, A2 => n8645, B1 => n811, B2 => 
                           n11891, ZN => n6968);
   U15516 : OAI22_X1 port map( A1 => n11940, A2 => n11892, B1 => n812, B2 => 
                           n11891, ZN => n6967);
   U15517 : OAI22_X1 port map( A1 => n11941, A2 => n11892, B1 => n813, B2 => 
                           n11891, ZN => n6966);
   U15518 : OAI22_X1 port map( A1 => n11942, A2 => n11892, B1 => n814, B2 => 
                           n11891, ZN => n6965);
   U15519 : OAI22_X1 port map( A1 => n11943, A2 => n11892, B1 => n815, B2 => 
                           n11891, ZN => n6964);
   U15520 : OAI22_X1 port map( A1 => n11944, A2 => n11892, B1 => n816, B2 => 
                           n11891, ZN => n6963);
   U15521 : OAI22_X1 port map( A1 => n11945, A2 => n8645, B1 => n817, B2 => 
                           n11891, ZN => n6962);
   U15522 : OAI22_X1 port map( A1 => n11946, A2 => n8645, B1 => n818, B2 => 
                           n11891, ZN => n6961);
   U15523 : OAI22_X1 port map( A1 => n11949, A2 => n8645, B1 => n819, B2 => 
                           n11891, ZN => n6960);
   U15524 : NAND2_X1 port map( A1 => n11893, A2 => n11913, ZN => n11894);
   U15525 : OAI22_X1 port map( A1 => n11916, A2 => n11896, B1 => n756, B2 => 
                           n11895, ZN => n6959);
   U15526 : OAI22_X1 port map( A1 => n11917, A2 => n11896, B1 => n757, B2 => 
                           n11895, ZN => n6958);
   U15527 : OAI22_X1 port map( A1 => n11918, A2 => n11896, B1 => n758, B2 => 
                           n11895, ZN => n6957);
   U15528 : OAI22_X1 port map( A1 => n11919, A2 => n11896, B1 => n759, B2 => 
                           n11895, ZN => n6956);
   U15529 : OAI22_X1 port map( A1 => n11920, A2 => n11896, B1 => n760, B2 => 
                           n11895, ZN => n6955);
   U15530 : OAI22_X1 port map( A1 => n11921, A2 => n11896, B1 => n761, B2 => 
                           n11895, ZN => n6954);
   U15531 : OAI22_X1 port map( A1 => n11922, A2 => n11896, B1 => n762, B2 => 
                           n11895, ZN => n6953);
   U15532 : OAI22_X1 port map( A1 => n11923, A2 => n11896, B1 => n763, B2 => 
                           n11895, ZN => n6952);
   U15533 : OAI22_X1 port map( A1 => n11924, A2 => n11896, B1 => n764, B2 => 
                           n11895, ZN => n6951);
   U15534 : OAI22_X1 port map( A1 => n11925, A2 => n11896, B1 => n765, B2 => 
                           n11895, ZN => n6950);
   U15535 : OAI22_X1 port map( A1 => n11926, A2 => n11896, B1 => n766, B2 => 
                           n11895, ZN => n6949);
   U15536 : OAI22_X1 port map( A1 => n11927, A2 => n11896, B1 => n767, B2 => 
                           n11895, ZN => n6948);
   U15537 : OAI22_X1 port map( A1 => n11928, A2 => n8646, B1 => n768, B2 => 
                           n11895, ZN => n6947);
   U15538 : OAI22_X1 port map( A1 => n11929, A2 => n8646, B1 => n769, B2 => 
                           n11895, ZN => n6946);
   U15539 : OAI22_X1 port map( A1 => n11930, A2 => n8646, B1 => n770, B2 => 
                           n11895, ZN => n6945);
   U15540 : OAI22_X1 port map( A1 => n11931, A2 => n8646, B1 => n771, B2 => 
                           n11895, ZN => n6944);
   U15541 : OAI22_X1 port map( A1 => n11932, A2 => n8646, B1 => n772, B2 => 
                           n11895, ZN => n6943);
   U15542 : OAI22_X1 port map( A1 => n11933, A2 => n8646, B1 => n773, B2 => 
                           n11895, ZN => n6942);
   U15543 : OAI22_X1 port map( A1 => n11934, A2 => n8646, B1 => n774, B2 => 
                           n11895, ZN => n6941);
   U15544 : OAI22_X1 port map( A1 => n11935, A2 => n8646, B1 => n775, B2 => 
                           n11895, ZN => n6940);
   U15545 : OAI22_X1 port map( A1 => n11936, A2 => n8646, B1 => n776, B2 => 
                           n11895, ZN => n6939);
   U15546 : OAI22_X1 port map( A1 => n11937, A2 => n8646, B1 => n777, B2 => 
                           n11895, ZN => n6938);
   U15547 : OAI22_X1 port map( A1 => n11938, A2 => n8646, B1 => n778, B2 => 
                           n11895, ZN => n6937);
   U15548 : OAI22_X1 port map( A1 => n11939, A2 => n8646, B1 => n779, B2 => 
                           n11895, ZN => n6936);
   U15549 : OAI22_X1 port map( A1 => n11940, A2 => n11896, B1 => n780, B2 => 
                           n11895, ZN => n6935);
   U15550 : OAI22_X1 port map( A1 => n11941, A2 => n11896, B1 => n781, B2 => 
                           n11895, ZN => n6934);
   U15551 : OAI22_X1 port map( A1 => n11942, A2 => n11896, B1 => n782, B2 => 
                           n11895, ZN => n6933);
   U15552 : OAI22_X1 port map( A1 => n11943, A2 => n11896, B1 => n783, B2 => 
                           n11895, ZN => n6932);
   U15553 : OAI22_X1 port map( A1 => n11944, A2 => n11896, B1 => n784, B2 => 
                           n11895, ZN => n6931);
   U15554 : OAI22_X1 port map( A1 => n11945, A2 => n8646, B1 => n785, B2 => 
                           n11895, ZN => n6930);
   U15555 : OAI22_X1 port map( A1 => n11946, A2 => n8646, B1 => n786, B2 => 
                           n11895, ZN => n6929);
   U15556 : OAI22_X1 port map( A1 => n11949, A2 => n8646, B1 => n787, B2 => 
                           n11895, ZN => n6928);
   U15557 : NAND2_X1 port map( A1 => n11897, A2 => n11913, ZN => n11898);
   U15558 : OAI22_X1 port map( A1 => n11916, A2 => n11900, B1 => n724, B2 => 
                           n11899, ZN => n6927);
   U15559 : OAI22_X1 port map( A1 => n11917, A2 => n11900, B1 => n725, B2 => 
                           n11899, ZN => n6926);
   U15560 : OAI22_X1 port map( A1 => n11918, A2 => n11900, B1 => n726, B2 => 
                           n11899, ZN => n6925);
   U15561 : OAI22_X1 port map( A1 => n11919, A2 => n11900, B1 => n727, B2 => 
                           n11899, ZN => n6924);
   U15562 : OAI22_X1 port map( A1 => n11920, A2 => n11900, B1 => n728, B2 => 
                           n11899, ZN => n6923);
   U15563 : OAI22_X1 port map( A1 => n11921, A2 => n11900, B1 => n729, B2 => 
                           n11899, ZN => n6922);
   U15564 : OAI22_X1 port map( A1 => n11922, A2 => n11900, B1 => n730, B2 => 
                           n11899, ZN => n6921);
   U15565 : OAI22_X1 port map( A1 => n11923, A2 => n11900, B1 => n731, B2 => 
                           n11899, ZN => n6920);
   U15566 : OAI22_X1 port map( A1 => n11924, A2 => n11900, B1 => n732, B2 => 
                           n11899, ZN => n6919);
   U15567 : OAI22_X1 port map( A1 => n11925, A2 => n11900, B1 => n733, B2 => 
                           n11899, ZN => n6918);
   U15568 : OAI22_X1 port map( A1 => n11926, A2 => n11900, B1 => n734, B2 => 
                           n11899, ZN => n6917);
   U15569 : OAI22_X1 port map( A1 => n11927, A2 => n11900, B1 => n735, B2 => 
                           n11899, ZN => n6916);
   U15570 : OAI22_X1 port map( A1 => n11928, A2 => n8647, B1 => n736, B2 => 
                           n11899, ZN => n6915);
   U15571 : OAI22_X1 port map( A1 => n11929, A2 => n8647, B1 => n737, B2 => 
                           n11899, ZN => n6914);
   U15572 : OAI22_X1 port map( A1 => n11930, A2 => n8647, B1 => n738, B2 => 
                           n11899, ZN => n6913);
   U15573 : OAI22_X1 port map( A1 => n11931, A2 => n8647, B1 => n739, B2 => 
                           n11899, ZN => n6912);
   U15574 : OAI22_X1 port map( A1 => n11932, A2 => n8647, B1 => n740, B2 => 
                           n11899, ZN => n6911);
   U15575 : OAI22_X1 port map( A1 => n11933, A2 => n8647, B1 => n741, B2 => 
                           n11899, ZN => n6910);
   U15576 : OAI22_X1 port map( A1 => n11934, A2 => n8647, B1 => n742, B2 => 
                           n11899, ZN => n6909);
   U15577 : OAI22_X1 port map( A1 => n11935, A2 => n8647, B1 => n743, B2 => 
                           n11899, ZN => n6908);
   U15578 : OAI22_X1 port map( A1 => n11936, A2 => n8647, B1 => n744, B2 => 
                           n11899, ZN => n6907);
   U15579 : OAI22_X1 port map( A1 => n11937, A2 => n8647, B1 => n745, B2 => 
                           n11899, ZN => n6906);
   U15580 : OAI22_X1 port map( A1 => n11938, A2 => n8647, B1 => n746, B2 => 
                           n11899, ZN => n6905);
   U15581 : OAI22_X1 port map( A1 => n11939, A2 => n8647, B1 => n747, B2 => 
                           n11899, ZN => n6904);
   U15582 : OAI22_X1 port map( A1 => n11940, A2 => n11900, B1 => n748, B2 => 
                           n11899, ZN => n6903);
   U15583 : OAI22_X1 port map( A1 => n11941, A2 => n11900, B1 => n749, B2 => 
                           n11899, ZN => n6902);
   U15584 : OAI22_X1 port map( A1 => n11942, A2 => n11900, B1 => n750, B2 => 
                           n11899, ZN => n6901);
   U15585 : OAI22_X1 port map( A1 => n11943, A2 => n11900, B1 => n751, B2 => 
                           n11899, ZN => n6900);
   U15586 : OAI22_X1 port map( A1 => n11944, A2 => n11900, B1 => n752, B2 => 
                           n11899, ZN => n6899);
   U15587 : OAI22_X1 port map( A1 => n11945, A2 => n8647, B1 => n753, B2 => 
                           n11899, ZN => n6898);
   U15588 : OAI22_X1 port map( A1 => n11946, A2 => n8647, B1 => n754, B2 => 
                           n11899, ZN => n6897);
   U15589 : OAI22_X1 port map( A1 => n11949, A2 => n8647, B1 => n755, B2 => 
                           n11899, ZN => n6896);
   U15590 : NAND2_X1 port map( A1 => n11901, A2 => n11913, ZN => n11902);
   U15591 : OAI22_X1 port map( A1 => n11916, A2 => n11904, B1 => n692, B2 => 
                           n11903, ZN => n6895);
   U15592 : OAI22_X1 port map( A1 => n11917, A2 => n11904, B1 => n693, B2 => 
                           n11903, ZN => n6894);
   U15593 : OAI22_X1 port map( A1 => n11918, A2 => n11904, B1 => n694, B2 => 
                           n11903, ZN => n6893);
   U15594 : OAI22_X1 port map( A1 => n11919, A2 => n11904, B1 => n695, B2 => 
                           n11903, ZN => n6892);
   U15595 : OAI22_X1 port map( A1 => n11920, A2 => n11904, B1 => n696, B2 => 
                           n11903, ZN => n6891);
   U15596 : OAI22_X1 port map( A1 => n11921, A2 => n11904, B1 => n697, B2 => 
                           n11903, ZN => n6890);
   U15597 : OAI22_X1 port map( A1 => n11922, A2 => n11904, B1 => n698, B2 => 
                           n11903, ZN => n6889);
   U15598 : OAI22_X1 port map( A1 => n11923, A2 => n11904, B1 => n699, B2 => 
                           n11903, ZN => n6888);
   U15599 : OAI22_X1 port map( A1 => n11924, A2 => n11904, B1 => n700, B2 => 
                           n11903, ZN => n6887);
   U15600 : OAI22_X1 port map( A1 => n11925, A2 => n11904, B1 => n701, B2 => 
                           n11903, ZN => n6886);
   U15601 : OAI22_X1 port map( A1 => n11926, A2 => n11904, B1 => n702, B2 => 
                           n11903, ZN => n6885);
   U15602 : OAI22_X1 port map( A1 => n11927, A2 => n11904, B1 => n703, B2 => 
                           n11903, ZN => n6884);
   U15603 : OAI22_X1 port map( A1 => n11928, A2 => n8648, B1 => n704, B2 => 
                           n11903, ZN => n6883);
   U15604 : OAI22_X1 port map( A1 => n11929, A2 => n8648, B1 => n705, B2 => 
                           n11903, ZN => n6882);
   U15605 : OAI22_X1 port map( A1 => n11930, A2 => n8648, B1 => n706, B2 => 
                           n11903, ZN => n6881);
   U15606 : OAI22_X1 port map( A1 => n11931, A2 => n8648, B1 => n707, B2 => 
                           n11903, ZN => n6880);
   U15607 : OAI22_X1 port map( A1 => n11932, A2 => n8648, B1 => n708, B2 => 
                           n11903, ZN => n6879);
   U15608 : OAI22_X1 port map( A1 => n11933, A2 => n8648, B1 => n709, B2 => 
                           n11903, ZN => n6878);
   U15609 : OAI22_X1 port map( A1 => n11934, A2 => n8648, B1 => n710, B2 => 
                           n11903, ZN => n6877);
   U15610 : OAI22_X1 port map( A1 => n11935, A2 => n8648, B1 => n711, B2 => 
                           n11903, ZN => n6876);
   U15611 : OAI22_X1 port map( A1 => n11936, A2 => n8648, B1 => n712, B2 => 
                           n11903, ZN => n6875);
   U15612 : OAI22_X1 port map( A1 => n11937, A2 => n8648, B1 => n713, B2 => 
                           n11903, ZN => n6874);
   U15613 : OAI22_X1 port map( A1 => n11938, A2 => n8648, B1 => n714, B2 => 
                           n11903, ZN => n6873);
   U15614 : OAI22_X1 port map( A1 => n11939, A2 => n8648, B1 => n715, B2 => 
                           n11903, ZN => n6872);
   U15615 : OAI22_X1 port map( A1 => n11940, A2 => n11904, B1 => n716, B2 => 
                           n11903, ZN => n6871);
   U15616 : OAI22_X1 port map( A1 => n11941, A2 => n11904, B1 => n717, B2 => 
                           n11903, ZN => n6870);
   U15617 : OAI22_X1 port map( A1 => n11942, A2 => n11904, B1 => n718, B2 => 
                           n11903, ZN => n6869);
   U15618 : OAI22_X1 port map( A1 => n11943, A2 => n11904, B1 => n719, B2 => 
                           n11903, ZN => n6868);
   U15619 : OAI22_X1 port map( A1 => n11944, A2 => n11904, B1 => n720, B2 => 
                           n11903, ZN => n6867);
   U15620 : OAI22_X1 port map( A1 => n11945, A2 => n8648, B1 => n721, B2 => 
                           n11903, ZN => n6866);
   U15621 : OAI22_X1 port map( A1 => n11946, A2 => n8648, B1 => n722, B2 => 
                           n11903, ZN => n6865);
   U15622 : OAI22_X1 port map( A1 => n11949, A2 => n8648, B1 => n723, B2 => 
                           n11903, ZN => n6864);
   U15623 : NAND2_X1 port map( A1 => n11905, A2 => n11913, ZN => n11906);
   U15624 : OAI22_X1 port map( A1 => n11916, A2 => n11908, B1 => n660, B2 => 
                           n11907, ZN => n6863);
   U15625 : OAI22_X1 port map( A1 => n11917, A2 => n11908, B1 => n661, B2 => 
                           n11907, ZN => n6862);
   U15626 : OAI22_X1 port map( A1 => n11918, A2 => n11908, B1 => n662, B2 => 
                           n11907, ZN => n6861);
   U15627 : OAI22_X1 port map( A1 => n11919, A2 => n11908, B1 => n663, B2 => 
                           n11907, ZN => n6860);
   U15628 : OAI22_X1 port map( A1 => n11920, A2 => n11908, B1 => n664, B2 => 
                           n11907, ZN => n6859);
   U15629 : OAI22_X1 port map( A1 => n11921, A2 => n11908, B1 => n665, B2 => 
                           n11907, ZN => n6858);
   U15630 : OAI22_X1 port map( A1 => n11922, A2 => n11908, B1 => n666, B2 => 
                           n11907, ZN => n6857);
   U15631 : OAI22_X1 port map( A1 => n11923, A2 => n11908, B1 => n667, B2 => 
                           n11907, ZN => n6856);
   U15632 : OAI22_X1 port map( A1 => n11924, A2 => n11908, B1 => n668, B2 => 
                           n11907, ZN => n6855);
   U15633 : OAI22_X1 port map( A1 => n11925, A2 => n11908, B1 => n669, B2 => 
                           n11907, ZN => n6854);
   U15634 : OAI22_X1 port map( A1 => n11926, A2 => n11908, B1 => n670, B2 => 
                           n11907, ZN => n6853);
   U15635 : OAI22_X1 port map( A1 => n11927, A2 => n11908, B1 => n671, B2 => 
                           n11907, ZN => n6852);
   U15636 : OAI22_X1 port map( A1 => n11928, A2 => n8649, B1 => n672, B2 => 
                           n11907, ZN => n6851);
   U15637 : OAI22_X1 port map( A1 => n11929, A2 => n8649, B1 => n673, B2 => 
                           n11907, ZN => n6850);
   U15638 : OAI22_X1 port map( A1 => n11930, A2 => n8649, B1 => n674, B2 => 
                           n11907, ZN => n6849);
   U15639 : OAI22_X1 port map( A1 => n11931, A2 => n8649, B1 => n675, B2 => 
                           n11907, ZN => n6848);
   U15640 : OAI22_X1 port map( A1 => n11932, A2 => n8649, B1 => n676, B2 => 
                           n11907, ZN => n6847);
   U15641 : OAI22_X1 port map( A1 => n11933, A2 => n8649, B1 => n677, B2 => 
                           n11907, ZN => n6846);
   U15642 : OAI22_X1 port map( A1 => n11934, A2 => n8649, B1 => n678, B2 => 
                           n11907, ZN => n6845);
   U15643 : OAI22_X1 port map( A1 => n11935, A2 => n8649, B1 => n679, B2 => 
                           n11907, ZN => n6844);
   U15644 : OAI22_X1 port map( A1 => n11936, A2 => n8649, B1 => n680, B2 => 
                           n11907, ZN => n6843);
   U15645 : OAI22_X1 port map( A1 => n11937, A2 => n8649, B1 => n681, B2 => 
                           n11907, ZN => n6842);
   U15646 : OAI22_X1 port map( A1 => n11938, A2 => n8649, B1 => n682, B2 => 
                           n11907, ZN => n6841);
   U15647 : OAI22_X1 port map( A1 => n11939, A2 => n8649, B1 => n683, B2 => 
                           n11907, ZN => n6840);
   U15648 : OAI22_X1 port map( A1 => n11940, A2 => n11908, B1 => n684, B2 => 
                           n11907, ZN => n6839);
   U15649 : OAI22_X1 port map( A1 => n11941, A2 => n11908, B1 => n685, B2 => 
                           n11907, ZN => n6838);
   U15650 : OAI22_X1 port map( A1 => n11942, A2 => n11908, B1 => n686, B2 => 
                           n11907, ZN => n6837);
   U15651 : OAI22_X1 port map( A1 => n11943, A2 => n11908, B1 => n687, B2 => 
                           n11907, ZN => n6836);
   U15652 : OAI22_X1 port map( A1 => n11944, A2 => n11908, B1 => n688, B2 => 
                           n11907, ZN => n6835);
   U15653 : OAI22_X1 port map( A1 => n11945, A2 => n8649, B1 => n689, B2 => 
                           n11907, ZN => n6834);
   U15654 : OAI22_X1 port map( A1 => n11946, A2 => n8649, B1 => n690, B2 => 
                           n11907, ZN => n6833);
   U15655 : OAI22_X1 port map( A1 => n11949, A2 => n8649, B1 => n691, B2 => 
                           n11907, ZN => n6832);
   U15656 : NAND2_X1 port map( A1 => n11909, A2 => n11913, ZN => n11910);
   U15657 : OAI22_X1 port map( A1 => n11916, A2 => n11912, B1 => n628, B2 => 
                           n11911, ZN => n6831);
   U15658 : OAI22_X1 port map( A1 => n11917, A2 => n11912, B1 => n629, B2 => 
                           n11911, ZN => n6830);
   U15659 : OAI22_X1 port map( A1 => n11918, A2 => n11912, B1 => n630, B2 => 
                           n11911, ZN => n6829);
   U15660 : OAI22_X1 port map( A1 => n11919, A2 => n11912, B1 => n631, B2 => 
                           n11911, ZN => n6828);
   U15661 : OAI22_X1 port map( A1 => n11920, A2 => n11912, B1 => n632, B2 => 
                           n11911, ZN => n6827);
   U15662 : OAI22_X1 port map( A1 => n11921, A2 => n11912, B1 => n633, B2 => 
                           n11911, ZN => n6826);
   U15663 : OAI22_X1 port map( A1 => n11922, A2 => n11912, B1 => n634, B2 => 
                           n11911, ZN => n6825);
   U15664 : OAI22_X1 port map( A1 => n11923, A2 => n11912, B1 => n635, B2 => 
                           n11911, ZN => n6824);
   U15665 : OAI22_X1 port map( A1 => n11924, A2 => n11912, B1 => n636, B2 => 
                           n11911, ZN => n6823);
   U15666 : OAI22_X1 port map( A1 => n11925, A2 => n11912, B1 => n637, B2 => 
                           n11911, ZN => n6822);
   U15667 : OAI22_X1 port map( A1 => n11926, A2 => n11912, B1 => n638, B2 => 
                           n11911, ZN => n6821);
   U15668 : OAI22_X1 port map( A1 => n11927, A2 => n11912, B1 => n639, B2 => 
                           n11911, ZN => n6820);
   U15669 : OAI22_X1 port map( A1 => n11928, A2 => n8650, B1 => n640, B2 => 
                           n11911, ZN => n6819);
   U15670 : OAI22_X1 port map( A1 => n11929, A2 => n8650, B1 => n641, B2 => 
                           n11911, ZN => n6818);
   U15671 : OAI22_X1 port map( A1 => n11930, A2 => n8650, B1 => n642, B2 => 
                           n11911, ZN => n6817);
   U15672 : OAI22_X1 port map( A1 => n11931, A2 => n8650, B1 => n643, B2 => 
                           n11911, ZN => n6816);
   U15673 : OAI22_X1 port map( A1 => n11932, A2 => n8650, B1 => n644, B2 => 
                           n11911, ZN => n6815);
   U15674 : OAI22_X1 port map( A1 => n11933, A2 => n8650, B1 => n645, B2 => 
                           n11911, ZN => n6814);
   U15675 : OAI22_X1 port map( A1 => n11934, A2 => n8650, B1 => n646, B2 => 
                           n11911, ZN => n6813);
   U15676 : OAI22_X1 port map( A1 => n11935, A2 => n8650, B1 => n647, B2 => 
                           n11911, ZN => n6812);
   U15677 : OAI22_X1 port map( A1 => n11936, A2 => n8650, B1 => n648, B2 => 
                           n11911, ZN => n6811);
   U15678 : OAI22_X1 port map( A1 => n11937, A2 => n8650, B1 => n649, B2 => 
                           n11911, ZN => n6810);
   U15679 : OAI22_X1 port map( A1 => n11938, A2 => n8650, B1 => n650, B2 => 
                           n11911, ZN => n6809);
   U15680 : OAI22_X1 port map( A1 => n11939, A2 => n8650, B1 => n651, B2 => 
                           n11911, ZN => n6808);
   U15681 : OAI22_X1 port map( A1 => n11940, A2 => n11912, B1 => n652, B2 => 
                           n11911, ZN => n6807);
   U15682 : OAI22_X1 port map( A1 => n11941, A2 => n11912, B1 => n653, B2 => 
                           n11911, ZN => n6806);
   U15683 : OAI22_X1 port map( A1 => n11942, A2 => n11912, B1 => n654, B2 => 
                           n11911, ZN => n6805);
   U15684 : OAI22_X1 port map( A1 => n11943, A2 => n11912, B1 => n655, B2 => 
                           n11911, ZN => n6804);
   U15685 : OAI22_X1 port map( A1 => n11944, A2 => n11912, B1 => n656, B2 => 
                           n11911, ZN => n6803);
   U15686 : OAI22_X1 port map( A1 => n11945, A2 => n8650, B1 => n657, B2 => 
                           n11911, ZN => n6802);
   U15687 : OAI22_X1 port map( A1 => n11946, A2 => n8650, B1 => n658, B2 => 
                           n11911, ZN => n6801);
   U15688 : OAI22_X1 port map( A1 => n11949, A2 => n8650, B1 => n659, B2 => 
                           n11911, ZN => n6800);
   U15689 : NAND2_X1 port map( A1 => n11914, A2 => n11913, ZN => n11915);
   U15690 : OAI22_X1 port map( A1 => n11916, A2 => n11948, B1 => n596, B2 => 
                           n11947, ZN => n6799);
   U15691 : OAI22_X1 port map( A1 => n11917, A2 => n11948, B1 => n597, B2 => 
                           n11947, ZN => n6798);
   U15692 : OAI22_X1 port map( A1 => n11918, A2 => n11948, B1 => n598, B2 => 
                           n11947, ZN => n6797);
   U15693 : OAI22_X1 port map( A1 => n11919, A2 => n11948, B1 => n599, B2 => 
                           n11947, ZN => n6796);
   U15694 : OAI22_X1 port map( A1 => n11920, A2 => n11948, B1 => n600, B2 => 
                           n11947, ZN => n6795);
   U15695 : OAI22_X1 port map( A1 => n11921, A2 => n11948, B1 => n601, B2 => 
                           n11947, ZN => n6794);
   U15696 : OAI22_X1 port map( A1 => n11922, A2 => n11948, B1 => n602, B2 => 
                           n11947, ZN => n6793);
   U15697 : OAI22_X1 port map( A1 => n11923, A2 => n11948, B1 => n603, B2 => 
                           n11947, ZN => n6792);
   U15698 : OAI22_X1 port map( A1 => n11924, A2 => n11948, B1 => n604, B2 => 
                           n11947, ZN => n6791);
   U15699 : OAI22_X1 port map( A1 => n11925, A2 => n11948, B1 => n605, B2 => 
                           n11947, ZN => n6790);
   U15700 : OAI22_X1 port map( A1 => n11926, A2 => n11948, B1 => n606, B2 => 
                           n11947, ZN => n6789);
   U15701 : OAI22_X1 port map( A1 => n11927, A2 => n11948, B1 => n607, B2 => 
                           n11947, ZN => n6788);
   U15702 : OAI22_X1 port map( A1 => n11928, A2 => n8651, B1 => n608, B2 => 
                           n11947, ZN => n6787);
   U15703 : OAI22_X1 port map( A1 => n11929, A2 => n8651, B1 => n609, B2 => 
                           n11947, ZN => n6786);
   U15704 : OAI22_X1 port map( A1 => n11930, A2 => n8651, B1 => n610, B2 => 
                           n11947, ZN => n6785);
   U15705 : OAI22_X1 port map( A1 => n11931, A2 => n8651, B1 => n611, B2 => 
                           n11947, ZN => n6784);
   U15706 : OAI22_X1 port map( A1 => n11932, A2 => n8651, B1 => n612, B2 => 
                           n11947, ZN => n6783);
   U15707 : OAI22_X1 port map( A1 => n11933, A2 => n8651, B1 => n613, B2 => 
                           n11947, ZN => n6782);
   U15708 : OAI22_X1 port map( A1 => n11934, A2 => n8651, B1 => n614, B2 => 
                           n11947, ZN => n6781);
   U15709 : OAI22_X1 port map( A1 => n11935, A2 => n8651, B1 => n615, B2 => 
                           n11947, ZN => n6780);
   U15710 : OAI22_X1 port map( A1 => n11936, A2 => n8651, B1 => n616, B2 => 
                           n11947, ZN => n6779);
   U15711 : OAI22_X1 port map( A1 => n11937, A2 => n8651, B1 => n617, B2 => 
                           n11947, ZN => n6778);
   U15712 : OAI22_X1 port map( A1 => n11938, A2 => n8651, B1 => n618, B2 => 
                           n11947, ZN => n6777);
   U15713 : OAI22_X1 port map( A1 => n11939, A2 => n8651, B1 => n619, B2 => 
                           n11947, ZN => n6776);
   U15714 : OAI22_X1 port map( A1 => n11940, A2 => n11948, B1 => n620, B2 => 
                           n11947, ZN => n6775);
   U15715 : OAI22_X1 port map( A1 => n11941, A2 => n11948, B1 => n621, B2 => 
                           n11947, ZN => n6774);
   U15716 : OAI22_X1 port map( A1 => n11942, A2 => n11948, B1 => n622, B2 => 
                           n11947, ZN => n6773);
   U15717 : OAI22_X1 port map( A1 => n11943, A2 => n11948, B1 => n623, B2 => 
                           n11947, ZN => n6772);
   U15718 : OAI22_X1 port map( A1 => n11944, A2 => n11948, B1 => n624, B2 => 
                           n11947, ZN => n6771);
   U15719 : OAI22_X1 port map( A1 => n11945, A2 => n8651, B1 => n625, B2 => 
                           n11947, ZN => n6770);
   U15720 : OAI22_X1 port map( A1 => n11946, A2 => n8651, B1 => n626, B2 => 
                           n11947, ZN => n6769);
   U15721 : OAI22_X1 port map( A1 => n11949, A2 => n8651, B1 => n627, B2 => 
                           n11947, ZN => n6768);
   U15722 : AOI22_X1 port map( A1 => i_RD1_0_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_A_0_port, ZN => n3383);
   U15723 : AOI22_X1 port map( A1 => i_RD1_1_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_A_1_port, ZN => n11951);
   U15724 : INV_X1 port map( A => n11951, ZN => n6735);
   U15725 : AOI22_X1 port map( A1 => i_RD1_2_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_A_2_port, ZN => n3382);
   U15726 : AOI22_X1 port map( A1 => i_RD1_3_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_A_3_port, ZN => n11952);
   U15727 : INV_X1 port map( A => n11952, ZN => n6734);
   U15728 : AOI22_X1 port map( A1 => i_RD1_4_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_A_4_port, ZN => n3381);
   U15729 : AOI22_X1 port map( A1 => i_RD1_5_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_A_5_port, ZN => n3380);
   U15730 : AOI22_X1 port map( A1 => i_RD1_6_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_A_6_port, ZN => n3379);
   U15731 : AOI22_X1 port map( A1 => i_RD1_7_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_A_7_port, ZN => n3378);
   U15732 : AOI22_X1 port map( A1 => i_RD1_8_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_A_8_port, ZN => n11953);
   U15733 : INV_X1 port map( A => n11953, ZN => n6733);
   U15734 : AOI22_X1 port map( A1 => i_RD1_9_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_A_9_port, ZN => n3377);
   U15735 : AOI22_X1 port map( A1 => i_RD1_10_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_10_port, ZN => n3376);
   U15736 : AOI22_X1 port map( A1 => i_RD1_11_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_11_port, ZN => n3375);
   U15737 : AOI22_X1 port map( A1 => i_RD1_12_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_12_port, ZN => n3374);
   U15738 : AOI22_X1 port map( A1 => i_RD1_13_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_13_port, ZN => n11954);
   U15739 : INV_X1 port map( A => n11954, ZN => n6732);
   U15740 : AOI22_X1 port map( A1 => i_RD1_14_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_14_port, ZN => n11955);
   U15741 : INV_X1 port map( A => n11955, ZN => n6731);
   U15742 : AOI22_X1 port map( A1 => i_RD1_15_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_15_port, ZN => n3373);
   U15743 : AOI22_X1 port map( A1 => i_RD1_16_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_16_port, ZN => n3372);
   U15744 : AOI22_X1 port map( A1 => i_RD1_17_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_17_port, ZN => n3371);
   U15745 : AOI22_X1 port map( A1 => i_RD1_18_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_18_port, ZN => n3370);
   U15746 : AOI22_X1 port map( A1 => i_RD1_19_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_19_port, ZN => n3369);
   U15747 : AOI22_X1 port map( A1 => i_RD1_21_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_21_port, ZN => n3368);
   U15748 : AOI22_X1 port map( A1 => i_RD1_22_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_22_port, ZN => n3367);
   U15749 : AOI22_X1 port map( A1 => i_RD1_23_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_23_port, ZN => n3366);
   U15750 : AOI22_X1 port map( A1 => i_RD1_24_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_24_port, ZN => n3365);
   U15751 : AOI22_X1 port map( A1 => i_RD1_25_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_25_port, ZN => n3364);
   U15752 : AOI22_X1 port map( A1 => i_RD1_26_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_26_port, ZN => n3363);
   U15753 : AOI22_X1 port map( A1 => i_RD1_27_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_27_port, ZN => n3362);
   U15754 : AOI22_X1 port map( A1 => i_RD1_28_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_28_port, ZN => n3361);
   U15755 : AOI22_X1 port map( A1 => i_RD1_29_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_29_port, ZN => n3360);
   U15756 : AOI22_X1 port map( A1 => i_RD1_30_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_30_port, ZN => n3359);
   U15757 : AOI22_X1 port map( A1 => i_RD1_31_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_A_31_port, ZN => n3358);
   U15758 : OR2_X1 port map( A1 => RST, A2 => n11956, ZN => n3357);
   U15759 : OR2_X1 port map( A1 => RST, A2 => n11957, ZN => n3356);
   U15760 : OR2_X1 port map( A1 => RST, A2 => n11958, ZN => n3355);
   U15761 : OR2_X1 port map( A1 => RST, A2 => n11959, ZN => n3354);
   U15762 : OR2_X1 port map( A1 => RST, A2 => n11960, ZN => n3353);
   U15763 : OR2_X1 port map( A1 => RST, A2 => n11961, ZN => n3352);
   U15764 : OR2_X1 port map( A1 => RST, A2 => n11962, ZN => n3351);
   U15765 : OR2_X1 port map( A1 => RST, A2 => n11963, ZN => n3349);
   U15766 : OR2_X1 port map( A1 => RST, A2 => n11964, ZN => n3348);
   U15767 : OR2_X1 port map( A1 => RST, A2 => n11965, ZN => n3346);
   U15768 : OR2_X1 port map( A1 => RST, A2 => n11966, ZN => n3344);
   U15769 : OR2_X1 port map( A1 => RST, A2 => n11967, ZN => n3343);
   U15770 : OR2_X1 port map( A1 => RST, A2 => n11968, ZN => n3334);
   U15771 : OR2_X1 port map( A1 => RST, A2 => n11969, ZN => n3333);
   U15772 : OR2_X1 port map( A1 => RST, A2 => n11970, ZN => n3331);
   U15773 : OR2_X1 port map( A1 => RST, A2 => n11971, ZN => n3329);
   U15774 : NOR2_X1 port map( A1 => n544, A2 => n543, ZN => n11973);
   U15775 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_2_port, A2 => 
                           n11973, ZN => n11975);
   U15776 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_4_port, A2 => 
                           n11976, ZN => n11978);
   U15777 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_6_port, A2 => 
                           n11979, ZN => n11981);
   U15778 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_8_port, A2 => 
                           n11982, ZN => n11984);
   U15779 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_10_port, A2 => 
                           n11985, ZN => n11987);
   U15780 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_12_port, A2 => 
                           n11988, ZN => n11990);
   U15781 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_14_port, A2 => 
                           n11991, ZN => n11993);
   U15782 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_16_port, A2 => 
                           n11994, ZN => n11996);
   U15783 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_18_port, A2 => 
                           n11997, ZN => n11999);
   U15784 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_20_port, A2 => 
                           n12000, ZN => n12002);
   U15785 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_22_port, A2 => 
                           n12003, ZN => n12005);
   U15786 : NOR2_X1 port map( A1 => n566, A2 => n12005, ZN => n12006);
   U15787 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_24_port, A2 => 
                           n12006, ZN => n12008);
   U15788 : NOR2_X1 port map( A1 => n568, A2 => n12008, ZN => n12009);
   U15789 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_26_port, A2 => 
                           n12009, ZN => n12012);
   U15790 : NOR2_X1 port map( A1 => n570, A2 => n12012, ZN => n12011);
   U15791 : INV_X1 port map( A => n12011, ZN => n12013);
   U15792 : NOR2_X1 port map( A1 => n571, A2 => n12013, ZN => n12014);
   U15793 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_29_port, A2 => 
                           n12014, ZN => n12016);
   U15794 : NOR2_X1 port map( A1 => n572, A2 => n12016, ZN => n12015);
   U15795 : OAI21_X1 port map( B1 => DECODEhw_i_tickcounter_31_port, B2 => 
                           n12015, A => n8691, ZN => n11972);
   U15796 : AOI21_X1 port map( B1 => DECODEhw_i_tickcounter_31_port, B2 => 
                           n12015, A => n11972, ZN => n7153);
   U15797 : AND2_X1 port map( A1 => n8689, A2 => n543, ZN => n7152);
   U15798 : AOI211_X1 port map( C1 => n543, C2 => n544, A => RST, B => n11973, 
                           ZN => n7151);
   U15799 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_2_port, C2 => 
                           n11973, A => n11975, B => n8698, ZN => n11974);
   U15800 : AOI211_X1 port map( C1 => n546, C2 => n11975, A => RST, B => n11976
                           , ZN => n7149);
   U15801 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_4_port, C2 => 
                           n11976, A => n11978, B => n8692, ZN => n11977);
   U15802 : INV_X1 port map( A => n11977, ZN => n7148);
   U15803 : AOI211_X1 port map( C1 => n548, C2 => n11978, A => RST, B => n11979
                           , ZN => n7147);
   U15804 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_6_port, C2 => 
                           n11979, A => n11981, B => n8688, ZN => n11980);
   U15805 : INV_X1 port map( A => n11980, ZN => n7146);
   U15806 : AOI211_X1 port map( C1 => n550, C2 => n11981, A => RST, B => n11982
                           , ZN => n7145);
   U15807 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_8_port, C2 => 
                           n11982, A => n11984, B => n8692, ZN => n11983);
   U15808 : INV_X1 port map( A => n11983, ZN => n7144);
   U15809 : AOI211_X1 port map( C1 => n552, C2 => n11984, A => RST, B => n11985
                           , ZN => n7143);
   U15810 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_10_port, C2 => 
                           n11985, A => n11987, B => n8692, ZN => n11986);
   U15811 : INV_X1 port map( A => n11986, ZN => n7142);
   U15812 : AOI211_X1 port map( C1 => n554, C2 => n11987, A => RST, B => n11988
                           , ZN => n7141);
   U15813 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_12_port, C2 => 
                           n11988, A => n11990, B => n8689, ZN => n11989);
   U15814 : INV_X1 port map( A => n11989, ZN => n7140);
   U15815 : AOI211_X1 port map( C1 => n556, C2 => n11990, A => RST, B => n11991
                           , ZN => n7139);
   U15816 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_14_port, C2 => 
                           n11991, A => n11993, B => n8692, ZN => n11992);
   U15817 : INV_X1 port map( A => n11992, ZN => n7138);
   U15818 : AOI211_X1 port map( C1 => n558, C2 => n11993, A => RST, B => n11994
                           , ZN => n7137);
   U15819 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_16_port, C2 => 
                           n11994, A => n11996, B => n8697, ZN => n11995);
   U15820 : INV_X1 port map( A => n11995, ZN => n7136);
   U15821 : AOI211_X1 port map( C1 => n560, C2 => n11996, A => RST, B => n11997
                           , ZN => n7135);
   U15822 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_18_port, C2 => 
                           n11997, A => n11999, B => n8695, ZN => n11998);
   U15823 : INV_X1 port map( A => n11998, ZN => n7134);
   U15824 : AOI211_X1 port map( C1 => n562, C2 => n11999, A => RST, B => n12000
                           , ZN => n7133);
   U15825 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_20_port, C2 => 
                           n12000, A => n12002, B => n8692, ZN => n12001);
   U15826 : INV_X1 port map( A => n12001, ZN => n7132);
   U15827 : AOI211_X1 port map( C1 => n564, C2 => n12002, A => RST, B => n12003
                           , ZN => n7131);
   U15828 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_22_port, C2 => 
                           n12003, A => n12005, B => n8688, ZN => n12004);
   U15829 : INV_X1 port map( A => n12004, ZN => n7130);
   U15830 : AOI211_X1 port map( C1 => n566, C2 => n12005, A => RST, B => n12006
                           , ZN => n7129);
   U15831 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_24_port, C2 => 
                           n12006, A => n12008, B => n8697, ZN => n12007);
   U15832 : INV_X1 port map( A => n12007, ZN => n7128);
   U15833 : AOI211_X1 port map( C1 => n568, C2 => n12008, A => RST, B => n12009
                           , ZN => n7127);
   U15834 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_26_port, C2 => 
                           n12009, A => n12012, B => n8692, ZN => n12010);
   U15835 : INV_X1 port map( A => n12010, ZN => n7126);
   U15836 : AOI211_X1 port map( C1 => n570, C2 => n12012, A => RST, B => n12011
                           , ZN => n7125);
   U15837 : AOI211_X1 port map( C1 => n571, C2 => n12013, A => RST, B => n12014
                           , ZN => n7124);
   U15838 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_29_port, C2 => 
                           n12014, A => n12016, B => n8690, ZN => n3280);
   U15839 : AOI211_X1 port map( C1 => n572, C2 => n12016, A => RST, B => n12015
                           , ZN => n7123);
   U15840 : AOI22_X1 port map( A1 => n8652, A2 => 
                           DataPath_RF_bus_reg_dataout_31_port, B1 => n12017, 
                           B2 => n8653, ZN => n3274);
   U15841 : INV_X1 port map( A => IRAM_DATA(26), ZN => n12019);
   U15842 : INV_X1 port map( A => IRAM_READY, ZN => n12020);
   U15843 : INV_X1 port map( A => IRAM_DATA(30), ZN => n12021);
   U15844 : AOI22_X1 port map( A1 => n10857, A2 => CU_I_CW_ID_6_port, B1 => 
                           n10851, B2 => CU_I_CW_EX_6_port, ZN => n2992);
   U15845 : AOI22_X1 port map( A1 => n10857, A2 => CU_I_CW_ID_0_port, B1 => 
                           n10851, B2 => CU_I_CW_EX_0_port, ZN => n2962);
   U15846 : AOI22_X1 port map( A1 => n10857, A2 => CU_I_CW_ID_1_port, B1 => 
                           n10851, B2 => CU_I_CW_EX_1_port, ZN => n2961);
   U15847 : AOI22_X1 port map( A1 => n10857, A2 => CU_I_CW_ID_2_port, B1 => 
                           n10851, B2 => CU_I_CW_EX_2_port, ZN => n2960);
   U15848 : AOI22_X1 port map( A1 => n10857, A2 => CU_I_CW_ID_3_port, B1 => 
                           n10851, B2 => CU_I_CW_EX_3_port, ZN => n2959);
   U15849 : AOI22_X1 port map( A1 => n10857, A2 => CU_I_CW_ID_4_port, B1 => 
                           n10851, B2 => CU_I_CW_EX_4_port, ZN => n2958);
   U15850 : AOI22_X1 port map( A1 => n10857, A2 => CU_I_CW_ID_5_port, B1 => 
                           n10851, B2 => CU_I_CW_EX_5_port, ZN => n2957);
   U15851 : AOI22_X1 port map( A1 => n10857, A2 => CU_I_CW_EX_0_port, B1 => 
                           n10851, B2 => CU_I_CW_MEM_0_port, ZN => n2956);
   U15852 : AOI22_X1 port map( A1 => n10857, A2 => CU_I_CW_EX_1_port, B1 => 
                           n10851, B2 => CU_I_CW_MEM_1_port, ZN => n2955);
   U15853 : OAI21_X1 port map( B1 => n7768, B2 => CU_I_CW_EX_2_port, A => n8695
                           , ZN => n2953);
   U15854 : NAND2_X1 port map( A1 => IR_1_port, A2 => IR_2_port, ZN => n12029);
   U15855 : NAND2_X1 port map( A1 => IR_2_port, A2 => n210, ZN => n12025);
   U15856 : AOI22_X1 port map( A1 => n8062, A2 => n10850, B1 => i_ALU_OP_0_port
                           , B2 => n10851, ZN => n12023);
   U15857 : OAI211_X1 port map( C1 => n12024, C2 => n12027, A => n10849, B => 
                           n12023, ZN => n7087);
   U15858 : NOR2_X1 port map( A1 => IR_1_port, A2 => IR_2_port, ZN => n12028);
   U15859 : INV_X1 port map( A => CU_I_CW_ID_16, ZN => n12030);
   U15860 : NAND2_X1 port map( A1 => n10857, A2 => CU_I_CW_ID_17, ZN => n12031)
                           ;
   U15861 : OAI21_X1 port map( B1 => n12032, B2 => n8674, A => n12031, ZN => 
                           n7077);
   U15862 : AOI22_X1 port map( A1 => n10857, A2 => CU_I_CW_ID_18, B1 => 
                           CU_I_CW_EX_18, B2 => n10851, ZN => n2887);
   U15863 : AOI22_X1 port map( A1 => n10848, A2 => 
                           DataPath_i_PIPLIN_WRB1_0_port, B1 => n7764, B2 => 
                           DataPath_i_PIPLIN_WRB2_0_port, ZN => n2886);
   U15864 : AOI22_X1 port map( A1 => n10848, A2 => 
                           DataPath_i_PIPLIN_WRB1_1_port, B1 => n7764, B2 => 
                           DataPath_i_PIPLIN_WRB2_1_port, ZN => n2885);
   U15865 : AOI22_X1 port map( A1 => n10848, A2 => 
                           DataPath_i_PIPLIN_WRB1_2_port, B1 => n7782, B2 => 
                           DataPath_i_PIPLIN_WRB2_2_port, ZN => n2884);
   U15866 : AOI22_X1 port map( A1 => n10848, A2 => 
                           DataPath_i_PIPLIN_WRB1_3_port, B1 => n7764, B2 => 
                           DataPath_i_PIPLIN_WRB2_3_port, ZN => n2883);
   U15867 : AOI22_X1 port map( A1 => n10848, A2 => 
                           DataPath_i_PIPLIN_WRB1_4_port, B1 => n7764, B2 => 
                           DataPath_i_PIPLIN_WRB2_4_port, ZN => n2882);
   U15868 : AOI22_X1 port map( A1 => CU_I_CW_ID_22, A2 => n10857, B1 => n10851,
                           B2 => CU_I_unsigned_1, ZN => n2876);
   U15869 : AOI22_X1 port map( A1 => n10857, A2 => CU_I_unsigned_1, B1 => 
                           i_UNSIG_SIGN_N, B2 => n10851, ZN => n2874);
   U15870 : AOI22_X1 port map( A1 => i_RD2_0_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_B_0_port, ZN => n2873);
   U15871 : AOI22_X1 port map( A1 => i_RD2_1_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_B_1_port, ZN => n2872);
   U15872 : AOI22_X1 port map( A1 => i_RD2_2_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_B_2_port, ZN => n2871);
   U15873 : AOI22_X1 port map( A1 => i_RD2_3_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_B_3_port, ZN => n2870);
   U15874 : AOI22_X1 port map( A1 => i_RD2_4_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_B_4_port, ZN => n2869);
   U15875 : AOI22_X1 port map( A1 => i_RD2_5_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_B_5_port, ZN => n2868);
   U15876 : AOI22_X1 port map( A1 => i_RD2_6_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_B_6_port, ZN => n12033);
   U15877 : INV_X1 port map( A => n12033, ZN => n7076);
   U15878 : AOI22_X1 port map( A1 => i_RD2_7_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_B_7_port, ZN => n2867);
   U15879 : AOI22_X1 port map( A1 => i_RD2_8_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_B_8_port, ZN => n2866);
   U15880 : AOI22_X1 port map( A1 => i_RD2_9_port, A2 => n10872, B1 => n10871, 
                           B2 => DataPath_i_PIPLIN_B_9_port, ZN => n2865);
   U15881 : AOI22_X1 port map( A1 => i_RD2_10_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_10_port, ZN => n2864);
   U15882 : AOI22_X1 port map( A1 => i_RD2_11_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_11_port, ZN => n2863);
   U15883 : AOI22_X1 port map( A1 => i_RD2_12_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_12_port, ZN => n2862);
   U15884 : AOI22_X1 port map( A1 => i_RD2_13_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_13_port, ZN => n2861);
   U15885 : AOI22_X1 port map( A1 => i_RD2_14_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_14_port, ZN => n2860);
   U15886 : AOI22_X1 port map( A1 => i_RD2_15_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_15_port, ZN => n2859);
   U15887 : AOI22_X1 port map( A1 => i_RD2_16_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_16_port, ZN => n12034);
   U15888 : INV_X1 port map( A => n12034, ZN => n7075);
   U15889 : AOI22_X1 port map( A1 => i_RD2_17_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_17_port, ZN => n2858);
   U15890 : AOI22_X1 port map( A1 => i_RD2_18_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_18_port, ZN => n2857);
   U15891 : AOI22_X1 port map( A1 => i_RD2_19_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_19_port, ZN => n2856);
   U15892 : AOI22_X1 port map( A1 => i_RD2_20_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_20_port, ZN => n2855);
   U15893 : AOI22_X1 port map( A1 => i_RD2_21_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_21_port, ZN => n2854);
   U15894 : AOI22_X1 port map( A1 => i_RD2_22_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_22_port, ZN => n2853);
   U15895 : AOI22_X1 port map( A1 => i_RD2_23_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_23_port, ZN => n2852);
   U15896 : AOI22_X1 port map( A1 => i_RD2_24_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_24_port, ZN => n2851);
   U15897 : AOI22_X1 port map( A1 => i_RD2_25_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_25_port, ZN => n2850);
   U15898 : AOI22_X1 port map( A1 => i_RD2_26_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_26_port, ZN => n2849);
   U15899 : AOI22_X1 port map( A1 => i_RD2_27_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_27_port, ZN => n2848);
   U15900 : AOI22_X1 port map( A1 => i_RD2_28_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_28_port, ZN => n2847);
   U15901 : AOI22_X1 port map( A1 => i_RD2_29_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_29_port, ZN => n2846);
   U15902 : AOI22_X1 port map( A1 => i_RD2_30_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_30_port, ZN => n2845);
   U15903 : AOI22_X1 port map( A1 => i_RD2_31_port, A2 => n10872, B1 => n10871,
                           B2 => DataPath_i_PIPLIN_B_31_port, ZN => n2844);
   U15904 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_0_port, 
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_0_port, ZN => n2843);
   U15905 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_1_port, 
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_1_port, ZN => n2842);
   U15906 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_2_port, 
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_2_port, ZN => n2841);
   U15907 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_3_port, 
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_3_port, ZN => n2840);
   U15908 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_4_port, 
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_4_port, ZN => n2839);
   U15909 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_5_port, 
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_5_port, ZN => n2838);
   U15910 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_6_port, 
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_6_port, ZN => n12035)
                           ;
   U15911 : INV_X1 port map( A => n12035, ZN => n7074);
   U15912 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_7_port, 
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_7_port, ZN => n2837);
   U15913 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_8_port, 
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_8_port, ZN => n2836);
   U15914 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_9_port, 
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_9_port, ZN => n2835);
   U15915 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_10_port,
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_10_port, ZN => n2834)
                           ;
   U15916 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_11_port,
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_11_port, ZN => n2833)
                           ;
   U15917 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_12_port,
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_12_port, ZN => n2832)
                           ;
   U15918 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_13_port,
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_13_port, ZN => n2831)
                           ;
   U15919 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_14_port,
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_14_port, ZN => n2830)
                           ;
   U15920 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_15_port,
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_15_port, ZN => n2829)
                           ;
   U15921 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_16_port,
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_16_port, ZN => n2828)
                           ;
   U15922 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_17_port,
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_17_port, ZN => n2827)
                           ;
   U15923 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_18_port,
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_18_port, ZN => n2826)
                           ;
   U15924 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_19_port,
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_19_port, ZN => n2825)
                           ;
   U15925 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_20_port,
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_20_port, ZN => n2824)
                           ;
   U15926 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_21_port,
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_21_port, ZN => n2823)
                           ;
   U15927 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_22_port,
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_22_port, ZN => n2822)
                           ;
   U15928 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_23_port,
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_23_port, ZN => n2821)
                           ;
   U15929 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_24_port,
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_24_port, ZN => n2820)
                           ;
   U15930 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_25_port,
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_25_port, ZN => n2819)
                           ;
   U15931 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_26_port,
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_26_port, ZN => n2818)
                           ;
   U15932 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_27_port,
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_27_port, ZN => n2817)
                           ;
   U15933 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_28_port,
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_28_port, ZN => n2816)
                           ;
   U15934 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_29_port,
                           B1 => n7782, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_29_port, ZN => n2815)
                           ;
   U15935 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_30_port,
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_30_port, ZN => n2814)
                           ;
   U15936 : AOI22_X1 port map( A1 => n10848, A2 => DataPath_i_PIPLIN_B_31_port,
                           B1 => n7764, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_31_port, ZN => n2813)
                           ;
   U15937 : NOR2_X1 port map( A1 => n12043, A2 => n12042, ZN => n12041);
   U15938 : AOI22_X1 port map( A1 => DataPath_RF_c_win_1_port, A2 => n12042, B1
                           => DataPath_RF_c_win_0_port, B2 => n12041, ZN => 
                           n12036);
   U15939 : OAI211_X1 port map( C1 => n8441, C2 => n12037, A => n12036, B => 
                           n8694, ZN => n7073);
   U15940 : NOR2_X1 port map( A1 => RST, A2 => n12038, ZN => n7072);
   U15941 : AOI222_X1 port map( A1 => DataPath_RF_c_win_3_port, A2 => n12042, 
                           B1 => DataPath_RF_c_win_2_port, B2 => n12041, C1 => 
                           DataPath_RF_c_win_1_port, C2 => n12043, ZN => n12039
                           );
   U15942 : NOR2_X1 port map( A1 => RST, A2 => n12039, ZN => n7071);
   U15943 : AOI222_X1 port map( A1 => DataPath_RF_c_win_3_port, A2 => n12041, 
                           B1 => n12043, B2 => DataPath_RF_c_win_2_port, C1 => 
                           n8678, C2 => n12042, ZN => n12040);
   U15944 : NOR2_X1 port map( A1 => RST, A2 => n12040, ZN => n7070);
   U15945 : AOI222_X1 port map( A1 => DataPath_RF_c_win_3_port, A2 => n12043, 
                           B1 => n12042, B2 => DataPath_RF_c_win_0_port, C1 => 
                           n8678, C2 => n12041, ZN => n12044);
   U15946 : NOR2_X1 port map( A1 => RST, A2 => n12044, ZN => n7069);
   U15947 : NAND2_X1 port map( A1 => n12208, A2 => n10846, ZN => n12049);
   U15948 : AOI21_X1 port map( B1 => n10852, B2 => n12047, A => n12208, ZN => 
                           n12055);
   U15949 : INV_X1 port map( A => n12049, ZN => n12054);
   U15950 : NOR2_X1 port map( A1 => n12055, A2 => n12054, ZN => n12053);
   U15951 : AOI22_X1 port map( A1 => DataPath_RF_c_swin_0_port, A2 => n12053, 
                           B1 => n12055, B2 => DataPath_RF_c_swin_4_port, ZN =>
                           n12048);
   U15952 : OAI211_X1 port map( C1 => n821, C2 => n12049, A => n12048, B => 
                           n8691, ZN => n7066);
   U15953 : AOI222_X1 port map( A1 => DataPath_RF_c_swin_1_port, A2 => n12053, 
                           B1 => DataPath_RF_c_swin_0_port, B2 => n12055, C1 =>
                           DataPath_RF_c_swin_2_port, C2 => n12054, ZN => 
                           n12050);
   U15954 : NOR2_X1 port map( A1 => RST, A2 => n12050, ZN => n7065);
   U15955 : AOI222_X1 port map( A1 => DataPath_RF_c_swin_2_port, A2 => n12053, 
                           B1 => DataPath_RF_c_swin_1_port, B2 => n12055, C1 =>
                           DataPath_RF_c_swin_3_port, C2 => n12054, ZN => 
                           n12051);
   U15956 : NOR2_X1 port map( A1 => RST, A2 => n12051, ZN => n7064);
   U15957 : AOI222_X1 port map( A1 => DataPath_RF_c_swin_2_port, A2 => n12055, 
                           B1 => DataPath_RF_c_swin_3_port, B2 => n12053, C1 =>
                           DataPath_RF_c_swin_4_port, C2 => n12054, ZN => 
                           n12052);
   U15958 : NOR2_X1 port map( A1 => RST, A2 => n12052, ZN => n7063);
   U15959 : AOI222_X1 port map( A1 => DataPath_RF_c_swin_3_port, A2 => n12055, 
                           B1 => DataPath_RF_c_swin_0_port, B2 => n12054, C1 =>
                           DataPath_RF_c_swin_4_port, C2 => n12053, ZN => 
                           n12056);
   U15960 : NOR2_X1 port map( A1 => RST, A2 => n12056, ZN => n7062);
   U15961 : AOI221_X1 port map( B1 => n12059, B2 => n10844, C1 => n12058, C2 =>
                           n10844, A => RST, ZN => n7061);
   U15962 : INV_X1 port map( A => i_RD1_1_port, ZN => n12060);
   U15963 : INV_X1 port map( A => i_RD1_8_port, ZN => n12062);
   U15964 : OAI21_X1 port map( B1 => n12062, B2 => n8549, A => n12061, ZN => 
                           n7051);
   U15965 : OAI21_X1 port map( B1 => n7759, B2 => n12064, A => n12063, ZN => 
                           n7050);
   U15966 : OAI21_X1 port map( B1 => n12067, B2 => n7759, A => n12066, ZN => 
                           n7041);
   U15967 : OAI21_X1 port map( B1 => n7759, B2 => n12069, A => n12068, ZN => 
                           n7040);
   U15968 : NOR2_X1 port map( A1 => n8319, A2 => n368, ZN => n12074);
   U15969 : NAND2_X1 port map( A1 => n8681, A2 => n368, ZN => n12088);
   U15970 : NOR2_X1 port map( A1 => n8319, A2 => n12091, ZN => n12072);
   U15971 : NOR2_X1 port map( A1 => n8681, A2 => n368, ZN => n12071);
   U15972 : INV_X1 port map( A => n12071, ZN => n12073);
   U15973 : NOR2_X1 port map( A1 => n12074, A2 => n12071, ZN => n12085);
   U15974 : NAND2_X1 port map( A1 => n8300, A2 => n12087, ZN => n12081);
   U15975 : INV_X1 port map( A => n12081, ZN => n12082);
   U15976 : INV_X1 port map( A => n12085, ZN => n12086);
   U15977 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_0_port, B1 => 
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_0_port, ZN => 
                           n2318);
   U15978 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_1_port, B1 => 
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_1_port, ZN => 
                           n2317);
   U15979 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_2_port, B1 => 
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_2_port, ZN => 
                           n2316);
   U15980 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_3_port, B1 => 
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_3_port, ZN => 
                           n2315);
   U15981 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_4_port, B1 => 
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_4_port, ZN => 
                           n2314);
   U15982 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_5_port, B1 => 
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_5_port, ZN => 
                           n2313);
   U15983 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_6_port, B1 => 
                           n12204, B2 => DataPath_i_REG_LDSTR_OUT_6_port, ZN =>
                           n2312);
   U15984 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_7_port, B1 => 
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_7_port, ZN => 
                           n2311);
   U15985 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_8_port, B1 => 
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_8_port, ZN => 
                           n2310);
   U15986 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_9_port, B1 => 
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_9_port, ZN => 
                           n2309);
   U15987 : AOI22_X1 port map( A1 => n8670, A2 => DRAM_DATA_OUT_10_port, B1 => 
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_10_port, ZN =>
                           n2308);
   U15988 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_11_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_11_port, ZN =>
                           n2307);
   U15989 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_12_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_12_port, ZN =>
                           n2306);
   U15990 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_13_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_13_port, ZN =>
                           n2305);
   U15991 : AOI22_X1 port map( A1 => n8670, A2 => DRAM_DATA_OUT_14_port, B1 => 
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_14_port, ZN =>
                           n2304);
   U15992 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_15_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_15_port, ZN =>
                           n2303);
   U15993 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_16_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_16_port, ZN =>
                           n2302);
   U15994 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_17_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_17_port, ZN =>
                           n2301);
   U15995 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_18_port, B1 =>
                           n12204, B2 => DataPath_i_REG_LDSTR_OUT_18_port, ZN 
                           => n2300);
   U15996 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_19_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_19_port, ZN =>
                           n2299);
   U15997 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_20_port, B1 =>
                           n12204, B2 => DataPath_i_REG_LDSTR_OUT_20_port, ZN 
                           => n2298);
   U15998 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_21_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_21_port, ZN =>
                           n2297);
   U15999 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_22_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_22_port, ZN =>
                           n2296);
   U16000 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_23_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_23_port, ZN =>
                           n2295);
   U16001 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_24_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_24_port, ZN =>
                           n2294);
   U16002 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_25_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_25_port, ZN =>
                           n2293);
   U16003 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_26_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_26_port, ZN =>
                           n2292);
   U16004 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_27_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_27_port, ZN =>
                           n2291);
   U16005 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_28_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_28_port, ZN =>
                           n2290);
   U16006 : AOI22_X1 port map( A1 => n8670, A2 => DRAM_DATA_OUT_29_port, B1 => 
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_29_port, ZN =>
                           n2289);
   U16007 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_30_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_30_port, ZN =>
                           n2288);
   U16008 : AOI22_X1 port map( A1 => n12203, A2 => DRAM_DATA_OUT_31_port, B1 =>
                           n7765, B2 => DataPath_i_REG_LDSTR_OUT_31_port, ZN =>
                           n2287);
   U16009 : NAND3_X1 port map( A1 => n12077, A2 => n12076, A3 => n12075, ZN => 
                           n12078);
   U16010 : AOI222_X1 port map( A1 => n12079, A2 => n10841, B1 => n7764, B2 => 
                           DRAM_ADDRESS_2_port, C1 => n12078, C2 => n10840, ZN 
                           => n2260);
   U16011 : NAND2_X1 port map( A1 => i_ALU_OP_3_port, A2 => n10869, ZN => 
                           n12090);
   U16012 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_0_port, A2 => 
                           n7765, B1 => n12203, B2 => n8388, ZN => n1258);
   U16013 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_1_port, A2 => 
                           n12204, B1 => n12203, B2 => n8376, ZN => n1257);
   U16014 : AOI22_X1 port map( A1 => n8670, A2 => DRAM_ADDRESS_2_port, B1 => 
                           n7765, B2 => DataPath_i_REG_MEM_ALUOUT_2_port, ZN =>
                           n1256);
   U16015 : AOI22_X1 port map( A1 => DRAM_ADDRESS_3_port, A2 => n8670, B1 => 
                           n7765, B2 => DataPath_i_REG_MEM_ALUOUT_3_port, ZN =>
                           n1255);
   U16016 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_4_port, A2 => 
                           n7765, B1 => n12203, B2 => DRAM_ADDRESS_4_port, ZN 
                           => n1254);
   U16017 : AOI22_X1 port map( A1 => n8670, A2 => DRAM_ADDRESS_5_port, B1 => 
                           n7765, B2 => DataPath_i_REG_MEM_ALUOUT_5_port, ZN =>
                           n1253);
   U16018 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_6_port, A2 => 
                           n12204, B1 => n12203, B2 => DRAM_ADDRESS_6_port, ZN 
                           => n1252);
   U16019 : AOI22_X1 port map( A1 => DRAM_ADDRESS_7_port, A2 => n8670, B1 => 
                           n7765, B2 => DataPath_i_REG_MEM_ALUOUT_7_port, ZN =>
                           n1251);
   U16020 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_8_port, A2 => 
                           n12204, B1 => n8670, B2 => DRAM_ADDRESS_8_port, ZN 
                           => n1250);
   U16021 : AOI22_X1 port map( A1 => DRAM_ADDRESS_9_port, A2 => n8670, B1 => 
                           n7765, B2 => DataPath_i_REG_MEM_ALUOUT_9_port, ZN =>
                           n1249);
   U16022 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_10_port, A2 => 
                           n7765, B1 => n8670, B2 => DRAM_ADDRESS_10_port, ZN 
                           => n1248);
   U16023 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_11_port, A2 => 
                           n7765, B1 => n8670, B2 => DRAM_ADDRESS_11_port, ZN 
                           => n1247);
   U16024 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_12_port, A2 => 
                           n7765, B1 => n8670, B2 => DRAM_ADDRESS_12_port, ZN 
                           => n1246);
   U16025 : AOI22_X1 port map( A1 => DRAM_ADDRESS_13_port, A2 => n8670, B1 => 
                           n7765, B2 => DataPath_i_REG_MEM_ALUOUT_13_port, ZN 
                           => n1245);
   U16026 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_14_port, A2 => 
                           n12204, B1 => n8670, B2 => DRAM_ADDRESS_14_port, ZN 
                           => n1244);
   U16027 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_15_port, A2 => 
                           n7765, B1 => n12203, B2 => DRAM_ADDRESS_15_port, ZN 
                           => n1243);
   U16028 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_16_port, A2 => 
                           n12204, B1 => n8670, B2 => DRAM_ADDRESS_16_port, ZN 
                           => n1242);
   U16029 : AOI22_X1 port map( A1 => DRAM_ADDRESS_17_port, A2 => n8670, B1 => 
                           n7765, B2 => DataPath_i_REG_MEM_ALUOUT_17_port, ZN 
                           => n1241);
   U16030 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_18_port, A2 => 
                           n12204, B1 => n8670, B2 => DRAM_ADDRESS_18_port, ZN 
                           => n1240);
   U16031 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_19_port, A2 => 
                           n12204, B1 => n8670, B2 => DRAM_ADDRESS_19_port, ZN 
                           => n1239);
   U16032 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_20_port, A2 => 
                           n7765, B1 => n12203, B2 => DRAM_ADDRESS_20_port, ZN 
                           => n1238);
   U16033 : AOI22_X1 port map( A1 => DRAM_ADDRESS_21_port, A2 => n8670, B1 => 
                           n7765, B2 => DataPath_i_REG_MEM_ALUOUT_21_port, ZN 
                           => n1237);
   U16034 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_22_port, A2 => 
                           n7765, B1 => n8670, B2 => DRAM_ADDRESS_22_port, ZN 
                           => n1236);
   U16035 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_23_port, A2 => 
                           n7765, B1 => n8670, B2 => DRAM_ADDRESS_23_port, ZN 
                           => n1235);
   U16036 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_24_port, A2 => 
                           n7765, B1 => n12203, B2 => DRAM_ADDRESS_24_port, ZN 
                           => n1234);
   U16037 : AOI22_X1 port map( A1 => DRAM_ADDRESS_25_port, A2 => n8670, B1 => 
                           n7765, B2 => DataPath_i_REG_MEM_ALUOUT_25_port, ZN 
                           => n1233);
   U16038 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_26_port, A2 => 
                           n7765, B1 => n12203, B2 => DRAM_ADDRESS_26_port, ZN 
                           => n1232);
   U16039 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_27_port, A2 => 
                           n7765, B1 => n12203, B2 => DRAM_ADDRESS_27_port, ZN 
                           => n1231);
   U16040 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_28_port, A2 => 
                           n7765, B1 => n12203, B2 => DRAM_ADDRESS_28_port, ZN 
                           => n1230);
   U16041 : AOI22_X1 port map( A1 => DRAM_ADDRESS_29_port, A2 => n8670, B1 => 
                           n7765, B2 => DataPath_i_REG_MEM_ALUOUT_29_port, ZN 
                           => n1229);
   U16042 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_30_port, A2 => 
                           n7765, B1 => n12203, B2 => DRAM_ADDRESS_30_port, ZN 
                           => n1228);
   U16043 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_31_port, A2 => 
                           n7765, B1 => n12203, B2 => DRAM_ADDRESS_31_port, ZN 
                           => n1225);
   U16044 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2528_port, B1 => n12106,
                           B2 => n12122, ZN => n1221);
   U16045 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2529_port, B1 => n12106,
                           B2 => n12123, ZN => n1220);
   U16046 : AOI22_X1 port map( A1 => n12108, A2 => 
                           DataPath_RF_bus_reg_dataout_2530_port, B1 => n12106,
                           B2 => n12124, ZN => n1219);
   U16047 : AOI22_X1 port map( A1 => n12108, A2 => 
                           DataPath_RF_bus_reg_dataout_2531_port, B1 => n12106,
                           B2 => n12125, ZN => n1218);
   U16048 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2532_port, B1 => n12106,
                           B2 => n12126, ZN => n1217);
   U16049 : OAI22_X1 port map( A1 => n12108, A2 => n12182, B1 => 
                           DataPath_RF_bus_reg_dataout_2533_port, B2 => n12107,
                           ZN => n1216);
   U16050 : AOI22_X1 port map( A1 => n12108, A2 => 
                           DataPath_RF_bus_reg_dataout_2534_port, B1 => n12106,
                           B2 => n12128, ZN => n1215);
   U16051 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2535_port, B1 => n12106,
                           B2 => n12129, ZN => n1214);
   U16052 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2536_port, B1 => n12106,
                           B2 => n12130, ZN => n1213);
   U16053 : AOI22_X1 port map( A1 => n12108, A2 => 
                           DataPath_RF_bus_reg_dataout_2537_port, B1 => n12106,
                           B2 => n12131, ZN => n1212);
   U16054 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2538_port, B1 => n12106,
                           B2 => n12132, ZN => n1211);
   U16055 : AOI22_X1 port map( A1 => n12108, A2 => 
                           DataPath_RF_bus_reg_dataout_2539_port, B1 => n12106,
                           B2 => n12133, ZN => n1210);
   U16056 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2540_port, B1 => n12106,
                           B2 => n12134, ZN => n1209);
   U16057 : AOI22_X1 port map( A1 => n12108, A2 => 
                           DataPath_RF_bus_reg_dataout_2541_port, B1 => n12106,
                           B2 => n12135, ZN => n1208);
   U16058 : OAI22_X1 port map( A1 => n12108, A2 => n12191, B1 => 
                           DataPath_RF_bus_reg_dataout_2542_port, B2 => n12107,
                           ZN => n1207);
   U16059 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2543_port, B1 => n12106,
                           B2 => n12136, ZN => n1206);
   U16060 : OAI22_X1 port map( A1 => n12108, A2 => n12159, B1 => 
                           DataPath_RF_bus_reg_dataout_2544_port, B2 => n12107,
                           ZN => n1205);
   U16061 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2545_port, B1 => n12106,
                           B2 => n12137, ZN => n1204);
   U16062 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2546_port, B1 => n12106,
                           B2 => n12138, ZN => n1203);
   U16063 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2547_port, B1 => n12106,
                           B2 => n12139, ZN => n1202);
   U16064 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2548_port, B1 => n12106,
                           B2 => n12101, ZN => n1201);
   U16065 : OAI22_X1 port map( A1 => n12108, A2 => n12164, B1 => 
                           DataPath_RF_bus_reg_dataout_2549_port, B2 => n12107,
                           ZN => n1200);
   U16066 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2550_port, B1 => n12106,
                           B2 => n12142, ZN => n1199);
   U16067 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2551_port, A2 
                           => n8654, B1 => n12166, B2 => n12107, ZN => n1198);
   U16068 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2552_port, B1 => n12106,
                           B2 => n12144, ZN => n1197);
   U16069 : OAI22_X1 port map( A1 => n12108, A2 => n12168, B1 => 
                           DataPath_RF_bus_reg_dataout_2553_port, B2 => n12107,
                           ZN => n1196);
   U16070 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2554_port, A2 
                           => n8654, B1 => n12169, B2 => n12107, ZN => n1195);
   U16071 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2555_port, B1 => n12106,
                           B2 => n12148, ZN => n1194);
   U16072 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2556_port, B1 => n12106,
                           B2 => n12149, ZN => n1193);
   U16073 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2557_port, B1 => n12106,
                           B2 => n12150, ZN => n1192);
   U16074 : AOI22_X1 port map( A1 => n8654, A2 => 
                           DataPath_RF_bus_reg_dataout_2558_port, B1 => n12106,
                           B2 => n12151, ZN => n1191);
   U16075 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2559_port, A2 
                           => n8654, B1 => n12107, B2 => n12175, ZN => n1188);
   U16076 : OAI22_X1 port map( A1 => n12177, A2 => n8656, B1 => 
                           DataPath_RF_bus_reg_dataout_2496_port, B2 => n8655, 
                           ZN => n1184);
   U16077 : OAI22_X1 port map( A1 => n12111, A2 => n12178, B1 => 
                           DataPath_RF_bus_reg_dataout_2497_port, B2 => n8655, 
                           ZN => n1183);
   U16078 : OAI22_X1 port map( A1 => n8656, A2 => n12179, B1 => 
                           DataPath_RF_bus_reg_dataout_2498_port, B2 => n12110,
                           ZN => n1182);
   U16079 : OAI22_X1 port map( A1 => n8656, A2 => n12180, B1 => 
                           DataPath_RF_bus_reg_dataout_2499_port, B2 => n12110,
                           ZN => n1181);
   U16080 : OAI22_X1 port map( A1 => n8656, A2 => n12181, B1 => 
                           DataPath_RF_bus_reg_dataout_2500_port, B2 => n12110,
                           ZN => n1180);
   U16081 : OAI22_X1 port map( A1 => n12182, A2 => n12111, B1 => 
                           DataPath_RF_bus_reg_dataout_2501_port, B2 => n12110,
                           ZN => n1179);
   U16082 : OAI22_X1 port map( A1 => n8656, A2 => n12183, B1 => 
                           DataPath_RF_bus_reg_dataout_2502_port, B2 => n12110,
                           ZN => n1178);
   U16083 : OAI22_X1 port map( A1 => n12111, A2 => n12184, B1 => 
                           DataPath_RF_bus_reg_dataout_2503_port, B2 => n8655, 
                           ZN => n1177);
   U16084 : OAI22_X1 port map( A1 => n8656, A2 => n12185, B1 => 
                           DataPath_RF_bus_reg_dataout_2504_port, B2 => n12110,
                           ZN => n1176);
   U16085 : OAI22_X1 port map( A1 => n8656, A2 => n12186, B1 => 
                           DataPath_RF_bus_reg_dataout_2505_port, B2 => n12110,
                           ZN => n1175);
   U16086 : OAI22_X1 port map( A1 => n12111, A2 => n12187, B1 => 
                           DataPath_RF_bus_reg_dataout_2506_port, B2 => n12110,
                           ZN => n1174);
   U16087 : OAI22_X1 port map( A1 => n12111, A2 => n12188, B1 => 
                           DataPath_RF_bus_reg_dataout_2507_port, B2 => n8655, 
                           ZN => n1173);
   U16088 : OAI22_X1 port map( A1 => n8656, A2 => n12189, B1 => 
                           DataPath_RF_bus_reg_dataout_2508_port, B2 => n12110,
                           ZN => n1172);
   U16089 : OAI22_X1 port map( A1 => n12111, A2 => n12190, B1 => 
                           DataPath_RF_bus_reg_dataout_2509_port, B2 => n8655, 
                           ZN => n1171);
   U16090 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2510_port, A2 
                           => n8656, B1 => n12191, B2 => n8655, ZN => n1170);
   U16091 : OAI22_X1 port map( A1 => n8656, A2 => n12192, B1 => 
                           DataPath_RF_bus_reg_dataout_2511_port, B2 => n8655, 
                           ZN => n1169);
   U16092 : OAI22_X1 port map( A1 => n12159, A2 => n8656, B1 => 
                           DataPath_RF_bus_reg_dataout_2512_port, B2 => n12110,
                           ZN => n1168);
   U16093 : OAI22_X1 port map( A1 => n8656, A2 => n12160, B1 => 
                           DataPath_RF_bus_reg_dataout_2513_port, B2 => n8655, 
                           ZN => n1167);
   U16094 : OAI22_X1 port map( A1 => n8656, A2 => n12161, B1 => 
                           DataPath_RF_bus_reg_dataout_2514_port, B2 => n8655, 
                           ZN => n1166);
   U16095 : OAI22_X1 port map( A1 => n12111, A2 => n12162, B1 => 
                           DataPath_RF_bus_reg_dataout_2515_port, B2 => n8655, 
                           ZN => n1165);
   U16096 : OAI22_X1 port map( A1 => n8656, A2 => n12163, B1 => 
                           DataPath_RF_bus_reg_dataout_2516_port, B2 => n8655, 
                           ZN => n1164);
   U16097 : OAI22_X1 port map( A1 => n12164, A2 => n12111, B1 => 
                           DataPath_RF_bus_reg_dataout_2517_port, B2 => n8655, 
                           ZN => n1163);
   U16098 : OAI22_X1 port map( A1 => n8656, A2 => n12165, B1 => 
                           DataPath_RF_bus_reg_dataout_2518_port, B2 => n8655, 
                           ZN => n1162);
   U16099 : OAI22_X1 port map( A1 => n12166, A2 => n12111, B1 => 
                           DataPath_RF_bus_reg_dataout_2519_port, B2 => n8655, 
                           ZN => n1161);
   U16100 : OAI22_X1 port map( A1 => n8656, A2 => n12167, B1 => 
                           DataPath_RF_bus_reg_dataout_2520_port, B2 => n8655, 
                           ZN => n1160);
   U16101 : OAI22_X1 port map( A1 => n12168, A2 => n12111, B1 => 
                           DataPath_RF_bus_reg_dataout_2521_port, B2 => n8655, 
                           ZN => n1159);
   U16102 : OAI22_X1 port map( A1 => n12169, A2 => n12111, B1 => 
                           DataPath_RF_bus_reg_dataout_2522_port, B2 => n8655, 
                           ZN => n1158);
   U16103 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2523_port, A2 
                           => n8656, B1 => n12170, B2 => n8655, ZN => n1157);
   U16104 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2524_port, A2 
                           => n8656, B1 => n12171, B2 => n8655, ZN => n1156);
   U16105 : OAI22_X1 port map( A1 => n8656, A2 => n12172, B1 => 
                           DataPath_RF_bus_reg_dataout_2525_port, B2 => n8655, 
                           ZN => n1155);
   U16106 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2526_port, A2 
                           => n8656, B1 => n12173, B2 => n8655, ZN => n1154);
   U16107 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2527_port, A2 
                           => n8656, B1 => n12175, B2 => n8655, ZN => n1151);
   U16108 : AOI22_X1 port map( A1 => n12177, A2 => n8657, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2464_port, ZN => n1147);
   U16109 : AOI22_X1 port map( A1 => n12178, A2 => n8657, B1 => n12114, B2 => 
                           DataPath_RF_bus_reg_dataout_2465_port, ZN => n1146);
   U16110 : AOI22_X1 port map( A1 => n12179, A2 => n8657, B1 => n12114, B2 => 
                           DataPath_RF_bus_reg_dataout_2466_port, ZN => n1145);
   U16111 : AOI22_X1 port map( A1 => n12180, A2 => n8657, B1 => n12114, B2 => 
                           DataPath_RF_bus_reg_dataout_2467_port, ZN => n1144);
   U16112 : AOI22_X1 port map( A1 => n12181, A2 => n8657, B1 => n12114, B2 => 
                           DataPath_RF_bus_reg_dataout_2468_port, ZN => n1143);
   U16113 : AOI22_X1 port map( A1 => n12182, A2 => n8657, B1 => n12114, B2 => 
                           DataPath_RF_bus_reg_dataout_2469_port, ZN => n1142);
   U16114 : AOI22_X1 port map( A1 => n12183, A2 => n8657, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2470_port, ZN => n1141);
   U16115 : AOI22_X1 port map( A1 => n12184, A2 => n8657, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2471_port, ZN => n1140);
   U16116 : AOI22_X1 port map( A1 => n12185, A2 => n8657, B1 => n12114, B2 => 
                           DataPath_RF_bus_reg_dataout_2472_port, ZN => n1139);
   U16117 : AOI22_X1 port map( A1 => n12186, A2 => n8657, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2473_port, ZN => n1138);
   U16118 : AOI22_X1 port map( A1 => n12187, A2 => n12113, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2474_port, ZN => n1137);
   U16119 : AOI22_X1 port map( A1 => n12188, A2 => n8657, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2475_port, ZN => n1136);
   U16120 : AOI22_X1 port map( A1 => n12189, A2 => n8657, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2476_port, ZN => n1135);
   U16121 : AOI22_X1 port map( A1 => n12190, A2 => n8657, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2477_port, ZN => n1134);
   U16122 : OAI22_X1 port map( A1 => n8658, A2 => n12191, B1 => 
                           DataPath_RF_bus_reg_dataout_2478_port, B2 => n8657, 
                           ZN => n1133);
   U16123 : AOI22_X1 port map( A1 => n12192, A2 => n8657, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2479_port, ZN => n1132);
   U16124 : AOI22_X1 port map( A1 => n12159, A2 => n8657, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2480_port, ZN => n1131);
   U16125 : AOI22_X1 port map( A1 => n12160, A2 => n12113, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2481_port, ZN => n1130);
   U16126 : AOI22_X1 port map( A1 => n12161, A2 => n12113, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2482_port, ZN => n1129);
   U16127 : AOI22_X1 port map( A1 => n12162, A2 => n8657, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2483_port, ZN => n1128);
   U16128 : AOI22_X1 port map( A1 => n12163, A2 => n12113, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2484_port, ZN => n1127);
   U16129 : AOI22_X1 port map( A1 => n12164, A2 => n12113, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2485_port, ZN => n1126);
   U16130 : AOI22_X1 port map( A1 => n12165, A2 => n8657, B1 => n12114, B2 => 
                           DataPath_RF_bus_reg_dataout_2486_port, ZN => n1125);
   U16131 : AOI22_X1 port map( A1 => n12166, A2 => n8657, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2487_port, ZN => n1124);
   U16132 : AOI22_X1 port map( A1 => n12167, A2 => n12113, B1 => n12114, B2 => 
                           DataPath_RF_bus_reg_dataout_2488_port, ZN => n1123);
   U16133 : AOI22_X1 port map( A1 => n12168, A2 => n12113, B1 => n12114, B2 => 
                           DataPath_RF_bus_reg_dataout_2489_port, ZN => n1122);
   U16134 : AOI22_X1 port map( A1 => n12169, A2 => n8657, B1 => n12114, B2 => 
                           DataPath_RF_bus_reg_dataout_2490_port, ZN => n1121);
   U16135 : AOI22_X1 port map( A1 => n12170, A2 => n12113, B1 => n12114, B2 => 
                           DataPath_RF_bus_reg_dataout_2491_port, ZN => n1120);
   U16136 : AOI22_X1 port map( A1 => n12171, A2 => n8657, B1 => n12114, B2 => 
                           DataPath_RF_bus_reg_dataout_2492_port, ZN => n1119);
   U16137 : AOI22_X1 port map( A1 => n12172, A2 => n12113, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2493_port, ZN => n1118);
   U16138 : AOI22_X1 port map( A1 => n12173, A2 => n12113, B1 => n8658, B2 => 
                           DataPath_RF_bus_reg_dataout_2494_port, ZN => n1117);
   U16139 : OAI22_X1 port map( A1 => n8658, A2 => n12175, B1 => 
                           DataPath_RF_bus_reg_dataout_2495_port, B2 => n8657, 
                           ZN => n1114);
   U16140 : OAI22_X1 port map( A1 => n12177, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2432_port, B2 => n8659, 
                           ZN => n1110);
   U16141 : OAI22_X1 port map( A1 => n12178, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2433_port, B2 => n8659, 
                           ZN => n1109);
   U16142 : OAI22_X1 port map( A1 => n12179, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2434_port, B2 => n12116,
                           ZN => n1108);
   U16143 : OAI22_X1 port map( A1 => n12180, A2 => n12117, B1 => 
                           DataPath_RF_bus_reg_dataout_2435_port, B2 => n12116,
                           ZN => n1107);
   U16144 : OAI22_X1 port map( A1 => n12181, A2 => n12117, B1 => 
                           DataPath_RF_bus_reg_dataout_2436_port, B2 => n12116,
                           ZN => n1106);
   U16145 : OAI22_X1 port map( A1 => n12182, A2 => n12117, B1 => 
                           DataPath_RF_bus_reg_dataout_2437_port, B2 => n12116,
                           ZN => n1105);
   U16146 : OAI22_X1 port map( A1 => n12183, A2 => n12117, B1 => 
                           DataPath_RF_bus_reg_dataout_2438_port, B2 => n12116,
                           ZN => n1104);
   U16147 : OAI22_X1 port map( A1 => n12184, A2 => n12117, B1 => 
                           DataPath_RF_bus_reg_dataout_2439_port, B2 => n12116,
                           ZN => n1103);
   U16148 : OAI22_X1 port map( A1 => n12185, A2 => n12117, B1 => 
                           DataPath_RF_bus_reg_dataout_2440_port, B2 => n12116,
                           ZN => n1102);
   U16149 : OAI22_X1 port map( A1 => n12186, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2441_port, B2 => n12116,
                           ZN => n1101);
   U16150 : OAI22_X1 port map( A1 => n12187, A2 => n12117, B1 => 
                           DataPath_RF_bus_reg_dataout_2442_port, B2 => n12116,
                           ZN => n1100);
   U16151 : OAI22_X1 port map( A1 => n12188, A2 => n12117, B1 => 
                           DataPath_RF_bus_reg_dataout_2443_port, B2 => n8659, 
                           ZN => n1099);
   U16152 : OAI22_X1 port map( A1 => n12189, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2444_port, B2 => n8659, 
                           ZN => n1098);
   U16153 : OAI22_X1 port map( A1 => n12190, A2 => n12117, B1 => 
                           DataPath_RF_bus_reg_dataout_2445_port, B2 => n8659, 
                           ZN => n1097);
   U16154 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2446_port, A2 
                           => n8660, B1 => n12191, B2 => n8659, ZN => n1096);
   U16155 : OAI22_X1 port map( A1 => n12192, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2447_port, B2 => n8659, 
                           ZN => n1095);
   U16156 : OAI22_X1 port map( A1 => n12159, A2 => n12117, B1 => 
                           DataPath_RF_bus_reg_dataout_2448_port, B2 => n12116,
                           ZN => n1094);
   U16157 : OAI22_X1 port map( A1 => n12160, A2 => n12117, B1 => 
                           DataPath_RF_bus_reg_dataout_2449_port, B2 => n8659, 
                           ZN => n1093);
   U16158 : OAI22_X1 port map( A1 => n12161, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2450_port, B2 => n8659, 
                           ZN => n1092);
   U16159 : OAI22_X1 port map( A1 => n12162, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2451_port, B2 => n8659, 
                           ZN => n1091);
   U16160 : OAI22_X1 port map( A1 => n12163, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2452_port, B2 => n8659, 
                           ZN => n1090);
   U16161 : OAI22_X1 port map( A1 => n12164, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2453_port, B2 => n8659, 
                           ZN => n1089);
   U16162 : OAI22_X1 port map( A1 => n12165, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2454_port, B2 => n8659, 
                           ZN => n1088);
   U16163 : OAI22_X1 port map( A1 => n12166, A2 => n12117, B1 => 
                           DataPath_RF_bus_reg_dataout_2455_port, B2 => n8659, 
                           ZN => n1087);
   U16164 : OAI22_X1 port map( A1 => n12167, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2456_port, B2 => n8659, 
                           ZN => n1086);
   U16165 : OAI22_X1 port map( A1 => n12168, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2457_port, B2 => n8659, 
                           ZN => n1085);
   U16166 : OAI22_X1 port map( A1 => n12169, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2458_port, B2 => n8659, 
                           ZN => n1084);
   U16167 : OAI22_X1 port map( A1 => n12170, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2459_port, B2 => n8659, 
                           ZN => n1083);
   U16168 : OAI22_X1 port map( A1 => n12171, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2460_port, B2 => n8659, 
                           ZN => n1082);
   U16169 : OAI22_X1 port map( A1 => n12172, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2461_port, B2 => n8659, 
                           ZN => n1081);
   U16170 : OAI22_X1 port map( A1 => n12173, A2 => n8660, B1 => 
                           DataPath_RF_bus_reg_dataout_2462_port, B2 => n8659, 
                           ZN => n1080);
   U16171 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2463_port, A2 
                           => n8660, B1 => n12175, B2 => n8659, ZN => n1077);
   U16172 : OAI22_X1 port map( A1 => n12177, A2 => n8662, B1 => 
                           DataPath_RF_bus_reg_dataout_2400_port, B2 => n12119,
                           ZN => n1073);
   U16173 : OAI22_X1 port map( A1 => n12178, A2 => n12120, B1 => 
                           DataPath_RF_bus_reg_dataout_2401_port, B2 => n12119,
                           ZN => n1072);
   U16174 : OAI22_X1 port map( A1 => n12179, A2 => n8662, B1 => 
                           DataPath_RF_bus_reg_dataout_2402_port, B2 => n12119,
                           ZN => n1071);
   U16175 : OAI22_X1 port map( A1 => n12180, A2 => n8662, B1 => 
                           DataPath_RF_bus_reg_dataout_2403_port, B2 => n12119,
                           ZN => n1070);
   U16176 : OAI22_X1 port map( A1 => n12181, A2 => n12120, B1 => 
                           DataPath_RF_bus_reg_dataout_2404_port, B2 => n8661, 
                           ZN => n1069);
   U16177 : AOI22_X1 port map( A1 => n12182, A2 => n8661, B1 => n8662, B2 => 
                           DataPath_RF_bus_reg_dataout_2405_port, ZN => n1068);
   U16178 : AOI22_X1 port map( A1 => n12183, A2 => n8661, B1 => n8662, B2 => 
                           DataPath_RF_bus_reg_dataout_2406_port, ZN => n1067);
   U16179 : AOI22_X1 port map( A1 => n12184, A2 => n8661, B1 => n8662, B2 => 
                           DataPath_RF_bus_reg_dataout_2407_port, ZN => n1066);
   U16180 : AOI22_X1 port map( A1 => n12185, A2 => n8661, B1 => n8662, B2 => 
                           DataPath_RF_bus_reg_dataout_2408_port, ZN => n1065);
   U16181 : AOI22_X1 port map( A1 => n12186, A2 => n12119, B1 => n8662, B2 => 
                           DataPath_RF_bus_reg_dataout_2409_port, ZN => n1064);
   U16182 : OAI22_X1 port map( A1 => n12187, A2 => n8662, B1 => 
                           DataPath_RF_bus_reg_dataout_2410_port, B2 => n12119,
                           ZN => n1063);
   U16183 : OAI22_X1 port map( A1 => n12188, A2 => n12120, B1 => 
                           DataPath_RF_bus_reg_dataout_2411_port, B2 => n8661, 
                           ZN => n1062);
   U16184 : AOI22_X1 port map( A1 => n12189, A2 => n8661, B1 => n8662, B2 => 
                           DataPath_RF_bus_reg_dataout_2412_port, ZN => n1061);
   U16185 : AOI22_X1 port map( A1 => n12190, A2 => n8661, B1 => n12120, B2 => 
                           DataPath_RF_bus_reg_dataout_2413_port, ZN => n1060);
   U16186 : OAI22_X1 port map( A1 => n8662, A2 => n12191, B1 => 
                           DataPath_RF_bus_reg_dataout_2414_port, B2 => n8661, 
                           ZN => n1059);
   U16187 : AOI22_X1 port map( A1 => n12192, A2 => n8661, B1 => n8662, B2 => 
                           DataPath_RF_bus_reg_dataout_2415_port, ZN => n1058);
   U16188 : AOI22_X1 port map( A1 => n12159, A2 => n8661, B1 => n8662, B2 => 
                           DataPath_RF_bus_reg_dataout_2416_port, ZN => n1057);
   U16189 : AOI22_X1 port map( A1 => n12160, A2 => n8661, B1 => n8662, B2 => 
                           DataPath_RF_bus_reg_dataout_2417_port, ZN => n1056);
   U16190 : OAI22_X1 port map( A1 => n12161, A2 => n12120, B1 => 
                           DataPath_RF_bus_reg_dataout_2418_port, B2 => n8661, 
                           ZN => n1055);
   U16191 : OAI22_X1 port map( A1 => n12162, A2 => n8662, B1 => 
                           DataPath_RF_bus_reg_dataout_2419_port, B2 => n12119,
                           ZN => n1054);
   U16192 : AOI22_X1 port map( A1 => n12163, A2 => n8661, B1 => n8662, B2 => 
                           DataPath_RF_bus_reg_dataout_2420_port, ZN => n1053);
   U16193 : OAI22_X1 port map( A1 => n12164, A2 => n12120, B1 => 
                           DataPath_RF_bus_reg_dataout_2421_port, B2 => n8661, 
                           ZN => n1052);
   U16194 : AOI22_X1 port map( A1 => n12165, A2 => n12119, B1 => n8662, B2 => 
                           DataPath_RF_bus_reg_dataout_2422_port, ZN => n1051);
   U16195 : AOI22_X1 port map( A1 => n12166, A2 => n8661, B1 => n12120, B2 => 
                           DataPath_RF_bus_reg_dataout_2423_port, ZN => n1050);
   U16196 : OAI22_X1 port map( A1 => n12167, A2 => n8662, B1 => 
                           DataPath_RF_bus_reg_dataout_2424_port, B2 => n12119,
                           ZN => n1049);
   U16197 : AOI22_X1 port map( A1 => n12168, A2 => n8661, B1 => n12120, B2 => 
                           DataPath_RF_bus_reg_dataout_2425_port, ZN => n1048);
   U16198 : AOI22_X1 port map( A1 => n12169, A2 => n8661, B1 => n12120, B2 => 
                           DataPath_RF_bus_reg_dataout_2426_port, ZN => n1047);
   U16199 : AOI22_X1 port map( A1 => n12170, A2 => n8661, B1 => n12120, B2 => 
                           DataPath_RF_bus_reg_dataout_2427_port, ZN => n1046);
   U16200 : AOI22_X1 port map( A1 => n12171, A2 => n8661, B1 => n12120, B2 => 
                           DataPath_RF_bus_reg_dataout_2428_port, ZN => n1045);
   U16201 : AOI22_X1 port map( A1 => n12172, A2 => n8661, B1 => n8662, B2 => 
                           DataPath_RF_bus_reg_dataout_2429_port, ZN => n1044);
   U16202 : OAI22_X1 port map( A1 => n12173, A2 => n8662, B1 => 
                           DataPath_RF_bus_reg_dataout_2430_port, B2 => n12119,
                           ZN => n1043);
   U16203 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2431_port, A2 
                           => n12120, B1 => n12175, B2 => n8661, ZN => n1040);
   U16204 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2368_port, A2 
                           => n8663, B1 => n12152, B2 => n12122, ZN => n1036);
   U16205 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2369_port, A2 
                           => n12154, B1 => n12152, B2 => n12123, ZN => n1035);
   U16206 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2370_port, A2 
                           => n8663, B1 => n12152, B2 => n12124, ZN => n1034);
   U16207 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2371_port, A2 
                           => n8663, B1 => n12152, B2 => n12125, ZN => n1033);
   U16208 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2372_port, A2 
                           => n8663, B1 => n12152, B2 => n12126, ZN => n1032);
   U16209 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2373_port, A2 
                           => n12154, B1 => n12152, B2 => n12127, ZN => n1031);
   U16210 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2374_port, A2 
                           => n8663, B1 => n12152, B2 => n12128, ZN => n1030);
   U16211 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2375_port, A2 
                           => n8663, B1 => n12152, B2 => n12129, ZN => n1029);
   U16212 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2376_port, A2 
                           => n8663, B1 => n12152, B2 => n12130, ZN => n1028);
   U16213 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2377_port, A2 
                           => n8663, B1 => n12152, B2 => n12131, ZN => n1027);
   U16214 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2378_port, A2 
                           => n8663, B1 => n12152, B2 => n12132, ZN => n1026);
   U16215 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2379_port, A2 
                           => n8663, B1 => n12152, B2 => n12133, ZN => n1025);
   U16216 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2380_port, A2 
                           => n8663, B1 => n12152, B2 => n12134, ZN => n1024);
   U16217 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2381_port, A2 
                           => n8663, B1 => n12152, B2 => n12135, ZN => n1023);
   U16218 : OAI22_X1 port map( A1 => n12154, A2 => n12191, B1 => 
                           DataPath_RF_bus_reg_dataout_2382_port, B2 => n12153,
                           ZN => n1022);
   U16219 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2383_port, A2 
                           => n8663, B1 => n12152, B2 => n12136, ZN => n1021);
   U16220 : OAI22_X1 port map( A1 => n12159, A2 => n12154, B1 => 
                           DataPath_RF_bus_reg_dataout_2384_port, B2 => n12153,
                           ZN => n1020);
   U16221 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2385_port, A2 
                           => n8663, B1 => n12152, B2 => n12137, ZN => n1019);
   U16222 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2386_port, A2 
                           => n12154, B1 => n12152, B2 => n12138, ZN => n1018);
   U16223 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2387_port, A2 
                           => n12154, B1 => n12152, B2 => n12139, ZN => n1017);
   U16224 : OAI22_X1 port map( A1 => n12163, A2 => n12154, B1 => 
                           DataPath_RF_bus_reg_dataout_2388_port, B2 => n12153,
                           ZN => n1016);
   U16225 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2389_port, A2 
                           => n12154, B1 => n12152, B2 => n12141, ZN => n1015);
   U16226 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2390_port, A2 
                           => n12154, B1 => n12152, B2 => n12142, ZN => n1014);
   U16227 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2391_port, A2 
                           => n8663, B1 => n12152, B2 => n12143, ZN => n1013);
   U16228 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2392_port, A2 
                           => n12154, B1 => n12152, B2 => n12144, ZN => n1012);
   U16229 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2393_port, A2 
                           => n8663, B1 => n12152, B2 => n12146, ZN => n1011);
   U16230 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2394_port, A2 
                           => n8663, B1 => n12152, B2 => n12147, ZN => n1010);
   U16231 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2395_port, A2 
                           => n8663, B1 => n12152, B2 => n12148, ZN => n1009);
   U16232 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2396_port, A2 
                           => n8663, B1 => n12152, B2 => n12149, ZN => n1008);
   U16233 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2397_port, A2 
                           => n8663, B1 => n12152, B2 => n12150, ZN => n1007);
   U16234 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2398_port, A2 
                           => n8663, B1 => n12152, B2 => n12151, ZN => n1006);
   U16235 : OAI22_X1 port map( A1 => n12154, A2 => n12175, B1 => 
                           DataPath_RF_bus_reg_dataout_2399_port, B2 => n12153,
                           ZN => n1003);
   U16236 : AOI22_X1 port map( A1 => n12177, A2 => n8664, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2336_port, ZN => n999);
   U16237 : AOI22_X1 port map( A1 => n12178, A2 => n8664, B1 => n12157, B2 => 
                           DataPath_RF_bus_reg_dataout_2337_port, ZN => n998);
   U16238 : AOI22_X1 port map( A1 => n12179, A2 => n8664, B1 => n12157, B2 => 
                           DataPath_RF_bus_reg_dataout_2338_port, ZN => n997);
   U16239 : AOI22_X1 port map( A1 => n12180, A2 => n8664, B1 => n12157, B2 => 
                           DataPath_RF_bus_reg_dataout_2339_port, ZN => n996);
   U16240 : AOI22_X1 port map( A1 => n12181, A2 => n8664, B1 => n12157, B2 => 
                           DataPath_RF_bus_reg_dataout_2340_port, ZN => n995);
   U16241 : AOI22_X1 port map( A1 => n12182, A2 => n8664, B1 => n12157, B2 => 
                           DataPath_RF_bus_reg_dataout_2341_port, ZN => n994);
   U16242 : AOI22_X1 port map( A1 => n12183, A2 => n8664, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2342_port, ZN => n993);
   U16243 : AOI22_X1 port map( A1 => n12184, A2 => n8664, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2343_port, ZN => n992);
   U16244 : AOI22_X1 port map( A1 => n12185, A2 => n8664, B1 => n12157, B2 => 
                           DataPath_RF_bus_reg_dataout_2344_port, ZN => n991);
   U16245 : AOI22_X1 port map( A1 => n12186, A2 => n8664, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2345_port, ZN => n990);
   U16246 : AOI22_X1 port map( A1 => n12187, A2 => n12156, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2346_port, ZN => n989);
   U16247 : AOI22_X1 port map( A1 => n12188, A2 => n8664, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2347_port, ZN => n988);
   U16248 : AOI22_X1 port map( A1 => n12189, A2 => n8664, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2348_port, ZN => n987);
   U16249 : AOI22_X1 port map( A1 => n12190, A2 => n8664, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2349_port, ZN => n986);
   U16250 : OAI22_X1 port map( A1 => n8665, A2 => n12191, B1 => 
                           DataPath_RF_bus_reg_dataout_2350_port, B2 => n8664, 
                           ZN => n985);
   U16251 : AOI22_X1 port map( A1 => n12192, A2 => n8664, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2351_port, ZN => n984);
   U16252 : AOI22_X1 port map( A1 => n12159, A2 => n8664, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2352_port, ZN => n983);
   U16253 : AOI22_X1 port map( A1 => n12160, A2 => n12156, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2353_port, ZN => n982);
   U16254 : AOI22_X1 port map( A1 => n12161, A2 => n12156, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2354_port, ZN => n981);
   U16255 : AOI22_X1 port map( A1 => n12162, A2 => n8664, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2355_port, ZN => n980);
   U16256 : AOI22_X1 port map( A1 => n12163, A2 => n12156, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2356_port, ZN => n979);
   U16257 : AOI22_X1 port map( A1 => n12164, A2 => n12156, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2357_port, ZN => n978);
   U16258 : AOI22_X1 port map( A1 => n12165, A2 => n8664, B1 => n12157, B2 => 
                           DataPath_RF_bus_reg_dataout_2358_port, ZN => n977);
   U16259 : AOI22_X1 port map( A1 => n12166, A2 => n8664, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2359_port, ZN => n976);
   U16260 : AOI22_X1 port map( A1 => n12167, A2 => n12156, B1 => n12157, B2 => 
                           DataPath_RF_bus_reg_dataout_2360_port, ZN => n975);
   U16261 : AOI22_X1 port map( A1 => n12168, A2 => n12156, B1 => n12157, B2 => 
                           DataPath_RF_bus_reg_dataout_2361_port, ZN => n974);
   U16262 : AOI22_X1 port map( A1 => n12169, A2 => n8664, B1 => n12157, B2 => 
                           DataPath_RF_bus_reg_dataout_2362_port, ZN => n973);
   U16263 : AOI22_X1 port map( A1 => n12170, A2 => n12156, B1 => n12157, B2 => 
                           DataPath_RF_bus_reg_dataout_2363_port, ZN => n972);
   U16264 : AOI22_X1 port map( A1 => n12171, A2 => n8664, B1 => n12157, B2 => 
                           DataPath_RF_bus_reg_dataout_2364_port, ZN => n971);
   U16265 : AOI22_X1 port map( A1 => n12172, A2 => n12156, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2365_port, ZN => n970);
   U16266 : AOI22_X1 port map( A1 => n12173, A2 => n12156, B1 => n8665, B2 => 
                           DataPath_RF_bus_reg_dataout_2366_port, ZN => n969);
   U16267 : OAI22_X1 port map( A1 => n8665, A2 => n12175, B1 => 
                           DataPath_RF_bus_reg_dataout_2367_port, B2 => n8664, 
                           ZN => n966);
   U16268 : OAI22_X1 port map( A1 => n12177, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2304_port, B2 => n8666, 
                           ZN => n962);
   U16269 : AOI22_X1 port map( A1 => n12178, A2 => n8666, B1 => n12176, B2 => 
                           DataPath_RF_bus_reg_dataout_2305_port, ZN => n961);
   U16270 : AOI22_X1 port map( A1 => n12179, A2 => n8666, B1 => n12176, B2 => 
                           DataPath_RF_bus_reg_dataout_2306_port, ZN => n960);
   U16271 : OAI22_X1 port map( A1 => n12180, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2307_port, B2 => n8666, 
                           ZN => n959);
   U16272 : OAI22_X1 port map( A1 => n12181, A2 => n12176, B1 => 
                           DataPath_RF_bus_reg_dataout_2308_port, B2 => n12174,
                           ZN => n958);
   U16273 : OAI22_X1 port map( A1 => n12182, A2 => n12176, B1 => 
                           DataPath_RF_bus_reg_dataout_2309_port, B2 => n12174,
                           ZN => n957);
   U16274 : OAI22_X1 port map( A1 => n12183, A2 => n12176, B1 => 
                           DataPath_RF_bus_reg_dataout_2310_port, B2 => n12174,
                           ZN => n956);
   U16275 : OAI22_X1 port map( A1 => n12184, A2 => n12176, B1 => 
                           DataPath_RF_bus_reg_dataout_2311_port, B2 => n12174,
                           ZN => n955);
   U16276 : OAI22_X1 port map( A1 => n12185, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2312_port, B2 => n12174,
                           ZN => n954);
   U16277 : OAI22_X1 port map( A1 => n12186, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2313_port, B2 => n12174,
                           ZN => n953);
   U16278 : OAI22_X1 port map( A1 => n12187, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2314_port, B2 => n12174,
                           ZN => n952);
   U16279 : OAI22_X1 port map( A1 => n12188, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2315_port, B2 => n12174,
                           ZN => n951);
   U16280 : OAI22_X1 port map( A1 => n12189, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2316_port, B2 => n8666, 
                           ZN => n950);
   U16281 : OAI22_X1 port map( A1 => n12190, A2 => n12176, B1 => 
                           DataPath_RF_bus_reg_dataout_2317_port, B2 => n8666, 
                           ZN => n949);
   U16282 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2318_port, A2 
                           => n8667, B1 => n12191, B2 => n8666, ZN => n948);
   U16283 : OAI22_X1 port map( A1 => n12192, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2319_port, B2 => n8666, 
                           ZN => n947);
   U16284 : OAI22_X1 port map( A1 => n12159, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2320_port, B2 => n12174,
                           ZN => n945);
   U16285 : OAI22_X1 port map( A1 => n12160, A2 => n12176, B1 => 
                           DataPath_RF_bus_reg_dataout_2321_port, B2 => n12174,
                           ZN => n943);
   U16286 : AOI22_X1 port map( A1 => n12161, A2 => n8666, B1 => n12176, B2 => 
                           DataPath_RF_bus_reg_dataout_2322_port, ZN => n941);
   U16287 : OAI22_X1 port map( A1 => n12162, A2 => n12176, B1 => 
                           DataPath_RF_bus_reg_dataout_2323_port, B2 => n8666, 
                           ZN => n939);
   U16288 : OAI22_X1 port map( A1 => n12163, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2324_port, B2 => n8666, 
                           ZN => n937);
   U16289 : OAI22_X1 port map( A1 => n12164, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2325_port, B2 => n8666, 
                           ZN => n935);
   U16290 : OAI22_X1 port map( A1 => n12165, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2326_port, B2 => n8666, 
                           ZN => n933);
   U16291 : OAI22_X1 port map( A1 => n12166, A2 => n12176, B1 => 
                           DataPath_RF_bus_reg_dataout_2327_port, B2 => n8666, 
                           ZN => n931);
   U16292 : OAI22_X1 port map( A1 => n12167, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2328_port, B2 => n8666, 
                           ZN => n929);
   U16293 : OAI22_X1 port map( A1 => n12168, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2329_port, B2 => n8666, 
                           ZN => n927);
   U16294 : OAI22_X1 port map( A1 => n12169, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2330_port, B2 => n8666, 
                           ZN => n925);
   U16295 : OAI22_X1 port map( A1 => n12170, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2331_port, B2 => n8666, 
                           ZN => n923);
   U16296 : OAI22_X1 port map( A1 => n12171, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2332_port, B2 => n8666, 
                           ZN => n921);
   U16297 : OAI22_X1 port map( A1 => n12172, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2333_port, B2 => n8666, 
                           ZN => n919);
   U16298 : OAI22_X1 port map( A1 => n12173, A2 => n8667, B1 => 
                           DataPath_RF_bus_reg_dataout_2334_port, B2 => n8666, 
                           ZN => n917);
   U16299 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2335_port, A2 
                           => n8667, B1 => n12175, B2 => n8666, ZN => n913);
   U16300 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2272_port, B1 => n12177,
                           B2 => n8669, ZN => n911);
   U16301 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2273_port, B1 => n12178,
                           B2 => n8669, ZN => n909);
   U16302 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2274_port, B1 => n12179,
                           B2 => n8669, ZN => n907);
   U16303 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2275_port, B1 => n12180,
                           B2 => n8669, ZN => n905);
   U16304 : AOI22_X1 port map( A1 => n12193, A2 => 
                           DataPath_RF_bus_reg_dataout_2276_port, B1 => n12181,
                           B2 => n8669, ZN => n903);
   U16305 : AOI22_X1 port map( A1 => n12193, A2 => 
                           DataPath_RF_bus_reg_dataout_2277_port, B1 => n12182,
                           B2 => n8669, ZN => n901);
   U16306 : AOI22_X1 port map( A1 => n12193, A2 => 
                           DataPath_RF_bus_reg_dataout_2278_port, B1 => n12183,
                           B2 => n8669, ZN => n899);
   U16307 : AOI22_X1 port map( A1 => n12193, A2 => 
                           DataPath_RF_bus_reg_dataout_2279_port, B1 => n12184,
                           B2 => n8669, ZN => n897);
   U16308 : AOI22_X1 port map( A1 => n12193, A2 => 
                           DataPath_RF_bus_reg_dataout_2280_port, B1 => n12185,
                           B2 => n8669, ZN => n895);
   U16309 : AOI22_X1 port map( A1 => n12193, A2 => 
                           DataPath_RF_bus_reg_dataout_2281_port, B1 => n12186,
                           B2 => n8669, ZN => n893);
   U16310 : AOI22_X1 port map( A1 => n12193, A2 => 
                           DataPath_RF_bus_reg_dataout_2282_port, B1 => n12187,
                           B2 => n8669, ZN => n891);
   U16311 : AOI22_X1 port map( A1 => n12193, A2 => 
                           DataPath_RF_bus_reg_dataout_2283_port, B1 => n12188,
                           B2 => n8669, ZN => n889);
   U16312 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2284_port, B1 => n12189,
                           B2 => n8669, ZN => n887);
   U16313 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2285_port, B1 => n12190,
                           B2 => n8669, ZN => n885);
   U16314 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2286_port, B1 => n12191,
                           B2 => n8669, ZN => n883);
   U16315 : AOI22_X1 port map( A1 => n8668, A2 => 
                           DataPath_RF_bus_reg_dataout_2287_port, B1 => n12192,
                           B2 => n8669, ZN => n879);
   U16316 : INV_X1 port map( A => n12194, ZN => DRAM_ISSUE);
   U16317 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => n10851, B1 => n10857, 
                           B2 => CU_I_CW_EX_5_port, ZN => n12195);
   U16318 : INV_X1 port map( A => n12195, ZN => n385);
   U16319 : AOI22_X1 port map( A1 => DATA_SIZE_1_port, A2 => n10851, B1 => 
                           n10857, B2 => CU_I_CW_EX_4_port, ZN => n12196);
   U16320 : INV_X1 port map( A => n12196, ZN => n384);
   U16321 : AOI22_X1 port map( A1 => DATA_SIZE_0_port, A2 => n10851, B1 => 
                           n10857, B2 => CU_I_CW_EX_3_port, ZN => n12197);
   U16322 : INV_X1 port map( A => n12197, ZN => n383);
   U16323 : AOI22_X1 port map( A1 => i_DATAMEM_WM, A2 => n10851, B1 => n10857, 
                           B2 => CU_I_CW_EX_6_port, ZN => n12198);
   U16324 : INV_X1 port map( A => n12198, ZN => n382);
   U16325 : AOI22_X1 port map( A1 => n8670, A2 => DataPath_i_PIPLIN_WRB2_4_port
                           , B1 => n7765, B2 => i_ADD_WB_4_port, ZN => n12199);
   U16326 : INV_X1 port map( A => n12199, ZN => n376);
   U16327 : AOI22_X1 port map( A1 => n8670, A2 => DataPath_i_PIPLIN_WRB2_3_port
                           , B1 => n7765, B2 => i_ADD_WB_3_port, ZN => n12200);
   U16328 : INV_X1 port map( A => n12200, ZN => n375);
   U16329 : AOI22_X1 port map( A1 => i_ADD_WB_2_port, A2 => n7765, B1 => n12203
                           , B2 => DataPath_i_PIPLIN_WRB2_2_port, ZN => n12201)
                           ;
   U16330 : INV_X1 port map( A => n12201, ZN => n374);
   U16331 : AOI22_X1 port map( A1 => i_ADD_WB_1_port, A2 => n7765, B1 => n12203
                           , B2 => DataPath_i_PIPLIN_WRB2_1_port, ZN => n12202)
                           ;
   U16332 : INV_X1 port map( A => n12202, ZN => n373);
   U16333 : AOI22_X1 port map( A1 => i_ADD_WB_0_port, A2 => n7765, B1 => n12203
                           , B2 => DataPath_i_PIPLIN_WRB2_0_port, ZN => n12205)
                           ;
   U16334 : INV_X1 port map( A => n12205, ZN => n372);
   IRAM_ISSUE <= '1';

end SYN_dlx_rtl;
