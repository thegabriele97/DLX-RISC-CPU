
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32.all;

entity mux_N32_M5_0 is

   port( S : in std_logic_vector (4 downto 0);  Q : in std_logic_vector (1023 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end mux_N32_M5_0;

architecture SYN_behav of mux_N32_M5_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687 : std_logic;

begin
   
   U2 : AOI22_X1 port map( A1 => n673, A2 => Q(509), B1 => n672, B2 => Q(573), 
                           ZN => n1);
   U3 : AOI22_X1 port map( A1 => n675, A2 => Q(669), B1 => n674, B2 => Q(477), 
                           ZN => n2);
   U4 : AOI22_X1 port map( A1 => n677, A2 => Q(381), B1 => n676, B2 => Q(317), 
                           ZN => n3);
   U5 : AOI22_X1 port map( A1 => n679, A2 => Q(413), B1 => n678, B2 => Q(285), 
                           ZN => n4);
   U6 : NAND4_X1 port map( A1 => n1, A2 => n2, A3 => n3, A4 => n4, ZN => n5);
   U7 : AOI22_X1 port map( A1 => n681, A2 => Q(349), B1 => n680, B2 => Q(445), 
                           ZN => n6);
   U8 : AOI22_X1 port map( A1 => n683, A2 => Q(253), B1 => n682, B2 => Q(157), 
                           ZN => n7);
   U9 : AOI22_X1 port map( A1 => n685, A2 => Q(93), B1 => n684, B2 => Q(189), 
                           ZN => n8);
   U10 : AOI22_X1 port map( A1 => n687, A2 => Q(221), B1 => n686, B2 => Q(61), 
                           ZN => n9);
   U11 : NAND4_X1 port map( A1 => n6, A2 => n7, A3 => n8, A4 => n9, ZN => n10);
   U12 : AOI22_X1 port map( A1 => n656, A2 => Q(1021), B1 => n655, B2 => Q(957)
                           , ZN => n11);
   U13 : AOI22_X1 port map( A1 => n658, A2 => Q(989), B1 => n657, B2 => Q(925),
                           ZN => n12);
   U14 : AOI222_X1 port map( A1 => n660, A2 => Q(829), B1 => n661, B2 => Q(125)
                           , C1 => n659, C2 => Q(765), ZN => n13);
   U15 : NAND3_X1 port map( A1 => n11, A2 => n12, A3 => n13, ZN => n14);
   U16 : AOI22_X1 port map( A1 => n663, A2 => Q(861), B1 => n662, B2 => Q(733),
                           ZN => n15);
   U17 : AOI22_X1 port map( A1 => n665, A2 => Q(797), B1 => n664, B2 => Q(893),
                           ZN => n16);
   U18 : NAND4_X1 port map( A1 => n635, A2 => n636, A3 => n15, A4 => n16, ZN =>
                           n17);
   U19 : OR4_X1 port map( A1 => n5, A2 => n10, A3 => n14, A4 => n17, ZN => 
                           Y(29));
   U20 : AOI22_X1 port map( A1 => n673, A2 => Q(499), B1 => n672, B2 => Q(563),
                           ZN => n18);
   U21 : AOI22_X1 port map( A1 => n675, A2 => Q(659), B1 => n674, B2 => Q(467),
                           ZN => n19);
   U22 : AOI22_X1 port map( A1 => n677, A2 => Q(371), B1 => n676, B2 => Q(307),
                           ZN => n20);
   U23 : AOI22_X1 port map( A1 => n679, A2 => Q(403), B1 => n678, B2 => Q(275),
                           ZN => n21);
   U24 : NAND4_X1 port map( A1 => n18, A2 => n19, A3 => n20, A4 => n21, ZN => 
                           n22);
   U25 : AOI22_X1 port map( A1 => n681, A2 => Q(339), B1 => n680, B2 => Q(435),
                           ZN => n23);
   U26 : AOI22_X1 port map( A1 => n683, A2 => Q(243), B1 => n682, B2 => Q(147),
                           ZN => n24);
   U27 : AOI22_X1 port map( A1 => n685, A2 => Q(83), B1 => n684, B2 => Q(179), 
                           ZN => n25);
   U28 : AOI22_X1 port map( A1 => n687, A2 => Q(211), B1 => n686, B2 => Q(51), 
                           ZN => n26);
   U29 : NAND4_X1 port map( A1 => n23, A2 => n24, A3 => n25, A4 => n26, ZN => 
                           n27);
   U30 : AOI22_X1 port map( A1 => n656, A2 => Q(1011), B1 => n655, B2 => Q(947)
                           , ZN => n28);
   U31 : AOI22_X1 port map( A1 => n658, A2 => Q(979), B1 => n657, B2 => Q(915),
                           ZN => n29);
   U32 : AOI222_X1 port map( A1 => n660, A2 => Q(819), B1 => n661, B2 => Q(115)
                           , C1 => n659, C2 => Q(755), ZN => n30);
   U33 : NAND3_X1 port map( A1 => n28, A2 => n29, A3 => n30, ZN => n31);
   U34 : AOI22_X1 port map( A1 => n663, A2 => Q(851), B1 => n662, B2 => Q(723),
                           ZN => n32);
   U35 : AOI22_X1 port map( A1 => n665, A2 => Q(787), B1 => n664, B2 => Q(883),
                           ZN => n33);
   U36 : NAND4_X1 port map( A1 => n613, A2 => n614, A3 => n32, A4 => n33, ZN =>
                           n34);
   U37 : OR4_X1 port map( A1 => n22, A2 => n27, A3 => n31, A4 => n34, ZN => 
                           Y(19));
   U38 : AOI22_X1 port map( A1 => n673, A2 => Q(498), B1 => n672, B2 => Q(562),
                           ZN => n35);
   U39 : AOI22_X1 port map( A1 => n675, A2 => Q(658), B1 => n674, B2 => Q(466),
                           ZN => n36);
   U40 : AOI22_X1 port map( A1 => n677, A2 => Q(370), B1 => n676, B2 => Q(306),
                           ZN => n37);
   U41 : AOI22_X1 port map( A1 => n679, A2 => Q(402), B1 => n678, B2 => Q(274),
                           ZN => n38);
   U42 : NAND4_X1 port map( A1 => n35, A2 => n36, A3 => n37, A4 => n38, ZN => 
                           n39);
   U43 : AOI22_X1 port map( A1 => n681, A2 => Q(338), B1 => n680, B2 => Q(434),
                           ZN => n40);
   U44 : AOI22_X1 port map( A1 => n683, A2 => Q(242), B1 => n682, B2 => Q(146),
                           ZN => n41);
   U45 : AOI22_X1 port map( A1 => n685, A2 => Q(82), B1 => n684, B2 => Q(178), 
                           ZN => n42);
   U46 : AOI22_X1 port map( A1 => n687, A2 => Q(210), B1 => n686, B2 => Q(50), 
                           ZN => n43);
   U47 : NAND4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n44);
   U48 : AOI22_X1 port map( A1 => n656, A2 => Q(1010), B1 => n655, B2 => Q(946)
                           , ZN => n45);
   U49 : AOI22_X1 port map( A1 => n658, A2 => Q(978), B1 => n657, B2 => Q(914),
                           ZN => n46);
   U50 : AOI222_X1 port map( A1 => n660, A2 => Q(818), B1 => n661, B2 => Q(114)
                           , C1 => n659, C2 => Q(754), ZN => n47);
   U51 : NAND3_X1 port map( A1 => n45, A2 => n46, A3 => n47, ZN => n48);
   U52 : AOI22_X1 port map( A1 => n663, A2 => Q(850), B1 => n662, B2 => Q(722),
                           ZN => n49);
   U53 : AOI22_X1 port map( A1 => n665, A2 => Q(786), B1 => n664, B2 => Q(882),
                           ZN => n50);
   U54 : NAND4_X1 port map( A1 => n611, A2 => n612, A3 => n49, A4 => n50, ZN =>
                           n51);
   U55 : OR4_X1 port map( A1 => n39, A2 => n44, A3 => n48, A4 => n51, ZN => 
                           Y(18));
   U56 : AOI22_X1 port map( A1 => n673, A2 => Q(497), B1 => n672, B2 => Q(561),
                           ZN => n52);
   U57 : AOI22_X1 port map( A1 => n675, A2 => Q(657), B1 => n674, B2 => Q(465),
                           ZN => n53);
   U58 : AOI22_X1 port map( A1 => n677, A2 => Q(369), B1 => n676, B2 => Q(305),
                           ZN => n54);
   U59 : AOI22_X1 port map( A1 => n679, A2 => Q(401), B1 => n678, B2 => Q(273),
                           ZN => n55);
   U60 : NAND4_X1 port map( A1 => n52, A2 => n53, A3 => n54, A4 => n55, ZN => 
                           n56);
   U61 : AOI22_X1 port map( A1 => n681, A2 => Q(337), B1 => n680, B2 => Q(433),
                           ZN => n57);
   U62 : AOI22_X1 port map( A1 => n683, A2 => Q(241), B1 => n682, B2 => Q(145),
                           ZN => n58);
   U63 : AOI22_X1 port map( A1 => n685, A2 => Q(81), B1 => n684, B2 => Q(177), 
                           ZN => n59);
   U64 : AOI22_X1 port map( A1 => n687, A2 => Q(209), B1 => n686, B2 => Q(49), 
                           ZN => n60);
   U65 : NAND4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           n61);
   U66 : AOI22_X1 port map( A1 => n656, A2 => Q(1009), B1 => n655, B2 => Q(945)
                           , ZN => n62);
   U67 : AOI22_X1 port map( A1 => n658, A2 => Q(977), B1 => n657, B2 => Q(913),
                           ZN => n63);
   U68 : AOI222_X1 port map( A1 => n660, A2 => Q(817), B1 => n661, B2 => Q(113)
                           , C1 => n659, C2 => Q(753), ZN => n64);
   U69 : NAND3_X1 port map( A1 => n62, A2 => n63, A3 => n64, ZN => n65);
   U70 : AOI22_X1 port map( A1 => n663, A2 => Q(849), B1 => n662, B2 => Q(721),
                           ZN => n66);
   U71 : AOI22_X1 port map( A1 => n665, A2 => Q(785), B1 => n664, B2 => Q(881),
                           ZN => n67);
   U72 : NAND4_X1 port map( A1 => n609, A2 => n610, A3 => n66, A4 => n67, ZN =>
                           n68);
   U73 : OR4_X1 port map( A1 => n56, A2 => n61, A3 => n65, A4 => n68, ZN => 
                           Y(17));
   U74 : AOI22_X1 port map( A1 => n673, A2 => Q(496), B1 => n672, B2 => Q(560),
                           ZN => n69);
   U75 : AOI22_X1 port map( A1 => n675, A2 => Q(656), B1 => n674, B2 => Q(464),
                           ZN => n70);
   U76 : AOI22_X1 port map( A1 => n677, A2 => Q(368), B1 => n676, B2 => Q(304),
                           ZN => n71);
   U77 : AOI22_X1 port map( A1 => n679, A2 => Q(400), B1 => n678, B2 => Q(272),
                           ZN => n72);
   U78 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           n73);
   U79 : AOI22_X1 port map( A1 => n681, A2 => Q(336), B1 => n680, B2 => Q(432),
                           ZN => n74);
   U80 : AOI22_X1 port map( A1 => n683, A2 => Q(240), B1 => n682, B2 => Q(144),
                           ZN => n75);
   U81 : AOI22_X1 port map( A1 => n685, A2 => Q(80), B1 => n684, B2 => Q(176), 
                           ZN => n76);
   U82 : AOI22_X1 port map( A1 => n687, A2 => Q(208), B1 => n686, B2 => Q(48), 
                           ZN => n77);
   U83 : NAND4_X1 port map( A1 => n74, A2 => n75, A3 => n76, A4 => n77, ZN => 
                           n78);
   U84 : AOI22_X1 port map( A1 => n656, A2 => Q(1008), B1 => n655, B2 => Q(944)
                           , ZN => n79);
   U85 : AOI22_X1 port map( A1 => n658, A2 => Q(976), B1 => n657, B2 => Q(912),
                           ZN => n80);
   U86 : AOI222_X1 port map( A1 => n660, A2 => Q(816), B1 => n661, B2 => Q(112)
                           , C1 => n659, C2 => Q(752), ZN => n81);
   U87 : NAND3_X1 port map( A1 => n79, A2 => n80, A3 => n81, ZN => n82);
   U88 : AOI22_X1 port map( A1 => n663, A2 => Q(848), B1 => n662, B2 => Q(720),
                           ZN => n83);
   U89 : AOI22_X1 port map( A1 => n665, A2 => Q(784), B1 => n664, B2 => Q(880),
                           ZN => n84);
   U90 : NAND4_X1 port map( A1 => n607, A2 => n608, A3 => n83, A4 => n84, ZN =>
                           n85);
   U91 : OR4_X1 port map( A1 => n73, A2 => n78, A3 => n82, A4 => n85, ZN => 
                           Y(16));
   U92 : AOI22_X1 port map( A1 => n673, A2 => Q(495), B1 => n672, B2 => Q(559),
                           ZN => n86);
   U93 : AOI22_X1 port map( A1 => n675, A2 => Q(655), B1 => n674, B2 => Q(463),
                           ZN => n87);
   U94 : AOI22_X1 port map( A1 => n677, A2 => Q(367), B1 => n676, B2 => Q(303),
                           ZN => n88);
   U95 : AOI22_X1 port map( A1 => n679, A2 => Q(399), B1 => n678, B2 => Q(271),
                           ZN => n89);
   U96 : NAND4_X1 port map( A1 => n86, A2 => n87, A3 => n88, A4 => n89, ZN => 
                           n90);
   U97 : AOI22_X1 port map( A1 => n681, A2 => Q(335), B1 => n680, B2 => Q(431),
                           ZN => n91);
   U98 : AOI22_X1 port map( A1 => n683, A2 => Q(239), B1 => n682, B2 => Q(143),
                           ZN => n92);
   U99 : AOI22_X1 port map( A1 => n685, A2 => Q(79), B1 => n684, B2 => Q(175), 
                           ZN => n93);
   U100 : AOI22_X1 port map( A1 => n687, A2 => Q(207), B1 => n686, B2 => Q(47),
                           ZN => n94);
   U101 : NAND4_X1 port map( A1 => n91, A2 => n92, A3 => n93, A4 => n94, ZN => 
                           n95);
   U102 : AOI22_X1 port map( A1 => n656, A2 => Q(1007), B1 => n655, B2 => 
                           Q(943), ZN => n96);
   U103 : AOI22_X1 port map( A1 => n658, A2 => Q(975), B1 => n657, B2 => Q(911)
                           , ZN => n97);
   U104 : AOI222_X1 port map( A1 => n660, A2 => Q(815), B1 => n661, B2 => 
                           Q(111), C1 => n659, C2 => Q(751), ZN => n98);
   U105 : NAND3_X1 port map( A1 => n96, A2 => n97, A3 => n98, ZN => n99);
   U106 : AOI22_X1 port map( A1 => n663, A2 => Q(847), B1 => n662, B2 => Q(719)
                           , ZN => n100);
   U107 : AOI22_X1 port map( A1 => n665, A2 => Q(783), B1 => n664, B2 => Q(879)
                           , ZN => n101);
   U108 : NAND4_X1 port map( A1 => n605, A2 => n606, A3 => n100, A4 => n101, ZN
                           => n102);
   U109 : OR4_X1 port map( A1 => n90, A2 => n95, A3 => n99, A4 => n102, ZN => 
                           Y(15));
   U110 : AOI22_X1 port map( A1 => n673, A2 => Q(494), B1 => n672, B2 => Q(558)
                           , ZN => n103);
   U111 : AOI22_X1 port map( A1 => n675, A2 => Q(654), B1 => n674, B2 => Q(462)
                           , ZN => n104);
   U112 : AOI22_X1 port map( A1 => n677, A2 => Q(366), B1 => n676, B2 => Q(302)
                           , ZN => n105);
   U113 : AOI22_X1 port map( A1 => n679, A2 => Q(398), B1 => n678, B2 => Q(270)
                           , ZN => n106);
   U114 : NAND4_X1 port map( A1 => n103, A2 => n104, A3 => n105, A4 => n106, ZN
                           => n107);
   U115 : AOI22_X1 port map( A1 => n681, A2 => Q(334), B1 => n680, B2 => Q(430)
                           , ZN => n108);
   U116 : AOI22_X1 port map( A1 => n683, A2 => Q(238), B1 => n682, B2 => Q(142)
                           , ZN => n109);
   U117 : AOI22_X1 port map( A1 => n685, A2 => Q(78), B1 => n684, B2 => Q(174),
                           ZN => n110);
   U118 : AOI22_X1 port map( A1 => n687, A2 => Q(206), B1 => n686, B2 => Q(46),
                           ZN => n111);
   U119 : NAND4_X1 port map( A1 => n108, A2 => n109, A3 => n110, A4 => n111, ZN
                           => n112);
   U120 : AOI22_X1 port map( A1 => n656, A2 => Q(1006), B1 => n655, B2 => 
                           Q(942), ZN => n113);
   U121 : AOI22_X1 port map( A1 => n658, A2 => Q(974), B1 => n657, B2 => Q(910)
                           , ZN => n114);
   U122 : AOI222_X1 port map( A1 => n660, A2 => Q(814), B1 => n661, B2 => 
                           Q(110), C1 => n659, C2 => Q(750), ZN => n115);
   U123 : NAND3_X1 port map( A1 => n113, A2 => n114, A3 => n115, ZN => n116);
   U124 : AOI22_X1 port map( A1 => n663, A2 => Q(846), B1 => n662, B2 => Q(718)
                           , ZN => n117);
   U125 : AOI22_X1 port map( A1 => n665, A2 => Q(782), B1 => n664, B2 => Q(878)
                           , ZN => n118);
   U126 : NAND4_X1 port map( A1 => n603, A2 => n604, A3 => n117, A4 => n118, ZN
                           => n119);
   U127 : OR4_X1 port map( A1 => n107, A2 => n112, A3 => n116, A4 => n119, ZN 
                           => Y(14));
   U128 : AOI22_X1 port map( A1 => n673, A2 => Q(493), B1 => n672, B2 => Q(557)
                           , ZN => n120);
   U129 : AOI22_X1 port map( A1 => n675, A2 => Q(653), B1 => n674, B2 => Q(461)
                           , ZN => n121);
   U130 : AOI22_X1 port map( A1 => n677, A2 => Q(365), B1 => n676, B2 => Q(301)
                           , ZN => n122);
   U131 : AOI22_X1 port map( A1 => n679, A2 => Q(397), B1 => n678, B2 => Q(269)
                           , ZN => n123);
   U132 : NAND4_X1 port map( A1 => n120, A2 => n121, A3 => n122, A4 => n123, ZN
                           => n124);
   U133 : AOI22_X1 port map( A1 => n681, A2 => Q(333), B1 => n680, B2 => Q(429)
                           , ZN => n125);
   U134 : AOI22_X1 port map( A1 => n683, A2 => Q(237), B1 => n682, B2 => Q(141)
                           , ZN => n126);
   U135 : AOI22_X1 port map( A1 => n685, A2 => Q(77), B1 => n684, B2 => Q(173),
                           ZN => n127);
   U136 : AOI22_X1 port map( A1 => n687, A2 => Q(205), B1 => n686, B2 => Q(45),
                           ZN => n128);
   U137 : NAND4_X1 port map( A1 => n125, A2 => n126, A3 => n127, A4 => n128, ZN
                           => n129);
   U138 : AOI22_X1 port map( A1 => n656, A2 => Q(1005), B1 => n655, B2 => 
                           Q(941), ZN => n130);
   U139 : AOI22_X1 port map( A1 => n658, A2 => Q(973), B1 => n657, B2 => Q(909)
                           , ZN => n131);
   U140 : AOI222_X1 port map( A1 => n660, A2 => Q(813), B1 => n661, B2 => 
                           Q(109), C1 => n659, C2 => Q(749), ZN => n132);
   U141 : NAND3_X1 port map( A1 => n130, A2 => n131, A3 => n132, ZN => n133);
   U142 : AOI22_X1 port map( A1 => n663, A2 => Q(845), B1 => n662, B2 => Q(717)
                           , ZN => n134);
   U143 : AOI22_X1 port map( A1 => n665, A2 => Q(781), B1 => n664, B2 => Q(877)
                           , ZN => n135);
   U144 : NAND4_X1 port map( A1 => n601, A2 => n602, A3 => n134, A4 => n135, ZN
                           => n136);
   U145 : OR4_X1 port map( A1 => n124, A2 => n129, A3 => n133, A4 => n136, ZN 
                           => Y(13));
   U146 : AOI22_X1 port map( A1 => n673, A2 => Q(492), B1 => n672, B2 => Q(556)
                           , ZN => n137);
   U147 : AOI22_X1 port map( A1 => n675, A2 => Q(652), B1 => n674, B2 => Q(460)
                           , ZN => n138);
   U148 : AOI22_X1 port map( A1 => n677, A2 => Q(364), B1 => n676, B2 => Q(300)
                           , ZN => n139);
   U149 : AOI22_X1 port map( A1 => n679, A2 => Q(396), B1 => n678, B2 => Q(268)
                           , ZN => n140);
   U150 : NAND4_X1 port map( A1 => n137, A2 => n138, A3 => n139, A4 => n140, ZN
                           => n141);
   U151 : AOI22_X1 port map( A1 => n681, A2 => Q(332), B1 => n680, B2 => Q(428)
                           , ZN => n142);
   U152 : AOI22_X1 port map( A1 => n683, A2 => Q(236), B1 => n682, B2 => Q(140)
                           , ZN => n143);
   U153 : AOI22_X1 port map( A1 => n685, A2 => Q(76), B1 => n684, B2 => Q(172),
                           ZN => n144);
   U154 : AOI22_X1 port map( A1 => n687, A2 => Q(204), B1 => n686, B2 => Q(44),
                           ZN => n145);
   U155 : NAND4_X1 port map( A1 => n142, A2 => n143, A3 => n144, A4 => n145, ZN
                           => n146);
   U156 : AOI22_X1 port map( A1 => n656, A2 => Q(1004), B1 => n655, B2 => 
                           Q(940), ZN => n147);
   U157 : AOI22_X1 port map( A1 => n658, A2 => Q(972), B1 => n657, B2 => Q(908)
                           , ZN => n148);
   U158 : AOI222_X1 port map( A1 => n660, A2 => Q(812), B1 => n661, B2 => 
                           Q(108), C1 => n659, C2 => Q(748), ZN => n149);
   U159 : NAND3_X1 port map( A1 => n147, A2 => n148, A3 => n149, ZN => n150);
   U160 : AOI22_X1 port map( A1 => n663, A2 => Q(844), B1 => n662, B2 => Q(716)
                           , ZN => n151);
   U161 : AOI22_X1 port map( A1 => n665, A2 => Q(780), B1 => n664, B2 => Q(876)
                           , ZN => n152);
   U162 : NAND4_X1 port map( A1 => n599, A2 => n600, A3 => n151, A4 => n152, ZN
                           => n153);
   U163 : OR4_X1 port map( A1 => n141, A2 => n146, A3 => n150, A4 => n153, ZN 
                           => Y(12));
   U164 : AOI22_X1 port map( A1 => n561, A2 => Q(511), B1 => n560, B2 => Q(575)
                           , ZN => n154);
   U165 : AOI22_X1 port map( A1 => n563, A2 => Q(671), B1 => n562, B2 => Q(479)
                           , ZN => n155);
   U166 : AOI22_X1 port map( A1 => n565, A2 => Q(383), B1 => n564, B2 => Q(319)
                           , ZN => n156);
   U167 : AOI22_X1 port map( A1 => n567, A2 => Q(415), B1 => n566, B2 => Q(287)
                           , ZN => n157);
   U168 : NAND4_X1 port map( A1 => n154, A2 => n155, A3 => n156, A4 => n157, ZN
                           => n158);
   U169 : AOI22_X1 port map( A1 => n569, A2 => Q(351), B1 => n568, B2 => Q(447)
                           , ZN => n159);
   U170 : AOI22_X1 port map( A1 => n571, A2 => Q(255), B1 => n570, B2 => Q(159)
                           , ZN => n160);
   U171 : AOI22_X1 port map( A1 => n573, A2 => Q(95), B1 => n572, B2 => Q(191),
                           ZN => n161);
   U172 : AOI22_X1 port map( A1 => n575, A2 => Q(223), B1 => n574, B2 => Q(63),
                           ZN => n162);
   U173 : NAND4_X1 port map( A1 => n159, A2 => n160, A3 => n161, A4 => n162, ZN
                           => n163);
   U174 : AOI22_X1 port map( A1 => n546, A2 => Q(1023), B1 => n545, B2 => 
                           Q(959), ZN => n164);
   U175 : AOI22_X1 port map( A1 => n548, A2 => Q(991), B1 => n547, B2 => Q(927)
                           , ZN => n165);
   U176 : AOI222_X1 port map( A1 => n550, A2 => Q(831), B1 => n551, B2 => 
                           Q(127), C1 => n549, C2 => Q(767), ZN => n166);
   U177 : NAND3_X1 port map( A1 => n164, A2 => n165, A3 => n166, ZN => n167);
   U178 : AOI22_X1 port map( A1 => n553, A2 => Q(863), B1 => n552, B2 => Q(735)
                           , ZN => n168);
   U179 : AOI22_X1 port map( A1 => n555, A2 => Q(799), B1 => n554, B2 => Q(895)
                           , ZN => n169);
   U180 : NAND4_X1 port map( A1 => n641, A2 => n642, A3 => n168, A4 => n169, ZN
                           => n170);
   U181 : OR4_X1 port map( A1 => n158, A2 => n163, A3 => n167, A4 => n170, ZN 
                           => Y(31));
   U182 : AOI22_X1 port map( A1 => n561, A2 => Q(510), B1 => n560, B2 => Q(574)
                           , ZN => n171);
   U183 : AOI22_X1 port map( A1 => n563, A2 => Q(670), B1 => n562, B2 => Q(478)
                           , ZN => n172);
   U184 : AOI22_X1 port map( A1 => n565, A2 => Q(382), B1 => n564, B2 => Q(318)
                           , ZN => n173);
   U185 : AOI22_X1 port map( A1 => n567, A2 => Q(414), B1 => n566, B2 => Q(286)
                           , ZN => n174);
   U186 : NAND4_X1 port map( A1 => n171, A2 => n172, A3 => n173, A4 => n174, ZN
                           => n175);
   U187 : AOI22_X1 port map( A1 => n569, A2 => Q(350), B1 => n568, B2 => Q(446)
                           , ZN => n176);
   U188 : AOI22_X1 port map( A1 => n571, A2 => Q(254), B1 => n570, B2 => Q(158)
                           , ZN => n177);
   U189 : AOI22_X1 port map( A1 => n573, A2 => Q(94), B1 => n572, B2 => Q(190),
                           ZN => n178);
   U190 : AOI22_X1 port map( A1 => n575, A2 => Q(222), B1 => n574, B2 => Q(62),
                           ZN => n179);
   U191 : NAND4_X1 port map( A1 => n176, A2 => n177, A3 => n178, A4 => n179, ZN
                           => n180);
   U192 : AOI22_X1 port map( A1 => n546, A2 => Q(1022), B1 => n545, B2 => 
                           Q(958), ZN => n181);
   U193 : AOI22_X1 port map( A1 => n548, A2 => Q(990), B1 => n547, B2 => Q(926)
                           , ZN => n182);
   U194 : AOI222_X1 port map( A1 => n550, A2 => Q(830), B1 => n551, B2 => 
                           Q(126), C1 => n549, C2 => Q(766), ZN => n183);
   U195 : NAND3_X1 port map( A1 => n181, A2 => n182, A3 => n183, ZN => n184);
   U196 : AOI22_X1 port map( A1 => n553, A2 => Q(862), B1 => n552, B2 => Q(734)
                           , ZN => n185);
   U197 : AOI22_X1 port map( A1 => n555, A2 => Q(798), B1 => n554, B2 => Q(894)
                           , ZN => n186);
   U198 : NAND4_X1 port map( A1 => n639, A2 => n640, A3 => n185, A4 => n186, ZN
                           => n187);
   U199 : OR4_X1 port map( A1 => n175, A2 => n180, A3 => n184, A4 => n187, ZN 
                           => Y(30));
   U200 : AOI22_X1 port map( A1 => n561, A2 => Q(508), B1 => n560, B2 => Q(572)
                           , ZN => n188);
   U201 : AOI22_X1 port map( A1 => n563, A2 => Q(668), B1 => n562, B2 => Q(476)
                           , ZN => n189);
   U202 : AOI22_X1 port map( A1 => n565, A2 => Q(380), B1 => n564, B2 => Q(316)
                           , ZN => n190);
   U203 : AOI22_X1 port map( A1 => n567, A2 => Q(412), B1 => n566, B2 => Q(284)
                           , ZN => n191);
   U204 : NAND4_X1 port map( A1 => n188, A2 => n189, A3 => n190, A4 => n191, ZN
                           => n192);
   U205 : AOI22_X1 port map( A1 => n569, A2 => Q(348), B1 => n568, B2 => Q(444)
                           , ZN => n193);
   U206 : AOI22_X1 port map( A1 => n571, A2 => Q(252), B1 => n570, B2 => Q(156)
                           , ZN => n194);
   U207 : AOI22_X1 port map( A1 => n573, A2 => Q(92), B1 => n572, B2 => Q(188),
                           ZN => n195);
   U208 : AOI22_X1 port map( A1 => n575, A2 => Q(220), B1 => n574, B2 => Q(60),
                           ZN => n196);
   U209 : NAND4_X1 port map( A1 => n193, A2 => n194, A3 => n195, A4 => n196, ZN
                           => n197);
   U210 : AOI22_X1 port map( A1 => n546, A2 => Q(1020), B1 => n545, B2 => 
                           Q(956), ZN => n198);
   U211 : AOI22_X1 port map( A1 => n548, A2 => Q(988), B1 => n547, B2 => Q(924)
                           , ZN => n199);
   U212 : AOI222_X1 port map( A1 => n550, A2 => Q(828), B1 => n551, B2 => 
                           Q(124), C1 => n549, C2 => Q(764), ZN => n200);
   U213 : NAND3_X1 port map( A1 => n198, A2 => n199, A3 => n200, ZN => n201);
   U214 : AOI22_X1 port map( A1 => n553, A2 => Q(860), B1 => n552, B2 => Q(732)
                           , ZN => n202);
   U215 : AOI22_X1 port map( A1 => n555, A2 => Q(796), B1 => n554, B2 => Q(892)
                           , ZN => n203);
   U216 : NAND4_X1 port map( A1 => n633, A2 => n634, A3 => n202, A4 => n203, ZN
                           => n204);
   U217 : OR4_X1 port map( A1 => n192, A2 => n197, A3 => n201, A4 => n204, ZN 
                           => Y(28));
   U218 : AOI22_X1 port map( A1 => n561, A2 => Q(507), B1 => n560, B2 => Q(571)
                           , ZN => n205);
   U219 : AOI22_X1 port map( A1 => n563, A2 => Q(667), B1 => n562, B2 => Q(475)
                           , ZN => n206);
   U220 : AOI22_X1 port map( A1 => n565, A2 => Q(379), B1 => n564, B2 => Q(315)
                           , ZN => n207);
   U221 : AOI22_X1 port map( A1 => n567, A2 => Q(411), B1 => n566, B2 => Q(283)
                           , ZN => n208);
   U222 : NAND4_X1 port map( A1 => n205, A2 => n206, A3 => n207, A4 => n208, ZN
                           => n209);
   U223 : AOI22_X1 port map( A1 => n569, A2 => Q(347), B1 => n568, B2 => Q(443)
                           , ZN => n210);
   U224 : AOI22_X1 port map( A1 => n571, A2 => Q(251), B1 => n570, B2 => Q(155)
                           , ZN => n211);
   U225 : AOI22_X1 port map( A1 => n573, A2 => Q(91), B1 => n572, B2 => Q(187),
                           ZN => n212);
   U226 : AOI22_X1 port map( A1 => n575, A2 => Q(219), B1 => n574, B2 => Q(59),
                           ZN => n213);
   U227 : NAND4_X1 port map( A1 => n210, A2 => n211, A3 => n212, A4 => n213, ZN
                           => n214);
   U228 : AOI22_X1 port map( A1 => n546, A2 => Q(1019), B1 => n545, B2 => 
                           Q(955), ZN => n215);
   U229 : AOI22_X1 port map( A1 => n548, A2 => Q(987), B1 => n547, B2 => Q(923)
                           , ZN => n216);
   U230 : AOI222_X1 port map( A1 => n550, A2 => Q(827), B1 => n551, B2 => 
                           Q(123), C1 => n549, C2 => Q(763), ZN => n217);
   U231 : NAND3_X1 port map( A1 => n215, A2 => n216, A3 => n217, ZN => n218);
   U232 : AOI22_X1 port map( A1 => n553, A2 => Q(859), B1 => n552, B2 => Q(731)
                           , ZN => n219);
   U233 : AOI22_X1 port map( A1 => n555, A2 => Q(795), B1 => n554, B2 => Q(891)
                           , ZN => n220);
   U234 : NAND4_X1 port map( A1 => n631, A2 => n632, A3 => n219, A4 => n220, ZN
                           => n221);
   U235 : OR4_X1 port map( A1 => n209, A2 => n214, A3 => n218, A4 => n221, ZN 
                           => Y(27));
   U236 : AOI22_X1 port map( A1 => n561, A2 => Q(506), B1 => n560, B2 => Q(570)
                           , ZN => n222);
   U237 : AOI22_X1 port map( A1 => n563, A2 => Q(666), B1 => n562, B2 => Q(474)
                           , ZN => n223);
   U238 : AOI22_X1 port map( A1 => n565, A2 => Q(378), B1 => n564, B2 => Q(314)
                           , ZN => n224);
   U239 : AOI22_X1 port map( A1 => n567, A2 => Q(410), B1 => n566, B2 => Q(282)
                           , ZN => n225);
   U240 : NAND4_X1 port map( A1 => n222, A2 => n223, A3 => n224, A4 => n225, ZN
                           => n226);
   U241 : AOI22_X1 port map( A1 => n569, A2 => Q(346), B1 => n568, B2 => Q(442)
                           , ZN => n227);
   U242 : AOI22_X1 port map( A1 => n571, A2 => Q(250), B1 => n570, B2 => Q(154)
                           , ZN => n228);
   U243 : AOI22_X1 port map( A1 => n573, A2 => Q(90), B1 => n572, B2 => Q(186),
                           ZN => n229);
   U244 : AOI22_X1 port map( A1 => n575, A2 => Q(218), B1 => n574, B2 => Q(58),
                           ZN => n230);
   U245 : NAND4_X1 port map( A1 => n227, A2 => n228, A3 => n229, A4 => n230, ZN
                           => n231);
   U246 : AOI22_X1 port map( A1 => n546, A2 => Q(1018), B1 => n545, B2 => 
                           Q(954), ZN => n232);
   U247 : AOI22_X1 port map( A1 => n548, A2 => Q(986), B1 => n547, B2 => Q(922)
                           , ZN => n233);
   U248 : AOI222_X1 port map( A1 => n550, A2 => Q(826), B1 => n551, B2 => 
                           Q(122), C1 => n549, C2 => Q(762), ZN => n234);
   U249 : NAND3_X1 port map( A1 => n232, A2 => n233, A3 => n234, ZN => n235);
   U250 : AOI22_X1 port map( A1 => n553, A2 => Q(858), B1 => n552, B2 => Q(730)
                           , ZN => n236);
   U251 : AOI22_X1 port map( A1 => n555, A2 => Q(794), B1 => n554, B2 => Q(890)
                           , ZN => n237);
   U252 : NAND4_X1 port map( A1 => n629, A2 => n630, A3 => n236, A4 => n237, ZN
                           => n238);
   U253 : OR4_X1 port map( A1 => n226, A2 => n231, A3 => n235, A4 => n238, ZN 
                           => Y(26));
   U254 : AOI22_X1 port map( A1 => n561, A2 => Q(505), B1 => n560, B2 => Q(569)
                           , ZN => n239);
   U255 : AOI22_X1 port map( A1 => n563, A2 => Q(665), B1 => n562, B2 => Q(473)
                           , ZN => n240);
   U256 : AOI22_X1 port map( A1 => n565, A2 => Q(377), B1 => n564, B2 => Q(313)
                           , ZN => n241);
   U257 : AOI22_X1 port map( A1 => n567, A2 => Q(409), B1 => n566, B2 => Q(281)
                           , ZN => n242);
   U258 : NAND4_X1 port map( A1 => n239, A2 => n240, A3 => n241, A4 => n242, ZN
                           => n243);
   U259 : AOI22_X1 port map( A1 => n569, A2 => Q(345), B1 => n568, B2 => Q(441)
                           , ZN => n244);
   U260 : AOI22_X1 port map( A1 => n571, A2 => Q(249), B1 => n570, B2 => Q(153)
                           , ZN => n245);
   U261 : AOI22_X1 port map( A1 => n573, A2 => Q(89), B1 => n572, B2 => Q(185),
                           ZN => n246);
   U262 : AOI22_X1 port map( A1 => n575, A2 => Q(217), B1 => n574, B2 => Q(57),
                           ZN => n247);
   U263 : NAND4_X1 port map( A1 => n244, A2 => n245, A3 => n246, A4 => n247, ZN
                           => n248);
   U264 : AOI22_X1 port map( A1 => n546, A2 => Q(1017), B1 => n545, B2 => 
                           Q(953), ZN => n249);
   U265 : AOI22_X1 port map( A1 => n548, A2 => Q(985), B1 => n547, B2 => Q(921)
                           , ZN => n250);
   U266 : AOI222_X1 port map( A1 => n550, A2 => Q(825), B1 => n551, B2 => 
                           Q(121), C1 => n549, C2 => Q(761), ZN => n251);
   U267 : NAND3_X1 port map( A1 => n249, A2 => n250, A3 => n251, ZN => n252);
   U268 : AOI22_X1 port map( A1 => n553, A2 => Q(857), B1 => n552, B2 => Q(729)
                           , ZN => n253);
   U269 : AOI22_X1 port map( A1 => n555, A2 => Q(793), B1 => n554, B2 => Q(889)
                           , ZN => n254);
   U270 : NAND4_X1 port map( A1 => n627, A2 => n628, A3 => n253, A4 => n254, ZN
                           => n255);
   U271 : OR4_X1 port map( A1 => n243, A2 => n248, A3 => n252, A4 => n255, ZN 
                           => Y(25));
   U272 : AOI22_X1 port map( A1 => n561, A2 => Q(504), B1 => n560, B2 => Q(568)
                           , ZN => n256);
   U273 : AOI22_X1 port map( A1 => n563, A2 => Q(664), B1 => n562, B2 => Q(472)
                           , ZN => n257);
   U274 : AOI22_X1 port map( A1 => n565, A2 => Q(376), B1 => n564, B2 => Q(312)
                           , ZN => n258);
   U275 : AOI22_X1 port map( A1 => n567, A2 => Q(408), B1 => n566, B2 => Q(280)
                           , ZN => n259);
   U276 : NAND4_X1 port map( A1 => n256, A2 => n257, A3 => n258, A4 => n259, ZN
                           => n260);
   U277 : AOI22_X1 port map( A1 => n569, A2 => Q(344), B1 => n568, B2 => Q(440)
                           , ZN => n261);
   U278 : AOI22_X1 port map( A1 => n571, A2 => Q(248), B1 => n570, B2 => Q(152)
                           , ZN => n262);
   U279 : AOI22_X1 port map( A1 => n573, A2 => Q(88), B1 => n572, B2 => Q(184),
                           ZN => n263);
   U280 : AOI22_X1 port map( A1 => n575, A2 => Q(216), B1 => n574, B2 => Q(56),
                           ZN => n264);
   U281 : NAND4_X1 port map( A1 => n261, A2 => n262, A3 => n263, A4 => n264, ZN
                           => n265);
   U282 : AOI22_X1 port map( A1 => n546, A2 => Q(1016), B1 => n545, B2 => 
                           Q(952), ZN => n266);
   U283 : AOI22_X1 port map( A1 => n548, A2 => Q(984), B1 => n547, B2 => Q(920)
                           , ZN => n267);
   U284 : AOI222_X1 port map( A1 => n550, A2 => Q(824), B1 => n551, B2 => 
                           Q(120), C1 => n549, C2 => Q(760), ZN => n268);
   U285 : NAND3_X1 port map( A1 => n266, A2 => n267, A3 => n268, ZN => n269);
   U286 : AOI22_X1 port map( A1 => n553, A2 => Q(856), B1 => n552, B2 => Q(728)
                           , ZN => n270);
   U287 : AOI22_X1 port map( A1 => n555, A2 => Q(792), B1 => n554, B2 => Q(888)
                           , ZN => n271);
   U288 : NAND4_X1 port map( A1 => n625, A2 => n626, A3 => n270, A4 => n271, ZN
                           => n272);
   U289 : OR4_X1 port map( A1 => n260, A2 => n265, A3 => n269, A4 => n272, ZN 
                           => Y(24));
   U290 : AOI22_X1 port map( A1 => n561, A2 => Q(503), B1 => n560, B2 => Q(567)
                           , ZN => n273);
   U291 : AOI22_X1 port map( A1 => n563, A2 => Q(663), B1 => n562, B2 => Q(471)
                           , ZN => n274);
   U292 : AOI22_X1 port map( A1 => n565, A2 => Q(375), B1 => n564, B2 => Q(311)
                           , ZN => n275);
   U293 : AOI22_X1 port map( A1 => n567, A2 => Q(407), B1 => n566, B2 => Q(279)
                           , ZN => n276);
   U294 : NAND4_X1 port map( A1 => n273, A2 => n274, A3 => n275, A4 => n276, ZN
                           => n277);
   U295 : AOI22_X1 port map( A1 => n569, A2 => Q(343), B1 => n568, B2 => Q(439)
                           , ZN => n278);
   U296 : AOI22_X1 port map( A1 => n571, A2 => Q(247), B1 => n570, B2 => Q(151)
                           , ZN => n279);
   U297 : AOI22_X1 port map( A1 => n573, A2 => Q(87), B1 => n572, B2 => Q(183),
                           ZN => n280);
   U298 : AOI22_X1 port map( A1 => n575, A2 => Q(215), B1 => n574, B2 => Q(55),
                           ZN => n281);
   U299 : NAND4_X1 port map( A1 => n278, A2 => n279, A3 => n280, A4 => n281, ZN
                           => n282);
   U300 : AOI22_X1 port map( A1 => n546, A2 => Q(1015), B1 => n545, B2 => 
                           Q(951), ZN => n283);
   U301 : AOI22_X1 port map( A1 => n548, A2 => Q(983), B1 => n547, B2 => Q(919)
                           , ZN => n284);
   U302 : AOI222_X1 port map( A1 => n550, A2 => Q(823), B1 => n551, B2 => 
                           Q(119), C1 => n549, C2 => Q(759), ZN => n285);
   U303 : NAND3_X1 port map( A1 => n283, A2 => n284, A3 => n285, ZN => n286);
   U304 : AOI22_X1 port map( A1 => n553, A2 => Q(855), B1 => n552, B2 => Q(727)
                           , ZN => n287);
   U305 : AOI22_X1 port map( A1 => n555, A2 => Q(791), B1 => n554, B2 => Q(887)
                           , ZN => n288);
   U306 : NAND4_X1 port map( A1 => n623, A2 => n624, A3 => n287, A4 => n288, ZN
                           => n289);
   U307 : OR4_X1 port map( A1 => n277, A2 => n282, A3 => n286, A4 => n289, ZN 
                           => Y(23));
   U308 : AOI22_X1 port map( A1 => n561, A2 => Q(502), B1 => n560, B2 => Q(566)
                           , ZN => n290);
   U309 : AOI22_X1 port map( A1 => n563, A2 => Q(662), B1 => n562, B2 => Q(470)
                           , ZN => n291);
   U310 : AOI22_X1 port map( A1 => n565, A2 => Q(374), B1 => n564, B2 => Q(310)
                           , ZN => n292);
   U311 : AOI22_X1 port map( A1 => n567, A2 => Q(406), B1 => n566, B2 => Q(278)
                           , ZN => n293);
   U312 : NAND4_X1 port map( A1 => n290, A2 => n291, A3 => n292, A4 => n293, ZN
                           => n294);
   U313 : AOI22_X1 port map( A1 => n569, A2 => Q(342), B1 => n568, B2 => Q(438)
                           , ZN => n295);
   U314 : AOI22_X1 port map( A1 => n571, A2 => Q(246), B1 => n570, B2 => Q(150)
                           , ZN => n296);
   U315 : AOI22_X1 port map( A1 => n573, A2 => Q(86), B1 => n572, B2 => Q(182),
                           ZN => n297);
   U316 : AOI22_X1 port map( A1 => n575, A2 => Q(214), B1 => n574, B2 => Q(54),
                           ZN => n298);
   U317 : NAND4_X1 port map( A1 => n295, A2 => n296, A3 => n297, A4 => n298, ZN
                           => n299);
   U318 : AOI22_X1 port map( A1 => n546, A2 => Q(1014), B1 => n545, B2 => 
                           Q(950), ZN => n300);
   U319 : AOI22_X1 port map( A1 => n548, A2 => Q(982), B1 => n547, B2 => Q(918)
                           , ZN => n301);
   U320 : AOI222_X1 port map( A1 => n550, A2 => Q(822), B1 => n551, B2 => 
                           Q(118), C1 => n549, C2 => Q(758), ZN => n302);
   U321 : NAND3_X1 port map( A1 => n300, A2 => n301, A3 => n302, ZN => n303);
   U322 : AOI22_X1 port map( A1 => n553, A2 => Q(854), B1 => n552, B2 => Q(726)
                           , ZN => n304);
   U323 : AOI22_X1 port map( A1 => n555, A2 => Q(790), B1 => n554, B2 => Q(886)
                           , ZN => n305);
   U324 : NAND4_X1 port map( A1 => n621, A2 => n622, A3 => n304, A4 => n305, ZN
                           => n306);
   U325 : OR4_X1 port map( A1 => n294, A2 => n299, A3 => n303, A4 => n306, ZN 
                           => Y(22));
   U326 : AOI22_X1 port map( A1 => n561, A2 => Q(501), B1 => n560, B2 => Q(565)
                           , ZN => n307);
   U327 : AOI22_X1 port map( A1 => n563, A2 => Q(661), B1 => n562, B2 => Q(469)
                           , ZN => n308);
   U328 : AOI22_X1 port map( A1 => n565, A2 => Q(373), B1 => n564, B2 => Q(309)
                           , ZN => n309);
   U329 : AOI22_X1 port map( A1 => n567, A2 => Q(405), B1 => n566, B2 => Q(277)
                           , ZN => n310);
   U330 : NAND4_X1 port map( A1 => n307, A2 => n308, A3 => n309, A4 => n310, ZN
                           => n311);
   U331 : AOI22_X1 port map( A1 => n569, A2 => Q(341), B1 => n568, B2 => Q(437)
                           , ZN => n312);
   U332 : AOI22_X1 port map( A1 => n571, A2 => Q(245), B1 => n570, B2 => Q(149)
                           , ZN => n313);
   U333 : AOI22_X1 port map( A1 => n573, A2 => Q(85), B1 => n572, B2 => Q(181),
                           ZN => n314);
   U334 : AOI22_X1 port map( A1 => n575, A2 => Q(213), B1 => n574, B2 => Q(53),
                           ZN => n315);
   U335 : NAND4_X1 port map( A1 => n312, A2 => n313, A3 => n314, A4 => n315, ZN
                           => n316);
   U336 : AOI22_X1 port map( A1 => n546, A2 => Q(1013), B1 => n545, B2 => 
                           Q(949), ZN => n317);
   U337 : AOI22_X1 port map( A1 => n548, A2 => Q(981), B1 => n547, B2 => Q(917)
                           , ZN => n318);
   U338 : AOI222_X1 port map( A1 => n550, A2 => Q(821), B1 => n551, B2 => 
                           Q(117), C1 => n549, C2 => Q(757), ZN => n319);
   U339 : NAND3_X1 port map( A1 => n317, A2 => n318, A3 => n319, ZN => n320);
   U340 : AOI22_X1 port map( A1 => n553, A2 => Q(853), B1 => n552, B2 => Q(725)
                           , ZN => n321);
   U341 : AOI22_X1 port map( A1 => n555, A2 => Q(789), B1 => n554, B2 => Q(885)
                           , ZN => n322);
   U342 : NAND4_X1 port map( A1 => n619, A2 => n620, A3 => n321, A4 => n322, ZN
                           => n323);
   U343 : OR4_X1 port map( A1 => n311, A2 => n316, A3 => n320, A4 => n323, ZN 
                           => Y(21));
   U344 : AOI22_X1 port map( A1 => n561, A2 => Q(500), B1 => n560, B2 => Q(564)
                           , ZN => n324);
   U345 : AOI22_X1 port map( A1 => n563, A2 => Q(660), B1 => n562, B2 => Q(468)
                           , ZN => n325);
   U346 : AOI22_X1 port map( A1 => n565, A2 => Q(372), B1 => n564, B2 => Q(308)
                           , ZN => n326);
   U347 : AOI22_X1 port map( A1 => n567, A2 => Q(404), B1 => n566, B2 => Q(276)
                           , ZN => n327);
   U348 : NAND4_X1 port map( A1 => n324, A2 => n325, A3 => n326, A4 => n327, ZN
                           => n328);
   U349 : AOI22_X1 port map( A1 => n569, A2 => Q(340), B1 => n568, B2 => Q(436)
                           , ZN => n329);
   U350 : AOI22_X1 port map( A1 => n571, A2 => Q(244), B1 => n570, B2 => Q(148)
                           , ZN => n330);
   U351 : AOI22_X1 port map( A1 => n573, A2 => Q(84), B1 => n572, B2 => Q(180),
                           ZN => n331);
   U352 : AOI22_X1 port map( A1 => n575, A2 => Q(212), B1 => n574, B2 => Q(52),
                           ZN => n332);
   U353 : NAND4_X1 port map( A1 => n329, A2 => n330, A3 => n331, A4 => n332, ZN
                           => n333);
   U354 : AOI22_X1 port map( A1 => n546, A2 => Q(1012), B1 => n545, B2 => 
                           Q(948), ZN => n334);
   U355 : AOI22_X1 port map( A1 => n548, A2 => Q(980), B1 => n547, B2 => Q(916)
                           , ZN => n335);
   U356 : AOI222_X1 port map( A1 => n550, A2 => Q(820), B1 => n551, B2 => 
                           Q(116), C1 => n549, C2 => Q(756), ZN => n336);
   U357 : NAND3_X1 port map( A1 => n334, A2 => n335, A3 => n336, ZN => n337);
   U358 : AOI22_X1 port map( A1 => n553, A2 => Q(852), B1 => n552, B2 => Q(724)
                           , ZN => n338);
   U359 : AOI22_X1 port map( A1 => n555, A2 => Q(788), B1 => n554, B2 => Q(884)
                           , ZN => n339);
   U360 : NAND4_X1 port map( A1 => n617, A2 => n618, A3 => n338, A4 => n339, ZN
                           => n340);
   U361 : OR4_X1 port map( A1 => n328, A2 => n333, A3 => n337, A4 => n340, ZN 
                           => Y(20));
   U362 : AOI22_X1 port map( A1 => n673, A2 => Q(491), B1 => n672, B2 => Q(555)
                           , ZN => n341);
   U363 : AOI22_X1 port map( A1 => n675, A2 => Q(651), B1 => n674, B2 => Q(459)
                           , ZN => n342);
   U364 : AOI22_X1 port map( A1 => n677, A2 => Q(363), B1 => n676, B2 => Q(299)
                           , ZN => n343);
   U365 : AOI22_X1 port map( A1 => n679, A2 => Q(395), B1 => n678, B2 => Q(267)
                           , ZN => n344);
   U366 : NAND4_X1 port map( A1 => n341, A2 => n342, A3 => n343, A4 => n344, ZN
                           => n345);
   U367 : AOI22_X1 port map( A1 => n681, A2 => Q(331), B1 => n680, B2 => Q(427)
                           , ZN => n346);
   U368 : AOI22_X1 port map( A1 => n683, A2 => Q(235), B1 => n682, B2 => Q(139)
                           , ZN => n347);
   U369 : AOI22_X1 port map( A1 => n685, A2 => Q(75), B1 => n684, B2 => Q(171),
                           ZN => n348);
   U370 : AOI22_X1 port map( A1 => n687, A2 => Q(203), B1 => n686, B2 => Q(43),
                           ZN => n349);
   U371 : NAND4_X1 port map( A1 => n346, A2 => n347, A3 => n348, A4 => n349, ZN
                           => n350);
   U372 : AOI22_X1 port map( A1 => n656, A2 => Q(1003), B1 => n655, B2 => 
                           Q(939), ZN => n351);
   U373 : AOI22_X1 port map( A1 => n658, A2 => Q(971), B1 => n657, B2 => Q(907)
                           , ZN => n352);
   U374 : AOI222_X1 port map( A1 => n660, A2 => Q(811), B1 => n661, B2 => 
                           Q(107), C1 => n659, C2 => Q(747), ZN => n353);
   U375 : NAND3_X1 port map( A1 => n351, A2 => n352, A3 => n353, ZN => n354);
   U376 : AOI22_X1 port map( A1 => n663, A2 => Q(843), B1 => n662, B2 => Q(715)
                           , ZN => n355);
   U377 : AOI22_X1 port map( A1 => n665, A2 => Q(779), B1 => n664, B2 => Q(875)
                           , ZN => n356);
   U378 : NAND4_X1 port map( A1 => n597, A2 => n598, A3 => n355, A4 => n356, ZN
                           => n357);
   U379 : OR4_X1 port map( A1 => n345, A2 => n350, A3 => n354, A4 => n357, ZN 
                           => Y(11));
   U380 : AOI22_X1 port map( A1 => n561, A2 => Q(490), B1 => n560, B2 => Q(554)
                           , ZN => n358);
   U381 : AOI22_X1 port map( A1 => n563, A2 => Q(650), B1 => n562, B2 => Q(458)
                           , ZN => n359);
   U382 : AOI22_X1 port map( A1 => n565, A2 => Q(362), B1 => n564, B2 => Q(298)
                           , ZN => n360);
   U383 : AOI22_X1 port map( A1 => n567, A2 => Q(394), B1 => n566, B2 => Q(266)
                           , ZN => n361);
   U384 : NAND4_X1 port map( A1 => n358, A2 => n359, A3 => n360, A4 => n361, ZN
                           => n362);
   U385 : AOI22_X1 port map( A1 => n569, A2 => Q(330), B1 => n568, B2 => Q(426)
                           , ZN => n363);
   U386 : AOI22_X1 port map( A1 => n571, A2 => Q(234), B1 => n570, B2 => Q(138)
                           , ZN => n364);
   U387 : AOI22_X1 port map( A1 => n573, A2 => Q(74), B1 => n572, B2 => Q(170),
                           ZN => n365);
   U388 : AOI22_X1 port map( A1 => n575, A2 => Q(202), B1 => n574, B2 => Q(42),
                           ZN => n366);
   U389 : NAND4_X1 port map( A1 => n363, A2 => n364, A3 => n365, A4 => n366, ZN
                           => n367);
   U390 : AOI22_X1 port map( A1 => n546, A2 => Q(1002), B1 => n545, B2 => 
                           Q(938), ZN => n368);
   U391 : AOI22_X1 port map( A1 => n548, A2 => Q(970), B1 => n547, B2 => Q(906)
                           , ZN => n369);
   U392 : AOI222_X1 port map( A1 => n550, A2 => Q(810), B1 => n551, B2 => 
                           Q(106), C1 => n549, C2 => Q(746), ZN => n370);
   U393 : NAND3_X1 port map( A1 => n368, A2 => n369, A3 => n370, ZN => n371);
   U394 : AOI22_X1 port map( A1 => n553, A2 => Q(842), B1 => n552, B2 => Q(714)
                           , ZN => n372);
   U395 : AOI22_X1 port map( A1 => n555, A2 => Q(778), B1 => n554, B2 => Q(874)
                           , ZN => n373);
   U396 : NAND4_X1 port map( A1 => n595, A2 => n596, A3 => n372, A4 => n373, ZN
                           => n374);
   U397 : OR4_X1 port map( A1 => n362, A2 => n367, A3 => n371, A4 => n374, ZN 
                           => Y(10));
   U398 : AOI22_X1 port map( A1 => n561, A2 => Q(489), B1 => n560, B2 => Q(553)
                           , ZN => n375);
   U399 : AOI22_X1 port map( A1 => n563, A2 => Q(649), B1 => n562, B2 => Q(457)
                           , ZN => n376);
   U400 : AOI22_X1 port map( A1 => n565, A2 => Q(361), B1 => n564, B2 => Q(297)
                           , ZN => n377);
   U401 : AOI22_X1 port map( A1 => n567, A2 => Q(393), B1 => n566, B2 => Q(265)
                           , ZN => n378);
   U402 : NAND4_X1 port map( A1 => n375, A2 => n376, A3 => n377, A4 => n378, ZN
                           => n379);
   U403 : AOI22_X1 port map( A1 => n569, A2 => Q(329), B1 => n568, B2 => Q(425)
                           , ZN => n380);
   U404 : AOI22_X1 port map( A1 => n571, A2 => Q(233), B1 => n570, B2 => Q(137)
                           , ZN => n381);
   U405 : AOI22_X1 port map( A1 => n573, A2 => Q(73), B1 => n572, B2 => Q(169),
                           ZN => n382);
   U406 : AOI22_X1 port map( A1 => n575, A2 => Q(201), B1 => n574, B2 => Q(41),
                           ZN => n383);
   U407 : NAND4_X1 port map( A1 => n380, A2 => n381, A3 => n382, A4 => n383, ZN
                           => n384);
   U408 : AOI22_X1 port map( A1 => n546, A2 => Q(1001), B1 => n545, B2 => 
                           Q(937), ZN => n385);
   U409 : AOI22_X1 port map( A1 => n548, A2 => Q(969), B1 => n547, B2 => Q(905)
                           , ZN => n386);
   U410 : AOI222_X1 port map( A1 => n550, A2 => Q(809), B1 => n551, B2 => 
                           Q(105), C1 => n549, C2 => Q(745), ZN => n387);
   U411 : NAND3_X1 port map( A1 => n385, A2 => n386, A3 => n387, ZN => n388);
   U412 : AOI22_X1 port map( A1 => n553, A2 => Q(841), B1 => n552, B2 => Q(713)
                           , ZN => n389);
   U413 : AOI22_X1 port map( A1 => n555, A2 => Q(777), B1 => n554, B2 => Q(873)
                           , ZN => n390);
   U414 : NAND4_X1 port map( A1 => n670, A2 => n671, A3 => n389, A4 => n390, ZN
                           => n391);
   U415 : OR4_X1 port map( A1 => n379, A2 => n384, A3 => n388, A4 => n391, ZN 
                           => Y(9));
   U416 : AOI22_X1 port map( A1 => n561, A2 => Q(488), B1 => n560, B2 => Q(552)
                           , ZN => n392);
   U417 : AOI22_X1 port map( A1 => n563, A2 => Q(648), B1 => n562, B2 => Q(456)
                           , ZN => n393);
   U418 : AOI22_X1 port map( A1 => n565, A2 => Q(360), B1 => n564, B2 => Q(296)
                           , ZN => n394);
   U419 : AOI22_X1 port map( A1 => n567, A2 => Q(392), B1 => n566, B2 => Q(264)
                           , ZN => n395);
   U420 : NAND4_X1 port map( A1 => n392, A2 => n393, A3 => n394, A4 => n395, ZN
                           => n396);
   U421 : AOI22_X1 port map( A1 => n569, A2 => Q(328), B1 => n568, B2 => Q(424)
                           , ZN => n397);
   U422 : AOI22_X1 port map( A1 => n571, A2 => Q(232), B1 => n570, B2 => Q(136)
                           , ZN => n398);
   U423 : AOI22_X1 port map( A1 => n573, A2 => Q(72), B1 => n572, B2 => Q(168),
                           ZN => n399);
   U424 : AOI22_X1 port map( A1 => n575, A2 => Q(200), B1 => n574, B2 => Q(40),
                           ZN => n400);
   U425 : NAND4_X1 port map( A1 => n397, A2 => n398, A3 => n399, A4 => n400, ZN
                           => n401);
   U426 : AOI22_X1 port map( A1 => n546, A2 => Q(1000), B1 => n545, B2 => 
                           Q(936), ZN => n402);
   U427 : AOI22_X1 port map( A1 => n548, A2 => Q(968), B1 => n547, B2 => Q(904)
                           , ZN => n403);
   U428 : AOI222_X1 port map( A1 => n550, A2 => Q(808), B1 => n551, B2 => 
                           Q(104), C1 => n549, C2 => Q(744), ZN => n404);
   U429 : NAND3_X1 port map( A1 => n402, A2 => n403, A3 => n404, ZN => n405);
   U430 : AOI22_X1 port map( A1 => n553, A2 => Q(840), B1 => n552, B2 => Q(712)
                           , ZN => n406);
   U431 : AOI22_X1 port map( A1 => n555, A2 => Q(776), B1 => n554, B2 => Q(872)
                           , ZN => n407);
   U432 : NAND4_X1 port map( A1 => n653, A2 => n654, A3 => n406, A4 => n407, ZN
                           => n408);
   U433 : OR4_X1 port map( A1 => n396, A2 => n401, A3 => n405, A4 => n408, ZN 
                           => Y(8));
   U434 : AOI22_X1 port map( A1 => n561, A2 => Q(487), B1 => n560, B2 => Q(551)
                           , ZN => n409);
   U435 : AOI22_X1 port map( A1 => n563, A2 => Q(647), B1 => n562, B2 => Q(455)
                           , ZN => n410);
   U436 : AOI22_X1 port map( A1 => n565, A2 => Q(359), B1 => n564, B2 => Q(295)
                           , ZN => n411);
   U437 : AOI22_X1 port map( A1 => n567, A2 => Q(391), B1 => n566, B2 => Q(263)
                           , ZN => n412);
   U438 : NAND4_X1 port map( A1 => n409, A2 => n410, A3 => n411, A4 => n412, ZN
                           => n413);
   U439 : AOI22_X1 port map( A1 => n569, A2 => Q(327), B1 => n568, B2 => Q(423)
                           , ZN => n414);
   U440 : AOI22_X1 port map( A1 => n571, A2 => Q(231), B1 => n570, B2 => Q(135)
                           , ZN => n415);
   U441 : AOI22_X1 port map( A1 => n573, A2 => Q(71), B1 => n572, B2 => Q(167),
                           ZN => n416);
   U442 : AOI22_X1 port map( A1 => n575, A2 => Q(199), B1 => n574, B2 => Q(39),
                           ZN => n417);
   U443 : NAND4_X1 port map( A1 => n414, A2 => n415, A3 => n416, A4 => n417, ZN
                           => n418);
   U444 : AOI22_X1 port map( A1 => n546, A2 => Q(999), B1 => n545, B2 => Q(935)
                           , ZN => n419);
   U445 : AOI22_X1 port map( A1 => n548, A2 => Q(967), B1 => n547, B2 => Q(903)
                           , ZN => n420);
   U446 : AOI222_X1 port map( A1 => n550, A2 => Q(807), B1 => n551, B2 => 
                           Q(103), C1 => n549, C2 => Q(743), ZN => n421);
   U447 : NAND3_X1 port map( A1 => n419, A2 => n420, A3 => n421, ZN => n422);
   U448 : AOI22_X1 port map( A1 => n553, A2 => Q(839), B1 => n552, B2 => Q(711)
                           , ZN => n423);
   U449 : AOI22_X1 port map( A1 => n555, A2 => Q(775), B1 => n554, B2 => Q(871)
                           , ZN => n424);
   U450 : NAND4_X1 port map( A1 => n651, A2 => n652, A3 => n423, A4 => n424, ZN
                           => n425);
   U451 : OR4_X1 port map( A1 => n413, A2 => n418, A3 => n422, A4 => n425, ZN 
                           => Y(7));
   U452 : AOI22_X1 port map( A1 => n561, A2 => Q(486), B1 => n560, B2 => Q(550)
                           , ZN => n426);
   U453 : AOI22_X1 port map( A1 => n563, A2 => Q(646), B1 => n562, B2 => Q(454)
                           , ZN => n427);
   U454 : AOI22_X1 port map( A1 => n565, A2 => Q(358), B1 => n564, B2 => Q(294)
                           , ZN => n428);
   U455 : AOI22_X1 port map( A1 => n567, A2 => Q(390), B1 => n566, B2 => Q(262)
                           , ZN => n429);
   U456 : NAND4_X1 port map( A1 => n426, A2 => n427, A3 => n428, A4 => n429, ZN
                           => n430);
   U457 : AOI22_X1 port map( A1 => n569, A2 => Q(326), B1 => n568, B2 => Q(422)
                           , ZN => n431);
   U458 : AOI22_X1 port map( A1 => n571, A2 => Q(230), B1 => n570, B2 => Q(134)
                           , ZN => n432);
   U459 : AOI22_X1 port map( A1 => n573, A2 => Q(70), B1 => n572, B2 => Q(166),
                           ZN => n433);
   U460 : AOI22_X1 port map( A1 => n575, A2 => Q(198), B1 => n574, B2 => Q(38),
                           ZN => n434);
   U461 : NAND4_X1 port map( A1 => n431, A2 => n432, A3 => n433, A4 => n434, ZN
                           => n435);
   U462 : AOI22_X1 port map( A1 => n546, A2 => Q(998), B1 => n545, B2 => Q(934)
                           , ZN => n436);
   U463 : AOI22_X1 port map( A1 => n548, A2 => Q(966), B1 => n547, B2 => Q(902)
                           , ZN => n437);
   U464 : AOI222_X1 port map( A1 => n550, A2 => Q(806), B1 => n551, B2 => 
                           Q(102), C1 => n549, C2 => Q(742), ZN => n438);
   U465 : NAND3_X1 port map( A1 => n436, A2 => n437, A3 => n438, ZN => n439);
   U466 : AOI22_X1 port map( A1 => n553, A2 => Q(838), B1 => n552, B2 => Q(710)
                           , ZN => n440);
   U467 : AOI22_X1 port map( A1 => n555, A2 => Q(774), B1 => n554, B2 => Q(870)
                           , ZN => n441);
   U468 : NAND4_X1 port map( A1 => n649, A2 => n650, A3 => n440, A4 => n441, ZN
                           => n442);
   U469 : OR4_X1 port map( A1 => n430, A2 => n435, A3 => n439, A4 => n442, ZN 
                           => Y(6));
   U470 : AOI22_X1 port map( A1 => n561, A2 => Q(485), B1 => n560, B2 => Q(549)
                           , ZN => n443);
   U471 : AOI22_X1 port map( A1 => n563, A2 => Q(645), B1 => n562, B2 => Q(453)
                           , ZN => n444);
   U472 : AOI22_X1 port map( A1 => n565, A2 => Q(357), B1 => n564, B2 => Q(293)
                           , ZN => n445);
   U473 : AOI22_X1 port map( A1 => n567, A2 => Q(389), B1 => n566, B2 => Q(261)
                           , ZN => n446);
   U474 : NAND4_X1 port map( A1 => n443, A2 => n444, A3 => n445, A4 => n446, ZN
                           => n447);
   U475 : AOI22_X1 port map( A1 => n569, A2 => Q(325), B1 => n568, B2 => Q(421)
                           , ZN => n448);
   U476 : AOI22_X1 port map( A1 => n571, A2 => Q(229), B1 => n570, B2 => Q(133)
                           , ZN => n449);
   U477 : AOI22_X1 port map( A1 => n573, A2 => Q(69), B1 => n572, B2 => Q(165),
                           ZN => n450);
   U478 : AOI22_X1 port map( A1 => n575, A2 => Q(197), B1 => n574, B2 => Q(37),
                           ZN => n451);
   U479 : NAND4_X1 port map( A1 => n448, A2 => n449, A3 => n450, A4 => n451, ZN
                           => n452);
   U480 : AOI22_X1 port map( A1 => n546, A2 => Q(997), B1 => n545, B2 => Q(933)
                           , ZN => n453);
   U481 : AOI22_X1 port map( A1 => n548, A2 => Q(965), B1 => n547, B2 => Q(901)
                           , ZN => n454);
   U482 : AOI222_X1 port map( A1 => n550, A2 => Q(805), B1 => n551, B2 => 
                           Q(101), C1 => n549, C2 => Q(741), ZN => n455);
   U483 : NAND3_X1 port map( A1 => n453, A2 => n454, A3 => n455, ZN => n456);
   U484 : AOI22_X1 port map( A1 => n553, A2 => Q(837), B1 => n552, B2 => Q(709)
                           , ZN => n457);
   U485 : AOI22_X1 port map( A1 => n555, A2 => Q(773), B1 => n554, B2 => Q(869)
                           , ZN => n458);
   U486 : NAND4_X1 port map( A1 => n647, A2 => n648, A3 => n457, A4 => n458, ZN
                           => n459);
   U487 : OR4_X1 port map( A1 => n447, A2 => n452, A3 => n456, A4 => n459, ZN 
                           => Y(5));
   U488 : AOI22_X1 port map( A1 => n561, A2 => Q(484), B1 => n560, B2 => Q(548)
                           , ZN => n460);
   U489 : AOI22_X1 port map( A1 => n563, A2 => Q(644), B1 => n562, B2 => Q(452)
                           , ZN => n461);
   U490 : AOI22_X1 port map( A1 => n565, A2 => Q(356), B1 => n564, B2 => Q(292)
                           , ZN => n462);
   U491 : AOI22_X1 port map( A1 => n567, A2 => Q(388), B1 => n566, B2 => Q(260)
                           , ZN => n463);
   U492 : NAND4_X1 port map( A1 => n460, A2 => n461, A3 => n462, A4 => n463, ZN
                           => n464);
   U493 : AOI22_X1 port map( A1 => n569, A2 => Q(324), B1 => n568, B2 => Q(420)
                           , ZN => n465);
   U494 : AOI22_X1 port map( A1 => n571, A2 => Q(228), B1 => n570, B2 => Q(132)
                           , ZN => n466);
   U495 : AOI22_X1 port map( A1 => n573, A2 => Q(68), B1 => n572, B2 => Q(164),
                           ZN => n467);
   U496 : AOI22_X1 port map( A1 => n575, A2 => Q(196), B1 => n574, B2 => Q(36),
                           ZN => n468);
   U497 : NAND4_X1 port map( A1 => n465, A2 => n466, A3 => n467, A4 => n468, ZN
                           => n469);
   U498 : AOI22_X1 port map( A1 => n546, A2 => Q(996), B1 => n545, B2 => Q(932)
                           , ZN => n470);
   U499 : AOI22_X1 port map( A1 => n548, A2 => Q(964), B1 => n547, B2 => Q(900)
                           , ZN => n471);
   U500 : AOI222_X1 port map( A1 => n550, A2 => Q(804), B1 => n551, B2 => 
                           Q(100), C1 => n549, C2 => Q(740), ZN => n472);
   U501 : NAND3_X1 port map( A1 => n470, A2 => n471, A3 => n472, ZN => n473);
   U502 : AOI22_X1 port map( A1 => n553, A2 => Q(836), B1 => n552, B2 => Q(708)
                           , ZN => n474);
   U503 : AOI22_X1 port map( A1 => n555, A2 => Q(772), B1 => n554, B2 => Q(868)
                           , ZN => n475);
   U504 : NAND4_X1 port map( A1 => n645, A2 => n646, A3 => n474, A4 => n475, ZN
                           => n476);
   U505 : OR4_X1 port map( A1 => n464, A2 => n469, A3 => n473, A4 => n476, ZN 
                           => Y(4));
   U506 : AOI22_X1 port map( A1 => n561, A2 => Q(483), B1 => n560, B2 => Q(547)
                           , ZN => n477);
   U507 : AOI22_X1 port map( A1 => n563, A2 => Q(643), B1 => n562, B2 => Q(451)
                           , ZN => n478);
   U508 : AOI22_X1 port map( A1 => n565, A2 => Q(355), B1 => n564, B2 => Q(291)
                           , ZN => n479);
   U509 : AOI22_X1 port map( A1 => n567, A2 => Q(387), B1 => n566, B2 => Q(259)
                           , ZN => n480);
   U510 : NAND4_X1 port map( A1 => n477, A2 => n478, A3 => n479, A4 => n480, ZN
                           => n481);
   U511 : AOI22_X1 port map( A1 => n569, A2 => Q(323), B1 => n568, B2 => Q(419)
                           , ZN => n482);
   U512 : AOI22_X1 port map( A1 => n571, A2 => Q(227), B1 => n570, B2 => Q(131)
                           , ZN => n483);
   U513 : AOI22_X1 port map( A1 => n573, A2 => Q(67), B1 => n572, B2 => Q(163),
                           ZN => n484);
   U514 : AOI22_X1 port map( A1 => n575, A2 => Q(195), B1 => n574, B2 => Q(35),
                           ZN => n485);
   U515 : NAND4_X1 port map( A1 => n482, A2 => n483, A3 => n484, A4 => n485, ZN
                           => n486);
   U516 : AOI22_X1 port map( A1 => n546, A2 => Q(995), B1 => n545, B2 => Q(931)
                           , ZN => n487);
   U517 : AOI22_X1 port map( A1 => n548, A2 => Q(963), B1 => n547, B2 => Q(899)
                           , ZN => n488);
   U518 : AOI222_X1 port map( A1 => n550, A2 => Q(803), B1 => n551, B2 => Q(99)
                           , C1 => n549, C2 => Q(739), ZN => n489);
   U519 : NAND3_X1 port map( A1 => n487, A2 => n488, A3 => n489, ZN => n490);
   U520 : AOI22_X1 port map( A1 => n553, A2 => Q(835), B1 => n552, B2 => Q(707)
                           , ZN => n491);
   U521 : AOI22_X1 port map( A1 => n555, A2 => Q(771), B1 => n554, B2 => Q(867)
                           , ZN => n492);
   U522 : NAND4_X1 port map( A1 => n643, A2 => n644, A3 => n491, A4 => n492, ZN
                           => n493);
   U523 : OR4_X1 port map( A1 => n481, A2 => n486, A3 => n490, A4 => n493, ZN 
                           => Y(3));
   U524 : AOI22_X1 port map( A1 => n561, A2 => Q(482), B1 => n560, B2 => Q(546)
                           , ZN => n494);
   U525 : AOI22_X1 port map( A1 => n563, A2 => Q(642), B1 => n562, B2 => Q(450)
                           , ZN => n495);
   U526 : AOI22_X1 port map( A1 => n565, A2 => Q(354), B1 => n564, B2 => Q(290)
                           , ZN => n496);
   U527 : AOI22_X1 port map( A1 => n567, A2 => Q(386), B1 => n566, B2 => Q(258)
                           , ZN => n497);
   U528 : NAND4_X1 port map( A1 => n494, A2 => n495, A3 => n496, A4 => n497, ZN
                           => n498);
   U529 : AOI22_X1 port map( A1 => n569, A2 => Q(322), B1 => n568, B2 => Q(418)
                           , ZN => n499);
   U530 : AOI22_X1 port map( A1 => n571, A2 => Q(226), B1 => n570, B2 => Q(130)
                           , ZN => n500);
   U531 : AOI22_X1 port map( A1 => n573, A2 => Q(66), B1 => n572, B2 => Q(162),
                           ZN => n501);
   U532 : AOI22_X1 port map( A1 => n575, A2 => Q(194), B1 => n574, B2 => Q(34),
                           ZN => n502);
   U533 : NAND4_X1 port map( A1 => n499, A2 => n500, A3 => n501, A4 => n502, ZN
                           => n503);
   U534 : AOI22_X1 port map( A1 => n546, A2 => Q(994), B1 => n545, B2 => Q(930)
                           , ZN => n504);
   U535 : AOI22_X1 port map( A1 => n548, A2 => Q(962), B1 => n547, B2 => Q(898)
                           , ZN => n505);
   U536 : AOI222_X1 port map( A1 => n550, A2 => Q(802), B1 => n551, B2 => Q(98)
                           , C1 => n549, C2 => Q(738), ZN => n506);
   U537 : NAND3_X1 port map( A1 => n504, A2 => n505, A3 => n506, ZN => n507);
   U538 : AOI22_X1 port map( A1 => n553, A2 => Q(834), B1 => n552, B2 => Q(706)
                           , ZN => n508);
   U539 : AOI22_X1 port map( A1 => n555, A2 => Q(770), B1 => n554, B2 => Q(866)
                           , ZN => n509);
   U540 : NAND4_X1 port map( A1 => n637, A2 => n638, A3 => n508, A4 => n509, ZN
                           => n510);
   U541 : OR4_X1 port map( A1 => n498, A2 => n503, A3 => n507, A4 => n510, ZN 
                           => Y(2));
   U542 : AOI22_X1 port map( A1 => n561, A2 => Q(481), B1 => n560, B2 => Q(545)
                           , ZN => n511);
   U543 : AOI22_X1 port map( A1 => n563, A2 => Q(641), B1 => n562, B2 => Q(449)
                           , ZN => n512);
   U544 : AOI22_X1 port map( A1 => n565, A2 => Q(353), B1 => n564, B2 => Q(289)
                           , ZN => n513);
   U545 : AOI22_X1 port map( A1 => n567, A2 => Q(385), B1 => n566, B2 => Q(257)
                           , ZN => n514);
   U546 : NAND4_X1 port map( A1 => n511, A2 => n512, A3 => n513, A4 => n514, ZN
                           => n515);
   U547 : AOI22_X1 port map( A1 => n569, A2 => Q(321), B1 => n568, B2 => Q(417)
                           , ZN => n516);
   U548 : AOI22_X1 port map( A1 => n571, A2 => Q(225), B1 => n570, B2 => Q(129)
                           , ZN => n517);
   U549 : AOI22_X1 port map( A1 => n573, A2 => Q(65), B1 => n572, B2 => Q(161),
                           ZN => n518);
   U550 : AOI22_X1 port map( A1 => n575, A2 => Q(193), B1 => n574, B2 => Q(33),
                           ZN => n519);
   U551 : NAND4_X1 port map( A1 => n516, A2 => n517, A3 => n518, A4 => n519, ZN
                           => n520);
   U552 : AOI22_X1 port map( A1 => n546, A2 => Q(993), B1 => n545, B2 => Q(929)
                           , ZN => n521);
   U553 : AOI22_X1 port map( A1 => n548, A2 => Q(961), B1 => n547, B2 => Q(897)
                           , ZN => n522);
   U554 : AOI222_X1 port map( A1 => n550, A2 => Q(801), B1 => n551, B2 => Q(97)
                           , C1 => n549, C2 => Q(737), ZN => n523);
   U555 : NAND3_X1 port map( A1 => n521, A2 => n522, A3 => n523, ZN => n524);
   U556 : AOI22_X1 port map( A1 => n553, A2 => Q(833), B1 => n552, B2 => Q(705)
                           , ZN => n525);
   U557 : AOI22_X1 port map( A1 => n555, A2 => Q(769), B1 => n554, B2 => Q(865)
                           , ZN => n526);
   U558 : NAND4_X1 port map( A1 => n615, A2 => n616, A3 => n525, A4 => n526, ZN
                           => n527);
   U559 : OR4_X1 port map( A1 => n515, A2 => n520, A3 => n524, A4 => n527, ZN 
                           => Y(1));
   U560 : AOI22_X1 port map( A1 => n561, A2 => Q(480), B1 => n560, B2 => Q(544)
                           , ZN => n528);
   U561 : AOI22_X1 port map( A1 => n563, A2 => Q(640), B1 => n562, B2 => Q(448)
                           , ZN => n529);
   U562 : AOI22_X1 port map( A1 => n565, A2 => Q(352), B1 => n564, B2 => Q(288)
                           , ZN => n530);
   U563 : AOI22_X1 port map( A1 => n567, A2 => Q(384), B1 => n566, B2 => Q(256)
                           , ZN => n531);
   U564 : NAND4_X1 port map( A1 => n528, A2 => n529, A3 => n530, A4 => n531, ZN
                           => n532);
   U565 : AOI22_X1 port map( A1 => n569, A2 => Q(320), B1 => n568, B2 => Q(416)
                           , ZN => n533);
   U566 : AOI22_X1 port map( A1 => n571, A2 => Q(224), B1 => n570, B2 => Q(128)
                           , ZN => n534);
   U567 : AOI22_X1 port map( A1 => n573, A2 => Q(64), B1 => n572, B2 => Q(160),
                           ZN => n535);
   U568 : AOI22_X1 port map( A1 => n575, A2 => Q(192), B1 => n574, B2 => Q(32),
                           ZN => n536);
   U569 : NAND4_X1 port map( A1 => n533, A2 => n534, A3 => n535, A4 => n536, ZN
                           => n537);
   U570 : AOI22_X1 port map( A1 => n546, A2 => Q(992), B1 => n545, B2 => Q(928)
                           , ZN => n538);
   U571 : AOI22_X1 port map( A1 => n548, A2 => Q(960), B1 => n547, B2 => Q(896)
                           , ZN => n539);
   U572 : AOI222_X1 port map( A1 => n550, A2 => Q(800), B1 => n551, B2 => Q(96)
                           , C1 => n549, C2 => Q(736), ZN => n540);
   U573 : NAND3_X1 port map( A1 => n538, A2 => n539, A3 => n540, ZN => n541);
   U574 : AOI22_X1 port map( A1 => n553, A2 => Q(832), B1 => n552, B2 => Q(704)
                           , ZN => n542);
   U575 : AOI22_X1 port map( A1 => n555, A2 => Q(768), B1 => n554, B2 => Q(864)
                           , ZN => n543);
   U576 : NAND4_X1 port map( A1 => n580, A2 => n581, A3 => n542, A4 => n543, ZN
                           => n544);
   U577 : OR4_X1 port map( A1 => n532, A2 => n537, A3 => n541, A4 => n544, ZN 
                           => Y(0));
   U578 : BUF_X1 port map( A => n686, Z => n574);
   U579 : BUF_X1 port map( A => n687, Z => n575);
   U580 : BUF_X1 port map( A => n684, Z => n572);
   U581 : BUF_X1 port map( A => n685, Z => n573);
   U582 : BUF_X1 port map( A => n682, Z => n570);
   U583 : BUF_X1 port map( A => n683, Z => n571);
   U584 : BUF_X1 port map( A => n680, Z => n568);
   U585 : BUF_X1 port map( A => n681, Z => n569);
   U586 : BUF_X1 port map( A => n678, Z => n566);
   U587 : BUF_X1 port map( A => n679, Z => n567);
   U588 : BUF_X1 port map( A => n676, Z => n564);
   U589 : BUF_X1 port map( A => n677, Z => n565);
   U590 : BUF_X1 port map( A => n674, Z => n562);
   U591 : BUF_X1 port map( A => n675, Z => n563);
   U592 : BUF_X1 port map( A => n672, Z => n560);
   U593 : BUF_X1 port map( A => n673, Z => n561);
   U594 : BUF_X1 port map( A => n668, Z => n558);
   U595 : BUF_X1 port map( A => n669, Z => n559);
   U596 : BUF_X1 port map( A => n666, Z => n556);
   U597 : BUF_X1 port map( A => n667, Z => n557);
   U598 : BUF_X1 port map( A => n664, Z => n554);
   U599 : BUF_X1 port map( A => n665, Z => n555);
   U600 : BUF_X1 port map( A => n662, Z => n552);
   U601 : BUF_X1 port map( A => n663, Z => n553);
   U602 : BUF_X1 port map( A => n661, Z => n551);
   U603 : BUF_X1 port map( A => n659, Z => n549);
   U604 : BUF_X1 port map( A => n660, Z => n550);
   U605 : OR2_X1 port map( A1 => S(1), A2 => S(2), ZN => n593);
   U606 : BUF_X1 port map( A => n657, Z => n547);
   U607 : BUF_X1 port map( A => n658, Z => n548);
   U608 : BUF_X1 port map( A => n655, Z => n545);
   U609 : OR2_X1 port map( A1 => n576, A2 => S(1), ZN => n590);
   U610 : BUF_X1 port map( A => n656, Z => n546);
   U611 : NAND2_X1 port map( A1 => S(1), A2 => S(2), ZN => n592);
   U612 : NAND3_X1 port map( A1 => S(3), A2 => S(4), A3 => S(0), ZN => n579);
   U613 : NOR2_X1 port map( A1 => n592, A2 => n579, ZN => n656);
   U614 : INV_X1 port map( A => S(2), ZN => n576);
   U615 : NOR2_X1 port map( A1 => n579, A2 => n590, ZN => n655);
   U616 : INV_X1 port map( A => S(0), ZN => n577);
   U617 : NAND3_X1 port map( A1 => S(4), A2 => S(3), A3 => n577, ZN => n578);
   U618 : NOR2_X1 port map( A1 => n592, A2 => n578, ZN => n658);
   U619 : NOR2_X1 port map( A1 => n590, A2 => n578, ZN => n657);
   U620 : NOR2_X1 port map( A1 => n579, A2 => n593, ZN => n660);
   U621 : INV_X1 port map( A => S(3), ZN => n587);
   U622 : NAND3_X1 port map( A1 => S(4), A2 => S(0), A3 => n587, ZN => n583);
   U623 : NOR2_X1 port map( A1 => n592, A2 => n583, ZN => n659);
   U624 : NAND2_X1 port map( A1 => S(1), A2 => n576, ZN => n589);
   U625 : INV_X1 port map( A => S(4), ZN => n582);
   U626 : NAND3_X1 port map( A1 => S(0), A2 => n587, A3 => n582, ZN => n594);
   U627 : NOR2_X1 port map( A1 => n589, A2 => n594, ZN => n661);
   U628 : NOR2_X1 port map( A1 => n589, A2 => n578, ZN => n663);
   U629 : NAND3_X1 port map( A1 => S(4), A2 => n587, A3 => n577, ZN => n584);
   U630 : NOR2_X1 port map( A1 => n592, A2 => n584, ZN => n662);
   U631 : NOR2_X1 port map( A1 => n578, A2 => n593, ZN => n665);
   U632 : NOR2_X1 port map( A1 => n589, A2 => n579, ZN => n664);
   U633 : NOR2_X1 port map( A1 => n590, A2 => n583, ZN => n667);
   U634 : NOR2_X1 port map( A1 => n589, A2 => n584, ZN => n666);
   U635 : AOI22_X1 port map( A1 => n557, A2 => Q(672), B1 => n556, B2 => Q(576)
                           , ZN => n581);
   U636 : NOR2_X1 port map( A1 => n593, A2 => n584, ZN => n669);
   U637 : NOR2_X1 port map( A1 => n589, A2 => n583, ZN => n668);
   U638 : AOI22_X1 port map( A1 => n559, A2 => Q(512), B1 => n558, B2 => Q(608)
                           , ZN => n580);
   U639 : NAND3_X1 port map( A1 => S(3), A2 => S(0), A3 => n582, ZN => n586);
   U640 : NOR2_X1 port map( A1 => n592, A2 => n586, ZN => n673);
   U641 : NOR2_X1 port map( A1 => n593, A2 => n583, ZN => n672);
   U642 : NOR2_X1 port map( A1 => n590, A2 => n584, ZN => n675);
   U643 : NOR2_X1 port map( A1 => S(4), A2 => S(0), ZN => n588);
   U644 : NAND2_X1 port map( A1 => S(3), A2 => n588, ZN => n585);
   U645 : NOR2_X1 port map( A1 => n592, A2 => n585, ZN => n674);
   U646 : NOR2_X1 port map( A1 => n589, A2 => n586, ZN => n677);
   U647 : NOR2_X1 port map( A1 => n593, A2 => n586, ZN => n676);
   U648 : NOR2_X1 port map( A1 => n590, A2 => n585, ZN => n679);
   U649 : NOR2_X1 port map( A1 => n593, A2 => n585, ZN => n678);
   U650 : NOR2_X1 port map( A1 => n589, A2 => n585, ZN => n681);
   U651 : NOR2_X1 port map( A1 => n590, A2 => n586, ZN => n680);
   U652 : NOR2_X1 port map( A1 => n594, A2 => n592, ZN => n683);
   U653 : NAND2_X1 port map( A1 => n588, A2 => n587, ZN => n591);
   U654 : NOR2_X1 port map( A1 => n590, A2 => n591, ZN => n682);
   U655 : NOR2_X1 port map( A1 => n589, A2 => n591, ZN => n685);
   U656 : NOR2_X1 port map( A1 => n594, A2 => n590, ZN => n684);
   U657 : NOR2_X1 port map( A1 => n592, A2 => n591, ZN => n687);
   U658 : NOR2_X1 port map( A1 => n594, A2 => n593, ZN => n686);
   U659 : AOI22_X1 port map( A1 => n557, A2 => Q(682), B1 => n556, B2 => Q(586)
                           , ZN => n596);
   U660 : AOI22_X1 port map( A1 => n559, A2 => Q(522), B1 => n558, B2 => Q(618)
                           , ZN => n595);
   U661 : AOI22_X1 port map( A1 => n667, A2 => Q(683), B1 => n666, B2 => Q(587)
                           , ZN => n598);
   U662 : AOI22_X1 port map( A1 => n669, A2 => Q(523), B1 => n668, B2 => Q(619)
                           , ZN => n597);
   U663 : AOI22_X1 port map( A1 => n667, A2 => Q(684), B1 => n666, B2 => Q(588)
                           , ZN => n600);
   U664 : AOI22_X1 port map( A1 => n669, A2 => Q(524), B1 => n668, B2 => Q(620)
                           , ZN => n599);
   U665 : AOI22_X1 port map( A1 => n667, A2 => Q(685), B1 => n666, B2 => Q(589)
                           , ZN => n602);
   U666 : AOI22_X1 port map( A1 => n669, A2 => Q(525), B1 => n668, B2 => Q(621)
                           , ZN => n601);
   U667 : AOI22_X1 port map( A1 => n667, A2 => Q(686), B1 => n666, B2 => Q(590)
                           , ZN => n604);
   U668 : AOI22_X1 port map( A1 => n669, A2 => Q(526), B1 => n668, B2 => Q(622)
                           , ZN => n603);
   U669 : AOI22_X1 port map( A1 => n667, A2 => Q(687), B1 => n666, B2 => Q(591)
                           , ZN => n606);
   U670 : AOI22_X1 port map( A1 => n669, A2 => Q(527), B1 => n668, B2 => Q(623)
                           , ZN => n605);
   U671 : AOI22_X1 port map( A1 => n667, A2 => Q(688), B1 => n666, B2 => Q(592)
                           , ZN => n608);
   U672 : AOI22_X1 port map( A1 => n669, A2 => Q(528), B1 => n668, B2 => Q(624)
                           , ZN => n607);
   U673 : AOI22_X1 port map( A1 => n667, A2 => Q(689), B1 => n666, B2 => Q(593)
                           , ZN => n610);
   U674 : AOI22_X1 port map( A1 => n669, A2 => Q(529), B1 => n668, B2 => Q(625)
                           , ZN => n609);
   U675 : AOI22_X1 port map( A1 => n667, A2 => Q(690), B1 => n666, B2 => Q(594)
                           , ZN => n612);
   U676 : AOI22_X1 port map( A1 => n669, A2 => Q(530), B1 => n668, B2 => Q(626)
                           , ZN => n611);
   U677 : AOI22_X1 port map( A1 => n667, A2 => Q(691), B1 => n666, B2 => Q(595)
                           , ZN => n614);
   U678 : AOI22_X1 port map( A1 => n669, A2 => Q(531), B1 => n668, B2 => Q(627)
                           , ZN => n613);
   U679 : AOI22_X1 port map( A1 => n557, A2 => Q(673), B1 => n556, B2 => Q(577)
                           , ZN => n616);
   U680 : AOI22_X1 port map( A1 => n559, A2 => Q(513), B1 => n558, B2 => Q(609)
                           , ZN => n615);
   U681 : AOI22_X1 port map( A1 => n557, A2 => Q(692), B1 => n556, B2 => Q(596)
                           , ZN => n618);
   U682 : AOI22_X1 port map( A1 => n559, A2 => Q(532), B1 => n558, B2 => Q(628)
                           , ZN => n617);
   U683 : AOI22_X1 port map( A1 => n557, A2 => Q(693), B1 => n556, B2 => Q(597)
                           , ZN => n620);
   U684 : AOI22_X1 port map( A1 => n559, A2 => Q(533), B1 => n558, B2 => Q(629)
                           , ZN => n619);
   U685 : AOI22_X1 port map( A1 => n557, A2 => Q(694), B1 => n556, B2 => Q(598)
                           , ZN => n622);
   U686 : AOI22_X1 port map( A1 => n559, A2 => Q(534), B1 => n558, B2 => Q(630)
                           , ZN => n621);
   U687 : AOI22_X1 port map( A1 => n557, A2 => Q(695), B1 => n556, B2 => Q(599)
                           , ZN => n624);
   U688 : AOI22_X1 port map( A1 => n559, A2 => Q(535), B1 => n558, B2 => Q(631)
                           , ZN => n623);
   U689 : AOI22_X1 port map( A1 => n557, A2 => Q(696), B1 => n556, B2 => Q(600)
                           , ZN => n626);
   U690 : AOI22_X1 port map( A1 => n559, A2 => Q(536), B1 => n558, B2 => Q(632)
                           , ZN => n625);
   U691 : AOI22_X1 port map( A1 => n557, A2 => Q(697), B1 => n556, B2 => Q(601)
                           , ZN => n628);
   U692 : AOI22_X1 port map( A1 => n559, A2 => Q(537), B1 => n558, B2 => Q(633)
                           , ZN => n627);
   U693 : AOI22_X1 port map( A1 => n557, A2 => Q(698), B1 => n556, B2 => Q(602)
                           , ZN => n630);
   U694 : AOI22_X1 port map( A1 => n559, A2 => Q(538), B1 => n558, B2 => Q(634)
                           , ZN => n629);
   U695 : AOI22_X1 port map( A1 => n557, A2 => Q(699), B1 => n556, B2 => Q(603)
                           , ZN => n632);
   U696 : AOI22_X1 port map( A1 => n559, A2 => Q(539), B1 => n558, B2 => Q(635)
                           , ZN => n631);
   U697 : AOI22_X1 port map( A1 => n557, A2 => Q(700), B1 => n556, B2 => Q(604)
                           , ZN => n634);
   U698 : AOI22_X1 port map( A1 => n559, A2 => Q(540), B1 => n558, B2 => Q(636)
                           , ZN => n633);
   U699 : AOI22_X1 port map( A1 => n667, A2 => Q(701), B1 => n666, B2 => Q(605)
                           , ZN => n636);
   U700 : AOI22_X1 port map( A1 => n669, A2 => Q(541), B1 => n668, B2 => Q(637)
                           , ZN => n635);
   U701 : AOI22_X1 port map( A1 => n557, A2 => Q(674), B1 => n556, B2 => Q(578)
                           , ZN => n638);
   U702 : AOI22_X1 port map( A1 => n559, A2 => Q(514), B1 => n558, B2 => Q(610)
                           , ZN => n637);
   U703 : AOI22_X1 port map( A1 => n557, A2 => Q(702), B1 => n556, B2 => Q(606)
                           , ZN => n640);
   U704 : AOI22_X1 port map( A1 => n559, A2 => Q(542), B1 => n558, B2 => Q(638)
                           , ZN => n639);
   U705 : AOI22_X1 port map( A1 => n557, A2 => Q(703), B1 => n556, B2 => Q(607)
                           , ZN => n642);
   U706 : AOI22_X1 port map( A1 => n559, A2 => Q(543), B1 => n558, B2 => Q(639)
                           , ZN => n641);
   U707 : AOI22_X1 port map( A1 => n557, A2 => Q(675), B1 => n556, B2 => Q(579)
                           , ZN => n644);
   U708 : AOI22_X1 port map( A1 => n559, A2 => Q(515), B1 => n558, B2 => Q(611)
                           , ZN => n643);
   U709 : AOI22_X1 port map( A1 => n557, A2 => Q(676), B1 => n556, B2 => Q(580)
                           , ZN => n646);
   U710 : AOI22_X1 port map( A1 => n559, A2 => Q(516), B1 => n558, B2 => Q(612)
                           , ZN => n645);
   U711 : AOI22_X1 port map( A1 => n557, A2 => Q(677), B1 => n556, B2 => Q(581)
                           , ZN => n648);
   U712 : AOI22_X1 port map( A1 => n559, A2 => Q(517), B1 => n558, B2 => Q(613)
                           , ZN => n647);
   U713 : AOI22_X1 port map( A1 => n557, A2 => Q(678), B1 => n556, B2 => Q(582)
                           , ZN => n650);
   U714 : AOI22_X1 port map( A1 => n559, A2 => Q(518), B1 => n558, B2 => Q(614)
                           , ZN => n649);
   U715 : AOI22_X1 port map( A1 => n557, A2 => Q(679), B1 => n556, B2 => Q(583)
                           , ZN => n652);
   U716 : AOI22_X1 port map( A1 => n559, A2 => Q(519), B1 => n558, B2 => Q(615)
                           , ZN => n651);
   U717 : AOI22_X1 port map( A1 => n557, A2 => Q(680), B1 => n556, B2 => Q(584)
                           , ZN => n654);
   U718 : AOI22_X1 port map( A1 => n559, A2 => Q(520), B1 => n558, B2 => Q(616)
                           , ZN => n653);
   U719 : AOI22_X1 port map( A1 => n557, A2 => Q(681), B1 => n556, B2 => Q(585)
                           , ZN => n671);
   U720 : AOI22_X1 port map( A1 => n559, A2 => Q(521), B1 => n558, B2 => Q(617)
                           , ZN => n670);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32.all;

entity select_block_NBIT_DATA32_N8_F5 is

   port( regs : in std_logic_vector (2559 downto 0);  win : in std_logic_vector
         (4 downto 0);  curr_proc_regs : out std_logic_vector (767 downto 0));

end select_block_NBIT_DATA32_N8_F5;

architecture SYN_behav of select_block_NBIT_DATA32_N8_F5 is

   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X16
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, 
      n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46
      , n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, 
      n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, 
      n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, 
      n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, 
      n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, 
      n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, 
      n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, 
      n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, 
      n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, 
      n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
      n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, 
      n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, 
      n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, 
      n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
      n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, 
      n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, 
      n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, 
      n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, 
      n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, 
      n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, 
      n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, 
      n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, 
      n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, 
      n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, 
      n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, 
      n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, 
      n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, 
      n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, 
      n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, 
      n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, 
      n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, 
      n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, 
      n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, 
      n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, 
      n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, 
      n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, 
      n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, 
      n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, 
      n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, 
      n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, 
      n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, 
      n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, 
      n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, 
      n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, 
      n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, 
      n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, 
      n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, 
      n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, 
      n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
      n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, 
      n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
      n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, 
      n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, 
      n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
      n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
      n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, 
      n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, 
      n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, 
      n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, 
      n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, 
      n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, 
      n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, 
      n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, 
      n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, 
      n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, 
      n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, 
      n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, 
      n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, 
      n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, 
      n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, 
      n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, 
      n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, 
      n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, 
      n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, 
      n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, 
      n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, 
      n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, 
      n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, 
      n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, 
      n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, 
      n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, 
      n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, 
      n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, 
      n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, 
      n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, 
      n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, 
      n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, 
      n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, 
      n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, 
      n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, 
      n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, 
      n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, 
      n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, 
      n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, 
      n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
      n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, 
      n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, 
      n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, 
      n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, 
      n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, 
      n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, 
      n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, 
      n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, 
      n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, 
      n2193, n2194, n2195, n2196, n2197, n2198, n2199 : std_logic;

begin
   
   U2 : CLKBUF_X3 port map( A => n2195, Z => n73);
   U3 : BUF_X1 port map( A => n67, Z => n1);
   U4 : BUF_X1 port map( A => n64, Z => n6);
   U5 : CLKBUF_X2 port map( A => n2195, Z => n16);
   U6 : BUF_X1 port map( A => n2185, Z => n67);
   U7 : BUF_X1 port map( A => n2185, Z => n65);
   U8 : INV_X2 port map( A => n2112, ZN => n2);
   U9 : BUF_X4 port map( A => n2195, Z => n68);
   U10 : CLKBUF_X3 port map( A => n2195, Z => n71);
   U11 : BUF_X1 port map( A => n101, Z => n15);
   U12 : INV_X1 port map( A => n2199, ZN => n18);
   U13 : NAND3_X2 port map( A1 => n119, A2 => win(0), A3 => n118, ZN => n2112);
   U14 : CLKBUF_X3 port map( A => n2195, Z => n3);
   U15 : NAND3_X2 port map( A1 => n117, A2 => n115, A3 => win(2), ZN => n2199);
   U16 : INV_X2 port map( A => n115, ZN => n4);
   U17 : INV_X2 port map( A => n64, ZN => n5);
   U18 : BUF_X2 port map( A => n64, Z => n47);
   U19 : INV_X2 port map( A => n2112, ZN => n7);
   U20 : INV_X2 port map( A => n64, ZN => n8);
   U21 : BUF_X2 port map( A => n77, Z => n9);
   U22 : INV_X2 port map( A => n2185, ZN => n10);
   U23 : BUF_X2 port map( A => n68, Z => n76);
   U24 : BUF_X2 port map( A => n2112, Z => n21);
   U25 : BUF_X2 port map( A => n78, Z => n11);
   U26 : BUF_X2 port map( A => n2112, Z => n22);
   U27 : BUF_X2 port map( A => n68, Z => n12);
   U28 : BUF_X2 port map( A => n102, Z => n100);
   U29 : NAND2_X2 port map( A1 => n119, A2 => win(1), ZN => n2185);
   U30 : BUF_X2 port map( A => n73, Z => n13);
   U31 : INV_X2 port map( A => n102, ZN => n14);
   U32 : INV_X2 port map( A => n102, ZN => n17);
   U33 : BUF_X16 port map( A => win(4), Z => n116);
   U34 : INV_X2 port map( A => n115, ZN => n19);
   U35 : BUF_X1 port map( A => n67, Z => n46);
   U36 : BUF_X1 port map( A => n2185, Z => n66);
   U37 : BUF_X1 port map( A => n68, Z => n78);
   U38 : INV_X1 port map( A => n64, ZN => n63);
   U39 : BUF_X1 port map( A => n73, Z => n77);
   U40 : INV_X1 port map( A => n115, ZN => n103);
   U41 : INV_X1 port map( A => win(4), ZN => n115);
   U42 : BUF_X1 port map( A => n101, Z => n99);
   U43 : BUF_X1 port map( A => n68, Z => n74);
   U44 : BUF_X1 port map( A => n73, Z => n70);
   U45 : BUF_X1 port map( A => n73, Z => n69);
   U46 : BUF_X1 port map( A => n68, Z => n75);
   U47 : BUF_X1 port map( A => n68, Z => n72);
   U48 : BUF_X1 port map( A => n2185, Z => n64);
   U49 : BUF_X1 port map( A => n2199, Z => n101);
   U50 : BUF_X1 port map( A => n2199, Z => n102);
   U51 : INV_X1 port map( A => n2112, ZN => n23);
   U52 : INV_X1 port map( A => n2112, ZN => n24);
   U53 : INV_X1 port map( A => n21, ZN => n25);
   U54 : INV_X1 port map( A => n2112, ZN => n26);
   U55 : INV_X1 port map( A => n2112, ZN => n27);
   U56 : INV_X1 port map( A => n2112, ZN => n28);
   U57 : INV_X1 port map( A => n2112, ZN => n29);
   U58 : INV_X1 port map( A => n2112, ZN => n30);
   U59 : INV_X1 port map( A => n2112, ZN => n31);
   U60 : INV_X1 port map( A => n2112, ZN => n32);
   U61 : INV_X1 port map( A => n2112, ZN => n33);
   U62 : INV_X1 port map( A => n2112, ZN => n34);
   U63 : INV_X1 port map( A => n2112, ZN => n35);
   U64 : INV_X1 port map( A => n2112, ZN => n36);
   U65 : INV_X1 port map( A => n2112, ZN => n37);
   U66 : INV_X1 port map( A => n2112, ZN => n38);
   U67 : INV_X1 port map( A => n2112, ZN => n39);
   U68 : INV_X1 port map( A => n2112, ZN => n40);
   U69 : INV_X1 port map( A => n2112, ZN => n41);
   U70 : INV_X1 port map( A => n2112, ZN => n42);
   U71 : INV_X1 port map( A => n2112, ZN => n43);
   U72 : INV_X1 port map( A => n2112, ZN => n44);
   U73 : INV_X1 port map( A => n2112, ZN => n45);
   U74 : INV_X1 port map( A => n47, ZN => n48);
   U75 : INV_X1 port map( A => n47, ZN => n49);
   U76 : INV_X1 port map( A => n47, ZN => n50);
   U77 : INV_X1 port map( A => n47, ZN => n51);
   U78 : INV_X1 port map( A => n2185, ZN => n52);
   U79 : INV_X1 port map( A => n2185, ZN => n53);
   U80 : INV_X1 port map( A => n2185, ZN => n54);
   U81 : INV_X1 port map( A => n2185, ZN => n55);
   U82 : INV_X1 port map( A => n2185, ZN => n56);
   U83 : INV_X1 port map( A => n2185, ZN => n57);
   U84 : INV_X1 port map( A => n2185, ZN => n58);
   U85 : INV_X1 port map( A => n2185, ZN => n59);
   U86 : INV_X1 port map( A => n2185, ZN => n60);
   U87 : INV_X1 port map( A => n2185, ZN => n61);
   U88 : INV_X1 port map( A => n2185, ZN => n62);
   U89 : INV_X1 port map( A => n2199, ZN => n79);
   U90 : INV_X1 port map( A => n2199, ZN => n80);
   U91 : INV_X1 port map( A => n2199, ZN => n81);
   U92 : INV_X1 port map( A => n2199, ZN => n82);
   U93 : INV_X1 port map( A => n2199, ZN => n83);
   U94 : INV_X1 port map( A => n2199, ZN => n84);
   U95 : INV_X1 port map( A => n2199, ZN => n85);
   U96 : INV_X1 port map( A => n2199, ZN => n86);
   U97 : INV_X1 port map( A => n2199, ZN => n87);
   U98 : INV_X1 port map( A => n2199, ZN => n88);
   U99 : INV_X1 port map( A => n102, ZN => n89);
   U100 : INV_X1 port map( A => n2199, ZN => n90);
   U101 : INV_X1 port map( A => n102, ZN => n91);
   U102 : INV_X1 port map( A => n2199, ZN => n92);
   U103 : INV_X1 port map( A => n102, ZN => n93);
   U104 : INV_X1 port map( A => n2199, ZN => n94);
   U105 : INV_X1 port map( A => n2199, ZN => n95);
   U106 : INV_X1 port map( A => n2199, ZN => n96);
   U107 : INV_X1 port map( A => n15, ZN => n97);
   U108 : INV_X1 port map( A => n2199, ZN => n98);
   U109 : INV_X1 port map( A => n115, ZN => n104);
   U110 : INV_X1 port map( A => n115, ZN => n105);
   U111 : INV_X1 port map( A => n115, ZN => n106);
   U112 : INV_X1 port map( A => n115, ZN => n107);
   U113 : INV_X1 port map( A => n115, ZN => n108);
   U114 : INV_X1 port map( A => n115, ZN => n109);
   U115 : INV_X1 port map( A => n115, ZN => n110);
   U116 : INV_X1 port map( A => n115, ZN => n111);
   U117 : INV_X1 port map( A => n115, ZN => n112);
   U118 : INV_X1 port map( A => n115, ZN => n113);
   U119 : INV_X1 port map( A => n115, ZN => n114);
   U120 : NOR3_X1 port map( A1 => win(3), A2 => n116, A3 => win(2), ZN => n119)
                           ;
   U121 : INV_X1 port map( A => regs(512), ZN => n1294);
   U122 : INV_X1 port map( A => win(3), ZN => n117);
   U123 : NOR2_X1 port map( A1 => n103, A2 => n117, ZN => n2195);
   U124 : AOI22_X1 port map( A1 => n116, A2 => regs(2048), B1 => n71, B2 => 
                           regs(1536), ZN => n121);
   U125 : INV_X1 port map( A => win(1), ZN => n118);
   U126 : AOI22_X1 port map( A1 => n94, A2 => regs(1024), B1 => n44, B2 => 
                           regs(0), ZN => n120);
   U127 : OAI211_X1 port map( C1 => n47, C2 => n1294, A => n121, B => n120, ZN 
                           => curr_proc_regs(0));
   U128 : INV_X1 port map( A => regs(1124), ZN => n1601);
   U129 : AOI22_X1 port map( A1 => n116, A2 => regs(2148), B1 => n71, B2 => 
                           regs(1636), ZN => n123);
   U130 : AOI22_X1 port map( A1 => n58, A2 => regs(612), B1 => n43, B2 => 
                           regs(100), ZN => n122);
   U131 : OAI211_X1 port map( C1 => n101, C2 => n1601, A => n123, B => n122, ZN
                           => curr_proc_regs(100));
   U132 : INV_X1 port map( A => regs(613), ZN => n1604);
   U133 : AOI22_X1 port map( A1 => n116, A2 => regs(2149), B1 => n71, B2 => 
                           regs(1637), ZN => n125);
   U134 : AOI22_X1 port map( A1 => n91, A2 => regs(1125), B1 => n44, B2 => 
                           regs(101), ZN => n124);
   U135 : OAI211_X1 port map( C1 => n47, C2 => n1604, A => n125, B => n124, ZN 
                           => curr_proc_regs(101));
   U136 : INV_X1 port map( A => regs(614), ZN => n1607);
   U137 : AOI22_X1 port map( A1 => n116, A2 => regs(2150), B1 => n71, B2 => 
                           regs(1638), ZN => n127);
   U138 : AOI22_X1 port map( A1 => n91, A2 => regs(1126), B1 => n43, B2 => 
                           regs(102), ZN => n126);
   U139 : OAI211_X1 port map( C1 => n47, C2 => n1607, A => n127, B => n126, ZN 
                           => curr_proc_regs(102));
   U140 : INV_X1 port map( A => regs(615), ZN => n1610);
   U141 : AOI22_X1 port map( A1 => n116, A2 => regs(2151), B1 => n71, B2 => 
                           regs(1639), ZN => n129);
   U142 : AOI22_X1 port map( A1 => n17, A2 => regs(1127), B1 => n43, B2 => 
                           regs(103), ZN => n128);
   U143 : OAI211_X1 port map( C1 => n47, C2 => n1610, A => n129, B => n128, ZN 
                           => curr_proc_regs(103));
   U144 : INV_X1 port map( A => regs(616), ZN => n1613);
   U145 : AOI22_X1 port map( A1 => n116, A2 => regs(2152), B1 => n71, B2 => 
                           regs(1640), ZN => n131);
   U146 : AOI22_X1 port map( A1 => n17, A2 => regs(1128), B1 => n43, B2 => 
                           regs(104), ZN => n130);
   U147 : OAI211_X1 port map( C1 => n47, C2 => n1613, A => n131, B => n130, ZN 
                           => curr_proc_regs(104));
   U148 : INV_X1 port map( A => regs(617), ZN => n1616);
   U149 : AOI22_X1 port map( A1 => n116, A2 => regs(2153), B1 => n71, B2 => 
                           regs(1641), ZN => n133);
   U150 : AOI22_X1 port map( A1 => n17, A2 => regs(1129), B1 => n43, B2 => 
                           regs(105), ZN => n132);
   U151 : OAI211_X1 port map( C1 => n47, C2 => n1616, A => n133, B => n132, ZN 
                           => curr_proc_regs(105));
   U152 : INV_X1 port map( A => regs(618), ZN => n1619);
   U153 : AOI22_X1 port map( A1 => n116, A2 => regs(2154), B1 => n71, B2 => 
                           regs(1642), ZN => n135);
   U154 : AOI22_X1 port map( A1 => n17, A2 => regs(1130), B1 => n43, B2 => 
                           regs(106), ZN => n134);
   U155 : OAI211_X1 port map( C1 => n47, C2 => n1619, A => n135, B => n134, ZN 
                           => curr_proc_regs(106));
   U156 : INV_X1 port map( A => regs(1131), ZN => n1622);
   U157 : AOI22_X1 port map( A1 => n116, A2 => regs(2155), B1 => n71, B2 => 
                           regs(1643), ZN => n137);
   U158 : AOI22_X1 port map( A1 => n8, A2 => regs(619), B1 => n43, B2 => 
                           regs(107), ZN => n136);
   U159 : OAI211_X1 port map( C1 => n101, C2 => n1622, A => n137, B => n136, ZN
                           => curr_proc_regs(107));
   U160 : INV_X1 port map( A => regs(620), ZN => n1628);
   U161 : AOI22_X1 port map( A1 => n116, A2 => regs(2156), B1 => n71, B2 => 
                           regs(1644), ZN => n139);
   U162 : AOI22_X1 port map( A1 => n81, A2 => regs(1132), B1 => n43, B2 => 
                           regs(108), ZN => n138);
   U163 : OAI211_X1 port map( C1 => n2185, C2 => n1628, A => n139, B => n138, 
                           ZN => curr_proc_regs(108));
   U164 : INV_X1 port map( A => regs(1133), ZN => n1631);
   U165 : AOI22_X1 port map( A1 => n116, A2 => regs(2157), B1 => n71, B2 => 
                           regs(1645), ZN => n141);
   U166 : AOI22_X1 port map( A1 => n49, A2 => regs(621), B1 => n43, B2 => 
                           regs(109), ZN => n140);
   U167 : OAI211_X1 port map( C1 => n101, C2 => n1631, A => n141, B => n140, ZN
                           => curr_proc_regs(109));
   U168 : INV_X1 port map( A => regs(522), ZN => n1323);
   U169 : AOI22_X1 port map( A1 => n116, A2 => regs(2058), B1 => n3, B2 => 
                           regs(1546), ZN => n143);
   U170 : AOI22_X1 port map( A1 => n17, A2 => regs(1034), B1 => n44, B2 => 
                           regs(10), ZN => n142);
   U171 : OAI211_X1 port map( C1 => n47, C2 => n1323, A => n143, B => n142, ZN 
                           => curr_proc_regs(10));
   U172 : INV_X1 port map( A => regs(622), ZN => n1634);
   U173 : AOI22_X1 port map( A1 => n116, A2 => regs(2158), B1 => n3, B2 => 
                           regs(1646), ZN => n145);
   U174 : AOI22_X1 port map( A1 => n17, A2 => regs(1134), B1 => n43, B2 => 
                           regs(110), ZN => n144);
   U175 : OAI211_X1 port map( C1 => n47, C2 => n1634, A => n145, B => n144, ZN 
                           => curr_proc_regs(110));
   U176 : INV_X1 port map( A => regs(623), ZN => n1637);
   U177 : AOI22_X1 port map( A1 => n116, A2 => regs(2159), B1 => n3, B2 => 
                           regs(1647), ZN => n147);
   U178 : AOI22_X1 port map( A1 => n17, A2 => regs(1135), B1 => n43, B2 => 
                           regs(111), ZN => n146);
   U179 : OAI211_X1 port map( C1 => n47, C2 => n1637, A => n147, B => n146, ZN 
                           => curr_proc_regs(111));
   U180 : INV_X1 port map( A => regs(624), ZN => n1640);
   U181 : AOI22_X1 port map( A1 => n116, A2 => regs(2160), B1 => n3, B2 => 
                           regs(1648), ZN => n149);
   U182 : AOI22_X1 port map( A1 => n18, A2 => regs(1136), B1 => n45, B2 => 
                           regs(112), ZN => n148);
   U183 : OAI211_X1 port map( C1 => n47, C2 => n1640, A => n149, B => n148, ZN 
                           => curr_proc_regs(112));
   U184 : INV_X1 port map( A => regs(625), ZN => n1643);
   U185 : AOI22_X1 port map( A1 => n116, A2 => regs(2161), B1 => n71, B2 => 
                           regs(1649), ZN => n151);
   U186 : AOI22_X1 port map( A1 => n17, A2 => regs(1137), B1 => n43, B2 => 
                           regs(113), ZN => n150);
   U187 : OAI211_X1 port map( C1 => n47, C2 => n1643, A => n151, B => n150, ZN 
                           => curr_proc_regs(113));
   U188 : INV_X1 port map( A => regs(626), ZN => n1646);
   U189 : AOI22_X1 port map( A1 => n116, A2 => regs(2162), B1 => n68, B2 => 
                           regs(1650), ZN => n153);
   U190 : AOI22_X1 port map( A1 => n17, A2 => regs(1138), B1 => n45, B2 => 
                           regs(114), ZN => n152);
   U191 : OAI211_X1 port map( C1 => n2185, C2 => n1646, A => n153, B => n152, 
                           ZN => curr_proc_regs(114));
   U192 : INV_X1 port map( A => regs(627), ZN => n1649);
   U193 : AOI22_X1 port map( A1 => n116, A2 => regs(2163), B1 => n73, B2 => 
                           regs(1651), ZN => n155);
   U194 : AOI22_X1 port map( A1 => n17, A2 => regs(1139), B1 => n44, B2 => 
                           regs(115), ZN => n154);
   U195 : OAI211_X1 port map( C1 => n47, C2 => n1649, A => n155, B => n154, ZN 
                           => curr_proc_regs(115));
   U196 : INV_X1 port map( A => regs(628), ZN => n1652);
   U197 : AOI22_X1 port map( A1 => n116, A2 => regs(2164), B1 => n16, B2 => 
                           regs(1652), ZN => n157);
   U198 : AOI22_X1 port map( A1 => n18, A2 => regs(1140), B1 => n44, B2 => 
                           regs(116), ZN => n156);
   U199 : OAI211_X1 port map( C1 => n47, C2 => n1652, A => n157, B => n156, ZN 
                           => curr_proc_regs(116));
   U200 : INV_X1 port map( A => regs(629), ZN => n1655);
   U201 : AOI22_X1 port map( A1 => n116, A2 => regs(2165), B1 => n16, B2 => 
                           regs(1653), ZN => n159);
   U202 : AOI22_X1 port map( A1 => n18, A2 => regs(1141), B1 => n45, B2 => 
                           regs(117), ZN => n158);
   U203 : OAI211_X1 port map( C1 => n47, C2 => n1655, A => n159, B => n158, ZN 
                           => curr_proc_regs(117));
   U204 : INV_X1 port map( A => regs(630), ZN => n1661);
   U205 : AOI22_X1 port map( A1 => n116, A2 => regs(2166), B1 => n9, B2 => 
                           regs(1654), ZN => n161);
   U206 : AOI22_X1 port map( A1 => n18, A2 => regs(1142), B1 => n43, B2 => 
                           regs(118), ZN => n160);
   U207 : OAI211_X1 port map( C1 => n47, C2 => n1661, A => n161, B => n160, ZN 
                           => curr_proc_regs(118));
   U208 : INV_X1 port map( A => regs(1143), ZN => n1664);
   U209 : AOI22_X1 port map( A1 => n116, A2 => regs(2167), B1 => n3, B2 => 
                           regs(1655), ZN => n163);
   U210 : AOI22_X1 port map( A1 => n49, A2 => regs(631), B1 => n45, B2 => 
                           regs(119), ZN => n162);
   U211 : OAI211_X1 port map( C1 => n101, C2 => n1664, A => n163, B => n162, ZN
                           => curr_proc_regs(119));
   U212 : INV_X1 port map( A => regs(523), ZN => n1326);
   U213 : AOI22_X1 port map( A1 => n116, A2 => regs(2059), B1 => n12, B2 => 
                           regs(1547), ZN => n165);
   U214 : AOI22_X1 port map( A1 => n18, A2 => regs(1035), B1 => n44, B2 => 
                           regs(11), ZN => n164);
   U215 : OAI211_X1 port map( C1 => n47, C2 => n1326, A => n165, B => n164, ZN 
                           => curr_proc_regs(11));
   U216 : INV_X1 port map( A => regs(1144), ZN => n1667);
   U217 : AOI22_X1 port map( A1 => n116, A2 => regs(2168), B1 => n12, B2 => 
                           regs(1656), ZN => n167);
   U218 : AOI22_X1 port map( A1 => n55, A2 => regs(632), B1 => n43, B2 => 
                           regs(120), ZN => n166);
   U219 : OAI211_X1 port map( C1 => n101, C2 => n1667, A => n167, B => n166, ZN
                           => curr_proc_regs(120));
   U220 : INV_X1 port map( A => regs(633), ZN => n1670);
   U221 : AOI22_X1 port map( A1 => n116, A2 => regs(2169), B1 => n12, B2 => 
                           regs(1657), ZN => n169);
   U222 : AOI22_X1 port map( A1 => n18, A2 => regs(1145), B1 => n45, B2 => 
                           regs(121), ZN => n168);
   U223 : OAI211_X1 port map( C1 => n47, C2 => n1670, A => n169, B => n168, ZN 
                           => curr_proc_regs(121));
   U224 : INV_X1 port map( A => regs(1146), ZN => n1673);
   U225 : AOI22_X1 port map( A1 => n116, A2 => regs(2170), B1 => n12, B2 => 
                           regs(1658), ZN => n171);
   U226 : AOI22_X1 port map( A1 => n57, A2 => regs(634), B1 => n44, B2 => 
                           regs(122), ZN => n170);
   U227 : OAI211_X1 port map( C1 => n101, C2 => n1673, A => n171, B => n170, ZN
                           => curr_proc_regs(122));
   U228 : INV_X1 port map( A => regs(635), ZN => n1676);
   U229 : AOI22_X1 port map( A1 => n116, A2 => regs(2171), B1 => n12, B2 => 
                           regs(1659), ZN => n173);
   U230 : AOI22_X1 port map( A1 => n17, A2 => regs(1147), B1 => n45, B2 => 
                           regs(123), ZN => n172);
   U231 : OAI211_X1 port map( C1 => n47, C2 => n1676, A => n173, B => n172, ZN 
                           => curr_proc_regs(123));
   U232 : INV_X1 port map( A => regs(1148), ZN => n1679);
   U233 : AOI22_X1 port map( A1 => n116, A2 => regs(2172), B1 => n12, B2 => 
                           regs(1660), ZN => n175);
   U234 : AOI22_X1 port map( A1 => n59, A2 => regs(636), B1 => n43, B2 => 
                           regs(124), ZN => n174);
   U235 : OAI211_X1 port map( C1 => n2199, C2 => n1679, A => n175, B => n174, 
                           ZN => curr_proc_regs(124));
   U236 : INV_X1 port map( A => regs(1149), ZN => n1682);
   U237 : AOI22_X1 port map( A1 => n116, A2 => regs(2173), B1 => n12, B2 => 
                           regs(1661), ZN => n177);
   U238 : AOI22_X1 port map( A1 => n61, A2 => regs(637), B1 => n45, B2 => 
                           regs(125), ZN => n176);
   U239 : OAI211_X1 port map( C1 => n101, C2 => n1682, A => n177, B => n176, ZN
                           => curr_proc_regs(125));
   U240 : INV_X1 port map( A => regs(1150), ZN => n1685);
   U241 : AOI22_X1 port map( A1 => n116, A2 => regs(2174), B1 => n12, B2 => 
                           regs(1662), ZN => n179);
   U242 : AOI22_X1 port map( A1 => n49, A2 => regs(638), B1 => n44, B2 => 
                           regs(126), ZN => n178);
   U243 : OAI211_X1 port map( C1 => n101, C2 => n1685, A => n179, B => n178, ZN
                           => curr_proc_regs(126));
   U244 : INV_X1 port map( A => regs(1151), ZN => n1688);
   U245 : AOI22_X1 port map( A1 => n116, A2 => regs(2175), B1 => n12, B2 => 
                           regs(1663), ZN => n181);
   U246 : AOI22_X1 port map( A1 => n50, A2 => regs(639), B1 => n44, B2 => 
                           regs(127), ZN => n180);
   U247 : OAI211_X1 port map( C1 => n101, C2 => n1688, A => n181, B => n180, ZN
                           => curr_proc_regs(127));
   U248 : INV_X1 port map( A => regs(1152), ZN => n1694);
   U249 : AOI22_X1 port map( A1 => n116, A2 => regs(2176), B1 => n12, B2 => 
                           regs(1664), ZN => n183);
   U250 : AOI22_X1 port map( A1 => n51, A2 => regs(640), B1 => n43, B2 => 
                           regs(128), ZN => n182);
   U251 : OAI211_X1 port map( C1 => n101, C2 => n1694, A => n183, B => n182, ZN
                           => curr_proc_regs(128));
   U252 : INV_X1 port map( A => regs(641), ZN => n1697);
   U253 : AOI22_X1 port map( A1 => n116, A2 => regs(2177), B1 => n12, B2 => 
                           regs(1665), ZN => n185);
   U254 : AOI22_X1 port map( A1 => n18, A2 => regs(1153), B1 => n45, B2 => 
                           regs(129), ZN => n184);
   U255 : OAI211_X1 port map( C1 => n47, C2 => n1697, A => n185, B => n184, ZN 
                           => curr_proc_regs(129));
   U256 : INV_X1 port map( A => regs(524), ZN => n1329);
   U257 : AOI22_X1 port map( A1 => n116, A2 => regs(2060), B1 => n13, B2 => 
                           regs(1548), ZN => n187);
   U258 : AOI22_X1 port map( A1 => n17, A2 => regs(1036), B1 => n44, B2 => 
                           regs(12), ZN => n186);
   U259 : OAI211_X1 port map( C1 => n47, C2 => n1329, A => n187, B => n186, ZN 
                           => curr_proc_regs(12));
   U260 : INV_X1 port map( A => regs(1154), ZN => n1700);
   U261 : AOI22_X1 port map( A1 => n116, A2 => regs(2178), B1 => n13, B2 => 
                           regs(1666), ZN => n189);
   U262 : AOI22_X1 port map( A1 => n48, A2 => regs(642), B1 => n44, B2 => 
                           regs(130), ZN => n188);
   U263 : OAI211_X1 port map( C1 => n101, C2 => n1700, A => n189, B => n188, ZN
                           => curr_proc_regs(130));
   U264 : INV_X1 port map( A => regs(1155), ZN => n1703);
   U265 : AOI22_X1 port map( A1 => n116, A2 => regs(2179), B1 => n13, B2 => 
                           regs(1667), ZN => n191);
   U266 : AOI22_X1 port map( A1 => n53, A2 => regs(643), B1 => n44, B2 => 
                           regs(131), ZN => n190);
   U267 : OAI211_X1 port map( C1 => n101, C2 => n1703, A => n191, B => n190, ZN
                           => curr_proc_regs(131));
   U268 : INV_X1 port map( A => regs(1156), ZN => n1706);
   U269 : AOI22_X1 port map( A1 => n116, A2 => regs(2180), B1 => n13, B2 => 
                           regs(1668), ZN => n193);
   U270 : AOI22_X1 port map( A1 => n52, A2 => regs(644), B1 => n44, B2 => 
                           regs(132), ZN => n192);
   U271 : OAI211_X1 port map( C1 => n101, C2 => n1706, A => n193, B => n192, ZN
                           => curr_proc_regs(132));
   U272 : INV_X1 port map( A => regs(1157), ZN => n1709);
   U273 : AOI22_X1 port map( A1 => n116, A2 => regs(2181), B1 => n13, B2 => 
                           regs(1669), ZN => n195);
   U274 : AOI22_X1 port map( A1 => n54, A2 => regs(645), B1 => n45, B2 => 
                           regs(133), ZN => n194);
   U275 : OAI211_X1 port map( C1 => n2199, C2 => n1709, A => n195, B => n194, 
                           ZN => curr_proc_regs(133));
   U276 : INV_X1 port map( A => regs(1158), ZN => n1712);
   U277 : AOI22_X1 port map( A1 => n116, A2 => regs(2182), B1 => n13, B2 => 
                           regs(1670), ZN => n197);
   U278 : AOI22_X1 port map( A1 => n49, A2 => regs(646), B1 => n44, B2 => 
                           regs(134), ZN => n196);
   U279 : OAI211_X1 port map( C1 => n101, C2 => n1712, A => n197, B => n196, ZN
                           => curr_proc_regs(134));
   U280 : INV_X1 port map( A => regs(647), ZN => n1715);
   U281 : AOI22_X1 port map( A1 => n116, A2 => regs(2183), B1 => n13, B2 => 
                           regs(1671), ZN => n199);
   U282 : AOI22_X1 port map( A1 => n17, A2 => regs(1159), B1 => n43, B2 => 
                           regs(135), ZN => n198);
   U283 : OAI211_X1 port map( C1 => n2185, C2 => n1715, A => n199, B => n198, 
                           ZN => curr_proc_regs(135));
   U284 : INV_X1 port map( A => regs(648), ZN => n1718);
   U285 : AOI22_X1 port map( A1 => n116, A2 => regs(2184), B1 => n13, B2 => 
                           regs(1672), ZN => n201);
   U286 : AOI22_X1 port map( A1 => n17, A2 => regs(1160), B1 => n45, B2 => 
                           regs(136), ZN => n200);
   U287 : OAI211_X1 port map( C1 => n47, C2 => n1718, A => n201, B => n200, ZN 
                           => curr_proc_regs(136));
   U288 : INV_X1 port map( A => regs(1161), ZN => n1721);
   U289 : AOI22_X1 port map( A1 => n116, A2 => regs(2185), B1 => n13, B2 => 
                           regs(1673), ZN => n203);
   U290 : AOI22_X1 port map( A1 => n49, A2 => regs(649), B1 => n44, B2 => 
                           regs(137), ZN => n202);
   U291 : OAI211_X1 port map( C1 => n2199, C2 => n1721, A => n203, B => n202, 
                           ZN => curr_proc_regs(137));
   U292 : INV_X1 port map( A => regs(650), ZN => n1727);
   U293 : AOI22_X1 port map( A1 => n116, A2 => regs(2186), B1 => n13, B2 => 
                           regs(1674), ZN => n205);
   U294 : AOI22_X1 port map( A1 => n17, A2 => regs(1162), B1 => n43, B2 => 
                           regs(138), ZN => n204);
   U295 : OAI211_X1 port map( C1 => n47, C2 => n1727, A => n205, B => n204, ZN 
                           => curr_proc_regs(138));
   U296 : INV_X1 port map( A => regs(1163), ZN => n1730);
   U297 : AOI22_X1 port map( A1 => n116, A2 => regs(2187), B1 => n13, B2 => 
                           regs(1675), ZN => n207);
   U298 : AOI22_X1 port map( A1 => n49, A2 => regs(651), B1 => n45, B2 => 
                           regs(139), ZN => n206);
   U299 : OAI211_X1 port map( C1 => n101, C2 => n1730, A => n207, B => n206, ZN
                           => curr_proc_regs(139));
   U300 : INV_X1 port map( A => regs(525), ZN => n1332);
   U301 : AOI22_X1 port map( A1 => n116, A2 => regs(2061), B1 => n71, B2 => 
                           regs(1549), ZN => n209);
   U302 : AOI22_X1 port map( A1 => n17, A2 => regs(1037), B1 => n45, B2 => 
                           regs(13), ZN => n208);
   U303 : OAI211_X1 port map( C1 => n47, C2 => n1332, A => n209, B => n208, ZN 
                           => curr_proc_regs(13));
   U304 : INV_X1 port map( A => regs(652), ZN => n1733);
   U305 : AOI22_X1 port map( A1 => n116, A2 => regs(2188), B1 => n12, B2 => 
                           regs(1676), ZN => n211);
   U306 : AOI22_X1 port map( A1 => n17, A2 => regs(1164), B1 => n45, B2 => 
                           regs(140), ZN => n210);
   U307 : OAI211_X1 port map( C1 => n47, C2 => n1733, A => n211, B => n210, ZN 
                           => curr_proc_regs(140));
   U308 : INV_X1 port map( A => regs(1165), ZN => n1736);
   U309 : AOI22_X1 port map( A1 => n116, A2 => regs(2189), B1 => n13, B2 => 
                           regs(1677), ZN => n213);
   U310 : AOI22_X1 port map( A1 => n49, A2 => regs(653), B1 => n45, B2 => 
                           regs(141), ZN => n212);
   U311 : OAI211_X1 port map( C1 => n2199, C2 => n1736, A => n213, B => n212, 
                           ZN => curr_proc_regs(141));
   U312 : INV_X1 port map( A => regs(654), ZN => n1739);
   U313 : AOI22_X1 port map( A1 => n116, A2 => regs(2190), B1 => n12, B2 => 
                           regs(1678), ZN => n215);
   U314 : AOI22_X1 port map( A1 => n17, A2 => regs(1166), B1 => n45, B2 => 
                           regs(142), ZN => n214);
   U315 : OAI211_X1 port map( C1 => n47, C2 => n1739, A => n215, B => n214, ZN 
                           => curr_proc_regs(142));
   U316 : INV_X1 port map( A => regs(1167), ZN => n1742);
   U317 : AOI22_X1 port map( A1 => n116, A2 => regs(2191), B1 => n71, B2 => 
                           regs(1679), ZN => n217);
   U318 : AOI22_X1 port map( A1 => n48, A2 => regs(655), B1 => n44, B2 => 
                           regs(143), ZN => n216);
   U319 : OAI211_X1 port map( C1 => n101, C2 => n1742, A => n217, B => n216, ZN
                           => curr_proc_regs(143));
   U320 : INV_X1 port map( A => regs(1168), ZN => n1745);
   U321 : AOI22_X1 port map( A1 => n116, A2 => regs(2192), B1 => n3, B2 => 
                           regs(1680), ZN => n219);
   U322 : AOI22_X1 port map( A1 => n48, A2 => regs(656), B1 => n44, B2 => 
                           regs(144), ZN => n218);
   U323 : OAI211_X1 port map( C1 => n102, C2 => n1745, A => n219, B => n218, ZN
                           => curr_proc_regs(144));
   U324 : INV_X1 port map( A => regs(657), ZN => n1748);
   U325 : AOI22_X1 port map( A1 => n116, A2 => regs(2193), B1 => n3, B2 => 
                           regs(1681), ZN => n221);
   U326 : AOI22_X1 port map( A1 => n95, A2 => regs(1169), B1 => n44, B2 => 
                           regs(145), ZN => n220);
   U327 : OAI211_X1 port map( C1 => n47, C2 => n1748, A => n221, B => n220, ZN 
                           => curr_proc_regs(145));
   U328 : INV_X1 port map( A => regs(1170), ZN => n1751);
   U329 : AOI22_X1 port map( A1 => n116, A2 => regs(2194), B1 => n12, B2 => 
                           regs(1682), ZN => n223);
   U330 : AOI22_X1 port map( A1 => n48, A2 => regs(658), B1 => n44, B2 => 
                           regs(146), ZN => n222);
   U331 : OAI211_X1 port map( C1 => n102, C2 => n1751, A => n223, B => n222, ZN
                           => curr_proc_regs(146));
   U332 : INV_X1 port map( A => regs(1171), ZN => n1754);
   U333 : AOI22_X1 port map( A1 => n116, A2 => regs(2195), B1 => n71, B2 => 
                           regs(1683), ZN => n225);
   U334 : AOI22_X1 port map( A1 => n48, A2 => regs(659), B1 => n44, B2 => 
                           regs(147), ZN => n224);
   U335 : OAI211_X1 port map( C1 => n99, C2 => n1754, A => n225, B => n224, ZN 
                           => curr_proc_regs(147));
   U336 : INV_X1 port map( A => regs(660), ZN => n1760);
   U337 : AOI22_X1 port map( A1 => n116, A2 => regs(2196), B1 => n12, B2 => 
                           regs(1684), ZN => n227);
   U338 : AOI22_X1 port map( A1 => n95, A2 => regs(1172), B1 => n44, B2 => 
                           regs(148), ZN => n226);
   U339 : OAI211_X1 port map( C1 => n47, C2 => n1760, A => n227, B => n226, ZN 
                           => curr_proc_regs(148));
   U340 : INV_X1 port map( A => regs(1173), ZN => n1763);
   U341 : AOI22_X1 port map( A1 => n116, A2 => regs(2197), B1 => n13, B2 => 
                           regs(1685), ZN => n229);
   U342 : AOI22_X1 port map( A1 => n48, A2 => regs(661), B1 => n44, B2 => 
                           regs(149), ZN => n228);
   U343 : OAI211_X1 port map( C1 => n102, C2 => n1763, A => n229, B => n228, ZN
                           => curr_proc_regs(149));
   U344 : INV_X1 port map( A => regs(1038), ZN => n1335);
   U345 : AOI22_X1 port map( A1 => n116, A2 => regs(2062), B1 => n12, B2 => 
                           regs(1550), ZN => n231);
   U346 : AOI22_X1 port map( A1 => n48, A2 => regs(526), B1 => n39, B2 => 
                           regs(14), ZN => n230);
   U347 : OAI211_X1 port map( C1 => n15, C2 => n1335, A => n231, B => n230, ZN 
                           => curr_proc_regs(14));
   U348 : INV_X1 port map( A => regs(1174), ZN => n1766);
   U349 : AOI22_X1 port map( A1 => n116, A2 => regs(2198), B1 => n69, B2 => 
                           regs(1686), ZN => n233);
   U350 : AOI22_X1 port map( A1 => n48, A2 => regs(662), B1 => n39, B2 => 
                           regs(150), ZN => n232);
   U351 : OAI211_X1 port map( C1 => n99, C2 => n1766, A => n233, B => n232, ZN 
                           => curr_proc_regs(150));
   U352 : INV_X1 port map( A => regs(1175), ZN => n1769);
   U353 : AOI22_X1 port map( A1 => n116, A2 => regs(2199), B1 => n71, B2 => 
                           regs(1687), ZN => n235);
   U354 : AOI22_X1 port map( A1 => n57, A2 => regs(663), B1 => n24, B2 => 
                           regs(151), ZN => n234);
   U355 : OAI211_X1 port map( C1 => n102, C2 => n1769, A => n235, B => n234, ZN
                           => curr_proc_regs(151));
   U356 : INV_X1 port map( A => regs(664), ZN => n1772);
   U357 : AOI22_X1 port map( A1 => n116, A2 => regs(2200), B1 => n71, B2 => 
                           regs(1688), ZN => n237);
   U358 : AOI22_X1 port map( A1 => n95, A2 => regs(1176), B1 => n23, B2 => 
                           regs(152), ZN => n236);
   U359 : OAI211_X1 port map( C1 => n47, C2 => n1772, A => n237, B => n236, ZN 
                           => curr_proc_regs(152));
   U360 : INV_X1 port map( A => regs(665), ZN => n1775);
   U361 : AOI22_X1 port map( A1 => n116, A2 => regs(2201), B1 => n68, B2 => 
                           regs(1689), ZN => n239);
   U362 : AOI22_X1 port map( A1 => n95, A2 => regs(1177), B1 => n45, B2 => 
                           regs(153), ZN => n238);
   U363 : OAI211_X1 port map( C1 => n47, C2 => n1775, A => n239, B => n238, ZN 
                           => curr_proc_regs(153));
   U364 : INV_X1 port map( A => regs(666), ZN => n1778);
   U365 : AOI22_X1 port map( A1 => n116, A2 => regs(2202), B1 => n12, B2 => 
                           regs(1690), ZN => n241);
   U366 : AOI22_X1 port map( A1 => n95, A2 => regs(1178), B1 => n45, B2 => 
                           regs(154), ZN => n240);
   U367 : OAI211_X1 port map( C1 => n47, C2 => n1778, A => n241, B => n240, ZN 
                           => curr_proc_regs(154));
   U368 : INV_X1 port map( A => regs(667), ZN => n1781);
   U369 : AOI22_X1 port map( A1 => n116, A2 => regs(2203), B1 => n13, B2 => 
                           regs(1691), ZN => n243);
   U370 : AOI22_X1 port map( A1 => n95, A2 => regs(1179), B1 => n45, B2 => 
                           regs(155), ZN => n242);
   U371 : OAI211_X1 port map( C1 => n47, C2 => n1781, A => n243, B => n242, ZN 
                           => curr_proc_regs(155));
   U372 : INV_X1 port map( A => regs(668), ZN => n1784);
   U373 : AOI22_X1 port map( A1 => n116, A2 => regs(2204), B1 => n12, B2 => 
                           regs(1692), ZN => n245);
   U374 : AOI22_X1 port map( A1 => n95, A2 => regs(1180), B1 => n45, B2 => 
                           regs(156), ZN => n244);
   U375 : OAI211_X1 port map( C1 => n1, C2 => n1784, A => n245, B => n244, ZN 
                           => curr_proc_regs(156));
   U376 : INV_X1 port map( A => regs(669), ZN => n1787);
   U377 : AOI22_X1 port map( A1 => n116, A2 => regs(2205), B1 => n69, B2 => 
                           regs(1693), ZN => n247);
   U378 : AOI22_X1 port map( A1 => n95, A2 => regs(1181), B1 => n45, B2 => 
                           regs(157), ZN => n246);
   U379 : OAI211_X1 port map( C1 => n1, C2 => n1787, A => n247, B => n246, ZN 
                           => curr_proc_regs(157));
   U380 : INV_X1 port map( A => regs(1182), ZN => n1793);
   U381 : AOI22_X1 port map( A1 => n116, A2 => regs(2206), B1 => n71, B2 => 
                           regs(1694), ZN => n249);
   U382 : AOI22_X1 port map( A1 => n59, A2 => regs(670), B1 => n45, B2 => 
                           regs(158), ZN => n248);
   U383 : OAI211_X1 port map( C1 => n2199, C2 => n1793, A => n249, B => n248, 
                           ZN => curr_proc_regs(158));
   U384 : INV_X1 port map( A => regs(1183), ZN => n1796);
   U385 : AOI22_X1 port map( A1 => n116, A2 => regs(2207), B1 => n71, B2 => 
                           regs(1695), ZN => n251);
   U386 : AOI22_X1 port map( A1 => n61, A2 => regs(671), B1 => n45, B2 => 
                           regs(159), ZN => n250);
   U387 : OAI211_X1 port map( C1 => n2199, C2 => n1796, A => n251, B => n250, 
                           ZN => curr_proc_regs(159));
   U388 : INV_X1 port map( A => regs(1039), ZN => n1338);
   U389 : AOI22_X1 port map( A1 => n116, A2 => regs(2063), B1 => n12, B2 => 
                           regs(1551), ZN => n253);
   U390 : AOI22_X1 port map( A1 => n56, A2 => regs(527), B1 => n24, B2 => 
                           regs(15), ZN => n252);
   U391 : OAI211_X1 port map( C1 => n2199, C2 => n1338, A => n253, B => n252, 
                           ZN => curr_proc_regs(15));
   U392 : INV_X1 port map( A => regs(1184), ZN => n1799);
   U393 : AOI22_X1 port map( A1 => n116, A2 => regs(2208), B1 => n13, B2 => 
                           regs(1696), ZN => n255);
   U394 : AOI22_X1 port map( A1 => n51, A2 => regs(672), B1 => n42, B2 => 
                           regs(160), ZN => n254);
   U395 : OAI211_X1 port map( C1 => n2199, C2 => n1799, A => n255, B => n254, 
                           ZN => curr_proc_regs(160));
   U396 : INV_X1 port map( A => regs(673), ZN => n1802);
   U397 : AOI22_X1 port map( A1 => n116, A2 => regs(2209), B1 => n12, B2 => 
                           regs(1697), ZN => n257);
   U398 : AOI22_X1 port map( A1 => n95, A2 => regs(1185), B1 => n39, B2 => 
                           regs(161), ZN => n256);
   U399 : OAI211_X1 port map( C1 => n1, C2 => n1802, A => n257, B => n256, ZN 
                           => curr_proc_regs(161));
   U400 : INV_X1 port map( A => regs(1186), ZN => n1805);
   U401 : AOI22_X1 port map( A1 => n116, A2 => regs(2210), B1 => n69, B2 => 
                           regs(1698), ZN => n259);
   U402 : AOI22_X1 port map( A1 => n50, A2 => regs(674), B1 => n24, B2 => 
                           regs(162), ZN => n258);
   U403 : OAI211_X1 port map( C1 => n2199, C2 => n1805, A => n259, B => n258, 
                           ZN => curr_proc_regs(162));
   U404 : INV_X1 port map( A => regs(1187), ZN => n1808);
   U405 : AOI22_X1 port map( A1 => n116, A2 => regs(2211), B1 => n71, B2 => 
                           regs(1699), ZN => n261);
   U406 : AOI22_X1 port map( A1 => n49, A2 => regs(675), B1 => n23, B2 => 
                           regs(163), ZN => n260);
   U407 : OAI211_X1 port map( C1 => n2199, C2 => n1808, A => n261, B => n260, 
                           ZN => curr_proc_regs(163));
   U408 : INV_X1 port map( A => regs(676), ZN => n1811);
   U409 : AOI22_X1 port map( A1 => n4, A2 => regs(2212), B1 => n71, B2 => 
                           regs(1700), ZN => n263);
   U410 : AOI22_X1 port map( A1 => n89, A2 => regs(1188), B1 => n24, B2 => 
                           regs(164), ZN => n262);
   U411 : OAI211_X1 port map( C1 => n1, C2 => n1811, A => n263, B => n262, ZN 
                           => curr_proc_regs(164));
   U412 : INV_X1 port map( A => regs(1189), ZN => n1814);
   U413 : AOI22_X1 port map( A1 => n19, A2 => regs(2213), B1 => n12, B2 => 
                           regs(1701), ZN => n265);
   U414 : AOI22_X1 port map( A1 => n53, A2 => regs(677), B1 => n42, B2 => 
                           regs(165), ZN => n264);
   U415 : OAI211_X1 port map( C1 => n2199, C2 => n1814, A => n265, B => n264, 
                           ZN => curr_proc_regs(165));
   U416 : INV_X1 port map( A => regs(678), ZN => n1817);
   U417 : AOI22_X1 port map( A1 => n19, A2 => regs(2214), B1 => n13, B2 => 
                           regs(1702), ZN => n267);
   U418 : AOI22_X1 port map( A1 => n91, A2 => regs(1190), B1 => n36, B2 => 
                           regs(166), ZN => n266);
   U419 : OAI211_X1 port map( C1 => n1, C2 => n1817, A => n267, B => n266, ZN 
                           => curr_proc_regs(166));
   U420 : INV_X1 port map( A => regs(679), ZN => n1820);
   U421 : AOI22_X1 port map( A1 => n19, A2 => regs(2215), B1 => n12, B2 => 
                           regs(1703), ZN => n269);
   U422 : AOI22_X1 port map( A1 => n17, A2 => regs(1191), B1 => n38, B2 => 
                           regs(167), ZN => n268);
   U423 : OAI211_X1 port map( C1 => n1, C2 => n1820, A => n269, B => n268, ZN 
                           => curr_proc_regs(167));
   U424 : INV_X1 port map( A => regs(680), ZN => n1826);
   U425 : AOI22_X1 port map( A1 => n19, A2 => regs(2216), B1 => n69, B2 => 
                           regs(1704), ZN => n271);
   U426 : AOI22_X1 port map( A1 => n93, A2 => regs(1192), B1 => n42, B2 => 
                           regs(168), ZN => n270);
   U427 : OAI211_X1 port map( C1 => n1, C2 => n1826, A => n271, B => n270, ZN 
                           => curr_proc_regs(168));
   U428 : INV_X1 port map( A => regs(1193), ZN => n1829);
   U429 : AOI22_X1 port map( A1 => n103, A2 => regs(2217), B1 => n71, B2 => 
                           regs(1705), ZN => n273);
   U430 : AOI22_X1 port map( A1 => n53, A2 => regs(681), B1 => n42, B2 => 
                           regs(169), ZN => n272);
   U431 : OAI211_X1 port map( C1 => n102, C2 => n1829, A => n273, B => n272, ZN
                           => curr_proc_regs(169));
   U432 : INV_X1 port map( A => regs(1040), ZN => n1341);
   U433 : AOI22_X1 port map( A1 => n103, A2 => regs(2064), B1 => n12, B2 => 
                           regs(1552), ZN => n275);
   U434 : AOI22_X1 port map( A1 => n53, A2 => regs(528), B1 => n26, B2 => 
                           regs(16), ZN => n274);
   U435 : OAI211_X1 port map( C1 => n99, C2 => n1341, A => n275, B => n274, ZN 
                           => curr_proc_regs(16));
   U436 : INV_X1 port map( A => regs(1194), ZN => n1832);
   U437 : AOI22_X1 port map( A1 => n19, A2 => regs(2218), B1 => n12, B2 => 
                           regs(1706), ZN => n277);
   U438 : AOI22_X1 port map( A1 => n53, A2 => regs(682), B1 => n26, B2 => 
                           regs(170), ZN => n276);
   U439 : OAI211_X1 port map( C1 => n99, C2 => n1832, A => n277, B => n276, ZN 
                           => curr_proc_regs(170));
   U440 : INV_X1 port map( A => regs(1195), ZN => n1835);
   U441 : AOI22_X1 port map( A1 => n103, A2 => regs(2219), B1 => n12, B2 => 
                           regs(1707), ZN => n279);
   U442 : AOI22_X1 port map( A1 => n53, A2 => regs(683), B1 => n28, B2 => 
                           regs(171), ZN => n278);
   U443 : OAI211_X1 port map( C1 => n99, C2 => n1835, A => n279, B => n278, ZN 
                           => curr_proc_regs(171));
   U444 : INV_X1 port map( A => regs(1196), ZN => n1838);
   U445 : AOI22_X1 port map( A1 => n4, A2 => regs(2220), B1 => n12, B2 => 
                           regs(1708), ZN => n281);
   U446 : AOI22_X1 port map( A1 => n53, A2 => regs(684), B1 => n27, B2 => 
                           regs(172), ZN => n280);
   U447 : OAI211_X1 port map( C1 => n102, C2 => n1838, A => n281, B => n280, ZN
                           => curr_proc_regs(172));
   U448 : INV_X1 port map( A => regs(1197), ZN => n1841);
   U449 : AOI22_X1 port map( A1 => n19, A2 => regs(2221), B1 => n12, B2 => 
                           regs(1709), ZN => n283);
   U450 : AOI22_X1 port map( A1 => n53, A2 => regs(685), B1 => n31, B2 => 
                           regs(173), ZN => n282);
   U451 : OAI211_X1 port map( C1 => n99, C2 => n1841, A => n283, B => n282, ZN 
                           => curr_proc_regs(173));
   U452 : INV_X1 port map( A => regs(686), ZN => n1844);
   U453 : AOI22_X1 port map( A1 => n4, A2 => regs(2222), B1 => n12, B2 => 
                           regs(1710), ZN => n285);
   U454 : AOI22_X1 port map( A1 => n17, A2 => regs(1198), B1 => n29, B2 => 
                           regs(174), ZN => n284);
   U455 : OAI211_X1 port map( C1 => n47, C2 => n1844, A => n285, B => n284, ZN 
                           => curr_proc_regs(174));
   U456 : INV_X1 port map( A => regs(687), ZN => n1847);
   U457 : AOI22_X1 port map( A1 => n19, A2 => regs(2223), B1 => n12, B2 => 
                           regs(1711), ZN => n287);
   U458 : AOI22_X1 port map( A1 => n89, A2 => regs(1199), B1 => n38, B2 => 
                           regs(175), ZN => n286);
   U459 : OAI211_X1 port map( C1 => n47, C2 => n1847, A => n287, B => n286, ZN 
                           => curr_proc_regs(175));
   U460 : INV_X1 port map( A => regs(1200), ZN => n1850);
   U461 : AOI22_X1 port map( A1 => n4, A2 => regs(2224), B1 => n12, B2 => 
                           regs(1712), ZN => n289);
   U462 : AOI22_X1 port map( A1 => n53, A2 => regs(688), B1 => n41, B2 => 
                           regs(176), ZN => n288);
   U463 : OAI211_X1 port map( C1 => n99, C2 => n1850, A => n289, B => n288, ZN 
                           => curr_proc_regs(176));
   U464 : INV_X1 port map( A => regs(689), ZN => n1853);
   U465 : AOI22_X1 port map( A1 => n4, A2 => regs(2225), B1 => n12, B2 => 
                           regs(1713), ZN => n291);
   U466 : AOI22_X1 port map( A1 => n89, A2 => regs(1201), B1 => n2, B2 => 
                           regs(177), ZN => n290);
   U467 : OAI211_X1 port map( C1 => n47, C2 => n1853, A => n291, B => n290, ZN 
                           => curr_proc_regs(177));
   U468 : INV_X1 port map( A => regs(1202), ZN => n1859);
   U469 : AOI22_X1 port map( A1 => n103, A2 => regs(2226), B1 => n12, B2 => 
                           regs(1714), ZN => n293);
   U470 : AOI22_X1 port map( A1 => n52, A2 => regs(690), B1 => n2, B2 => 
                           regs(178), ZN => n292);
   U471 : OAI211_X1 port map( C1 => n2199, C2 => n1859, A => n293, B => n292, 
                           ZN => curr_proc_regs(178));
   U472 : INV_X1 port map( A => regs(691), ZN => n1862);
   U473 : AOI22_X1 port map( A1 => n4, A2 => regs(2227), B1 => n12, B2 => 
                           regs(1715), ZN => n295);
   U474 : AOI22_X1 port map( A1 => n17, A2 => regs(1203), B1 => n7, B2 => 
                           regs(179), ZN => n294);
   U475 : OAI211_X1 port map( C1 => n47, C2 => n1862, A => n295, B => n294, ZN 
                           => curr_proc_regs(179));
   U476 : INV_X1 port map( A => regs(1041), ZN => n1344);
   U477 : AOI22_X1 port map( A1 => n19, A2 => regs(2065), B1 => n16, B2 => 
                           regs(1553), ZN => n297);
   U478 : AOI22_X1 port map( A1 => n52, A2 => regs(529), B1 => n29, B2 => 
                           regs(17), ZN => n296);
   U479 : OAI211_X1 port map( C1 => n100, C2 => n1344, A => n297, B => n296, ZN
                           => curr_proc_regs(17));
   U480 : INV_X1 port map( A => regs(692), ZN => n1865);
   U481 : AOI22_X1 port map( A1 => n19, A2 => regs(2228), B1 => n16, B2 => 
                           regs(1716), ZN => n299);
   U482 : AOI22_X1 port map( A1 => n91, A2 => regs(1204), B1 => n38, B2 => 
                           regs(180), ZN => n298);
   U483 : OAI211_X1 port map( C1 => n47, C2 => n1865, A => n299, B => n298, ZN 
                           => curr_proc_regs(180));
   U484 : INV_X1 port map( A => regs(693), ZN => n1868);
   U485 : AOI22_X1 port map( A1 => n4, A2 => regs(2229), B1 => n12, B2 => 
                           regs(1717), ZN => n301);
   U486 : AOI22_X1 port map( A1 => n92, A2 => regs(1205), B1 => n41, B2 => 
                           regs(181), ZN => n300);
   U487 : OAI211_X1 port map( C1 => n47, C2 => n1868, A => n301, B => n300, ZN 
                           => curr_proc_regs(181));
   U488 : INV_X1 port map( A => regs(694), ZN => n1871);
   U489 : AOI22_X1 port map( A1 => n103, A2 => regs(2230), B1 => n3, B2 => 
                           regs(1718), ZN => n303);
   U490 : AOI22_X1 port map( A1 => n17, A2 => regs(1206), B1 => n2, B2 => 
                           regs(182), ZN => n302);
   U491 : OAI211_X1 port map( C1 => n47, C2 => n1871, A => n303, B => n302, ZN 
                           => curr_proc_regs(182));
   U492 : INV_X1 port map( A => regs(695), ZN => n1874);
   U493 : AOI22_X1 port map( A1 => n19, A2 => regs(2231), B1 => n3, B2 => 
                           regs(1719), ZN => n305);
   U494 : AOI22_X1 port map( A1 => n17, A2 => regs(1207), B1 => n33, B2 => 
                           regs(183), ZN => n304);
   U495 : OAI211_X1 port map( C1 => n2185, C2 => n1874, A => n305, B => n304, 
                           ZN => curr_proc_regs(183));
   U496 : INV_X1 port map( A => regs(696), ZN => n1877);
   U497 : AOI22_X1 port map( A1 => n19, A2 => regs(2232), B1 => n71, B2 => 
                           regs(1720), ZN => n307);
   U498 : AOI22_X1 port map( A1 => n18, A2 => regs(1208), B1 => n30, B2 => 
                           regs(184), ZN => n306);
   U499 : OAI211_X1 port map( C1 => n47, C2 => n1877, A => n307, B => n306, ZN 
                           => curr_proc_regs(184));
   U500 : INV_X1 port map( A => regs(697), ZN => n1880);
   U501 : AOI22_X1 port map( A1 => n19, A2 => regs(2233), B1 => n68, B2 => 
                           regs(1721), ZN => n309);
   U502 : AOI22_X1 port map( A1 => n94, A2 => regs(1209), B1 => n32, B2 => 
                           regs(185), ZN => n308);
   U503 : OAI211_X1 port map( C1 => n2185, C2 => n1880, A => n309, B => n308, 
                           ZN => curr_proc_regs(185));
   U504 : INV_X1 port map( A => regs(1210), ZN => n1883);
   U505 : AOI22_X1 port map( A1 => n116, A2 => regs(2234), B1 => n73, B2 => 
                           regs(1722), ZN => n311);
   U506 : AOI22_X1 port map( A1 => n52, A2 => regs(698), B1 => n37, B2 => 
                           regs(186), ZN => n310);
   U507 : OAI211_X1 port map( C1 => n2199, C2 => n1883, A => n311, B => n310, 
                           ZN => curr_proc_regs(186));
   U508 : INV_X1 port map( A => regs(1211), ZN => n1886);
   U509 : AOI22_X1 port map( A1 => n4, A2 => regs(2235), B1 => n16, B2 => 
                           regs(1723), ZN => n313);
   U510 : AOI22_X1 port map( A1 => n59, A2 => regs(699), B1 => n40, B2 => 
                           regs(187), ZN => n312);
   U511 : OAI211_X1 port map( C1 => n100, C2 => n1886, A => n313, B => n312, ZN
                           => curr_proc_regs(187));
   U512 : INV_X1 port map( A => regs(700), ZN => n1895);
   U513 : AOI22_X1 port map( A1 => n19, A2 => regs(2236), B1 => n16, B2 => 
                           regs(1724), ZN => n315);
   U514 : AOI22_X1 port map( A1 => n95, A2 => regs(1212), B1 => n28, B2 => 
                           regs(188), ZN => n314);
   U515 : OAI211_X1 port map( C1 => n47, C2 => n1895, A => n315, B => n314, ZN 
                           => curr_proc_regs(188));
   U516 : INV_X1 port map( A => regs(701), ZN => n1898);
   U517 : AOI22_X1 port map( A1 => n103, A2 => regs(2237), B1 => n11, B2 => 
                           regs(1725), ZN => n317);
   U518 : AOI22_X1 port map( A1 => n91, A2 => regs(1213), B1 => n27, B2 => 
                           regs(189), ZN => n316);
   U519 : OAI211_X1 port map( C1 => n2185, C2 => n1898, A => n317, B => n316, 
                           ZN => curr_proc_regs(189));
   U520 : INV_X1 port map( A => regs(1042), ZN => n1349);
   U521 : AOI22_X1 port map( A1 => n4, A2 => regs(2066), B1 => n12, B2 => 
                           regs(1554), ZN => n319);
   U522 : AOI22_X1 port map( A1 => n57, A2 => regs(530), B1 => n40, B2 => 
                           regs(18), ZN => n318);
   U523 : OAI211_X1 port map( C1 => n2199, C2 => n1349, A => n319, B => n318, 
                           ZN => curr_proc_regs(18));
   U524 : INV_X1 port map( A => regs(702), ZN => n1901);
   U525 : AOI22_X1 port map( A1 => n19, A2 => regs(2238), B1 => n13, B2 => 
                           regs(1726), ZN => n321);
   U526 : AOI22_X1 port map( A1 => n89, A2 => regs(1214), B1 => n28, B2 => 
                           regs(190), ZN => n320);
   U527 : OAI211_X1 port map( C1 => n47, C2 => n1901, A => n321, B => n320, ZN 
                           => curr_proc_regs(190));
   U528 : INV_X1 port map( A => regs(703), ZN => n1904);
   U529 : AOI22_X1 port map( A1 => n19, A2 => regs(2239), B1 => n3, B2 => 
                           regs(1727), ZN => n323);
   U530 : AOI22_X1 port map( A1 => n93, A2 => regs(1215), B1 => n27, B2 => 
                           regs(191), ZN => n322);
   U531 : OAI211_X1 port map( C1 => n2185, C2 => n1904, A => n323, B => n322, 
                           ZN => curr_proc_regs(191));
   U532 : INV_X1 port map( A => regs(1216), ZN => n1907);
   U533 : AOI22_X1 port map( A1 => n19, A2 => regs(2240), B1 => n71, B2 => 
                           regs(1728), ZN => n325);
   U534 : AOI22_X1 port map( A1 => n55, A2 => regs(704), B1 => n26, B2 => 
                           regs(192), ZN => n324);
   U535 : OAI211_X1 port map( C1 => n100, C2 => n1907, A => n325, B => n324, ZN
                           => curr_proc_regs(192));
   U536 : INV_X1 port map( A => regs(1217), ZN => n1910);
   U537 : AOI22_X1 port map( A1 => n19, A2 => regs(2241), B1 => n12, B2 => 
                           regs(1729), ZN => n327);
   U538 : AOI22_X1 port map( A1 => n54, A2 => regs(705), B1 => n2, B2 => 
                           regs(193), ZN => n326);
   U539 : OAI211_X1 port map( C1 => n100, C2 => n1910, A => n327, B => n326, ZN
                           => curr_proc_regs(193));
   U540 : INV_X1 port map( A => regs(1218), ZN => n1913);
   U541 : AOI22_X1 port map( A1 => n116, A2 => regs(2242), B1 => n13, B2 => 
                           regs(1730), ZN => n329);
   U542 : AOI22_X1 port map( A1 => n52, A2 => regs(706), B1 => n29, B2 => 
                           regs(194), ZN => n328);
   U543 : OAI211_X1 port map( C1 => n15, C2 => n1913, A => n329, B => n328, ZN 
                           => curr_proc_regs(194));
   U544 : INV_X1 port map( A => regs(1219), ZN => n1916);
   U545 : AOI22_X1 port map( A1 => n19, A2 => regs(2243), B1 => n69, B2 => 
                           regs(1731), ZN => n331);
   U546 : AOI22_X1 port map( A1 => n53, A2 => regs(707), B1 => n31, B2 => 
                           regs(195), ZN => n330);
   U547 : OAI211_X1 port map( C1 => n15, C2 => n1916, A => n331, B => n330, ZN 
                           => curr_proc_regs(195));
   U548 : INV_X1 port map( A => regs(708), ZN => n1919);
   U549 : AOI22_X1 port map( A1 => n103, A2 => regs(2244), B1 => n71, B2 => 
                           regs(1732), ZN => n333);
   U550 : AOI22_X1 port map( A1 => n17, A2 => regs(1220), B1 => n31, B2 => 
                           regs(196), ZN => n332);
   U551 : OAI211_X1 port map( C1 => n65, C2 => n1919, A => n333, B => n332, ZN 
                           => curr_proc_regs(196));
   U552 : INV_X1 port map( A => regs(1221), ZN => n1922);
   U553 : AOI22_X1 port map( A1 => n4, A2 => regs(2245), B1 => n69, B2 => 
                           regs(1733), ZN => n335);
   U554 : AOI22_X1 port map( A1 => n54, A2 => regs(709), B1 => n29, B2 => 
                           regs(197), ZN => n334);
   U555 : OAI211_X1 port map( C1 => n15, C2 => n1922, A => n335, B => n334, ZN 
                           => curr_proc_regs(197));
   U556 : INV_X1 port map( A => regs(1222), ZN => n1928);
   U557 : AOI22_X1 port map( A1 => n19, A2 => regs(2246), B1 => n71, B2 => 
                           regs(1734), ZN => n337);
   U558 : AOI22_X1 port map( A1 => n48, A2 => regs(710), B1 => n2, B2 => 
                           regs(198), ZN => n336);
   U559 : OAI211_X1 port map( C1 => n15, C2 => n1928, A => n337, B => n336, ZN 
                           => curr_proc_regs(198));
   U560 : INV_X1 port map( A => regs(711), ZN => n1931);
   U561 : AOI22_X1 port map( A1 => n19, A2 => regs(2247), B1 => n12, B2 => 
                           regs(1735), ZN => n339);
   U562 : AOI22_X1 port map( A1 => n93, A2 => regs(1223), B1 => n31, B2 => 
                           regs(199), ZN => n338);
   U563 : OAI211_X1 port map( C1 => n66, C2 => n1931, A => n339, B => n338, ZN 
                           => curr_proc_regs(199));
   U564 : INV_X1 port map( A => regs(531), ZN => n1352);
   U565 : AOI22_X1 port map( A1 => n103, A2 => regs(2067), B1 => n71, B2 => 
                           regs(1555), ZN => n341);
   U566 : AOI22_X1 port map( A1 => n89, A2 => regs(1043), B1 => n42, B2 => 
                           regs(19), ZN => n340);
   U567 : OAI211_X1 port map( C1 => n2185, C2 => n1352, A => n341, B => n340, 
                           ZN => curr_proc_regs(19));
   U568 : INV_X1 port map( A => regs(513), ZN => n1297);
   U569 : AOI22_X1 port map( A1 => win(4), A2 => regs(2049), B1 => n12, B2 => 
                           regs(1537), ZN => n343);
   U570 : AOI22_X1 port map( A1 => n91, A2 => regs(1025), B1 => n42, B2 => 
                           regs(1), ZN => n342);
   U571 : OAI211_X1 port map( C1 => n2185, C2 => n1297, A => n343, B => n342, 
                           ZN => curr_proc_regs(1));
   U572 : INV_X1 port map( A => regs(1224), ZN => n1934);
   U573 : AOI22_X1 port map( A1 => n103, A2 => regs(2248), B1 => n12, B2 => 
                           regs(1736), ZN => n345);
   U574 : AOI22_X1 port map( A1 => n52, A2 => regs(712), B1 => n42, B2 => 
                           regs(200), ZN => n344);
   U575 : OAI211_X1 port map( C1 => n15, C2 => n1934, A => n345, B => n344, ZN 
                           => curr_proc_regs(200));
   U576 : INV_X1 port map( A => regs(1225), ZN => n1937);
   U577 : AOI22_X1 port map( A1 => n4, A2 => regs(2249), B1 => n69, B2 => 
                           regs(1737), ZN => n347);
   U578 : AOI22_X1 port map( A1 => n48, A2 => regs(713), B1 => n42, B2 => 
                           regs(201), ZN => n346);
   U579 : OAI211_X1 port map( C1 => n15, C2 => n1937, A => n347, B => n346, ZN 
                           => curr_proc_regs(201));
   U580 : INV_X1 port map( A => regs(714), ZN => n1940);
   U581 : AOI22_X1 port map( A1 => n19, A2 => regs(2250), B1 => n71, B2 => 
                           regs(1738), ZN => n349);
   U582 : AOI22_X1 port map( A1 => n93, A2 => regs(1226), B1 => n26, B2 => 
                           regs(202), ZN => n348);
   U583 : OAI211_X1 port map( C1 => n67, C2 => n1940, A => n349, B => n348, ZN 
                           => curr_proc_regs(202));
   U584 : INV_X1 port map( A => regs(715), ZN => n1943);
   U585 : AOI22_X1 port map( A1 => n103, A2 => regs(2251), B1 => n71, B2 => 
                           regs(1739), ZN => n351);
   U586 : AOI22_X1 port map( A1 => n17, A2 => regs(1227), B1 => n33, B2 => 
                           regs(203), ZN => n350);
   U587 : OAI211_X1 port map( C1 => n65, C2 => n1943, A => n351, B => n350, ZN 
                           => curr_proc_regs(203));
   U588 : INV_X1 port map( A => regs(1228), ZN => n1946);
   U589 : AOI22_X1 port map( A1 => n4, A2 => regs(2252), B1 => n16, B2 => 
                           regs(1740), ZN => n353);
   U590 : AOI22_X1 port map( A1 => n50, A2 => regs(716), B1 => n27, B2 => 
                           regs(204), ZN => n352);
   U591 : OAI211_X1 port map( C1 => n15, C2 => n1946, A => n353, B => n352, ZN 
                           => curr_proc_regs(204));
   U592 : INV_X1 port map( A => regs(1229), ZN => n1949);
   U593 : AOI22_X1 port map( A1 => n19, A2 => regs(2253), B1 => n69, B2 => 
                           regs(1741), ZN => n355);
   U594 : AOI22_X1 port map( A1 => n52, A2 => regs(717), B1 => n33, B2 => 
                           regs(205), ZN => n354);
   U595 : OAI211_X1 port map( C1 => n100, C2 => n1949, A => n355, B => n354, ZN
                           => curr_proc_regs(205));
   U596 : INV_X1 port map( A => regs(718), ZN => n1952);
   U597 : AOI22_X1 port map( A1 => n19, A2 => regs(2254), B1 => n16, B2 => 
                           regs(1742), ZN => n357);
   U598 : AOI22_X1 port map( A1 => n17, A2 => regs(1230), B1 => n30, B2 => 
                           regs(206), ZN => n356);
   U599 : OAI211_X1 port map( C1 => n2185, C2 => n1952, A => n357, B => n356, 
                           ZN => curr_proc_regs(206));
   U600 : INV_X1 port map( A => regs(719), ZN => n1955);
   U601 : AOI22_X1 port map( A1 => n116, A2 => regs(2255), B1 => n75, B2 => 
                           regs(1743), ZN => n359);
   U602 : AOI22_X1 port map( A1 => n96, A2 => regs(1231), B1 => n32, B2 => 
                           regs(207), ZN => n358);
   U603 : OAI211_X1 port map( C1 => n1, C2 => n1955, A => n359, B => n358, ZN 
                           => curr_proc_regs(207));
   U604 : INV_X1 port map( A => regs(1232), ZN => n1961);
   U605 : AOI22_X1 port map( A1 => n103, A2 => regs(2256), B1 => n12, B2 => 
                           regs(1744), ZN => n361);
   U606 : AOI22_X1 port map( A1 => n52, A2 => regs(720), B1 => n37, B2 => 
                           regs(208), ZN => n360);
   U607 : OAI211_X1 port map( C1 => n2199, C2 => n1961, A => n361, B => n360, 
                           ZN => curr_proc_regs(208));
   U608 : INV_X1 port map( A => regs(1233), ZN => n1964);
   U609 : AOI22_X1 port map( A1 => n4, A2 => regs(2257), B1 => n71, B2 => 
                           regs(1745), ZN => n363);
   U610 : AOI22_X1 port map( A1 => n52, A2 => regs(721), B1 => n29, B2 => 
                           regs(209), ZN => n362);
   U611 : OAI211_X1 port map( C1 => n100, C2 => n1964, A => n363, B => n362, ZN
                           => curr_proc_regs(209));
   U612 : INV_X1 port map( A => regs(1044), ZN => n1355);
   U613 : AOI22_X1 port map( A1 => n19, A2 => regs(2068), B1 => n13, B2 => 
                           regs(1556), ZN => n365);
   U614 : AOI22_X1 port map( A1 => n52, A2 => regs(532), B1 => n29, B2 => 
                           regs(20), ZN => n364);
   U615 : OAI211_X1 port map( C1 => n2199, C2 => n1355, A => n365, B => n364, 
                           ZN => curr_proc_regs(20));
   U616 : INV_X1 port map( A => regs(1234), ZN => n1967);
   U617 : AOI22_X1 port map( A1 => n19, A2 => regs(2258), B1 => n12, B2 => 
                           regs(1746), ZN => n367);
   U618 : AOI22_X1 port map( A1 => n52, A2 => regs(722), B1 => n38, B2 => 
                           regs(210), ZN => n366);
   U619 : OAI211_X1 port map( C1 => n100, C2 => n1967, A => n367, B => n366, ZN
                           => curr_proc_regs(210));
   U620 : INV_X1 port map( A => regs(1235), ZN => n1970);
   U621 : AOI22_X1 port map( A1 => n116, A2 => regs(2259), B1 => n69, B2 => 
                           regs(1747), ZN => n369);
   U622 : AOI22_X1 port map( A1 => n52, A2 => regs(723), B1 => n31, B2 => 
                           regs(211), ZN => n368);
   U623 : OAI211_X1 port map( C1 => n2199, C2 => n1970, A => n369, B => n368, 
                           ZN => curr_proc_regs(211));
   U624 : INV_X1 port map( A => regs(724), ZN => n1973);
   U625 : AOI22_X1 port map( A1 => n103, A2 => regs(2260), B1 => n71, B2 => 
                           regs(1748), ZN => n371);
   U626 : AOI22_X1 port map( A1 => n89, A2 => regs(1236), B1 => n42, B2 => 
                           regs(212), ZN => n370);
   U627 : OAI211_X1 port map( C1 => n65, C2 => n1973, A => n371, B => n370, ZN 
                           => curr_proc_regs(212));
   U628 : INV_X1 port map( A => regs(1237), ZN => n1976);
   U629 : AOI22_X1 port map( A1 => n116, A2 => regs(2261), B1 => n71, B2 => 
                           regs(1749), ZN => n373);
   U630 : AOI22_X1 port map( A1 => n52, A2 => regs(725), B1 => n42, B2 => 
                           regs(213), ZN => n372);
   U631 : OAI211_X1 port map( C1 => n100, C2 => n1976, A => n373, B => n372, ZN
                           => curr_proc_regs(213));
   U632 : INV_X1 port map( A => regs(1238), ZN => n1979);
   U633 : AOI22_X1 port map( A1 => n116, A2 => regs(2262), B1 => n73, B2 => 
                           regs(1750), ZN => n375);
   U634 : AOI22_X1 port map( A1 => n52, A2 => regs(726), B1 => n42, B2 => 
                           regs(214), ZN => n374);
   U635 : OAI211_X1 port map( C1 => n100, C2 => n1979, A => n375, B => n374, ZN
                           => curr_proc_regs(214));
   U636 : INV_X1 port map( A => regs(1239), ZN => n1982);
   U637 : AOI22_X1 port map( A1 => n116, A2 => regs(2263), B1 => n71, B2 => 
                           regs(1751), ZN => n377);
   U638 : AOI22_X1 port map( A1 => n53, A2 => regs(727), B1 => n42, B2 => 
                           regs(215), ZN => n376);
   U639 : OAI211_X1 port map( C1 => n100, C2 => n1982, A => n377, B => n376, ZN
                           => curr_proc_regs(215));
   U640 : INV_X1 port map( A => regs(1240), ZN => n1985);
   U641 : AOI22_X1 port map( A1 => n116, A2 => regs(2264), B1 => n68, B2 => 
                           regs(1752), ZN => n379);
   U642 : AOI22_X1 port map( A1 => n61, A2 => regs(728), B1 => n42, B2 => 
                           regs(216), ZN => n378);
   U643 : OAI211_X1 port map( C1 => n100, C2 => n1985, A => n379, B => n378, ZN
                           => curr_proc_regs(216));
   U644 : INV_X1 port map( A => regs(1241), ZN => n1988);
   U645 : AOI22_X1 port map( A1 => n116, A2 => regs(2265), B1 => n73, B2 => 
                           regs(1753), ZN => n381);
   U646 : AOI22_X1 port map( A1 => n53, A2 => regs(729), B1 => n42, B2 => 
                           regs(217), ZN => n380);
   U647 : OAI211_X1 port map( C1 => n100, C2 => n1988, A => n381, B => n380, ZN
                           => curr_proc_regs(217));
   U648 : INV_X1 port map( A => regs(1242), ZN => n1994);
   U649 : AOI22_X1 port map( A1 => n116, A2 => regs(2266), B1 => n71, B2 => 
                           regs(1754), ZN => n383);
   U650 : AOI22_X1 port map( A1 => n59, A2 => regs(730), B1 => n42, B2 => 
                           regs(218), ZN => n382);
   U651 : OAI211_X1 port map( C1 => n101, C2 => n1994, A => n383, B => n382, ZN
                           => curr_proc_regs(218));
   U652 : INV_X1 port map( A => regs(731), ZN => n1997);
   U653 : AOI22_X1 port map( A1 => n116, A2 => regs(2267), B1 => n69, B2 => 
                           regs(1755), ZN => n385);
   U654 : AOI22_X1 port map( A1 => n93, A2 => regs(1243), B1 => n26, B2 => 
                           regs(219), ZN => n384);
   U655 : OAI211_X1 port map( C1 => n2185, C2 => n1997, A => n385, B => n384, 
                           ZN => curr_proc_regs(219));
   U656 : INV_X1 port map( A => regs(533), ZN => n1358);
   U657 : AOI22_X1 port map( A1 => n116, A2 => regs(2069), B1 => n69, B2 => 
                           regs(1557), ZN => n387);
   U658 : AOI22_X1 port map( A1 => n17, A2 => regs(1045), B1 => n33, B2 => 
                           regs(21), ZN => n386);
   U659 : OAI211_X1 port map( C1 => n2185, C2 => n1358, A => n387, B => n386, 
                           ZN => curr_proc_regs(21));
   U660 : INV_X1 port map( A => regs(732), ZN => n2000);
   U661 : AOI22_X1 port map( A1 => n116, A2 => regs(2268), B1 => n69, B2 => 
                           regs(1756), ZN => n389);
   U662 : AOI22_X1 port map( A1 => n87, A2 => regs(1244), B1 => n30, B2 => 
                           regs(220), ZN => n388);
   U663 : OAI211_X1 port map( C1 => n2185, C2 => n2000, A => n389, B => n388, 
                           ZN => curr_proc_regs(220));
   U664 : INV_X1 port map( A => regs(1245), ZN => n2003);
   U665 : AOI22_X1 port map( A1 => n116, A2 => regs(2269), B1 => n69, B2 => 
                           regs(1757), ZN => n391);
   U666 : AOI22_X1 port map( A1 => n57, A2 => regs(733), B1 => n33, B2 => 
                           regs(221), ZN => n390);
   U667 : OAI211_X1 port map( C1 => n100, C2 => n2003, A => n391, B => n390, ZN
                           => curr_proc_regs(221));
   U668 : INV_X1 port map( A => regs(734), ZN => n2006);
   U669 : AOI22_X1 port map( A1 => n116, A2 => regs(2270), B1 => n69, B2 => 
                           regs(1758), ZN => n393);
   U670 : AOI22_X1 port map( A1 => n88, A2 => regs(1246), B1 => n7, B2 => 
                           regs(222), ZN => n392);
   U671 : OAI211_X1 port map( C1 => n2185, C2 => n2006, A => n393, B => n392, 
                           ZN => curr_proc_regs(222));
   U672 : INV_X1 port map( A => regs(735), ZN => n2009);
   U673 : AOI22_X1 port map( A1 => win(4), A2 => regs(2271), B1 => n69, B2 => 
                           regs(1759), ZN => n395);
   U674 : AOI22_X1 port map( A1 => n89, A2 => regs(1247), B1 => n7, B2 => 
                           regs(223), ZN => n394);
   U675 : OAI211_X1 port map( C1 => n2185, C2 => n2009, A => n395, B => n394, 
                           ZN => curr_proc_regs(223));
   U676 : INV_X1 port map( A => regs(1248), ZN => n2012);
   U677 : AOI22_X1 port map( A1 => n113, A2 => regs(2272), B1 => n69, B2 => 
                           regs(1760), ZN => n397);
   U678 : AOI22_X1 port map( A1 => n55, A2 => regs(736), B1 => n25, B2 => 
                           regs(224), ZN => n396);
   U679 : OAI211_X1 port map( C1 => n100, C2 => n2012, A => n397, B => n396, ZN
                           => curr_proc_regs(224));
   U680 : INV_X1 port map( A => regs(1249), ZN => n2015);
   U681 : AOI22_X1 port map( A1 => n114, A2 => regs(2273), B1 => n69, B2 => 
                           regs(1761), ZN => n399);
   U682 : AOI22_X1 port map( A1 => n54, A2 => regs(737), B1 => n29, B2 => 
                           regs(225), ZN => n398);
   U683 : OAI211_X1 port map( C1 => n99, C2 => n2015, A => n399, B => n398, ZN 
                           => curr_proc_regs(225));
   U684 : INV_X1 port map( A => regs(738), ZN => n2018);
   U685 : AOI22_X1 port map( A1 => n114, A2 => regs(2274), B1 => n69, B2 => 
                           regs(1762), ZN => n401);
   U686 : AOI22_X1 port map( A1 => n17, A2 => regs(1250), B1 => n29, B2 => 
                           regs(226), ZN => n400);
   U687 : OAI211_X1 port map( C1 => n1, C2 => n2018, A => n401, B => n400, ZN 
                           => curr_proc_regs(226));
   U688 : INV_X1 port map( A => regs(1251), ZN => n2021);
   U689 : AOI22_X1 port map( A1 => n113, A2 => regs(2275), B1 => n69, B2 => 
                           regs(1763), ZN => n403);
   U690 : AOI22_X1 port map( A1 => n52, A2 => regs(739), B1 => n7, B2 => 
                           regs(227), ZN => n402);
   U691 : OAI211_X1 port map( C1 => n99, C2 => n2021, A => n403, B => n402, ZN 
                           => curr_proc_regs(227));
   U692 : INV_X1 port map( A => regs(1252), ZN => n2027);
   U693 : AOI22_X1 port map( A1 => win(4), A2 => regs(2276), B1 => n69, B2 => 
                           regs(1764), ZN => n405);
   U694 : AOI22_X1 port map( A1 => n53, A2 => regs(740), B1 => n38, B2 => 
                           regs(228), ZN => n404);
   U695 : OAI211_X1 port map( C1 => n99, C2 => n2027, A => n405, B => n404, ZN 
                           => curr_proc_regs(228));
   U696 : INV_X1 port map( A => regs(1253), ZN => n2030);
   U697 : AOI22_X1 port map( A1 => n113, A2 => regs(2277), B1 => n13, B2 => 
                           regs(1765), ZN => n407);
   U698 : AOI22_X1 port map( A1 => n56, A2 => regs(741), B1 => n32, B2 => 
                           regs(229), ZN => n406);
   U699 : OAI211_X1 port map( C1 => n99, C2 => n2030, A => n407, B => n406, ZN 
                           => curr_proc_regs(229));
   U700 : INV_X1 port map( A => regs(534), ZN => n1361);
   U701 : AOI22_X1 port map( A1 => n114, A2 => regs(2070), B1 => n12, B2 => 
                           regs(1558), ZN => n409);
   U702 : AOI22_X1 port map( A1 => n94, A2 => regs(1046), B1 => n37, B2 => 
                           regs(22), ZN => n408);
   U703 : OAI211_X1 port map( C1 => n64, C2 => n1361, A => n409, B => n408, ZN 
                           => curr_proc_regs(22));
   U704 : INV_X1 port map( A => regs(1254), ZN => n2033);
   U705 : AOI22_X1 port map( A1 => win(4), A2 => regs(2278), B1 => n13, B2 => 
                           regs(1766), ZN => n411);
   U706 : AOI22_X1 port map( A1 => n48, A2 => regs(742), B1 => n40, B2 => 
                           regs(230), ZN => n410);
   U707 : OAI211_X1 port map( C1 => n99, C2 => n2033, A => n411, B => n410, ZN 
                           => curr_proc_regs(230));
   U708 : INV_X1 port map( A => regs(1255), ZN => n2036);
   U709 : AOI22_X1 port map( A1 => n114, A2 => regs(2279), B1 => n12, B2 => 
                           regs(1767), ZN => n413);
   U710 : AOI22_X1 port map( A1 => n57, A2 => regs(743), B1 => n28, B2 => 
                           regs(231), ZN => n412);
   U711 : OAI211_X1 port map( C1 => n99, C2 => n2036, A => n413, B => n412, ZN 
                           => curr_proc_regs(231));
   U712 : INV_X1 port map( A => regs(1256), ZN => n2039);
   U713 : AOI22_X1 port map( A1 => win(4), A2 => regs(2280), B1 => n69, B2 => 
                           regs(1768), ZN => n415);
   U714 : AOI22_X1 port map( A1 => n53, A2 => regs(744), B1 => n33, B2 => 
                           regs(232), ZN => n414);
   U715 : OAI211_X1 port map( C1 => n99, C2 => n2039, A => n415, B => n414, ZN 
                           => curr_proc_regs(232));
   U716 : INV_X1 port map( A => regs(1257), ZN => n2042);
   U717 : AOI22_X1 port map( A1 => n113, A2 => regs(2281), B1 => n71, B2 => 
                           regs(1769), ZN => n417);
   U718 : AOI22_X1 port map( A1 => n52, A2 => regs(745), B1 => n30, B2 => 
                           regs(233), ZN => n416);
   U719 : OAI211_X1 port map( C1 => n101, C2 => n2042, A => n417, B => n416, ZN
                           => curr_proc_regs(233));
   U720 : INV_X1 port map( A => regs(1258), ZN => n2045);
   U721 : AOI22_X1 port map( A1 => win(4), A2 => regs(2282), B1 => n69, B2 => 
                           regs(1770), ZN => n419);
   U722 : AOI22_X1 port map( A1 => n56, A2 => regs(746), B1 => n32, B2 => 
                           regs(234), ZN => n418);
   U723 : OAI211_X1 port map( C1 => n102, C2 => n2045, A => n419, B => n418, ZN
                           => curr_proc_regs(234));
   U724 : INV_X1 port map( A => regs(747), ZN => n2048);
   U725 : AOI22_X1 port map( A1 => n113, A2 => regs(2283), B1 => n3, B2 => 
                           regs(1771), ZN => n421);
   U726 : AOI22_X1 port map( A1 => n94, A2 => regs(1259), B1 => n37, B2 => 
                           regs(235), ZN => n420);
   U727 : OAI211_X1 port map( C1 => n65, C2 => n2048, A => n421, B => n420, ZN 
                           => curr_proc_regs(235));
   U728 : INV_X1 port map( A => regs(748), ZN => n2051);
   U729 : AOI22_X1 port map( A1 => n114, A2 => regs(2284), B1 => n12, B2 => 
                           regs(1772), ZN => n423);
   U730 : AOI22_X1 port map( A1 => n94, A2 => regs(1260), B1 => n40, B2 => 
                           regs(236), ZN => n422);
   U731 : OAI211_X1 port map( C1 => n1, C2 => n2051, A => n423, B => n422, ZN 
                           => curr_proc_regs(236));
   U732 : INV_X1 port map( A => regs(1261), ZN => n2054);
   U733 : AOI22_X1 port map( A1 => n114, A2 => regs(2285), B1 => n71, B2 => 
                           regs(1773), ZN => n425);
   U734 : AOI22_X1 port map( A1 => n61, A2 => regs(749), B1 => n28, B2 => 
                           regs(237), ZN => n424);
   U735 : OAI211_X1 port map( C1 => n101, C2 => n2054, A => n425, B => n424, ZN
                           => curr_proc_regs(237));
   U736 : INV_X1 port map( A => regs(750), ZN => n2060);
   U737 : AOI22_X1 port map( A1 => win(4), A2 => regs(2286), B1 => n3, B2 => 
                           regs(1774), ZN => n427);
   U738 : AOI22_X1 port map( A1 => n94, A2 => regs(1262), B1 => n27, B2 => 
                           regs(238), ZN => n426);
   U739 : OAI211_X1 port map( C1 => n67, C2 => n2060, A => n427, B => n426, ZN 
                           => curr_proc_regs(238));
   U740 : INV_X1 port map( A => regs(751), ZN => n2063);
   U741 : AOI22_X1 port map( A1 => n113, A2 => regs(2287), B1 => n71, B2 => 
                           regs(1775), ZN => n429);
   U742 : AOI22_X1 port map( A1 => n94, A2 => regs(1263), B1 => n40, B2 => 
                           regs(239), ZN => n428);
   U743 : OAI211_X1 port map( C1 => n65, C2 => n2063, A => n429, B => n428, ZN 
                           => curr_proc_regs(239));
   U744 : INV_X1 port map( A => regs(1047), ZN => n1364);
   U745 : AOI22_X1 port map( A1 => n114, A2 => regs(2071), B1 => n71, B2 => 
                           regs(1559), ZN => n431);
   U746 : AOI22_X1 port map( A1 => n59, A2 => regs(535), B1 => n33, B2 => 
                           regs(23), ZN => n430);
   U747 : OAI211_X1 port map( C1 => n100, C2 => n1364, A => n431, B => n430, ZN
                           => curr_proc_regs(23));
   U748 : INV_X1 port map( A => regs(1264), ZN => n2066);
   U749 : AOI22_X1 port map( A1 => win(4), A2 => regs(2288), B1 => n71, B2 => 
                           regs(1776), ZN => n433);
   U750 : AOI22_X1 port map( A1 => n57, A2 => regs(752), B1 => n30, B2 => 
                           regs(240), ZN => n432);
   U751 : OAI211_X1 port map( C1 => n100, C2 => n2066, A => n433, B => n432, ZN
                           => curr_proc_regs(240));
   U752 : INV_X1 port map( A => regs(753), ZN => n2069);
   U753 : AOI22_X1 port map( A1 => win(4), A2 => regs(2289), B1 => n71, B2 => 
                           regs(1777), ZN => n435);
   U754 : AOI22_X1 port map( A1 => n94, A2 => regs(1265), B1 => n32, B2 => 
                           regs(241), ZN => n434);
   U755 : OAI211_X1 port map( C1 => n46, C2 => n2069, A => n435, B => n434, ZN 
                           => curr_proc_regs(241));
   U756 : INV_X1 port map( A => regs(1266), ZN => n2072);
   U757 : AOI22_X1 port map( A1 => n113, A2 => regs(2290), B1 => n71, B2 => 
                           regs(1778), ZN => n437);
   U758 : AOI22_X1 port map( A1 => n55, A2 => regs(754), B1 => n27, B2 => 
                           regs(242), ZN => n436);
   U759 : OAI211_X1 port map( C1 => n102, C2 => n2072, A => n437, B => n436, ZN
                           => curr_proc_regs(242));
   U760 : INV_X1 port map( A => regs(755), ZN => n2075);
   U761 : AOI22_X1 port map( A1 => n113, A2 => regs(2291), B1 => n71, B2 => 
                           regs(1779), ZN => n439);
   U762 : AOI22_X1 port map( A1 => n94, A2 => regs(1267), B1 => n37, B2 => 
                           regs(243), ZN => n438);
   U763 : OAI211_X1 port map( C1 => n2185, C2 => n2075, A => n439, B => n438, 
                           ZN => curr_proc_regs(243));
   U764 : INV_X1 port map( A => regs(756), ZN => n2078);
   U765 : AOI22_X1 port map( A1 => n114, A2 => regs(2292), B1 => n71, B2 => 
                           regs(1780), ZN => n441);
   U766 : AOI22_X1 port map( A1 => n93, A2 => regs(1268), B1 => n32, B2 => 
                           regs(244), ZN => n440);
   U767 : OAI211_X1 port map( C1 => n2185, C2 => n2078, A => n441, B => n440, 
                           ZN => curr_proc_regs(244));
   U768 : INV_X1 port map( A => regs(1269), ZN => n2081);
   U769 : AOI22_X1 port map( A1 => win(4), A2 => regs(2293), B1 => n71, B2 => 
                           regs(1781), ZN => n443);
   U770 : AOI22_X1 port map( A1 => n54, A2 => regs(757), B1 => n37, B2 => 
                           regs(245), ZN => n442);
   U771 : OAI211_X1 port map( C1 => n100, C2 => n2081, A => n443, B => n442, ZN
                           => curr_proc_regs(245));
   U772 : INV_X1 port map( A => regs(1270), ZN => n2084);
   U773 : AOI22_X1 port map( A1 => n113, A2 => regs(2294), B1 => n71, B2 => 
                           regs(1782), ZN => n445);
   U774 : AOI22_X1 port map( A1 => n52, A2 => regs(758), B1 => n27, B2 => 
                           regs(246), ZN => n444);
   U775 : OAI211_X1 port map( C1 => n2199, C2 => n2084, A => n445, B => n444, 
                           ZN => curr_proc_regs(246));
   U776 : INV_X1 port map( A => regs(759), ZN => n2087);
   U777 : AOI22_X1 port map( A1 => n114, A2 => regs(2295), B1 => n71, B2 => 
                           regs(1783), ZN => n447);
   U778 : AOI22_X1 port map( A1 => n93, A2 => regs(1271), B1 => n33, B2 => 
                           regs(247), ZN => n446);
   U779 : OAI211_X1 port map( C1 => n6, C2 => n2087, A => n447, B => n446, ZN 
                           => curr_proc_regs(247));
   U780 : INV_X1 port map( A => regs(760), ZN => n2093);
   U781 : AOI22_X1 port map( A1 => win(4), A2 => regs(2296), B1 => n71, B2 => 
                           regs(1784), ZN => n449);
   U782 : AOI22_X1 port map( A1 => n93, A2 => regs(1272), B1 => n30, B2 => 
                           regs(248), ZN => n448);
   U783 : OAI211_X1 port map( C1 => n65, C2 => n2093, A => n449, B => n448, ZN 
                           => curr_proc_regs(248));
   U784 : INV_X1 port map( A => regs(761), ZN => n2096);
   U785 : AOI22_X1 port map( A1 => n113, A2 => regs(2297), B1 => n71, B2 => 
                           regs(1785), ZN => n451);
   U786 : AOI22_X1 port map( A1 => n93, A2 => regs(1273), B1 => n28, B2 => 
                           regs(249), ZN => n450);
   U787 : OAI211_X1 port map( C1 => n6, C2 => n2096, A => n451, B => n450, ZN 
                           => curr_proc_regs(249));
   U788 : INV_X1 port map( A => regs(536), ZN => n1367);
   U789 : AOI22_X1 port map( A1 => n114, A2 => regs(2072), B1 => n12, B2 => 
                           regs(1560), ZN => n453);
   U790 : AOI22_X1 port map( A1 => n93, A2 => regs(1048), B1 => n40, B2 => 
                           regs(24), ZN => n452);
   U791 : OAI211_X1 port map( C1 => n6, C2 => n1367, A => n453, B => n452, ZN 
                           => curr_proc_regs(24));
   U792 : INV_X1 port map( A => regs(762), ZN => n2099);
   U793 : AOI22_X1 port map( A1 => win(4), A2 => regs(2298), B1 => n13, B2 => 
                           regs(1786), ZN => n455);
   U794 : AOI22_X1 port map( A1 => n93, A2 => regs(1274), B1 => n33, B2 => 
                           regs(250), ZN => n454);
   U795 : OAI211_X1 port map( C1 => n66, C2 => n2099, A => n455, B => n454, ZN 
                           => curr_proc_regs(250));
   U796 : INV_X1 port map( A => regs(1275), ZN => n2102);
   U797 : AOI22_X1 port map( A1 => n113, A2 => regs(2299), B1 => n12, B2 => 
                           regs(1787), ZN => n457);
   U798 : AOI22_X1 port map( A1 => n51, A2 => regs(763), B1 => n30, B2 => 
                           regs(251), ZN => n456);
   U799 : OAI211_X1 port map( C1 => n2199, C2 => n2102, A => n457, B => n456, 
                           ZN => curr_proc_regs(251));
   U800 : INV_X1 port map( A => regs(1276), ZN => n2105);
   U801 : AOI22_X1 port map( A1 => n114, A2 => regs(2300), B1 => n69, B2 => 
                           regs(1788), ZN => n459);
   U802 : AOI22_X1 port map( A1 => n51, A2 => regs(764), B1 => n26, B2 => 
                           regs(252), ZN => n458);
   U803 : OAI211_X1 port map( C1 => n99, C2 => n2105, A => n459, B => n458, ZN 
                           => curr_proc_regs(252));
   U804 : INV_X1 port map( A => regs(765), ZN => n2108);
   U805 : AOI22_X1 port map( A1 => n114, A2 => regs(2301), B1 => n71, B2 => 
                           regs(1789), ZN => n461);
   U806 : AOI22_X1 port map( A1 => n93, A2 => regs(1277), B1 => n32, B2 => 
                           regs(253), ZN => n460);
   U807 : OAI211_X1 port map( C1 => n1, C2 => n2108, A => n461, B => n460, ZN 
                           => curr_proc_regs(253));
   U808 : INV_X1 port map( A => regs(766), ZN => n2111);
   U809 : AOI22_X1 port map( A1 => n114, A2 => regs(2302), B1 => n71, B2 => 
                           regs(1790), ZN => n463);
   U810 : AOI22_X1 port map( A1 => n93, A2 => regs(1278), B1 => n33, B2 => 
                           regs(254), ZN => n462);
   U811 : OAI211_X1 port map( C1 => n2185, C2 => n2111, A => n463, B => n462, 
                           ZN => curr_proc_regs(254));
   U812 : INV_X1 port map( A => regs(1279), ZN => n2115);
   U813 : AOI22_X1 port map( A1 => n114, A2 => regs(2303), B1 => n16, B2 => 
                           regs(1791), ZN => n465);
   U814 : AOI22_X1 port map( A1 => n51, A2 => regs(767), B1 => n30, B2 => 
                           regs(255), ZN => n464);
   U815 : OAI211_X1 port map( C1 => n15, C2 => n2115, A => n465, B => n464, ZN 
                           => curr_proc_regs(255));
   U816 : NAND2_X1 port map( A1 => regs(768), A2 => n62, ZN => n468);
   U817 : AOI22_X1 port map( A1 => n93, A2 => regs(1280), B1 => n26, B2 => 
                           regs(256), ZN => n467);
   U818 : AOI22_X1 port map( A1 => n114, A2 => regs(2304), B1 => n2195, B2 => 
                           regs(1792), ZN => n466);
   U819 : NAND3_X1 port map( A1 => n468, A2 => n467, A3 => n466, ZN => 
                           curr_proc_regs(256));
   U820 : NAND2_X1 port map( A1 => regs(1281), A2 => n18, ZN => n471);
   U821 : AOI22_X1 port map( A1 => n51, A2 => regs(769), B1 => n40, B2 => 
                           regs(257), ZN => n470);
   U822 : AOI22_X1 port map( A1 => n114, A2 => regs(2305), B1 => n72, B2 => 
                           regs(1793), ZN => n469);
   U823 : NAND3_X1 port map( A1 => n471, A2 => n470, A3 => n469, ZN => 
                           curr_proc_regs(257));
   U824 : NAND2_X1 port map( A1 => regs(1282), A2 => n17, ZN => n474);
   U825 : AOI22_X1 port map( A1 => n57, A2 => regs(770), B1 => n37, B2 => 
                           regs(258), ZN => n473);
   U826 : AOI22_X1 port map( A1 => n114, A2 => regs(2306), B1 => n3, B2 => 
                           regs(1794), ZN => n472);
   U827 : NAND3_X1 port map( A1 => n474, A2 => n473, A3 => n472, ZN => 
                           curr_proc_regs(258));
   U828 : NAND2_X1 port map( A1 => regs(1283), A2 => n17, ZN => n477);
   U829 : AOI22_X1 port map( A1 => n59, A2 => regs(771), B1 => n27, B2 => 
                           regs(259), ZN => n476);
   U830 : AOI22_X1 port map( A1 => n114, A2 => regs(2307), B1 => n70, B2 => 
                           regs(1795), ZN => n475);
   U831 : NAND3_X1 port map( A1 => n477, A2 => n476, A3 => n475, ZN => 
                           curr_proc_regs(259));
   U832 : INV_X1 port map( A => regs(1049), ZN => n1370);
   U833 : AOI22_X1 port map( A1 => n114, A2 => regs(2073), B1 => n70, B2 => 
                           regs(1561), ZN => n479);
   U834 : AOI22_X1 port map( A1 => n61, A2 => regs(537), B1 => n33, B2 => 
                           regs(25), ZN => n478);
   U835 : OAI211_X1 port map( C1 => n99, C2 => n1370, A => n479, B => n478, ZN 
                           => curr_proc_regs(25));
   U836 : NAND2_X1 port map( A1 => regs(1284), A2 => n93, ZN => n482);
   U837 : AOI22_X1 port map( A1 => n56, A2 => regs(772), B1 => n30, B2 => 
                           regs(260), ZN => n481);
   U838 : AOI22_X1 port map( A1 => n114, A2 => regs(2308), B1 => n70, B2 => 
                           regs(1796), ZN => n480);
   U839 : NAND3_X1 port map( A1 => n482, A2 => n481, A3 => n480, ZN => 
                           curr_proc_regs(260));
   U840 : NAND2_X1 port map( A1 => regs(1285), A2 => n18, ZN => n485);
   U841 : AOI22_X1 port map( A1 => n49, A2 => regs(773), B1 => n32, B2 => 
                           regs(261), ZN => n484);
   U842 : AOI22_X1 port map( A1 => n114, A2 => regs(2309), B1 => n70, B2 => 
                           regs(1797), ZN => n483);
   U843 : NAND3_X1 port map( A1 => n485, A2 => n484, A3 => n483, ZN => 
                           curr_proc_regs(261));
   U844 : NAND2_X1 port map( A1 => regs(1286), A2 => n91, ZN => n488);
   U845 : AOI22_X1 port map( A1 => n50, A2 => regs(774), B1 => n28, B2 => 
                           regs(262), ZN => n487);
   U846 : AOI22_X1 port map( A1 => n114, A2 => regs(2310), B1 => n70, B2 => 
                           regs(1798), ZN => n486);
   U847 : NAND3_X1 port map( A1 => n488, A2 => n487, A3 => n486, ZN => 
                           curr_proc_regs(262));
   U848 : NAND2_X1 port map( A1 => regs(775), A2 => n5, ZN => n491);
   U849 : AOI22_X1 port map( A1 => n92, A2 => regs(1287), B1 => n27, B2 => 
                           regs(263), ZN => n490);
   U850 : AOI22_X1 port map( A1 => win(4), A2 => regs(2311), B1 => n70, B2 => 
                           regs(1799), ZN => n489);
   U851 : NAND3_X1 port map( A1 => n491, A2 => n490, A3 => n489, ZN => 
                           curr_proc_regs(263));
   U852 : NAND2_X1 port map( A1 => regs(1288), A2 => n18, ZN => n494);
   U853 : AOI22_X1 port map( A1 => n51, A2 => regs(776), B1 => n26, B2 => 
                           regs(264), ZN => n493);
   U854 : AOI22_X1 port map( A1 => win(4), A2 => regs(2312), B1 => n70, B2 => 
                           regs(1800), ZN => n492);
   U855 : NAND3_X1 port map( A1 => n494, A2 => n493, A3 => n492, ZN => 
                           curr_proc_regs(264));
   U856 : NAND2_X1 port map( A1 => regs(1289), A2 => n89, ZN => n497);
   U857 : AOI22_X1 port map( A1 => n8, A2 => regs(777), B1 => n37, B2 => 
                           regs(265), ZN => n496);
   U858 : AOI22_X1 port map( A1 => win(4), A2 => regs(2313), B1 => n70, B2 => 
                           regs(1801), ZN => n495);
   U859 : NAND3_X1 port map( A1 => n497, A2 => n496, A3 => n495, ZN => 
                           curr_proc_regs(265));
   U860 : NAND2_X1 port map( A1 => regs(778), A2 => n5, ZN => n500);
   U861 : AOI22_X1 port map( A1 => n92, A2 => regs(1290), B1 => n30, B2 => 
                           regs(266), ZN => n499);
   U862 : AOI22_X1 port map( A1 => win(4), A2 => regs(2314), B1 => n70, B2 => 
                           regs(1802), ZN => n498);
   U863 : NAND3_X1 port map( A1 => n500, A2 => n499, A3 => n498, ZN => 
                           curr_proc_regs(266));
   U864 : NAND2_X1 port map( A1 => regs(779), A2 => n63, ZN => n503);
   U865 : AOI22_X1 port map( A1 => n92, A2 => regs(1291), B1 => n32, B2 => 
                           regs(267), ZN => n502);
   U866 : AOI22_X1 port map( A1 => n114, A2 => regs(2315), B1 => n70, B2 => 
                           regs(1803), ZN => n501);
   U867 : NAND3_X1 port map( A1 => n503, A2 => n502, A3 => n501, ZN => 
                           curr_proc_regs(267));
   U868 : NAND2_X1 port map( A1 => regs(780), A2 => n63, ZN => n506);
   U869 : AOI22_X1 port map( A1 => n92, A2 => regs(1292), B1 => n40, B2 => 
                           regs(268), ZN => n505);
   U870 : AOI22_X1 port map( A1 => n113, A2 => regs(2316), B1 => n70, B2 => 
                           regs(1804), ZN => n504);
   U871 : NAND3_X1 port map( A1 => n506, A2 => n505, A3 => n504, ZN => 
                           curr_proc_regs(268));
   U872 : NAND2_X1 port map( A1 => regs(781), A2 => n63, ZN => n509);
   U873 : AOI22_X1 port map( A1 => n92, A2 => regs(1293), B1 => n32, B2 => 
                           regs(269), ZN => n508);
   U874 : AOI22_X1 port map( A1 => n107, A2 => regs(2317), B1 => n73, B2 => 
                           regs(1805), ZN => n507);
   U875 : NAND3_X1 port map( A1 => n509, A2 => n508, A3 => n507, ZN => 
                           curr_proc_regs(269));
   U876 : INV_X1 port map( A => regs(1050), ZN => n1373);
   U877 : AOI22_X1 port map( A1 => n108, A2 => regs(2074), B1 => n73, B2 => 
                           regs(1562), ZN => n511);
   U878 : AOI22_X1 port map( A1 => n61, A2 => regs(538), B1 => n37, B2 => 
                           regs(26), ZN => n510);
   U879 : OAI211_X1 port map( C1 => n2199, C2 => n1373, A => n511, B => n510, 
                           ZN => curr_proc_regs(26));
   U880 : NAND2_X1 port map( A1 => regs(1294), A2 => n18, ZN => n514);
   U881 : AOI22_X1 port map( A1 => n8, A2 => regs(782), B1 => n40, B2 => 
                           regs(270), ZN => n513);
   U882 : AOI22_X1 port map( A1 => n109, A2 => regs(2318), B1 => n73, B2 => 
                           regs(1806), ZN => n512);
   U883 : NAND3_X1 port map( A1 => n514, A2 => n513, A3 => n512, ZN => 
                           curr_proc_regs(270));
   U884 : NAND2_X1 port map( A1 => regs(1295), A2 => n18, ZN => n517);
   U885 : AOI22_X1 port map( A1 => n52, A2 => regs(783), B1 => n28, B2 => 
                           regs(271), ZN => n516);
   U886 : AOI22_X1 port map( A1 => n104, A2 => regs(2319), B1 => n73, B2 => 
                           regs(1807), ZN => n515);
   U887 : NAND3_X1 port map( A1 => n517, A2 => n516, A3 => n515, ZN => 
                           curr_proc_regs(271));
   U888 : NAND2_X1 port map( A1 => regs(784), A2 => n5, ZN => n520);
   U889 : AOI22_X1 port map( A1 => n91, A2 => regs(1296), B1 => n28, B2 => 
                           regs(272), ZN => n519);
   U890 : AOI22_X1 port map( A1 => n4, A2 => regs(2320), B1 => n73, B2 => 
                           regs(1808), ZN => n518);
   U891 : NAND3_X1 port map( A1 => n520, A2 => n519, A3 => n518, ZN => 
                           curr_proc_regs(272));
   U892 : NAND2_X1 port map( A1 => regs(785), A2 => n63, ZN => n523);
   U893 : AOI22_X1 port map( A1 => n91, A2 => regs(1297), B1 => n27, B2 => 
                           regs(273), ZN => n522);
   U894 : AOI22_X1 port map( A1 => n116, A2 => regs(2321), B1 => n73, B2 => 
                           regs(1809), ZN => n521);
   U895 : NAND3_X1 port map( A1 => n523, A2 => n522, A3 => n521, ZN => 
                           curr_proc_regs(273));
   U896 : NAND2_X1 port map( A1 => regs(1298), A2 => n18, ZN => n526);
   U897 : AOI22_X1 port map( A1 => n8, A2 => regs(786), B1 => n26, B2 => 
                           regs(274), ZN => n525);
   U898 : AOI22_X1 port map( A1 => n116, A2 => regs(2322), B1 => n73, B2 => 
                           regs(1810), ZN => n524);
   U899 : NAND3_X1 port map( A1 => n526, A2 => n525, A3 => n524, ZN => 
                           curr_proc_regs(274));
   U900 : NAND2_X1 port map( A1 => regs(787), A2 => n5, ZN => n529);
   U901 : AOI22_X1 port map( A1 => n91, A2 => regs(1299), B1 => n28, B2 => 
                           regs(275), ZN => n528);
   U902 : AOI22_X1 port map( A1 => n116, A2 => regs(2323), B1 => n73, B2 => 
                           regs(1811), ZN => n527);
   U903 : NAND3_X1 port map( A1 => n529, A2 => n528, A3 => n527, ZN => 
                           curr_proc_regs(275));
   U904 : NAND2_X1 port map( A1 => regs(1300), A2 => n18, ZN => n532);
   U905 : AOI22_X1 port map( A1 => n53, A2 => regs(788), B1 => n32, B2 => 
                           regs(276), ZN => n531);
   U906 : AOI22_X1 port map( A1 => n116, A2 => regs(2324), B1 => n73, B2 => 
                           regs(1812), ZN => n530);
   U907 : NAND3_X1 port map( A1 => n532, A2 => n531, A3 => n530, ZN => 
                           curr_proc_regs(276));
   U908 : NAND2_X1 port map( A1 => regs(789), A2 => n5, ZN => n535);
   U909 : AOI22_X1 port map( A1 => n91, A2 => regs(1301), B1 => n37, B2 => 
                           regs(277), ZN => n534);
   U910 : AOI22_X1 port map( A1 => n116, A2 => regs(2325), B1 => n73, B2 => 
                           regs(1813), ZN => n533);
   U911 : NAND3_X1 port map( A1 => n535, A2 => n534, A3 => n533, ZN => 
                           curr_proc_regs(277));
   U912 : NAND2_X1 port map( A1 => regs(1302), A2 => n18, ZN => n538);
   U913 : AOI22_X1 port map( A1 => n49, A2 => regs(790), B1 => n37, B2 => 
                           regs(278), ZN => n537);
   U914 : AOI22_X1 port map( A1 => n116, A2 => regs(2326), B1 => n73, B2 => 
                           regs(1814), ZN => n536);
   U915 : NAND3_X1 port map( A1 => n538, A2 => n537, A3 => n536, ZN => 
                           curr_proc_regs(278));
   U916 : NAND2_X1 port map( A1 => regs(791), A2 => n5, ZN => n541);
   U917 : AOI22_X1 port map( A1 => n90, A2 => regs(1303), B1 => n38, B2 => 
                           regs(279), ZN => n540);
   U918 : AOI22_X1 port map( A1 => n116, A2 => regs(2327), B1 => n3, B2 => 
                           regs(1815), ZN => n539);
   U919 : NAND3_X1 port map( A1 => n541, A2 => n540, A3 => n539, ZN => 
                           curr_proc_regs(279));
   U920 : INV_X1 port map( A => regs(1051), ZN => n1376);
   U921 : AOI22_X1 port map( A1 => n116, A2 => regs(2075), B1 => n3, B2 => 
                           regs(1563), ZN => n543);
   U922 : AOI22_X1 port map( A1 => n8, A2 => regs(539), B1 => n7, B2 => 
                           regs(27), ZN => n542);
   U923 : OAI211_X1 port map( C1 => n2199, C2 => n1376, A => n543, B => n542, 
                           ZN => curr_proc_regs(27));
   U924 : NAND2_X1 port map( A1 => regs(792), A2 => n63, ZN => n546);
   U925 : AOI22_X1 port map( A1 => n90, A2 => regs(1304), B1 => n41, B2 => 
                           regs(280), ZN => n545);
   U926 : AOI22_X1 port map( A1 => n116, A2 => regs(2328), B1 => n71, B2 => 
                           regs(1816), ZN => n544);
   U927 : NAND3_X1 port map( A1 => n546, A2 => n545, A3 => n544, ZN => 
                           curr_proc_regs(280));
   U928 : NAND2_X1 port map( A1 => regs(793), A2 => n5, ZN => n549);
   U929 : AOI22_X1 port map( A1 => n90, A2 => regs(1305), B1 => n38, B2 => 
                           regs(281), ZN => n548);
   U930 : AOI22_X1 port map( A1 => n116, A2 => regs(2329), B1 => n71, B2 => 
                           regs(1817), ZN => n547);
   U931 : NAND3_X1 port map( A1 => n549, A2 => n548, A3 => n547, ZN => 
                           curr_proc_regs(281));
   U932 : NAND2_X1 port map( A1 => regs(1306), A2 => n18, ZN => n552);
   U933 : AOI22_X1 port map( A1 => n48, A2 => regs(794), B1 => n26, B2 => 
                           regs(282), ZN => n551);
   U934 : AOI22_X1 port map( A1 => n116, A2 => regs(2330), B1 => n68, B2 => 
                           regs(1818), ZN => n550);
   U935 : NAND3_X1 port map( A1 => n552, A2 => n551, A3 => n550, ZN => 
                           curr_proc_regs(282));
   U936 : NAND2_X1 port map( A1 => regs(1307), A2 => n18, ZN => n555);
   U937 : AOI22_X1 port map( A1 => n8, A2 => regs(795), B1 => n27, B2 => 
                           regs(283), ZN => n554);
   U938 : AOI22_X1 port map( A1 => n116, A2 => regs(2331), B1 => n73, B2 => 
                           regs(1819), ZN => n553);
   U939 : NAND3_X1 port map( A1 => n555, A2 => n554, A3 => n553, ZN => 
                           curr_proc_regs(283));
   U940 : NAND2_X1 port map( A1 => regs(1308), A2 => n18, ZN => n558);
   U941 : AOI22_X1 port map( A1 => n48, A2 => regs(796), B1 => n40, B2 => 
                           regs(284), ZN => n557);
   U942 : AOI22_X1 port map( A1 => n116, A2 => regs(2332), B1 => n73, B2 => 
                           regs(1820), ZN => n556);
   U943 : NAND3_X1 port map( A1 => n558, A2 => n557, A3 => n556, ZN => 
                           curr_proc_regs(284));
   U944 : NAND2_X1 port map( A1 => regs(797), A2 => n5, ZN => n561);
   U945 : AOI22_X1 port map( A1 => n90, A2 => regs(1309), B1 => n40, B2 => 
                           regs(285), ZN => n560);
   U946 : AOI22_X1 port map( A1 => n116, A2 => regs(2333), B1 => n73, B2 => 
                           regs(1821), ZN => n559);
   U947 : NAND3_X1 port map( A1 => n561, A2 => n560, A3 => n559, ZN => 
                           curr_proc_regs(285));
   U948 : NAND2_X1 port map( A1 => regs(798), A2 => n5, ZN => n564);
   U949 : AOI22_X1 port map( A1 => n90, A2 => regs(1310), B1 => n28, B2 => 
                           regs(286), ZN => n563);
   U950 : AOI22_X1 port map( A1 => n116, A2 => regs(2334), B1 => n16, B2 => 
                           regs(1822), ZN => n562);
   U951 : NAND3_X1 port map( A1 => n564, A2 => n563, A3 => n562, ZN => 
                           curr_proc_regs(286));
   U952 : NAND2_X1 port map( A1 => regs(1311), A2 => n14, ZN => n567);
   U953 : AOI22_X1 port map( A1 => n5, A2 => regs(799), B1 => n33, B2 => 
                           regs(287), ZN => n566);
   U954 : AOI22_X1 port map( A1 => n116, A2 => regs(2335), B1 => n16, B2 => 
                           regs(1823), ZN => n565);
   U955 : NAND3_X1 port map( A1 => n567, A2 => n566, A3 => n565, ZN => 
                           curr_proc_regs(287));
   U956 : NAND2_X1 port map( A1 => regs(800), A2 => n5, ZN => n570);
   U957 : AOI22_X1 port map( A1 => n89, A2 => regs(1312), B1 => n30, B2 => 
                           regs(288), ZN => n569);
   U958 : AOI22_X1 port map( A1 => n116, A2 => regs(2336), B1 => n12, B2 => 
                           regs(1824), ZN => n568);
   U959 : NAND3_X1 port map( A1 => n570, A2 => n569, A3 => n568, ZN => 
                           curr_proc_regs(288));
   U960 : NAND2_X1 port map( A1 => regs(801), A2 => n5, ZN => n573);
   U961 : AOI22_X1 port map( A1 => n91, A2 => regs(1313), B1 => n41, B2 => 
                           regs(289), ZN => n572);
   U962 : AOI22_X1 port map( A1 => n116, A2 => regs(2337), B1 => n72, B2 => 
                           regs(1825), ZN => n571);
   U963 : NAND3_X1 port map( A1 => n573, A2 => n572, A3 => n571, ZN => 
                           curr_proc_regs(289));
   U964 : INV_X1 port map( A => regs(540), ZN => n1381);
   U965 : AOI22_X1 port map( A1 => n116, A2 => regs(2076), B1 => n72, B2 => 
                           regs(1564), ZN => n575);
   U966 : AOI22_X1 port map( A1 => n89, A2 => regs(1052), B1 => n41, B2 => 
                           regs(28), ZN => n574);
   U967 : OAI211_X1 port map( C1 => n65, C2 => n1381, A => n575, B => n574, ZN 
                           => curr_proc_regs(28));
   U968 : NAND2_X1 port map( A1 => regs(802), A2 => n63, ZN => n578);
   U969 : AOI22_X1 port map( A1 => n90, A2 => regs(1314), B1 => n25, B2 => 
                           regs(290), ZN => n577);
   U970 : AOI22_X1 port map( A1 => n116, A2 => regs(2338), B1 => n72, B2 => 
                           regs(1826), ZN => n576);
   U971 : NAND3_X1 port map( A1 => n578, A2 => n577, A3 => n576, ZN => 
                           curr_proc_regs(290));
   U972 : NAND2_X1 port map( A1 => regs(803), A2 => n5, ZN => n581);
   U973 : AOI22_X1 port map( A1 => n90, A2 => regs(1315), B1 => n2, B2 => 
                           regs(291), ZN => n580);
   U974 : AOI22_X1 port map( A1 => n116, A2 => regs(2339), B1 => n72, B2 => 
                           regs(1827), ZN => n579);
   U975 : NAND3_X1 port map( A1 => n581, A2 => n580, A3 => n579, ZN => 
                           curr_proc_regs(291));
   U976 : NAND2_X1 port map( A1 => regs(804), A2 => n5, ZN => n584);
   U977 : AOI22_X1 port map( A1 => n90, A2 => regs(1316), B1 => n41, B2 => 
                           regs(292), ZN => n583);
   U978 : AOI22_X1 port map( A1 => n116, A2 => regs(2340), B1 => n72, B2 => 
                           regs(1828), ZN => n582);
   U979 : NAND3_X1 port map( A1 => n584, A2 => n583, A3 => n582, ZN => 
                           curr_proc_regs(292));
   U980 : NAND2_X1 port map( A1 => regs(1317), A2 => n14, ZN => n587);
   U981 : AOI22_X1 port map( A1 => n5, A2 => regs(805), B1 => n2, B2 => 
                           regs(293), ZN => n586);
   U982 : AOI22_X1 port map( A1 => n116, A2 => regs(2341), B1 => n72, B2 => 
                           regs(1829), ZN => n585);
   U983 : NAND3_X1 port map( A1 => n587, A2 => n586, A3 => n585, ZN => 
                           curr_proc_regs(293));
   U984 : NAND2_X1 port map( A1 => regs(806), A2 => n5, ZN => n590);
   U985 : AOI22_X1 port map( A1 => n90, A2 => regs(1318), B1 => n2, B2 => 
                           regs(294), ZN => n589);
   U986 : AOI22_X1 port map( A1 => n116, A2 => regs(2342), B1 => n72, B2 => 
                           regs(1830), ZN => n588);
   U987 : NAND3_X1 port map( A1 => n590, A2 => n589, A3 => n588, ZN => 
                           curr_proc_regs(294));
   U988 : NAND2_X1 port map( A1 => regs(1319), A2 => n14, ZN => n593);
   U989 : AOI22_X1 port map( A1 => n5, A2 => regs(807), B1 => n7, B2 => 
                           regs(295), ZN => n592);
   U990 : AOI22_X1 port map( A1 => n116, A2 => regs(2343), B1 => n72, B2 => 
                           regs(1831), ZN => n591);
   U991 : NAND3_X1 port map( A1 => n593, A2 => n592, A3 => n591, ZN => 
                           curr_proc_regs(295));
   U992 : NAND2_X1 port map( A1 => regs(808), A2 => n5, ZN => n596);
   U993 : AOI22_X1 port map( A1 => n90, A2 => regs(1320), B1 => n7, B2 => 
                           regs(296), ZN => n595);
   U994 : AOI22_X1 port map( A1 => n116, A2 => regs(2344), B1 => n72, B2 => 
                           regs(1832), ZN => n594);
   U995 : NAND3_X1 port map( A1 => n596, A2 => n595, A3 => n594, ZN => 
                           curr_proc_regs(296));
   U996 : NAND2_X1 port map( A1 => regs(809), A2 => n5, ZN => n599);
   U997 : AOI22_X1 port map( A1 => n90, A2 => regs(1321), B1 => n25, B2 => 
                           regs(297), ZN => n598);
   U998 : AOI22_X1 port map( A1 => n116, A2 => regs(2345), B1 => n72, B2 => 
                           regs(1833), ZN => n597);
   U999 : NAND3_X1 port map( A1 => n599, A2 => n598, A3 => n597, ZN => 
                           curr_proc_regs(297));
   U1000 : NAND2_X1 port map( A1 => regs(1322), A2 => n14, ZN => n602);
   U1001 : AOI22_X1 port map( A1 => n8, A2 => regs(810), B1 => n38, B2 => 
                           regs(298), ZN => n601);
   U1002 : AOI22_X1 port map( A1 => n116, A2 => regs(2346), B1 => n72, B2 => 
                           regs(1834), ZN => n600);
   U1003 : NAND3_X1 port map( A1 => n602, A2 => n601, A3 => n600, ZN => 
                           curr_proc_regs(298));
   U1004 : NAND2_X1 port map( A1 => regs(811), A2 => n5, ZN => n605);
   U1005 : AOI22_X1 port map( A1 => n91, A2 => regs(1323), B1 => n2, B2 => 
                           regs(299), ZN => n604);
   U1006 : AOI22_X1 port map( A1 => n116, A2 => regs(2347), B1 => n68, B2 => 
                           regs(1835), ZN => n603);
   U1007 : NAND3_X1 port map( A1 => n605, A2 => n604, A3 => n603, ZN => 
                           curr_proc_regs(299));
   U1008 : INV_X1 port map( A => regs(1053), ZN => n1384);
   U1009 : AOI22_X1 port map( A1 => n116, A2 => regs(2077), B1 => n71, B2 => 
                           regs(1565), ZN => n607);
   U1010 : AOI22_X1 port map( A1 => n50, A2 => regs(541), B1 => n2, B2 => 
                           regs(29), ZN => n606);
   U1011 : OAI211_X1 port map( C1 => n15, C2 => n1384, A => n607, B => n606, ZN
                           => curr_proc_regs(29));
   U1012 : INV_X1 port map( A => regs(514), ZN => n1300);
   U1013 : AOI22_X1 port map( A1 => n116, A2 => regs(2050), B1 => n73, B2 => 
                           regs(1538), ZN => n609);
   U1014 : AOI22_X1 port map( A1 => n91, A2 => regs(1026), B1 => n2, B2 => 
                           regs(2), ZN => n608);
   U1015 : OAI211_X1 port map( C1 => n67, C2 => n1300, A => n609, B => n608, ZN
                           => curr_proc_regs(2));
   U1016 : NAND2_X1 port map( A1 => regs(812), A2 => n5, ZN => n612);
   U1017 : AOI22_X1 port map( A1 => n91, A2 => regs(1324), B1 => n31, B2 => 
                           regs(300), ZN => n611);
   U1018 : AOI22_X1 port map( A1 => n116, A2 => regs(2348), B1 => n11, B2 => 
                           regs(1836), ZN => n610);
   U1019 : NAND3_X1 port map( A1 => n612, A2 => n611, A3 => n610, ZN => 
                           curr_proc_regs(300));
   U1020 : NAND2_X1 port map( A1 => regs(813), A2 => n5, ZN => n615);
   U1021 : AOI22_X1 port map( A1 => n91, A2 => regs(1325), B1 => n38, B2 => 
                           regs(301), ZN => n614);
   U1022 : AOI22_X1 port map( A1 => n116, A2 => regs(2349), B1 => n3, B2 => 
                           regs(1837), ZN => n613);
   U1023 : NAND3_X1 port map( A1 => n615, A2 => n614, A3 => n613, ZN => 
                           curr_proc_regs(301));
   U1024 : NAND2_X1 port map( A1 => regs(814), A2 => n5, ZN => n618);
   U1025 : AOI22_X1 port map( A1 => n91, A2 => regs(1326), B1 => n41, B2 => 
                           regs(302), ZN => n617);
   U1026 : AOI22_X1 port map( A1 => n116, A2 => regs(2350), B1 => n3, B2 => 
                           regs(1838), ZN => n616);
   U1027 : NAND3_X1 port map( A1 => n618, A2 => n617, A3 => n616, ZN => 
                           curr_proc_regs(302));
   U1028 : NAND2_X1 port map( A1 => regs(815), A2 => n5, ZN => n621);
   U1029 : AOI22_X1 port map( A1 => n91, A2 => regs(1327), B1 => n2, B2 => 
                           regs(303), ZN => n620);
   U1030 : AOI22_X1 port map( A1 => n116, A2 => regs(2351), B1 => n3, B2 => 
                           regs(1839), ZN => n619);
   U1031 : NAND3_X1 port map( A1 => n621, A2 => n620, A3 => n619, ZN => 
                           curr_proc_regs(303));
   U1032 : NAND2_X1 port map( A1 => regs(1328), A2 => n14, ZN => n624);
   U1033 : AOI22_X1 port map( A1 => n49, A2 => regs(816), B1 => n2, B2 => 
                           regs(304), ZN => n623);
   U1034 : AOI22_X1 port map( A1 => n116, A2 => regs(2352), B1 => n3, B2 => 
                           regs(1840), ZN => n622);
   U1035 : NAND3_X1 port map( A1 => n624, A2 => n623, A3 => n622, ZN => 
                           curr_proc_regs(304));
   U1036 : NAND2_X1 port map( A1 => regs(817), A2 => n63, ZN => n627);
   U1037 : AOI22_X1 port map( A1 => n91, A2 => regs(1329), B1 => n7, B2 => 
                           regs(305), ZN => n626);
   U1038 : AOI22_X1 port map( A1 => n116, A2 => regs(2353), B1 => n70, B2 => 
                           regs(1841), ZN => n625);
   U1039 : NAND3_X1 port map( A1 => n627, A2 => n626, A3 => n625, ZN => 
                           curr_proc_regs(305));
   U1040 : NAND2_X1 port map( A1 => regs(1330), A2 => n14, ZN => n630);
   U1041 : AOI22_X1 port map( A1 => n8, A2 => regs(818), B1 => n7, B2 => 
                           regs(306), ZN => n629);
   U1042 : AOI22_X1 port map( A1 => n116, A2 => regs(2354), B1 => n75, B2 => 
                           regs(1842), ZN => n628);
   U1043 : NAND3_X1 port map( A1 => n630, A2 => n629, A3 => n628, ZN => 
                           curr_proc_regs(306));
   U1044 : NAND2_X1 port map( A1 => regs(1331), A2 => n14, ZN => n633);
   U1045 : AOI22_X1 port map( A1 => n8, A2 => regs(819), B1 => n25, B2 => 
                           regs(307), ZN => n632);
   U1046 : AOI22_X1 port map( A1 => n116, A2 => regs(2355), B1 => n16, B2 => 
                           regs(1843), ZN => n631);
   U1047 : NAND3_X1 port map( A1 => n633, A2 => n632, A3 => n631, ZN => 
                           curr_proc_regs(307));
   U1048 : NAND2_X1 port map( A1 => regs(820), A2 => n5, ZN => n636);
   U1049 : AOI22_X1 port map( A1 => n92, A2 => regs(1332), B1 => n36, B2 => 
                           regs(308), ZN => n635);
   U1050 : AOI22_X1 port map( A1 => n116, A2 => regs(2356), B1 => n11, B2 => 
                           regs(1844), ZN => n634);
   U1051 : NAND3_X1 port map( A1 => n636, A2 => n635, A3 => n634, ZN => 
                           curr_proc_regs(308));
   U1052 : NAND2_X1 port map( A1 => regs(821), A2 => n5, ZN => n639);
   U1053 : AOI22_X1 port map( A1 => n92, A2 => regs(1333), B1 => n35, B2 => 
                           regs(309), ZN => n638);
   U1054 : AOI22_X1 port map( A1 => n116, A2 => regs(2357), B1 => n11, B2 => 
                           regs(1845), ZN => n637);
   U1055 : NAND3_X1 port map( A1 => n639, A2 => n638, A3 => n637, ZN => 
                           curr_proc_regs(309));
   U1056 : INV_X1 port map( A => regs(1054), ZN => n1387);
   U1057 : AOI22_X1 port map( A1 => n116, A2 => regs(2078), B1 => n11, B2 => 
                           regs(1566), ZN => n641);
   U1058 : AOI22_X1 port map( A1 => n56, A2 => regs(542), B1 => n34, B2 => 
                           regs(30), ZN => n640);
   U1059 : OAI211_X1 port map( C1 => n2199, C2 => n1387, A => n641, B => n640, 
                           ZN => curr_proc_regs(30));
   U1060 : NAND2_X1 port map( A1 => regs(822), A2 => n5, ZN => n644);
   U1061 : AOI22_X1 port map( A1 => n92, A2 => regs(1334), B1 => n39, B2 => 
                           regs(310), ZN => n643);
   U1062 : AOI22_X1 port map( A1 => n116, A2 => regs(2358), B1 => n11, B2 => 
                           regs(1846), ZN => n642);
   U1063 : NAND3_X1 port map( A1 => n644, A2 => n643, A3 => n642, ZN => 
                           curr_proc_regs(310));
   U1064 : NAND2_X1 port map( A1 => regs(823), A2 => n5, ZN => n647);
   U1065 : AOI22_X1 port map( A1 => n92, A2 => regs(1335), B1 => n41, B2 => 
                           regs(311), ZN => n646);
   U1066 : AOI22_X1 port map( A1 => n116, A2 => regs(2359), B1 => n11, B2 => 
                           regs(1847), ZN => n645);
   U1067 : NAND3_X1 port map( A1 => n647, A2 => n646, A3 => n645, ZN => 
                           curr_proc_regs(311));
   U1068 : NAND2_X1 port map( A1 => regs(824), A2 => n5, ZN => n650);
   U1069 : AOI22_X1 port map( A1 => n92, A2 => regs(1336), B1 => n2, B2 => 
                           regs(312), ZN => n649);
   U1070 : AOI22_X1 port map( A1 => n116, A2 => regs(2360), B1 => n11, B2 => 
                           regs(1848), ZN => n648);
   U1071 : NAND3_X1 port map( A1 => n650, A2 => n649, A3 => n648, ZN => 
                           curr_proc_regs(312));
   U1072 : NAND2_X1 port map( A1 => regs(1337), A2 => n14, ZN => n653);
   U1073 : AOI22_X1 port map( A1 => n8, A2 => regs(825), B1 => n2, B2 => 
                           regs(313), ZN => n652);
   U1074 : AOI22_X1 port map( A1 => n116, A2 => regs(2361), B1 => n11, B2 => 
                           regs(1849), ZN => n651);
   U1075 : NAND3_X1 port map( A1 => n653, A2 => n652, A3 => n651, ZN => 
                           curr_proc_regs(313));
   U1076 : NAND2_X1 port map( A1 => regs(826), A2 => n5, ZN => n656);
   U1077 : AOI22_X1 port map( A1 => n92, A2 => regs(1338), B1 => n7, B2 => 
                           regs(314), ZN => n655);
   U1078 : AOI22_X1 port map( A1 => n116, A2 => regs(2362), B1 => n11, B2 => 
                           regs(1850), ZN => n654);
   U1079 : NAND3_X1 port map( A1 => n656, A2 => n655, A3 => n654, ZN => 
                           curr_proc_regs(314));
   U1080 : NAND2_X1 port map( A1 => regs(1339), A2 => n85, ZN => n659);
   U1081 : AOI22_X1 port map( A1 => n8, A2 => regs(827), B1 => n7, B2 => 
                           regs(315), ZN => n658);
   U1082 : AOI22_X1 port map( A1 => n116, A2 => regs(2363), B1 => n11, B2 => 
                           regs(1851), ZN => n657);
   U1083 : NAND3_X1 port map( A1 => n659, A2 => n658, A3 => n657, ZN => 
                           curr_proc_regs(315));
   U1084 : NAND2_X1 port map( A1 => regs(1340), A2 => n84, ZN => n662);
   U1085 : AOI22_X1 port map( A1 => n55, A2 => regs(828), B1 => n25, B2 => 
                           regs(316), ZN => n661);
   U1086 : AOI22_X1 port map( A1 => n116, A2 => regs(2364), B1 => n11, B2 => 
                           regs(1852), ZN => n660);
   U1087 : NAND3_X1 port map( A1 => n662, A2 => n661, A3 => n660, ZN => 
                           curr_proc_regs(316));
   U1088 : NAND2_X1 port map( A1 => regs(1341), A2 => n94, ZN => n665);
   U1089 : AOI22_X1 port map( A1 => n8, A2 => regs(829), B1 => n2, B2 => 
                           regs(317), ZN => n664);
   U1090 : AOI22_X1 port map( A1 => n116, A2 => regs(2365), B1 => n11, B2 => 
                           regs(1853), ZN => n663);
   U1091 : NAND3_X1 port map( A1 => n665, A2 => n664, A3 => n663, ZN => 
                           curr_proc_regs(317));
   U1092 : NAND2_X1 port map( A1 => regs(1342), A2 => n82, ZN => n668);
   U1093 : AOI22_X1 port map( A1 => n8, A2 => regs(830), B1 => n29, B2 => 
                           regs(318), ZN => n667);
   U1094 : AOI22_X1 port map( A1 => n116, A2 => regs(2366), B1 => n68, B2 => 
                           regs(1854), ZN => n666);
   U1095 : NAND3_X1 port map( A1 => n668, A2 => n667, A3 => n666, ZN => 
                           curr_proc_regs(318));
   U1096 : NAND2_X1 port map( A1 => regs(831), A2 => n5, ZN => n671);
   U1097 : AOI22_X1 port map( A1 => n93, A2 => regs(1343), B1 => n38, B2 => 
                           regs(319), ZN => n670);
   U1098 : AOI22_X1 port map( A1 => n116, A2 => regs(2367), B1 => n68, B2 => 
                           regs(1855), ZN => n669);
   U1099 : NAND3_X1 port map( A1 => n671, A2 => n670, A3 => n669, ZN => 
                           curr_proc_regs(319));
   U1100 : INV_X1 port map( A => regs(543), ZN => n1390);
   U1101 : AOI22_X1 port map( A1 => n116, A2 => regs(2079), B1 => n68, B2 => 
                           regs(1567), ZN => n673);
   U1102 : AOI22_X1 port map( A1 => n93, A2 => regs(1055), B1 => n41, B2 => 
                           regs(31), ZN => n672);
   U1103 : OAI211_X1 port map( C1 => n2185, C2 => n1390, A => n673, B => n672, 
                           ZN => curr_proc_regs(31));
   U1104 : NAND2_X1 port map( A1 => regs(1344), A2 => n98, ZN => n676);
   U1105 : AOI22_X1 port map( A1 => n8, A2 => regs(832), B1 => n2, B2 => 
                           regs(320), ZN => n675);
   U1106 : AOI22_X1 port map( A1 => n116, A2 => regs(2368), B1 => n68, B2 => 
                           regs(1856), ZN => n674);
   U1107 : NAND3_X1 port map( A1 => n676, A2 => n675, A3 => n674, ZN => 
                           curr_proc_regs(320));
   U1108 : NAND2_X1 port map( A1 => regs(1345), A2 => n84, ZN => n679);
   U1109 : AOI22_X1 port map( A1 => n10, A2 => regs(833), B1 => n41, B2 => 
                           regs(321), ZN => n678);
   U1110 : AOI22_X1 port map( A1 => n116, A2 => regs(2369), B1 => n68, B2 => 
                           regs(1857), ZN => n677);
   U1111 : NAND3_X1 port map( A1 => n679, A2 => n678, A3 => n677, ZN => 
                           curr_proc_regs(321));
   U1112 : NAND2_X1 port map( A1 => regs(834), A2 => n62, ZN => n682);
   U1113 : AOI22_X1 port map( A1 => n94, A2 => regs(1346), B1 => n45, B2 => 
                           regs(322), ZN => n681);
   U1114 : AOI22_X1 port map( A1 => n116, A2 => regs(2370), B1 => n68, B2 => 
                           regs(1858), ZN => n680);
   U1115 : NAND3_X1 port map( A1 => n682, A2 => n681, A3 => n680, ZN => 
                           curr_proc_regs(322));
   U1116 : NAND2_X1 port map( A1 => regs(835), A2 => n53, ZN => n685);
   U1117 : AOI22_X1 port map( A1 => n94, A2 => regs(1347), B1 => n44, B2 => 
                           regs(323), ZN => n684);
   U1118 : AOI22_X1 port map( A1 => n116, A2 => regs(2371), B1 => n68, B2 => 
                           regs(1859), ZN => n683);
   U1119 : NAND3_X1 port map( A1 => n685, A2 => n684, A3 => n683, ZN => 
                           curr_proc_regs(323));
   U1120 : NAND2_X1 port map( A1 => regs(1348), A2 => n79, ZN => n688);
   U1121 : AOI22_X1 port map( A1 => n5, A2 => regs(836), B1 => n43, B2 => 
                           regs(324), ZN => n687);
   U1122 : AOI22_X1 port map( A1 => n116, A2 => regs(2372), B1 => n68, B2 => 
                           regs(1860), ZN => n686);
   U1123 : NAND3_X1 port map( A1 => n688, A2 => n687, A3 => n686, ZN => 
                           curr_proc_regs(324));
   U1124 : NAND2_X1 port map( A1 => regs(837), A2 => n10, ZN => n691);
   U1125 : AOI22_X1 port map( A1 => n94, A2 => regs(1349), B1 => n27, B2 => 
                           regs(325), ZN => n690);
   U1126 : AOI22_X1 port map( A1 => n116, A2 => regs(2373), B1 => n68, B2 => 
                           regs(1861), ZN => n689);
   U1127 : NAND3_X1 port map( A1 => n691, A2 => n690, A3 => n689, ZN => 
                           curr_proc_regs(325));
   U1128 : NAND2_X1 port map( A1 => regs(838), A2 => n55, ZN => n694);
   U1129 : AOI22_X1 port map( A1 => n94, A2 => regs(1350), B1 => n26, B2 => 
                           regs(326), ZN => n693);
   U1130 : AOI22_X1 port map( A1 => n116, A2 => regs(2374), B1 => n68, B2 => 
                           regs(1862), ZN => n692);
   U1131 : NAND3_X1 port map( A1 => n694, A2 => n693, A3 => n692, ZN => 
                           curr_proc_regs(326));
   U1132 : NAND2_X1 port map( A1 => regs(1351), A2 => n96, ZN => n697);
   U1133 : AOI22_X1 port map( A1 => n8, A2 => regs(839), B1 => n25, B2 => 
                           regs(327), ZN => n696);
   U1134 : AOI22_X1 port map( A1 => n116, A2 => regs(2375), B1 => n68, B2 => 
                           regs(1863), ZN => n695);
   U1135 : NAND3_X1 port map( A1 => n697, A2 => n696, A3 => n695, ZN => 
                           curr_proc_regs(327));
   U1136 : NAND2_X1 port map( A1 => regs(1352), A2 => n96, ZN => n700);
   U1137 : AOI22_X1 port map( A1 => n10, A2 => regs(840), B1 => n7, B2 => 
                           regs(328), ZN => n699);
   U1138 : AOI22_X1 port map( A1 => n116, A2 => regs(2376), B1 => n68, B2 => 
                           regs(1864), ZN => n698);
   U1139 : NAND3_X1 port map( A1 => n700, A2 => n699, A3 => n698, ZN => 
                           curr_proc_regs(328));
   U1140 : NAND2_X1 port map( A1 => regs(841), A2 => n5, ZN => n703);
   U1141 : AOI22_X1 port map( A1 => n93, A2 => regs(1353), B1 => n25, B2 => 
                           regs(329), ZN => n702);
   U1142 : AOI22_X1 port map( A1 => n116, A2 => regs(2377), B1 => n73, B2 => 
                           regs(1865), ZN => n701);
   U1143 : NAND3_X1 port map( A1 => n703, A2 => n702, A3 => n701, ZN => 
                           curr_proc_regs(329));
   U1144 : INV_X1 port map( A => regs(544), ZN => n1393);
   U1145 : AOI22_X1 port map( A1 => n116, A2 => regs(2080), B1 => n68, B2 => 
                           regs(1568), ZN => n705);
   U1146 : AOI22_X1 port map( A1 => n91, A2 => regs(1056), B1 => n7, B2 => 
                           regs(32), ZN => n704);
   U1147 : OAI211_X1 port map( C1 => n67, C2 => n1393, A => n705, B => n704, ZN
                           => curr_proc_regs(32));
   U1148 : NAND2_X1 port map( A1 => regs(1354), A2 => n96, ZN => n708);
   U1149 : AOI22_X1 port map( A1 => n49, A2 => regs(842), B1 => n7, B2 => 
                           regs(330), ZN => n707);
   U1150 : AOI22_X1 port map( A1 => n116, A2 => regs(2378), B1 => n73, B2 => 
                           regs(1866), ZN => n706);
   U1151 : NAND3_X1 port map( A1 => n708, A2 => n707, A3 => n706, ZN => 
                           curr_proc_regs(330));
   U1152 : NAND2_X1 port map( A1 => regs(843), A2 => n60, ZN => n711);
   U1153 : AOI22_X1 port map( A1 => n17, A2 => regs(1355), B1 => n7, B2 => 
                           regs(331), ZN => n710);
   U1154 : AOI22_X1 port map( A1 => n116, A2 => regs(2379), B1 => n68, B2 => 
                           regs(1867), ZN => n709);
   U1155 : NAND3_X1 port map( A1 => n711, A2 => n710, A3 => n709, ZN => 
                           curr_proc_regs(331));
   U1156 : NAND2_X1 port map( A1 => regs(1356), A2 => n14, ZN => n714);
   U1157 : AOI22_X1 port map( A1 => n49, A2 => regs(844), B1 => n7, B2 => 
                           regs(332), ZN => n713);
   U1158 : AOI22_X1 port map( A1 => n116, A2 => regs(2380), B1 => n73, B2 => 
                           regs(1868), ZN => n712);
   U1159 : NAND3_X1 port map( A1 => n714, A2 => n713, A3 => n712, ZN => 
                           curr_proc_regs(332));
   U1160 : NAND2_X1 port map( A1 => regs(845), A2 => n5, ZN => n717);
   U1161 : AOI22_X1 port map( A1 => n89, A2 => regs(1357), B1 => n25, B2 => 
                           regs(333), ZN => n716);
   U1162 : AOI22_X1 port map( A1 => n116, A2 => regs(2381), B1 => n68, B2 => 
                           regs(1869), ZN => n715);
   U1163 : NAND3_X1 port map( A1 => n717, A2 => n716, A3 => n715, ZN => 
                           curr_proc_regs(333));
   U1164 : NAND2_X1 port map( A1 => regs(846), A2 => n60, ZN => n720);
   U1165 : AOI22_X1 port map( A1 => n91, A2 => regs(1358), B1 => n7, B2 => 
                           regs(334), ZN => n719);
   U1166 : AOI22_X1 port map( A1 => n116, A2 => regs(2382), B1 => n73, B2 => 
                           regs(1870), ZN => n718);
   U1167 : NAND3_X1 port map( A1 => n720, A2 => n719, A3 => n718, ZN => 
                           curr_proc_regs(334));
   U1168 : NAND2_X1 port map( A1 => regs(847), A2 => n10, ZN => n723);
   U1169 : AOI22_X1 port map( A1 => n17, A2 => regs(1359), B1 => n2, B2 => 
                           regs(335), ZN => n722);
   U1170 : AOI22_X1 port map( A1 => n116, A2 => regs(2383), B1 => n68, B2 => 
                           regs(1871), ZN => n721);
   U1171 : NAND3_X1 port map( A1 => n723, A2 => n722, A3 => n721, ZN => 
                           curr_proc_regs(335));
   U1172 : NAND2_X1 port map( A1 => regs(1360), A2 => n95, ZN => n726);
   U1173 : AOI22_X1 port map( A1 => n52, A2 => regs(848), B1 => n7, B2 => 
                           regs(336), ZN => n725);
   U1174 : AOI22_X1 port map( A1 => n116, A2 => regs(2384), B1 => n73, B2 => 
                           regs(1872), ZN => n724);
   U1175 : NAND3_X1 port map( A1 => n726, A2 => n725, A3 => n724, ZN => 
                           curr_proc_regs(336));
   U1176 : NAND2_X1 port map( A1 => regs(849), A2 => n5, ZN => n729);
   U1177 : AOI22_X1 port map( A1 => n17, A2 => regs(1361), B1 => n31, B2 => 
                           regs(337), ZN => n728);
   U1178 : AOI22_X1 port map( A1 => n116, A2 => regs(2385), B1 => n68, B2 => 
                           regs(1873), ZN => n727);
   U1179 : NAND3_X1 port map( A1 => n729, A2 => n728, A3 => n727, ZN => 
                           curr_proc_regs(337));
   U1180 : NAND2_X1 port map( A1 => regs(1362), A2 => n92, ZN => n732);
   U1181 : AOI22_X1 port map( A1 => n50, A2 => regs(850), B1 => n43, B2 => 
                           regs(338), ZN => n731);
   U1182 : AOI22_X1 port map( A1 => n116, A2 => regs(2386), B1 => n73, B2 => 
                           regs(1874), ZN => n730);
   U1183 : NAND3_X1 port map( A1 => n732, A2 => n731, A3 => n730, ZN => 
                           curr_proc_regs(338));
   U1184 : NAND2_X1 port map( A1 => regs(1363), A2 => n96, ZN => n735);
   U1185 : AOI22_X1 port map( A1 => n50, A2 => regs(851), B1 => n43, B2 => 
                           regs(339), ZN => n734);
   U1186 : AOI22_X1 port map( A1 => n116, A2 => regs(2387), B1 => n72, B2 => 
                           regs(1875), ZN => n733);
   U1187 : NAND3_X1 port map( A1 => n735, A2 => n734, A3 => n733, ZN => 
                           curr_proc_regs(339));
   U1188 : INV_X1 port map( A => regs(1057), ZN => n1396);
   U1189 : AOI22_X1 port map( A1 => n116, A2 => regs(2081), B1 => n74, B2 => 
                           regs(1569), ZN => n737);
   U1190 : AOI22_X1 port map( A1 => n51, A2 => regs(545), B1 => n43, B2 => 
                           regs(33), ZN => n736);
   U1191 : OAI211_X1 port map( C1 => n15, C2 => n1396, A => n737, B => n736, ZN
                           => curr_proc_regs(33));
   U1192 : NAND2_X1 port map( A1 => regs(1364), A2 => n83, ZN => n740);
   U1193 : AOI22_X1 port map( A1 => n51, A2 => regs(852), B1 => n43, B2 => 
                           regs(340), ZN => n739);
   U1194 : AOI22_X1 port map( A1 => n116, A2 => regs(2388), B1 => n3, B2 => 
                           regs(1876), ZN => n738);
   U1195 : NAND3_X1 port map( A1 => n740, A2 => n739, A3 => n738, ZN => 
                           curr_proc_regs(340));
   U1196 : NAND2_X1 port map( A1 => regs(1365), A2 => n82, ZN => n743);
   U1197 : AOI22_X1 port map( A1 => n50, A2 => regs(853), B1 => n31, B2 => 
                           regs(341), ZN => n742);
   U1198 : AOI22_X1 port map( A1 => n116, A2 => regs(2389), B1 => n70, B2 => 
                           regs(1877), ZN => n741);
   U1199 : NAND3_X1 port map( A1 => n743, A2 => n742, A3 => n741, ZN => 
                           curr_proc_regs(341));
   U1200 : NAND2_X1 port map( A1 => regs(1366), A2 => n85, ZN => n746);
   U1201 : AOI22_X1 port map( A1 => n50, A2 => regs(854), B1 => n29, B2 => 
                           regs(342), ZN => n745);
   U1202 : AOI22_X1 port map( A1 => n116, A2 => regs(2390), B1 => n73, B2 => 
                           regs(1878), ZN => n744);
   U1203 : NAND3_X1 port map( A1 => n746, A2 => n745, A3 => n744, ZN => 
                           curr_proc_regs(342));
   U1204 : NAND2_X1 port map( A1 => regs(855), A2 => n5, ZN => n749);
   U1205 : AOI22_X1 port map( A1 => n93, A2 => regs(1367), B1 => n38, B2 => 
                           regs(343), ZN => n748);
   U1206 : AOI22_X1 port map( A1 => n116, A2 => regs(2391), B1 => n74, B2 => 
                           regs(1879), ZN => n747);
   U1207 : NAND3_X1 port map( A1 => n749, A2 => n748, A3 => n747, ZN => 
                           curr_proc_regs(343));
   U1208 : NAND2_X1 port map( A1 => regs(856), A2 => n5, ZN => n752);
   U1209 : AOI22_X1 port map( A1 => n89, A2 => regs(1368), B1 => n41, B2 => 
                           regs(344), ZN => n751);
   U1210 : AOI22_X1 port map( A1 => n116, A2 => regs(2392), B1 => n71, B2 => 
                           regs(1880), ZN => n750);
   U1211 : NAND3_X1 port map( A1 => n752, A2 => n751, A3 => n750, ZN => 
                           curr_proc_regs(344));
   U1212 : NAND2_X1 port map( A1 => regs(1369), A2 => n98, ZN => n755);
   U1213 : AOI22_X1 port map( A1 => n50, A2 => regs(857), B1 => n2, B2 => 
                           regs(345), ZN => n754);
   U1214 : AOI22_X1 port map( A1 => n116, A2 => regs(2393), B1 => n70, B2 => 
                           regs(1881), ZN => n753);
   U1215 : NAND3_X1 port map( A1 => n755, A2 => n754, A3 => n753, ZN => 
                           curr_proc_regs(345));
   U1216 : NAND2_X1 port map( A1 => regs(1370), A2 => n17, ZN => n758);
   U1217 : AOI22_X1 port map( A1 => n50, A2 => regs(858), B1 => n2, B2 => 
                           regs(346), ZN => n757);
   U1218 : AOI22_X1 port map( A1 => n116, A2 => regs(2394), B1 => n73, B2 => 
                           regs(1882), ZN => n756);
   U1219 : NAND3_X1 port map( A1 => n758, A2 => n757, A3 => n756, ZN => 
                           curr_proc_regs(346));
   U1220 : NAND2_X1 port map( A1 => regs(859), A2 => n63, ZN => n761);
   U1221 : AOI22_X1 port map( A1 => n17, A2 => regs(1371), B1 => n7, B2 => 
                           regs(347), ZN => n760);
   U1222 : AOI22_X1 port map( A1 => n116, A2 => regs(2395), B1 => n74, B2 => 
                           regs(1883), ZN => n759);
   U1223 : NAND3_X1 port map( A1 => n761, A2 => n760, A3 => n759, ZN => 
                           curr_proc_regs(347));
   U1224 : NAND2_X1 port map( A1 => regs(860), A2 => n63, ZN => n764);
   U1225 : AOI22_X1 port map( A1 => n17, A2 => regs(1372), B1 => n34, B2 => 
                           regs(348), ZN => n763);
   U1226 : AOI22_X1 port map( A1 => n116, A2 => regs(2396), B1 => n74, B2 => 
                           regs(1884), ZN => n762);
   U1227 : NAND3_X1 port map( A1 => n764, A2 => n763, A3 => n762, ZN => 
                           curr_proc_regs(348));
   U1228 : NAND2_X1 port map( A1 => regs(861), A2 => n55, ZN => n767);
   U1229 : AOI22_X1 port map( A1 => n17, A2 => regs(1373), B1 => n36, B2 => 
                           regs(349), ZN => n766);
   U1230 : AOI22_X1 port map( A1 => n116, A2 => regs(2397), B1 => n3, B2 => 
                           regs(1885), ZN => n765);
   U1231 : NAND3_X1 port map( A1 => n767, A2 => n766, A3 => n765, ZN => 
                           curr_proc_regs(349));
   U1232 : INV_X1 port map( A => regs(546), ZN => n1399);
   U1233 : AOI22_X1 port map( A1 => n116, A2 => regs(2082), B1 => n3, B2 => 
                           regs(1570), ZN => n769);
   U1234 : AOI22_X1 port map( A1 => n93, A2 => regs(1058), B1 => n34, B2 => 
                           regs(34), ZN => n768);
   U1235 : OAI211_X1 port map( C1 => n64, C2 => n1399, A => n769, B => n768, ZN
                           => curr_proc_regs(34));
   U1236 : NAND2_X1 port map( A1 => regs(862), A2 => n54, ZN => n772);
   U1237 : AOI22_X1 port map( A1 => n91, A2 => regs(1374), B1 => n36, B2 => 
                           regs(350), ZN => n771);
   U1238 : AOI22_X1 port map( A1 => n116, A2 => regs(2398), B1 => n70, B2 => 
                           regs(1886), ZN => n770);
   U1239 : NAND3_X1 port map( A1 => n772, A2 => n771, A3 => n770, ZN => 
                           curr_proc_regs(350));
   U1240 : NAND2_X1 port map( A1 => regs(863), A2 => n58, ZN => n775);
   U1241 : AOI22_X1 port map( A1 => n90, A2 => regs(1375), B1 => n33, B2 => 
                           regs(351), ZN => n774);
   U1242 : AOI22_X1 port map( A1 => n116, A2 => regs(2399), B1 => n73, B2 => 
                           regs(1887), ZN => n773);
   U1243 : NAND3_X1 port map( A1 => n775, A2 => n774, A3 => n773, ZN => 
                           curr_proc_regs(351));
   U1244 : NAND2_X1 port map( A1 => regs(864), A2 => n57, ZN => n778);
   U1245 : AOI22_X1 port map( A1 => n91, A2 => regs(1376), B1 => n33, B2 => 
                           regs(352), ZN => n777);
   U1246 : AOI22_X1 port map( A1 => n116, A2 => regs(2400), B1 => n74, B2 => 
                           regs(1888), ZN => n776);
   U1247 : NAND3_X1 port map( A1 => n778, A2 => n777, A3 => n776, ZN => 
                           curr_proc_regs(352));
   U1248 : NAND2_X1 port map( A1 => regs(1377), A2 => n82, ZN => n781);
   U1249 : AOI22_X1 port map( A1 => n51, A2 => regs(865), B1 => n33, B2 => 
                           regs(353), ZN => n780);
   U1250 : AOI22_X1 port map( A1 => n116, A2 => regs(2401), B1 => n73, B2 => 
                           regs(1889), ZN => n779);
   U1251 : NAND3_X1 port map( A1 => n781, A2 => n780, A3 => n779, ZN => 
                           curr_proc_regs(353));
   U1252 : NAND2_X1 port map( A1 => regs(866), A2 => n54, ZN => n784);
   U1253 : AOI22_X1 port map( A1 => n17, A2 => regs(1378), B1 => n33, B2 => 
                           regs(354), ZN => n783);
   U1254 : AOI22_X1 port map( A1 => n116, A2 => regs(2402), B1 => n70, B2 => 
                           regs(1890), ZN => n782);
   U1255 : NAND3_X1 port map( A1 => n784, A2 => n783, A3 => n782, ZN => 
                           curr_proc_regs(354));
   U1256 : NAND2_X1 port map( A1 => regs(867), A2 => n51, ZN => n787);
   U1257 : AOI22_X1 port map( A1 => n93, A2 => regs(1379), B1 => n33, B2 => 
                           regs(355), ZN => n786);
   U1258 : AOI22_X1 port map( A1 => n116, A2 => regs(2403), B1 => n70, B2 => 
                           regs(1891), ZN => n785);
   U1259 : NAND3_X1 port map( A1 => n787, A2 => n786, A3 => n785, ZN => 
                           curr_proc_regs(355));
   U1260 : NAND2_X1 port map( A1 => regs(868), A2 => n49, ZN => n790);
   U1261 : AOI22_X1 port map( A1 => n17, A2 => regs(1380), B1 => n33, B2 => 
                           regs(356), ZN => n789);
   U1262 : AOI22_X1 port map( A1 => n116, A2 => regs(2404), B1 => n73, B2 => 
                           regs(1892), ZN => n788);
   U1263 : NAND3_X1 port map( A1 => n790, A2 => n789, A3 => n788, ZN => 
                           curr_proc_regs(356));
   U1264 : NAND2_X1 port map( A1 => regs(869), A2 => n61, ZN => n793);
   U1265 : AOI22_X1 port map( A1 => n89, A2 => regs(1381), B1 => n33, B2 => 
                           regs(357), ZN => n792);
   U1266 : AOI22_X1 port map( A1 => n116, A2 => regs(2405), B1 => n74, B2 => 
                           regs(1893), ZN => n791);
   U1267 : NAND3_X1 port map( A1 => n793, A2 => n792, A3 => n791, ZN => 
                           curr_proc_regs(357));
   U1268 : NAND2_X1 port map( A1 => regs(870), A2 => n10, ZN => n796);
   U1269 : AOI22_X1 port map( A1 => n95, A2 => regs(1382), B1 => n34, B2 => 
                           regs(358), ZN => n795);
   U1270 : AOI22_X1 port map( A1 => n116, A2 => regs(2406), B1 => n73, B2 => 
                           regs(1894), ZN => n794);
   U1271 : NAND3_X1 port map( A1 => n796, A2 => n795, A3 => n794, ZN => 
                           curr_proc_regs(358));
   U1272 : NAND2_X1 port map( A1 => regs(871), A2 => n10, ZN => n799);
   U1273 : AOI22_X1 port map( A1 => n95, A2 => regs(1383), B1 => n36, B2 => 
                           regs(359), ZN => n798);
   U1274 : AOI22_X1 port map( A1 => n116, A2 => regs(2407), B1 => n16, B2 => 
                           regs(1895), ZN => n797);
   U1275 : NAND3_X1 port map( A1 => n799, A2 => n798, A3 => n797, ZN => 
                           curr_proc_regs(359));
   U1276 : INV_X1 port map( A => regs(1059), ZN => n1402);
   U1277 : AOI22_X1 port map( A1 => n116, A2 => regs(2083), B1 => n16, B2 => 
                           regs(1571), ZN => n801);
   U1278 : AOI22_X1 port map( A1 => n51, A2 => regs(547), B1 => n36, B2 => 
                           regs(35), ZN => n800);
   U1279 : OAI211_X1 port map( C1 => n2199, C2 => n1402, A => n801, B => n800, 
                           ZN => curr_proc_regs(35));
   U1280 : NAND2_X1 port map( A1 => regs(872), A2 => n10, ZN => n804);
   U1281 : AOI22_X1 port map( A1 => n17, A2 => regs(1384), B1 => n35, B2 => 
                           regs(360), ZN => n803);
   U1282 : AOI22_X1 port map( A1 => n116, A2 => regs(2408), B1 => n78, B2 => 
                           regs(1896), ZN => n802);
   U1283 : NAND3_X1 port map( A1 => n804, A2 => n803, A3 => n802, ZN => 
                           curr_proc_regs(360));
   U1284 : NAND2_X1 port map( A1 => regs(1385), A2 => n98, ZN => n807);
   U1285 : AOI22_X1 port map( A1 => n49, A2 => regs(873), B1 => n36, B2 => 
                           regs(361), ZN => n806);
   U1286 : AOI22_X1 port map( A1 => n116, A2 => regs(2409), B1 => n3, B2 => 
                           regs(1897), ZN => n805);
   U1287 : NAND3_X1 port map( A1 => n807, A2 => n806, A3 => n805, ZN => 
                           curr_proc_regs(361));
   U1288 : NAND2_X1 port map( A1 => regs(1386), A2 => n84, ZN => n810);
   U1289 : AOI22_X1 port map( A1 => n51, A2 => regs(874), B1 => n35, B2 => 
                           regs(362), ZN => n809);
   U1290 : AOI22_X1 port map( A1 => n116, A2 => regs(2410), B1 => n3, B2 => 
                           regs(1898), ZN => n808);
   U1291 : NAND3_X1 port map( A1 => n810, A2 => n809, A3 => n808, ZN => 
                           curr_proc_regs(362));
   U1292 : NAND2_X1 port map( A1 => regs(875), A2 => n60, ZN => n813);
   U1293 : AOI22_X1 port map( A1 => n17, A2 => regs(1387), B1 => n34, B2 => 
                           regs(363), ZN => n812);
   U1294 : AOI22_X1 port map( A1 => n116, A2 => regs(2411), B1 => n3, B2 => 
                           regs(1899), ZN => n811);
   U1295 : NAND3_X1 port map( A1 => n813, A2 => n812, A3 => n811, ZN => 
                           curr_proc_regs(363));
   U1296 : NAND2_X1 port map( A1 => regs(876), A2 => n10, ZN => n816);
   U1297 : AOI22_X1 port map( A1 => n18, A2 => regs(1388), B1 => n34, B2 => 
                           regs(364), ZN => n815);
   U1298 : AOI22_X1 port map( A1 => n116, A2 => regs(2412), B1 => n73, B2 => 
                           regs(1900), ZN => n814);
   U1299 : NAND3_X1 port map( A1 => n816, A2 => n815, A3 => n814, ZN => 
                           curr_proc_regs(364));
   U1300 : NAND2_X1 port map( A1 => regs(877), A2 => n62, ZN => n819);
   U1301 : AOI22_X1 port map( A1 => n18, A2 => regs(1389), B1 => n35, B2 => 
                           regs(365), ZN => n818);
   U1302 : AOI22_X1 port map( A1 => n116, A2 => regs(2413), B1 => n71, B2 => 
                           regs(1901), ZN => n817);
   U1303 : NAND3_X1 port map( A1 => n819, A2 => n818, A3 => n817, ZN => 
                           curr_proc_regs(365));
   U1304 : NAND2_X1 port map( A1 => regs(1390), A2 => n86, ZN => n822);
   U1305 : AOI22_X1 port map( A1 => n51, A2 => regs(878), B1 => n36, B2 => 
                           regs(366), ZN => n821);
   U1306 : AOI22_X1 port map( A1 => n116, A2 => regs(2414), B1 => n68, B2 => 
                           regs(1902), ZN => n820);
   U1307 : NAND3_X1 port map( A1 => n822, A2 => n821, A3 => n820, ZN => 
                           curr_proc_regs(366));
   U1308 : NAND2_X1 port map( A1 => regs(1391), A2 => n98, ZN => n825);
   U1309 : AOI22_X1 port map( A1 => n50, A2 => regs(879), B1 => n35, B2 => 
                           regs(367), ZN => n824);
   U1310 : AOI22_X1 port map( A1 => n116, A2 => regs(2415), B1 => n73, B2 => 
                           regs(1903), ZN => n823);
   U1311 : NAND3_X1 port map( A1 => n825, A2 => n824, A3 => n823, ZN => 
                           curr_proc_regs(367));
   U1312 : NAND2_X1 port map( A1 => regs(1392), A2 => n14, ZN => n828);
   U1313 : AOI22_X1 port map( A1 => n50, A2 => regs(880), B1 => n34, B2 => 
                           regs(368), ZN => n827);
   U1314 : AOI22_X1 port map( A1 => n116, A2 => regs(2416), B1 => n74, B2 => 
                           regs(1904), ZN => n826);
   U1315 : NAND3_X1 port map( A1 => n828, A2 => n827, A3 => n826, ZN => 
                           curr_proc_regs(368));
   U1316 : NAND2_X1 port map( A1 => regs(1393), A2 => n14, ZN => n831);
   U1317 : AOI22_X1 port map( A1 => n49, A2 => regs(881), B1 => n36, B2 => 
                           regs(369), ZN => n830);
   U1318 : AOI22_X1 port map( A1 => n116, A2 => regs(2417), B1 => n68, B2 => 
                           regs(1905), ZN => n829);
   U1319 : NAND3_X1 port map( A1 => n831, A2 => n830, A3 => n829, ZN => 
                           curr_proc_regs(369));
   U1320 : INV_X1 port map( A => regs(1060), ZN => n1405);
   U1321 : AOI22_X1 port map( A1 => n116, A2 => regs(2084), B1 => n73, B2 => 
                           regs(1572), ZN => n833);
   U1322 : AOI22_X1 port map( A1 => n56, A2 => regs(548), B1 => n35, B2 => 
                           regs(36), ZN => n832);
   U1323 : OAI211_X1 port map( C1 => n99, C2 => n1405, A => n833, B => n832, ZN
                           => curr_proc_regs(36));
   U1324 : NAND2_X1 port map( A1 => regs(1394), A2 => n14, ZN => n836);
   U1325 : AOI22_X1 port map( A1 => n50, A2 => regs(882), B1 => n34, B2 => 
                           regs(370), ZN => n835);
   U1326 : AOI22_X1 port map( A1 => n116, A2 => regs(2418), B1 => n73, B2 => 
                           regs(1906), ZN => n834);
   U1327 : NAND3_X1 port map( A1 => n836, A2 => n835, A3 => n834, ZN => 
                           curr_proc_regs(370));
   U1328 : NAND2_X1 port map( A1 => regs(883), A2 => n49, ZN => n839);
   U1329 : AOI22_X1 port map( A1 => n17, A2 => regs(1395), B1 => n35, B2 => 
                           regs(371), ZN => n838);
   U1330 : AOI22_X1 port map( A1 => n116, A2 => regs(2419), B1 => n70, B2 => 
                           regs(1907), ZN => n837);
   U1331 : NAND3_X1 port map( A1 => n839, A2 => n838, A3 => n837, ZN => 
                           curr_proc_regs(371));
   U1332 : NAND2_X1 port map( A1 => regs(1396), A2 => n14, ZN => n842);
   U1333 : AOI22_X1 port map( A1 => n50, A2 => regs(884), B1 => n36, B2 => 
                           regs(372), ZN => n841);
   U1334 : AOI22_X1 port map( A1 => n116, A2 => regs(2420), B1 => n74, B2 => 
                           regs(1908), ZN => n840);
   U1335 : NAND3_X1 port map( A1 => n842, A2 => n841, A3 => n840, ZN => 
                           curr_proc_regs(372));
   U1336 : NAND2_X1 port map( A1 => regs(885), A2 => n10, ZN => n845);
   U1337 : AOI22_X1 port map( A1 => n17, A2 => regs(1397), B1 => n35, B2 => 
                           regs(373), ZN => n844);
   U1338 : AOI22_X1 port map( A1 => n116, A2 => regs(2421), B1 => n16, B2 => 
                           regs(1909), ZN => n843);
   U1339 : NAND3_X1 port map( A1 => n845, A2 => n844, A3 => n843, ZN => 
                           curr_proc_regs(373));
   U1340 : NAND2_X1 port map( A1 => regs(886), A2 => n10, ZN => n848);
   U1341 : AOI22_X1 port map( A1 => n17, A2 => regs(1398), B1 => n34, B2 => 
                           regs(374), ZN => n847);
   U1342 : AOI22_X1 port map( A1 => n116, A2 => regs(2422), B1 => n74, B2 => 
                           regs(1910), ZN => n846);
   U1343 : NAND3_X1 port map( A1 => n848, A2 => n847, A3 => n846, ZN => 
                           curr_proc_regs(374));
   U1344 : NAND2_X1 port map( A1 => regs(887), A2 => n62, ZN => n851);
   U1345 : AOI22_X1 port map( A1 => n18, A2 => regs(1399), B1 => n34, B2 => 
                           regs(375), ZN => n850);
   U1346 : AOI22_X1 port map( A1 => n116, A2 => regs(2423), B1 => n16, B2 => 
                           regs(1911), ZN => n849);
   U1347 : NAND3_X1 port map( A1 => n851, A2 => n850, A3 => n849, ZN => 
                           curr_proc_regs(375));
   U1348 : NAND2_X1 port map( A1 => regs(1400), A2 => n14, ZN => n854);
   U1349 : AOI22_X1 port map( A1 => n49, A2 => regs(888), B1 => n36, B2 => 
                           regs(376), ZN => n853);
   U1350 : AOI22_X1 port map( A1 => n116, A2 => regs(2424), B1 => n70, B2 => 
                           regs(1912), ZN => n852);
   U1351 : NAND3_X1 port map( A1 => n854, A2 => n853, A3 => n852, ZN => 
                           curr_proc_regs(376));
   U1352 : NAND2_X1 port map( A1 => regs(889), A2 => n62, ZN => n857);
   U1353 : AOI22_X1 port map( A1 => n17, A2 => regs(1401), B1 => n35, B2 => 
                           regs(377), ZN => n856);
   U1354 : AOI22_X1 port map( A1 => n116, A2 => regs(2425), B1 => n70, B2 => 
                           regs(1913), ZN => n855);
   U1355 : NAND3_X1 port map( A1 => n857, A2 => n856, A3 => n855, ZN => 
                           curr_proc_regs(377));
   U1356 : NAND2_X1 port map( A1 => regs(890), A2 => n10, ZN => n860);
   U1357 : AOI22_X1 port map( A1 => n18, A2 => regs(1402), B1 => n34, B2 => 
                           regs(378), ZN => n859);
   U1358 : AOI22_X1 port map( A1 => n116, A2 => regs(2426), B1 => n16, B2 => 
                           regs(1914), ZN => n858);
   U1359 : NAND3_X1 port map( A1 => n860, A2 => n859, A3 => n858, ZN => 
                           curr_proc_regs(378));
   U1360 : NAND2_X1 port map( A1 => regs(1403), A2 => n14, ZN => n863);
   U1361 : AOI22_X1 port map( A1 => n51, A2 => regs(891), B1 => n34, B2 => 
                           regs(379), ZN => n862);
   U1362 : AOI22_X1 port map( A1 => n116, A2 => regs(2427), B1 => n16, B2 => 
                           regs(1915), ZN => n861);
   U1363 : NAND3_X1 port map( A1 => n863, A2 => n862, A3 => n861, ZN => 
                           curr_proc_regs(379));
   U1364 : INV_X1 port map( A => regs(549), ZN => n1408);
   U1365 : AOI22_X1 port map( A1 => n116, A2 => regs(2085), B1 => n9, B2 => 
                           regs(1573), ZN => n865);
   U1366 : AOI22_X1 port map( A1 => n93, A2 => regs(1061), B1 => n34, B2 => 
                           regs(37), ZN => n864);
   U1367 : OAI211_X1 port map( C1 => n2185, C2 => n1408, A => n865, B => n864, 
                           ZN => curr_proc_regs(37));
   U1368 : NAND2_X1 port map( A1 => regs(1404), A2 => n14, ZN => n868);
   U1369 : AOI22_X1 port map( A1 => n51, A2 => regs(892), B1 => n34, B2 => 
                           regs(380), ZN => n867);
   U1370 : AOI22_X1 port map( A1 => n116, A2 => regs(2428), B1 => n3, B2 => 
                           regs(1916), ZN => n866);
   U1371 : NAND3_X1 port map( A1 => n868, A2 => n867, A3 => n866, ZN => 
                           curr_proc_regs(380));
   U1372 : NAND2_X1 port map( A1 => regs(893), A2 => n54, ZN => n871);
   U1373 : AOI22_X1 port map( A1 => n89, A2 => regs(1405), B1 => n35, B2 => 
                           regs(381), ZN => n870);
   U1374 : AOI22_X1 port map( A1 => n116, A2 => regs(2429), B1 => n3, B2 => 
                           regs(1917), ZN => n869);
   U1375 : NAND3_X1 port map( A1 => n871, A2 => n870, A3 => n869, ZN => 
                           curr_proc_regs(381));
   U1376 : NAND2_X1 port map( A1 => regs(1406), A2 => n17, ZN => n874);
   U1377 : AOI22_X1 port map( A1 => n48, A2 => regs(894), B1 => n34, B2 => 
                           regs(382), ZN => n873);
   U1378 : AOI22_X1 port map( A1 => n116, A2 => regs(2430), B1 => n3, B2 => 
                           regs(1918), ZN => n872);
   U1379 : NAND3_X1 port map( A1 => n874, A2 => n873, A3 => n872, ZN => 
                           curr_proc_regs(382));
   U1380 : NAND2_X1 port map( A1 => regs(895), A2 => n59, ZN => n877);
   U1381 : AOI22_X1 port map( A1 => n82, A2 => regs(1407), B1 => n36, B2 => 
                           regs(383), ZN => n876);
   U1382 : AOI22_X1 port map( A1 => n116, A2 => regs(2431), B1 => n3, B2 => 
                           regs(1919), ZN => n875);
   U1383 : NAND3_X1 port map( A1 => n877, A2 => n876, A3 => n875, ZN => 
                           curr_proc_regs(383));
   U1384 : NAND2_X1 port map( A1 => regs(1408), A2 => n96, ZN => n880);
   U1385 : AOI22_X1 port map( A1 => n50, A2 => regs(896), B1 => n35, B2 => 
                           regs(384), ZN => n879);
   U1386 : AOI22_X1 port map( A1 => n116, A2 => regs(2432), B1 => n71, B2 => 
                           regs(1920), ZN => n878);
   U1387 : NAND3_X1 port map( A1 => n880, A2 => n879, A3 => n878, ZN => 
                           curr_proc_regs(384));
   U1388 : NAND2_X1 port map( A1 => regs(897), A2 => n63, ZN => n883);
   U1389 : AOI22_X1 port map( A1 => n82, A2 => regs(1409), B1 => n34, B2 => 
                           regs(385), ZN => n882);
   U1390 : AOI22_X1 port map( A1 => n116, A2 => regs(2433), B1 => n68, B2 => 
                           regs(1921), ZN => n881);
   U1391 : NAND3_X1 port map( A1 => n883, A2 => n882, A3 => n881, ZN => 
                           curr_proc_regs(385));
   U1392 : NAND2_X1 port map( A1 => regs(898), A2 => n63, ZN => n886);
   U1393 : AOI22_X1 port map( A1 => n82, A2 => regs(1410), B1 => n36, B2 => 
                           regs(386), ZN => n885);
   U1394 : AOI22_X1 port map( A1 => n116, A2 => regs(2434), B1 => n73, B2 => 
                           regs(1922), ZN => n884);
   U1395 : NAND3_X1 port map( A1 => n886, A2 => n885, A3 => n884, ZN => 
                           curr_proc_regs(386));
   U1396 : NAND2_X1 port map( A1 => regs(899), A2 => n63, ZN => n889);
   U1397 : AOI22_X1 port map( A1 => n82, A2 => regs(1411), B1 => n35, B2 => 
                           regs(387), ZN => n888);
   U1398 : AOI22_X1 port map( A1 => n116, A2 => regs(2435), B1 => n16, B2 => 
                           regs(1923), ZN => n887);
   U1399 : NAND3_X1 port map( A1 => n889, A2 => n888, A3 => n887, ZN => 
                           curr_proc_regs(387));
   U1400 : NAND2_X1 port map( A1 => regs(1412), A2 => n14, ZN => n892);
   U1401 : AOI22_X1 port map( A1 => n53, A2 => regs(900), B1 => n35, B2 => 
                           regs(388), ZN => n891);
   U1402 : AOI22_X1 port map( A1 => n116, A2 => regs(2436), B1 => n73, B2 => 
                           regs(1924), ZN => n890);
   U1403 : NAND3_X1 port map( A1 => n892, A2 => n891, A3 => n890, ZN => 
                           curr_proc_regs(388));
   U1404 : NAND2_X1 port map( A1 => regs(1413), A2 => n14, ZN => n895);
   U1405 : AOI22_X1 port map( A1 => n50, A2 => regs(901), B1 => n35, B2 => 
                           regs(389), ZN => n894);
   U1406 : AOI22_X1 port map( A1 => n116, A2 => regs(2437), B1 => n73, B2 => 
                           regs(1925), ZN => n893);
   U1407 : NAND3_X1 port map( A1 => n895, A2 => n894, A3 => n893, ZN => 
                           curr_proc_regs(389));
   U1408 : INV_X1 port map( A => regs(550), ZN => n1413);
   U1409 : AOI22_X1 port map( A1 => n116, A2 => regs(2086), B1 => n73, B2 => 
                           regs(1574), ZN => n897);
   U1410 : AOI22_X1 port map( A1 => n82, A2 => regs(1062), B1 => n35, B2 => 
                           regs(38), ZN => n896);
   U1411 : OAI211_X1 port map( C1 => n65, C2 => n1413, A => n897, B => n896, ZN
                           => curr_proc_regs(38));
   U1412 : NAND2_X1 port map( A1 => regs(1414), A2 => n97, ZN => n900);
   U1413 : AOI22_X1 port map( A1 => n49, A2 => regs(902), B1 => n35, B2 => 
                           regs(390), ZN => n899);
   U1414 : AOI22_X1 port map( A1 => n116, A2 => regs(2438), B1 => n16, B2 => 
                           regs(1926), ZN => n898);
   U1415 : NAND3_X1 port map( A1 => n900, A2 => n899, A3 => n898, ZN => 
                           curr_proc_regs(390));
   U1416 : NAND2_X1 port map( A1 => regs(903), A2 => n63, ZN => n903);
   U1417 : AOI22_X1 port map( A1 => n82, A2 => regs(1415), B1 => n34, B2 => 
                           regs(391), ZN => n902);
   U1418 : AOI22_X1 port map( A1 => n116, A2 => regs(2439), B1 => n73, B2 => 
                           regs(1927), ZN => n901);
   U1419 : NAND3_X1 port map( A1 => n903, A2 => n902, A3 => n901, ZN => 
                           curr_proc_regs(391));
   U1420 : NAND2_X1 port map( A1 => regs(904), A2 => n62, ZN => n906);
   U1421 : AOI22_X1 port map( A1 => n82, A2 => regs(1416), B1 => n34, B2 => 
                           regs(392), ZN => n905);
   U1422 : AOI22_X1 port map( A1 => n116, A2 => regs(2440), B1 => n16, B2 => 
                           regs(1928), ZN => n904);
   U1423 : NAND3_X1 port map( A1 => n906, A2 => n905, A3 => n904, ZN => 
                           curr_proc_regs(392));
   U1424 : NAND2_X1 port map( A1 => regs(905), A2 => n63, ZN => n909);
   U1425 : AOI22_X1 port map( A1 => n82, A2 => regs(1417), B1 => n34, B2 => 
                           regs(393), ZN => n908);
   U1426 : AOI22_X1 port map( A1 => n116, A2 => regs(2441), B1 => n73, B2 => 
                           regs(1929), ZN => n907);
   U1427 : NAND3_X1 port map( A1 => n909, A2 => n908, A3 => n907, ZN => 
                           curr_proc_regs(393));
   U1428 : NAND2_X1 port map( A1 => regs(1418), A2 => n14, ZN => n912);
   U1429 : AOI22_X1 port map( A1 => n61, A2 => regs(906), B1 => n34, B2 => 
                           regs(394), ZN => n911);
   U1430 : AOI22_X1 port map( A1 => n116, A2 => regs(2442), B1 => n74, B2 => 
                           regs(1930), ZN => n910);
   U1431 : NAND3_X1 port map( A1 => n912, A2 => n911, A3 => n910, ZN => 
                           curr_proc_regs(394));
   U1432 : NAND2_X1 port map( A1 => regs(907), A2 => n60, ZN => n915);
   U1433 : AOI22_X1 port map( A1 => n82, A2 => regs(1419), B1 => n34, B2 => 
                           regs(395), ZN => n914);
   U1434 : AOI22_X1 port map( A1 => n116, A2 => regs(2443), B1 => n3, B2 => 
                           regs(1931), ZN => n913);
   U1435 : NAND3_X1 port map( A1 => n915, A2 => n914, A3 => n913, ZN => 
                           curr_proc_regs(395));
   U1436 : NAND2_X1 port map( A1 => regs(908), A2 => n48, ZN => n918);
   U1437 : AOI22_X1 port map( A1 => n82, A2 => regs(1420), B1 => n34, B2 => 
                           regs(396), ZN => n917);
   U1438 : AOI22_X1 port map( A1 => n116, A2 => regs(2444), B1 => n73, B2 => 
                           regs(1932), ZN => n916);
   U1439 : NAND3_X1 port map( A1 => n918, A2 => n917, A3 => n916, ZN => 
                           curr_proc_regs(396));
   U1440 : NAND2_X1 port map( A1 => regs(909), A2 => n63, ZN => n921);
   U1441 : AOI22_X1 port map( A1 => n98, A2 => regs(1421), B1 => n34, B2 => 
                           regs(397), ZN => n920);
   U1442 : AOI22_X1 port map( A1 => n116, A2 => regs(2445), B1 => n3, B2 => 
                           regs(1933), ZN => n919);
   U1443 : NAND3_X1 port map( A1 => n921, A2 => n920, A3 => n919, ZN => 
                           curr_proc_regs(397));
   U1444 : NAND2_X1 port map( A1 => regs(910), A2 => n62, ZN => n924);
   U1445 : AOI22_X1 port map( A1 => n18, A2 => regs(1422), B1 => n36, B2 => 
                           regs(398), ZN => n923);
   U1446 : AOI22_X1 port map( A1 => n116, A2 => regs(2446), B1 => n74, B2 => 
                           regs(1934), ZN => n922);
   U1447 : NAND3_X1 port map( A1 => n924, A2 => n923, A3 => n922, ZN => 
                           curr_proc_regs(398));
   U1448 : NAND2_X1 port map( A1 => regs(1423), A2 => n14, ZN => n927);
   U1449 : AOI22_X1 port map( A1 => n60, A2 => regs(911), B1 => n36, B2 => 
                           regs(399), ZN => n926);
   U1450 : AOI22_X1 port map( A1 => n116, A2 => regs(2447), B1 => n74, B2 => 
                           regs(1935), ZN => n925);
   U1451 : NAND3_X1 port map( A1 => n927, A2 => n926, A3 => n925, ZN => 
                           curr_proc_regs(399));
   U1452 : INV_X1 port map( A => regs(551), ZN => n1416);
   U1453 : AOI22_X1 port map( A1 => n116, A2 => regs(2087), B1 => n74, B2 => 
                           regs(1575), ZN => n929);
   U1454 : AOI22_X1 port map( A1 => n90, A2 => regs(1063), B1 => n36, B2 => 
                           regs(39), ZN => n928);
   U1455 : OAI211_X1 port map( C1 => n6, C2 => n1416, A => n929, B => n928, ZN 
                           => curr_proc_regs(39));
   U1456 : INV_X1 port map( A => regs(515), ZN => n1303);
   U1457 : AOI22_X1 port map( A1 => n116, A2 => regs(2051), B1 => n74, B2 => 
                           regs(1539), ZN => n931);
   U1458 : AOI22_X1 port map( A1 => n80, A2 => regs(1027), B1 => n36, B2 => 
                           regs(3), ZN => n930);
   U1459 : OAI211_X1 port map( C1 => n2185, C2 => n1303, A => n931, B => n930, 
                           ZN => curr_proc_regs(3));
   U1460 : NAND2_X1 port map( A1 => regs(912), A2 => n63, ZN => n934);
   U1461 : AOI22_X1 port map( A1 => n96, A2 => regs(1424), B1 => n35, B2 => 
                           regs(400), ZN => n933);
   U1462 : AOI22_X1 port map( A1 => n116, A2 => regs(2448), B1 => n74, B2 => 
                           regs(1936), ZN => n932);
   U1463 : NAND3_X1 port map( A1 => n934, A2 => n933, A3 => n932, ZN => 
                           curr_proc_regs(400));
   U1464 : NAND2_X1 port map( A1 => regs(913), A2 => n58, ZN => n937);
   U1465 : AOI22_X1 port map( A1 => n96, A2 => regs(1425), B1 => n35, B2 => 
                           regs(401), ZN => n936);
   U1466 : AOI22_X1 port map( A1 => n116, A2 => regs(2449), B1 => n74, B2 => 
                           regs(1937), ZN => n935);
   U1467 : NAND3_X1 port map( A1 => n937, A2 => n936, A3 => n935, ZN => 
                           curr_proc_regs(401));
   U1468 : NAND2_X1 port map( A1 => regs(1426), A2 => n14, ZN => n940);
   U1469 : AOI22_X1 port map( A1 => n61, A2 => regs(914), B1 => n35, B2 => 
                           regs(402), ZN => n939);
   U1470 : AOI22_X1 port map( A1 => n116, A2 => regs(2450), B1 => n74, B2 => 
                           regs(1938), ZN => n938);
   U1471 : NAND3_X1 port map( A1 => n940, A2 => n939, A3 => n938, ZN => 
                           curr_proc_regs(402));
   U1472 : NAND2_X1 port map( A1 => regs(1427), A2 => n85, ZN => n943);
   U1473 : AOI22_X1 port map( A1 => n60, A2 => regs(915), B1 => n35, B2 => 
                           regs(403), ZN => n942);
   U1474 : AOI22_X1 port map( A1 => n116, A2 => regs(2451), B1 => n74, B2 => 
                           regs(1939), ZN => n941);
   U1475 : NAND3_X1 port map( A1 => n943, A2 => n942, A3 => n941, ZN => 
                           curr_proc_regs(403));
   U1476 : NAND2_X1 port map( A1 => regs(1428), A2 => n14, ZN => n946);
   U1477 : AOI22_X1 port map( A1 => n61, A2 => regs(916), B1 => n35, B2 => 
                           regs(404), ZN => n945);
   U1478 : AOI22_X1 port map( A1 => n116, A2 => regs(2452), B1 => n74, B2 => 
                           regs(1940), ZN => n944);
   U1479 : NAND3_X1 port map( A1 => n946, A2 => n945, A3 => n944, ZN => 
                           curr_proc_regs(404));
   U1480 : NAND2_X1 port map( A1 => regs(917), A2 => n63, ZN => n949);
   U1481 : AOI22_X1 port map( A1 => n95, A2 => regs(1429), B1 => n35, B2 => 
                           regs(405), ZN => n948);
   U1482 : AOI22_X1 port map( A1 => n116, A2 => regs(2453), B1 => n74, B2 => 
                           regs(1941), ZN => n947);
   U1483 : NAND3_X1 port map( A1 => n949, A2 => n948, A3 => n947, ZN => 
                           curr_proc_regs(405));
   U1484 : NAND2_X1 port map( A1 => regs(1430), A2 => n14, ZN => n952);
   U1485 : AOI22_X1 port map( A1 => n60, A2 => regs(918), B1 => n35, B2 => 
                           regs(406), ZN => n951);
   U1486 : AOI22_X1 port map( A1 => n116, A2 => regs(2454), B1 => n74, B2 => 
                           regs(1942), ZN => n950);
   U1487 : NAND3_X1 port map( A1 => n952, A2 => n951, A3 => n950, ZN => 
                           curr_proc_regs(406));
   U1488 : NAND2_X1 port map( A1 => regs(919), A2 => n62, ZN => n955);
   U1489 : AOI22_X1 port map( A1 => n81, A2 => regs(1431), B1 => n38, B2 => 
                           regs(407), ZN => n954);
   U1490 : AOI22_X1 port map( A1 => n116, A2 => regs(2455), B1 => n68, B2 => 
                           regs(1943), ZN => n953);
   U1491 : NAND3_X1 port map( A1 => n955, A2 => n954, A3 => n953, ZN => 
                           curr_proc_regs(407));
   U1492 : NAND2_X1 port map( A1 => regs(1432), A2 => n88, ZN => n958);
   U1493 : AOI22_X1 port map( A1 => n61, A2 => regs(920), B1 => n41, B2 => 
                           regs(408), ZN => n957);
   U1494 : AOI22_X1 port map( A1 => n116, A2 => regs(2456), B1 => n73, B2 => 
                           regs(1944), ZN => n956);
   U1495 : NAND3_X1 port map( A1 => n958, A2 => n957, A3 => n956, ZN => 
                           curr_proc_regs(408));
   U1496 : NAND2_X1 port map( A1 => regs(921), A2 => n10, ZN => n961);
   U1497 : AOI22_X1 port map( A1 => n81, A2 => regs(1433), B1 => n45, B2 => 
                           regs(409), ZN => n960);
   U1498 : AOI22_X1 port map( A1 => n116, A2 => regs(2457), B1 => n16, B2 => 
                           regs(1945), ZN => n959);
   U1499 : NAND3_X1 port map( A1 => n961, A2 => n960, A3 => n959, ZN => 
                           curr_proc_regs(409));
   U1500 : INV_X1 port map( A => regs(552), ZN => n1419);
   U1501 : AOI22_X1 port map( A1 => n116, A2 => regs(2088), B1 => n16, B2 => 
                           regs(1576), ZN => n963);
   U1502 : AOI22_X1 port map( A1 => n82, A2 => regs(1064), B1 => n44, B2 => 
                           regs(40), ZN => n962);
   U1503 : OAI211_X1 port map( C1 => n64, C2 => n1419, A => n963, B => n962, ZN
                           => curr_proc_regs(40));
   U1504 : NAND2_X1 port map( A1 => regs(1434), A2 => n79, ZN => n966);
   U1505 : AOI22_X1 port map( A1 => n8, A2 => regs(922), B1 => n36, B2 => 
                           regs(410), ZN => n965);
   U1506 : AOI22_X1 port map( A1 => n116, A2 => regs(2458), B1 => n69, B2 => 
                           regs(1946), ZN => n964);
   U1507 : NAND3_X1 port map( A1 => n966, A2 => n965, A3 => n964, ZN => 
                           curr_proc_regs(410));
   U1508 : NAND2_X1 port map( A1 => regs(1435), A2 => n84, ZN => n969);
   U1509 : AOI22_X1 port map( A1 => n8, A2 => regs(923), B1 => n36, B2 => 
                           regs(411), ZN => n968);
   U1510 : AOI22_X1 port map( A1 => n116, A2 => regs(2459), B1 => n3, B2 => 
                           regs(1947), ZN => n967);
   U1511 : NAND3_X1 port map( A1 => n969, A2 => n968, A3 => n967, ZN => 
                           curr_proc_regs(411));
   U1512 : NAND2_X1 port map( A1 => regs(924), A2 => n10, ZN => n972);
   U1513 : AOI22_X1 port map( A1 => n83, A2 => regs(1436), B1 => n36, B2 => 
                           regs(412), ZN => n971);
   U1514 : AOI22_X1 port map( A1 => n116, A2 => regs(2460), B1 => n3, B2 => 
                           regs(1948), ZN => n970);
   U1515 : NAND3_X1 port map( A1 => n972, A2 => n971, A3 => n970, ZN => 
                           curr_proc_regs(412));
   U1516 : NAND2_X1 port map( A1 => regs(1437), A2 => n86, ZN => n975);
   U1517 : AOI22_X1 port map( A1 => n57, A2 => regs(925), B1 => n36, B2 => 
                           regs(413), ZN => n974);
   U1518 : AOI22_X1 port map( A1 => n116, A2 => regs(2461), B1 => n3, B2 => 
                           regs(1949), ZN => n973);
   U1519 : NAND3_X1 port map( A1 => n975, A2 => n974, A3 => n973, ZN => 
                           curr_proc_regs(413));
   U1520 : NAND2_X1 port map( A1 => regs(1438), A2 => n80, ZN => n978);
   U1521 : AOI22_X1 port map( A1 => n61, A2 => regs(926), B1 => n36, B2 => 
                           regs(414), ZN => n977);
   U1522 : AOI22_X1 port map( A1 => n116, A2 => regs(2462), B1 => n71, B2 => 
                           regs(1950), ZN => n976);
   U1523 : NAND3_X1 port map( A1 => n978, A2 => n977, A3 => n976, ZN => 
                           curr_proc_regs(414));
   U1524 : NAND2_X1 port map( A1 => regs(927), A2 => n5, ZN => n981);
   U1525 : AOI22_X1 port map( A1 => n95, A2 => regs(1439), B1 => n36, B2 => 
                           regs(415), ZN => n980);
   U1526 : AOI22_X1 port map( A1 => n116, A2 => regs(2463), B1 => n71, B2 => 
                           regs(1951), ZN => n979);
   U1527 : NAND3_X1 port map( A1 => n981, A2 => n980, A3 => n979, ZN => 
                           curr_proc_regs(415));
   U1528 : NAND2_X1 port map( A1 => regs(1440), A2 => n95, ZN => n984);
   U1529 : AOI22_X1 port map( A1 => n61, A2 => regs(928), B1 => n36, B2 => 
                           regs(416), ZN => n983);
   U1530 : AOI22_X1 port map( A1 => n116, A2 => regs(2464), B1 => n68, B2 => 
                           regs(1952), ZN => n982);
   U1531 : NAND3_X1 port map( A1 => n984, A2 => n983, A3 => n982, ZN => 
                           curr_proc_regs(416));
   U1532 : NAND2_X1 port map( A1 => regs(929), A2 => n62, ZN => n987);
   U1533 : AOI22_X1 port map( A1 => n84, A2 => regs(1441), B1 => n24, B2 => 
                           regs(417), ZN => n986);
   U1534 : AOI22_X1 port map( A1 => n116, A2 => regs(2465), B1 => n16, B2 => 
                           regs(1953), ZN => n985);
   U1535 : NAND3_X1 port map( A1 => n987, A2 => n986, A3 => n985, ZN => 
                           curr_proc_regs(417));
   U1536 : NAND2_X1 port map( A1 => regs(1442), A2 => n91, ZN => n990);
   U1537 : AOI22_X1 port map( A1 => n62, A2 => regs(930), B1 => n23, B2 => 
                           regs(418), ZN => n989);
   U1538 : AOI22_X1 port map( A1 => n116, A2 => regs(2466), B1 => n77, B2 => 
                           regs(1954), ZN => n988);
   U1539 : NAND3_X1 port map( A1 => n990, A2 => n989, A3 => n988, ZN => 
                           curr_proc_regs(418));
   U1540 : NAND2_X1 port map( A1 => regs(1443), A2 => n85, ZN => n993);
   U1541 : AOI22_X1 port map( A1 => n61, A2 => regs(931), B1 => n24, B2 => 
                           regs(419), ZN => n992);
   U1542 : AOI22_X1 port map( A1 => n116, A2 => regs(2467), B1 => n3, B2 => 
                           regs(1955), ZN => n991);
   U1543 : NAND3_X1 port map( A1 => n993, A2 => n992, A3 => n991, ZN => 
                           curr_proc_regs(419));
   U1544 : INV_X1 port map( A => regs(1065), ZN => n1422);
   U1545 : AOI22_X1 port map( A1 => n116, A2 => regs(2089), B1 => n3, B2 => 
                           regs(1577), ZN => n995);
   U1546 : AOI22_X1 port map( A1 => n62, A2 => regs(553), B1 => n34, B2 => 
                           regs(41), ZN => n994);
   U1547 : OAI211_X1 port map( C1 => n15, C2 => n1422, A => n995, B => n994, ZN
                           => curr_proc_regs(41));
   U1548 : NAND2_X1 port map( A1 => regs(1444), A2 => n82, ZN => n998);
   U1549 : AOI22_X1 port map( A1 => n60, A2 => regs(932), B1 => n35, B2 => 
                           regs(420), ZN => n997);
   U1550 : AOI22_X1 port map( A1 => n116, A2 => regs(2468), B1 => n3, B2 => 
                           regs(1956), ZN => n996);
   U1551 : NAND3_X1 port map( A1 => n998, A2 => n997, A3 => n996, ZN => 
                           curr_proc_regs(420));
   U1552 : NAND2_X1 port map( A1 => regs(933), A2 => n10, ZN => n1001);
   U1553 : AOI22_X1 port map( A1 => n85, A2 => regs(1445), B1 => n34, B2 => 
                           regs(421), ZN => n1000);
   U1554 : AOI22_X1 port map( A1 => n116, A2 => regs(2469), B1 => n71, B2 => 
                           regs(1957), ZN => n999);
   U1555 : NAND3_X1 port map( A1 => n1001, A2 => n1000, A3 => n999, ZN => 
                           curr_proc_regs(421));
   U1556 : NAND2_X1 port map( A1 => regs(1446), A2 => n96, ZN => n1004);
   U1557 : AOI22_X1 port map( A1 => n62, A2 => regs(934), B1 => n39, B2 => 
                           regs(422), ZN => n1003);
   U1558 : AOI22_X1 port map( A1 => n116, A2 => regs(2470), B1 => n71, B2 => 
                           regs(1958), ZN => n1002);
   U1559 : NAND3_X1 port map( A1 => n1004, A2 => n1003, A3 => n1002, ZN => 
                           curr_proc_regs(422));
   U1560 : NAND2_X1 port map( A1 => regs(1447), A2 => n96, ZN => n1007);
   U1561 : AOI22_X1 port map( A1 => n61, A2 => regs(935), B1 => n24, B2 => 
                           regs(423), ZN => n1006);
   U1562 : AOI22_X1 port map( A1 => n116, A2 => regs(2471), B1 => n68, B2 => 
                           regs(1959), ZN => n1005);
   U1563 : NAND3_X1 port map( A1 => n1007, A2 => n1006, A3 => n1005, ZN => 
                           curr_proc_regs(423));
   U1564 : NAND2_X1 port map( A1 => regs(1448), A2 => n96, ZN => n1010);
   U1565 : AOI22_X1 port map( A1 => n54, A2 => regs(936), B1 => n23, B2 => 
                           regs(424), ZN => n1009);
   U1566 : AOI22_X1 port map( A1 => n116, A2 => regs(2472), B1 => n73, B2 => 
                           regs(1960), ZN => n1008);
   U1567 : NAND3_X1 port map( A1 => n1010, A2 => n1009, A3 => n1008, ZN => 
                           curr_proc_regs(424));
   U1568 : NAND2_X1 port map( A1 => regs(1449), A2 => n96, ZN => n1013);
   U1569 : AOI22_X1 port map( A1 => n52, A2 => regs(937), B1 => n25, B2 => 
                           regs(425), ZN => n1012);
   U1570 : AOI22_X1 port map( A1 => n116, A2 => regs(2473), B1 => n3, B2 => 
                           regs(1961), ZN => n1011);
   U1571 : NAND3_X1 port map( A1 => n1013, A2 => n1012, A3 => n1011, ZN => 
                           curr_proc_regs(425));
   U1572 : NAND2_X1 port map( A1 => regs(938), A2 => n10, ZN => n1016);
   U1573 : AOI22_X1 port map( A1 => n86, A2 => regs(1450), B1 => n42, B2 => 
                           regs(426), ZN => n1015);
   U1574 : AOI22_X1 port map( A1 => n116, A2 => regs(2474), B1 => n73, B2 => 
                           regs(1962), ZN => n1014);
   U1575 : NAND3_X1 port map( A1 => n1016, A2 => n1015, A3 => n1014, ZN => 
                           curr_proc_regs(426));
   U1576 : NAND2_X1 port map( A1 => regs(1451), A2 => n94, ZN => n1019);
   U1577 : AOI22_X1 port map( A1 => n53, A2 => regs(939), B1 => n28, B2 => 
                           regs(427), ZN => n1018);
   U1578 : AOI22_X1 port map( A1 => n116, A2 => regs(2475), B1 => n74, B2 => 
                           regs(1963), ZN => n1017);
   U1579 : NAND3_X1 port map( A1 => n1019, A2 => n1018, A3 => n1017, ZN => 
                           curr_proc_regs(427));
   U1580 : NAND2_X1 port map( A1 => regs(1452), A2 => n95, ZN => n1022);
   U1581 : AOI22_X1 port map( A1 => n55, A2 => regs(940), B1 => n27, B2 => 
                           regs(428), ZN => n1021);
   U1582 : AOI22_X1 port map( A1 => n116, A2 => regs(2476), B1 => n3, B2 => 
                           regs(1964), ZN => n1020);
   U1583 : NAND3_X1 port map( A1 => n1022, A2 => n1021, A3 => n1020, ZN => 
                           curr_proc_regs(428));
   U1584 : NAND2_X1 port map( A1 => regs(941), A2 => n56, ZN => n1025);
   U1585 : AOI22_X1 port map( A1 => n87, A2 => regs(1453), B1 => n26, B2 => 
                           regs(429), ZN => n1024);
   U1586 : AOI22_X1 port map( A1 => n116, A2 => regs(2477), B1 => n70, B2 => 
                           regs(1965), ZN => n1023);
   U1587 : NAND3_X1 port map( A1 => n1025, A2 => n1024, A3 => n1023, ZN => 
                           curr_proc_regs(429));
   U1588 : INV_X1 port map( A => regs(1066), ZN => n1425);
   U1589 : AOI22_X1 port map( A1 => n116, A2 => regs(2090), B1 => n70, B2 => 
                           regs(1578), ZN => n1027);
   U1590 : AOI22_X1 port map( A1 => n48, A2 => regs(554), B1 => n32, B2 => 
                           regs(42), ZN => n1026);
   U1591 : OAI211_X1 port map( C1 => n102, C2 => n1425, A => n1027, B => n1026,
                           ZN => curr_proc_regs(42));
   U1592 : NAND2_X1 port map( A1 => regs(942), A2 => n10, ZN => n1030);
   U1593 : AOI22_X1 port map( A1 => n88, A2 => regs(1454), B1 => n39, B2 => 
                           regs(430), ZN => n1029);
   U1594 : AOI22_X1 port map( A1 => n116, A2 => regs(2478), B1 => n70, B2 => 
                           regs(1966), ZN => n1028);
   U1595 : NAND3_X1 port map( A1 => n1030, A2 => n1029, A3 => n1028, ZN => 
                           curr_proc_regs(430));
   U1596 : NAND2_X1 port map( A1 => regs(1455), A2 => n90, ZN => n1033);
   U1597 : AOI22_X1 port map( A1 => n51, A2 => regs(943), B1 => n24, B2 => 
                           regs(431), ZN => n1032);
   U1598 : AOI22_X1 port map( A1 => n116, A2 => regs(2479), B1 => n74, B2 => 
                           regs(1967), ZN => n1031);
   U1599 : NAND3_X1 port map( A1 => n1033, A2 => n1032, A3 => n1031, ZN => 
                           curr_proc_regs(431));
   U1600 : NAND2_X1 port map( A1 => regs(1456), A2 => n94, ZN => n1036);
   U1601 : AOI22_X1 port map( A1 => n50, A2 => regs(944), B1 => n23, B2 => 
                           regs(432), ZN => n1035);
   U1602 : AOI22_X1 port map( A1 => n116, A2 => regs(2480), B1 => n73, B2 => 
                           regs(1968), ZN => n1034);
   U1603 : NAND3_X1 port map( A1 => n1036, A2 => n1035, A3 => n1034, ZN => 
                           curr_proc_regs(432));
   U1604 : NAND2_X1 port map( A1 => regs(945), A2 => n10, ZN => n1039);
   U1605 : AOI22_X1 port map( A1 => n88, A2 => regs(1457), B1 => n39, B2 => 
                           regs(433), ZN => n1038);
   U1606 : AOI22_X1 port map( A1 => n116, A2 => regs(2481), B1 => n71, B2 => 
                           regs(1969), ZN => n1037);
   U1607 : NAND3_X1 port map( A1 => n1039, A2 => n1038, A3 => n1037, ZN => 
                           curr_proc_regs(433));
   U1608 : NAND2_X1 port map( A1 => regs(1458), A2 => n95, ZN => n1042);
   U1609 : AOI22_X1 port map( A1 => n49, A2 => regs(946), B1 => n35, B2 => 
                           regs(434), ZN => n1041);
   U1610 : AOI22_X1 port map( A1 => n116, A2 => regs(2482), B1 => n73, B2 => 
                           regs(1970), ZN => n1040);
   U1611 : NAND3_X1 port map( A1 => n1042, A2 => n1041, A3 => n1040, ZN => 
                           curr_proc_regs(434));
   U1612 : NAND2_X1 port map( A1 => regs(947), A2 => n61, ZN => n1045);
   U1613 : AOI22_X1 port map( A1 => n87, A2 => regs(1459), B1 => n42, B2 => 
                           regs(435), ZN => n1044);
   U1614 : AOI22_X1 port map( A1 => n116, A2 => regs(2483), B1 => n70, B2 => 
                           regs(1971), ZN => n1043);
   U1615 : NAND3_X1 port map( A1 => n1045, A2 => n1044, A3 => n1043, ZN => 
                           curr_proc_regs(435));
   U1616 : NAND2_X1 port map( A1 => regs(948), A2 => n50, ZN => n1048);
   U1617 : AOI22_X1 port map( A1 => n81, A2 => regs(1460), B1 => n39, B2 => 
                           regs(436), ZN => n1047);
   U1618 : AOI22_X1 port map( A1 => n116, A2 => regs(2484), B1 => n74, B2 => 
                           regs(1972), ZN => n1046);
   U1619 : NAND3_X1 port map( A1 => n1048, A2 => n1047, A3 => n1046, ZN => 
                           curr_proc_regs(436));
   U1620 : NAND2_X1 port map( A1 => regs(1461), A2 => n84, ZN => n1051);
   U1621 : AOI22_X1 port map( A1 => n56, A2 => regs(949), B1 => n23, B2 => 
                           regs(437), ZN => n1050);
   U1622 : AOI22_X1 port map( A1 => n116, A2 => regs(2485), B1 => n75, B2 => 
                           regs(1973), ZN => n1049);
   U1623 : NAND3_X1 port map( A1 => n1051, A2 => n1050, A3 => n1049, ZN => 
                           curr_proc_regs(437));
   U1624 : NAND2_X1 port map( A1 => regs(1462), A2 => n93, ZN => n1054);
   U1625 : AOI22_X1 port map( A1 => n61, A2 => regs(950), B1 => n39, B2 => 
                           regs(438), ZN => n1053);
   U1626 : AOI22_X1 port map( A1 => n116, A2 => regs(2486), B1 => n68, B2 => 
                           regs(1974), ZN => n1052);
   U1627 : NAND3_X1 port map( A1 => n1054, A2 => n1053, A3 => n1052, ZN => 
                           curr_proc_regs(438));
   U1628 : NAND2_X1 port map( A1 => regs(951), A2 => n10, ZN => n1057);
   U1629 : AOI22_X1 port map( A1 => n83, A2 => regs(1463), B1 => n42, B2 => 
                           regs(439), ZN => n1056);
   U1630 : AOI22_X1 port map( A1 => n116, A2 => regs(2487), B1 => n68, B2 => 
                           regs(1975), ZN => n1055);
   U1631 : NAND3_X1 port map( A1 => n1057, A2 => n1056, A3 => n1055, ZN => 
                           curr_proc_regs(439));
   U1632 : INV_X1 port map( A => regs(1067), ZN => n1428);
   U1633 : AOI22_X1 port map( A1 => n116, A2 => regs(2091), B1 => n72, B2 => 
                           regs(1579), ZN => n1059);
   U1634 : AOI22_X1 port map( A1 => n51, A2 => regs(555), B1 => n23, B2 => 
                           regs(43), ZN => n1058);
   U1635 : OAI211_X1 port map( C1 => n2199, C2 => n1428, A => n1059, B => n1058
                           , ZN => curr_proc_regs(43));
   U1636 : NAND2_X1 port map( A1 => regs(952), A2 => n10, ZN => n1062);
   U1637 : AOI22_X1 port map( A1 => n98, A2 => regs(1464), B1 => n26, B2 => 
                           regs(440), ZN => n1061);
   U1638 : AOI22_X1 port map( A1 => n116, A2 => regs(2488), B1 => n75, B2 => 
                           regs(1976), ZN => n1060);
   U1639 : NAND3_X1 port map( A1 => n1062, A2 => n1061, A3 => n1060, ZN => 
                           curr_proc_regs(440));
   U1640 : NAND2_X1 port map( A1 => regs(1465), A2 => n14, ZN => n1065);
   U1641 : AOI22_X1 port map( A1 => n54, A2 => regs(953), B1 => n30, B2 => 
                           regs(441), ZN => n1064);
   U1642 : AOI22_X1 port map( A1 => n116, A2 => regs(2489), B1 => n68, B2 => 
                           regs(1977), ZN => n1063);
   U1643 : NAND3_X1 port map( A1 => n1065, A2 => n1064, A3 => n1063, ZN => 
                           curr_proc_regs(441));
   U1644 : NAND2_X1 port map( A1 => regs(954), A2 => n10, ZN => n1068);
   U1645 : AOI22_X1 port map( A1 => n81, A2 => regs(1466), B1 => n33, B2 => 
                           regs(442), ZN => n1067);
   U1646 : AOI22_X1 port map( A1 => n116, A2 => regs(2490), B1 => n68, B2 => 
                           regs(1978), ZN => n1066);
   U1647 : NAND3_X1 port map( A1 => n1068, A2 => n1067, A3 => n1066, ZN => 
                           curr_proc_regs(442));
   U1648 : NAND2_X1 port map( A1 => regs(955), A2 => n10, ZN => n1071);
   U1649 : AOI22_X1 port map( A1 => n81, A2 => regs(1467), B1 => n30, B2 => 
                           regs(443), ZN => n1070);
   U1650 : AOI22_X1 port map( A1 => n116, A2 => regs(2491), B1 => n72, B2 => 
                           regs(1979), ZN => n1069);
   U1651 : NAND3_X1 port map( A1 => n1071, A2 => n1070, A3 => n1069, ZN => 
                           curr_proc_regs(443));
   U1652 : NAND2_X1 port map( A1 => regs(956), A2 => n10, ZN => n1074);
   U1653 : AOI22_X1 port map( A1 => n81, A2 => regs(1468), B1 => n32, B2 => 
                           regs(444), ZN => n1073);
   U1654 : AOI22_X1 port map( A1 => n116, A2 => regs(2492), B1 => n75, B2 => 
                           regs(1980), ZN => n1072);
   U1655 : NAND3_X1 port map( A1 => n1074, A2 => n1073, A3 => n1072, ZN => 
                           curr_proc_regs(444));
   U1656 : NAND2_X1 port map( A1 => regs(957), A2 => n10, ZN => n1077);
   U1657 : AOI22_X1 port map( A1 => n81, A2 => regs(1469), B1 => n37, B2 => 
                           regs(445), ZN => n1076);
   U1658 : AOI22_X1 port map( A1 => n109, A2 => regs(2493), B1 => n68, B2 => 
                           regs(1981), ZN => n1075);
   U1659 : NAND3_X1 port map( A1 => n1077, A2 => n1076, A3 => n1075, ZN => 
                           curr_proc_regs(445));
   U1660 : NAND2_X1 port map( A1 => regs(1470), A2 => n14, ZN => n1080);
   U1661 : AOI22_X1 port map( A1 => n54, A2 => regs(958), B1 => n40, B2 => 
                           regs(446), ZN => n1079);
   U1662 : AOI22_X1 port map( A1 => n104, A2 => regs(2494), B1 => n68, B2 => 
                           regs(1982), ZN => n1078);
   U1663 : NAND3_X1 port map( A1 => n1080, A2 => n1079, A3 => n1078, ZN => 
                           curr_proc_regs(446));
   U1664 : NAND2_X1 port map( A1 => regs(959), A2 => n10, ZN => n1083);
   U1665 : AOI22_X1 port map( A1 => n81, A2 => regs(1471), B1 => n32, B2 => 
                           regs(447), ZN => n1082);
   U1666 : AOI22_X1 port map( A1 => n105, A2 => regs(2495), B1 => n68, B2 => 
                           regs(1983), ZN => n1081);
   U1667 : NAND3_X1 port map( A1 => n1083, A2 => n1082, A3 => n1081, ZN => 
                           curr_proc_regs(447));
   U1668 : NAND2_X1 port map( A1 => regs(960), A2 => n10, ZN => n1086);
   U1669 : AOI22_X1 port map( A1 => n81, A2 => regs(1472), B1 => n37, B2 => 
                           regs(448), ZN => n1085);
   U1670 : AOI22_X1 port map( A1 => n106, A2 => regs(2496), B1 => n68, B2 => 
                           regs(1984), ZN => n1084);
   U1671 : NAND3_X1 port map( A1 => n1086, A2 => n1085, A3 => n1084, ZN => 
                           curr_proc_regs(448));
   U1672 : NAND2_X1 port map( A1 => regs(961), A2 => n48, ZN => n1089);
   U1673 : AOI22_X1 port map( A1 => n81, A2 => regs(1473), B1 => n40, B2 => 
                           regs(449), ZN => n1088);
   U1674 : AOI22_X1 port map( A1 => n112, A2 => regs(2497), B1 => n72, B2 => 
                           regs(1985), ZN => n1087);
   U1675 : NAND3_X1 port map( A1 => n1089, A2 => n1088, A3 => n1087, ZN => 
                           curr_proc_regs(449));
   U1676 : INV_X1 port map( A => regs(556), ZN => n1431);
   U1677 : AOI22_X1 port map( A1 => n111, A2 => regs(2092), B1 => n72, B2 => 
                           regs(1580), ZN => n1091);
   U1678 : AOI22_X1 port map( A1 => n81, A2 => regs(1068), B1 => n28, B2 => 
                           regs(44), ZN => n1090);
   U1679 : OAI211_X1 port map( C1 => n66, C2 => n1431, A => n1091, B => n1090, 
                           ZN => curr_proc_regs(44));
   U1680 : NAND2_X1 port map( A1 => regs(962), A2 => n10, ZN => n1094);
   U1681 : AOI22_X1 port map( A1 => n81, A2 => regs(1474), B1 => n23, B2 => 
                           regs(450), ZN => n1093);
   U1682 : AOI22_X1 port map( A1 => n116, A2 => regs(2498), B1 => n75, B2 => 
                           regs(1986), ZN => n1092);
   U1683 : NAND3_X1 port map( A1 => n1094, A2 => n1093, A3 => n1092, ZN => 
                           curr_proc_regs(450));
   U1684 : NAND2_X1 port map( A1 => regs(1475), A2 => n17, ZN => n1097);
   U1685 : AOI22_X1 port map( A1 => n54, A2 => regs(963), B1 => n42, B2 => 
                           regs(451), ZN => n1096);
   U1686 : AOI22_X1 port map( A1 => n116, A2 => regs(2499), B1 => n68, B2 => 
                           regs(1987), ZN => n1095);
   U1687 : NAND3_X1 port map( A1 => n1097, A2 => n1096, A3 => n1095, ZN => 
                           curr_proc_regs(451));
   U1688 : NAND2_X1 port map( A1 => regs(1476), A2 => n14, ZN => n1100);
   U1689 : AOI22_X1 port map( A1 => n54, A2 => regs(964), B1 => n43, B2 => 
                           regs(452), ZN => n1099);
   U1690 : AOI22_X1 port map( A1 => n116, A2 => regs(2500), B1 => n68, B2 => 
                           regs(1988), ZN => n1098);
   U1691 : NAND3_X1 port map( A1 => n1100, A2 => n1099, A3 => n1098, ZN => 
                           curr_proc_regs(452));
   U1692 : NAND2_X1 port map( A1 => regs(1477), A2 => n98, ZN => n1103);
   U1693 : AOI22_X1 port map( A1 => n54, A2 => regs(965), B1 => n24, B2 => 
                           regs(453), ZN => n1102);
   U1694 : AOI22_X1 port map( A1 => n116, A2 => regs(2501), B1 => n75, B2 => 
                           regs(1989), ZN => n1101);
   U1695 : NAND3_X1 port map( A1 => n1103, A2 => n1102, A3 => n1101, ZN => 
                           curr_proc_regs(453));
   U1696 : NAND2_X1 port map( A1 => regs(1478), A2 => n97, ZN => n1106);
   U1697 : AOI22_X1 port map( A1 => n54, A2 => regs(966), B1 => n42, B2 => 
                           regs(454), ZN => n1105);
   U1698 : AOI22_X1 port map( A1 => n116, A2 => regs(2502), B1 => n72, B2 => 
                           regs(1990), ZN => n1104);
   U1699 : NAND3_X1 port map( A1 => n1106, A2 => n1105, A3 => n1104, ZN => 
                           curr_proc_regs(454));
   U1700 : NAND2_X1 port map( A1 => regs(967), A2 => n10, ZN => n1109);
   U1701 : AOI22_X1 port map( A1 => n81, A2 => regs(1479), B1 => n39, B2 => 
                           regs(455), ZN => n1108);
   U1702 : AOI22_X1 port map( A1 => n116, A2 => regs(2503), B1 => n75, B2 => 
                           regs(1991), ZN => n1107);
   U1703 : NAND3_X1 port map( A1 => n1109, A2 => n1108, A3 => n1107, ZN => 
                           curr_proc_regs(455));
   U1704 : NAND2_X1 port map( A1 => regs(968), A2 => n58, ZN => n1112);
   U1705 : AOI22_X1 port map( A1 => n81, A2 => regs(1480), B1 => n24, B2 => 
                           regs(456), ZN => n1111);
   U1706 : AOI22_X1 port map( A1 => n116, A2 => regs(2504), B1 => n68, B2 => 
                           regs(1992), ZN => n1110);
   U1707 : NAND3_X1 port map( A1 => n1112, A2 => n1111, A3 => n1110, ZN => 
                           curr_proc_regs(456));
   U1708 : NAND2_X1 port map( A1 => regs(1481), A2 => n81, ZN => n1115);
   U1709 : AOI22_X1 port map( A1 => n54, A2 => regs(969), B1 => n2, B2 => 
                           regs(457), ZN => n1114);
   U1710 : AOI22_X1 port map( A1 => n116, A2 => regs(2505), B1 => n75, B2 => 
                           regs(1993), ZN => n1113);
   U1711 : NAND3_X1 port map( A1 => n1115, A2 => n1114, A3 => n1113, ZN => 
                           curr_proc_regs(457));
   U1712 : NAND2_X1 port map( A1 => regs(1482), A2 => n80, ZN => n1118);
   U1713 : AOI22_X1 port map( A1 => n54, A2 => regs(970), B1 => n7, B2 => 
                           regs(458), ZN => n1117);
   U1714 : AOI22_X1 port map( A1 => n116, A2 => regs(2506), B1 => n75, B2 => 
                           regs(1994), ZN => n1116);
   U1715 : NAND3_X1 port map( A1 => n1118, A2 => n1117, A3 => n1116, ZN => 
                           curr_proc_regs(458));
   U1716 : NAND2_X1 port map( A1 => regs(1483), A2 => n79, ZN => n1121);
   U1717 : AOI22_X1 port map( A1 => n54, A2 => regs(971), B1 => n7, B2 => 
                           regs(459), ZN => n1120);
   U1718 : AOI22_X1 port map( A1 => n116, A2 => regs(2507), B1 => n75, B2 => 
                           regs(1995), ZN => n1119);
   U1719 : NAND3_X1 port map( A1 => n1121, A2 => n1120, A3 => n1119, ZN => 
                           curr_proc_regs(459));
   U1720 : INV_X1 port map( A => regs(557), ZN => n1434);
   U1721 : AOI22_X1 port map( A1 => n116, A2 => regs(2093), B1 => n75, B2 => 
                           regs(1581), ZN => n1123);
   U1722 : AOI22_X1 port map( A1 => n80, A2 => regs(1069), B1 => n25, B2 => 
                           regs(45), ZN => n1122);
   U1723 : OAI211_X1 port map( C1 => n65, C2 => n1434, A => n1123, B => n1122, 
                           ZN => curr_proc_regs(45));
   U1724 : NAND2_X1 port map( A1 => regs(1484), A2 => n83, ZN => n1126);
   U1725 : AOI22_X1 port map( A1 => n54, A2 => regs(972), B1 => n37, B2 => 
                           regs(460), ZN => n1125);
   U1726 : AOI22_X1 port map( A1 => n116, A2 => regs(2508), B1 => n75, B2 => 
                           regs(1996), ZN => n1124);
   U1727 : NAND3_X1 port map( A1 => n1126, A2 => n1125, A3 => n1124, ZN => 
                           curr_proc_regs(460));
   U1728 : NAND2_X1 port map( A1 => regs(973), A2 => n10, ZN => n1129);
   U1729 : AOI22_X1 port map( A1 => n80, A2 => regs(1485), B1 => n40, B2 => 
                           regs(461), ZN => n1128);
   U1730 : AOI22_X1 port map( A1 => n107, A2 => regs(2509), B1 => n75, B2 => 
                           regs(1997), ZN => n1127);
   U1731 : NAND3_X1 port map( A1 => n1129, A2 => n1128, A3 => n1127, ZN => 
                           curr_proc_regs(461));
   U1732 : NAND2_X1 port map( A1 => regs(974), A2 => n57, ZN => n1132);
   U1733 : AOI22_X1 port map( A1 => n80, A2 => regs(1486), B1 => n28, B2 => 
                           regs(462), ZN => n1131);
   U1734 : AOI22_X1 port map( A1 => n108, A2 => regs(2510), B1 => n75, B2 => 
                           regs(1998), ZN => n1130);
   U1735 : NAND3_X1 port map( A1 => n1132, A2 => n1131, A3 => n1130, ZN => 
                           curr_proc_regs(462));
   U1736 : NAND2_X1 port map( A1 => regs(975), A2 => n59, ZN => n1135);
   U1737 : AOI22_X1 port map( A1 => n80, A2 => regs(1487), B1 => n27, B2 => 
                           regs(463), ZN => n1134);
   U1738 : AOI22_X1 port map( A1 => n109, A2 => regs(2511), B1 => n75, B2 => 
                           regs(1999), ZN => n1133);
   U1739 : NAND3_X1 port map( A1 => n1135, A2 => n1134, A3 => n1133, ZN => 
                           curr_proc_regs(463));
   U1740 : NAND2_X1 port map( A1 => regs(1488), A2 => n90, ZN => n1138);
   U1741 : AOI22_X1 port map( A1 => n55, A2 => regs(976), B1 => n26, B2 => 
                           regs(464), ZN => n1137);
   U1742 : AOI22_X1 port map( A1 => n109, A2 => regs(2512), B1 => n75, B2 => 
                           regs(2000), ZN => n1136);
   U1743 : NAND3_X1 port map( A1 => n1138, A2 => n1137, A3 => n1136, ZN => 
                           curr_proc_regs(464));
   U1744 : NAND2_X1 port map( A1 => regs(977), A2 => n56, ZN => n1141);
   U1745 : AOI22_X1 port map( A1 => n80, A2 => regs(1489), B1 => n33, B2 => 
                           regs(465), ZN => n1140);
   U1746 : AOI22_X1 port map( A1 => n108, A2 => regs(2513), B1 => n75, B2 => 
                           regs(2001), ZN => n1139);
   U1747 : NAND3_X1 port map( A1 => n1141, A2 => n1140, A3 => n1139, ZN => 
                           curr_proc_regs(465));
   U1748 : NAND2_X1 port map( A1 => regs(1490), A2 => n94, ZN => n1144);
   U1749 : AOI22_X1 port map( A1 => n50, A2 => regs(978), B1 => n30, B2 => 
                           regs(466), ZN => n1143);
   U1750 : AOI22_X1 port map( A1 => n107, A2 => regs(2514), B1 => n75, B2 => 
                           regs(2002), ZN => n1142);
   U1751 : NAND3_X1 port map( A1 => n1144, A2 => n1143, A3 => n1142, ZN => 
                           curr_proc_regs(466));
   U1752 : NAND2_X1 port map( A1 => regs(979), A2 => n50, ZN => n1147);
   U1753 : AOI22_X1 port map( A1 => n80, A2 => regs(1491), B1 => n37, B2 => 
                           regs(467), ZN => n1146);
   U1754 : AOI22_X1 port map( A1 => n108, A2 => regs(2515), B1 => n75, B2 => 
                           regs(2003), ZN => n1145);
   U1755 : NAND3_X1 port map( A1 => n1147, A2 => n1146, A3 => n1145, ZN => 
                           curr_proc_regs(467));
   U1756 : NAND2_X1 port map( A1 => regs(1492), A2 => n92, ZN => n1150);
   U1757 : AOI22_X1 port map( A1 => n49, A2 => regs(980), B1 => n37, B2 => 
                           regs(468), ZN => n1149);
   U1758 : AOI22_X1 port map( A1 => n109, A2 => regs(2516), B1 => n68, B2 => 
                           regs(2004), ZN => n1148);
   U1759 : NAND3_X1 port map( A1 => n1150, A2 => n1149, A3 => n1148, ZN => 
                           curr_proc_regs(468));
   U1760 : NAND2_X1 port map( A1 => regs(981), A2 => n62, ZN => n1153);
   U1761 : AOI22_X1 port map( A1 => n80, A2 => regs(1493), B1 => n37, B2 => 
                           regs(469), ZN => n1152);
   U1762 : AOI22_X1 port map( A1 => n107, A2 => regs(2517), B1 => n68, B2 => 
                           regs(2005), ZN => n1151);
   U1763 : NAND3_X1 port map( A1 => n1153, A2 => n1152, A3 => n1151, ZN => 
                           curr_proc_regs(469));
   U1764 : INV_X1 port map( A => regs(558), ZN => n1437);
   U1765 : AOI22_X1 port map( A1 => n109, A2 => regs(2094), B1 => n68, B2 => 
                           regs(1582), ZN => n1155);
   U1766 : AOI22_X1 port map( A1 => n80, A2 => regs(1070), B1 => n37, B2 => 
                           regs(46), ZN => n1154);
   U1767 : OAI211_X1 port map( C1 => n1, C2 => n1437, A => n1155, B => n1154, 
                           ZN => curr_proc_regs(46));
   U1768 : NAND2_X1 port map( A1 => regs(982), A2 => n58, ZN => n1158);
   U1769 : AOI22_X1 port map( A1 => n80, A2 => regs(1494), B1 => n25, B2 => 
                           regs(470), ZN => n1157);
   U1770 : AOI22_X1 port map( A1 => n107, A2 => regs(2518), B1 => n68, B2 => 
                           regs(2006), ZN => n1156);
   U1771 : NAND3_X1 port map( A1 => n1158, A2 => n1157, A3 => n1156, ZN => 
                           curr_proc_regs(470));
   U1772 : NAND2_X1 port map( A1 => regs(1495), A2 => n92, ZN => n1161);
   U1773 : AOI22_X1 port map( A1 => n56, A2 => regs(983), B1 => n25, B2 => 
                           regs(471), ZN => n1160);
   U1774 : AOI22_X1 port map( A1 => n108, A2 => regs(2519), B1 => n72, B2 => 
                           regs(2007), ZN => n1159);
   U1775 : NAND3_X1 port map( A1 => n1161, A2 => n1160, A3 => n1159, ZN => 
                           curr_proc_regs(471));
   U1776 : NAND2_X1 port map( A1 => regs(1496), A2 => n90, ZN => n1164);
   U1777 : AOI22_X1 port map( A1 => n61, A2 => regs(984), B1 => n31, B2 => 
                           regs(472), ZN => n1163);
   U1778 : AOI22_X1 port map( A1 => n107, A2 => regs(2520), B1 => n75, B2 => 
                           regs(2008), ZN => n1162);
   U1779 : NAND3_X1 port map( A1 => n1164, A2 => n1163, A3 => n1162, ZN => 
                           curr_proc_regs(472));
   U1780 : NAND2_X1 port map( A1 => regs(985), A2 => n10, ZN => n1167);
   U1781 : AOI22_X1 port map( A1 => n80, A2 => regs(1497), B1 => n29, B2 => 
                           regs(473), ZN => n1166);
   U1782 : AOI22_X1 port map( A1 => n108, A2 => regs(2521), B1 => n68, B2 => 
                           regs(2009), ZN => n1165);
   U1783 : NAND3_X1 port map( A1 => n1167, A2 => n1166, A3 => n1165, ZN => 
                           curr_proc_regs(473));
   U1784 : NAND2_X1 port map( A1 => regs(986), A2 => n10, ZN => n1170);
   U1785 : AOI22_X1 port map( A1 => n80, A2 => regs(1498), B1 => n38, B2 => 
                           regs(474), ZN => n1169);
   U1786 : AOI22_X1 port map( A1 => n109, A2 => regs(2522), B1 => n68, B2 => 
                           regs(2010), ZN => n1168);
   U1787 : NAND3_X1 port map( A1 => n1170, A2 => n1169, A3 => n1168, ZN => 
                           curr_proc_regs(474));
   U1788 : NAND2_X1 port map( A1 => regs(1499), A2 => n96, ZN => n1173);
   U1789 : AOI22_X1 port map( A1 => n59, A2 => regs(987), B1 => n41, B2 => 
                           regs(475), ZN => n1172);
   U1790 : AOI22_X1 port map( A1 => n109, A2 => regs(2523), B1 => n68, B2 => 
                           regs(2011), ZN => n1171);
   U1791 : NAND3_X1 port map( A1 => n1173, A2 => n1172, A3 => n1171, ZN => 
                           curr_proc_regs(475));
   U1792 : NAND2_X1 port map( A1 => regs(1500), A2 => n96, ZN => n1176);
   U1793 : AOI22_X1 port map( A1 => n57, A2 => regs(988), B1 => n2, B2 => 
                           regs(476), ZN => n1175);
   U1794 : AOI22_X1 port map( A1 => n107, A2 => regs(2524), B1 => n72, B2 => 
                           regs(2012), ZN => n1174);
   U1795 : NAND3_X1 port map( A1 => n1176, A2 => n1175, A3 => n1174, ZN => 
                           curr_proc_regs(476));
   U1796 : NAND2_X1 port map( A1 => regs(989), A2 => n60, ZN => n1179);
   U1797 : AOI22_X1 port map( A1 => n80, A2 => regs(1501), B1 => n38, B2 => 
                           regs(477), ZN => n1178);
   U1798 : AOI22_X1 port map( A1 => n108, A2 => regs(2525), B1 => n72, B2 => 
                           regs(2013), ZN => n1177);
   U1799 : NAND3_X1 port map( A1 => n1179, A2 => n1178, A3 => n1177, ZN => 
                           curr_proc_regs(477));
   U1800 : NAND2_X1 port map( A1 => regs(990), A2 => n51, ZN => n1182);
   U1801 : AOI22_X1 port map( A1 => n81, A2 => regs(1502), B1 => n38, B2 => 
                           regs(478), ZN => n1181);
   U1802 : AOI22_X1 port map( A1 => n109, A2 => regs(2526), B1 => n75, B2 => 
                           regs(2014), ZN => n1180);
   U1803 : NAND3_X1 port map( A1 => n1182, A2 => n1181, A3 => n1180, ZN => 
                           curr_proc_regs(478));
   U1804 : NAND2_X1 port map( A1 => regs(991), A2 => n62, ZN => n1185);
   U1805 : AOI22_X1 port map( A1 => n87, A2 => regs(1503), B1 => n38, B2 => 
                           regs(479), ZN => n1184);
   U1806 : AOI22_X1 port map( A1 => n107, A2 => regs(2527), B1 => n68, B2 => 
                           regs(2015), ZN => n1183);
   U1807 : NAND3_X1 port map( A1 => n1185, A2 => n1184, A3 => n1183, ZN => 
                           curr_proc_regs(479));
   U1808 : INV_X1 port map( A => regs(559), ZN => n1440);
   U1809 : AOI22_X1 port map( A1 => n107, A2 => regs(2095), B1 => n68, B2 => 
                           regs(1583), ZN => n1187);
   U1810 : AOI22_X1 port map( A1 => n87, A2 => regs(1071), B1 => n38, B2 => 
                           regs(47), ZN => n1186);
   U1811 : OAI211_X1 port map( C1 => n64, C2 => n1440, A => n1187, B => n1186, 
                           ZN => curr_proc_regs(47));
   U1812 : NAND2_X1 port map( A1 => regs(992), A2 => n52, ZN => n1190);
   U1813 : AOI22_X1 port map( A1 => n88, A2 => regs(1504), B1 => n37, B2 => 
                           regs(480), ZN => n1189);
   U1814 : AOI22_X1 port map( A1 => n108, A2 => regs(2528), B1 => n68, B2 => 
                           regs(2016), ZN => n1188);
   U1815 : NAND3_X1 port map( A1 => n1190, A2 => n1189, A3 => n1188, ZN => 
                           curr_proc_regs(480));
   U1816 : NAND2_X1 port map( A1 => regs(1505), A2 => n96, ZN => n1193);
   U1817 : AOI22_X1 port map( A1 => n55, A2 => regs(993), B1 => n37, B2 => 
                           regs(481), ZN => n1192);
   U1818 : AOI22_X1 port map( A1 => n108, A2 => regs(2529), B1 => n72, B2 => 
                           regs(2017), ZN => n1191);
   U1819 : NAND3_X1 port map( A1 => n1193, A2 => n1192, A3 => n1191, ZN => 
                           curr_proc_regs(481));
   U1820 : NAND2_X1 port map( A1 => regs(1506), A2 => n96, ZN => n1196);
   U1821 : AOI22_X1 port map( A1 => n54, A2 => regs(994), B1 => n37, B2 => 
                           regs(482), ZN => n1195);
   U1822 : AOI22_X1 port map( A1 => n109, A2 => regs(2530), B1 => n75, B2 => 
                           regs(2018), ZN => n1194);
   U1823 : NAND3_X1 port map( A1 => n1196, A2 => n1195, A3 => n1194, ZN => 
                           curr_proc_regs(482));
   U1824 : NAND2_X1 port map( A1 => regs(995), A2 => n5, ZN => n1199);
   U1825 : AOI22_X1 port map( A1 => n94, A2 => regs(1507), B1 => n37, B2 => 
                           regs(483), ZN => n1198);
   U1826 : AOI22_X1 port map( A1 => n107, A2 => regs(2531), B1 => n72, B2 => 
                           regs(2019), ZN => n1197);
   U1827 : NAND3_X1 port map( A1 => n1199, A2 => n1198, A3 => n1197, ZN => 
                           curr_proc_regs(483));
   U1828 : NAND2_X1 port map( A1 => regs(996), A2 => n63, ZN => n1202);
   U1829 : AOI22_X1 port map( A1 => n98, A2 => regs(1508), B1 => n37, B2 => 
                           regs(484), ZN => n1201);
   U1830 : AOI22_X1 port map( A1 => n108, A2 => regs(2532), B1 => n75, B2 => 
                           regs(2020), ZN => n1200);
   U1831 : NAND3_X1 port map( A1 => n1202, A2 => n1201, A3 => n1200, ZN => 
                           curr_proc_regs(484));
   U1832 : NAND2_X1 port map( A1 => regs(997), A2 => n63, ZN => n1205);
   U1833 : AOI22_X1 port map( A1 => n96, A2 => regs(1509), B1 => n37, B2 => 
                           regs(485), ZN => n1204);
   U1834 : AOI22_X1 port map( A1 => n109, A2 => regs(2533), B1 => n68, B2 => 
                           regs(2021), ZN => n1203);
   U1835 : NAND3_X1 port map( A1 => n1205, A2 => n1204, A3 => n1203, ZN => 
                           curr_proc_regs(485));
   U1836 : NAND2_X1 port map( A1 => regs(998), A2 => n5, ZN => n1208);
   U1837 : AOI22_X1 port map( A1 => n79, A2 => regs(1510), B1 => n37, B2 => 
                           regs(486), ZN => n1207);
   U1838 : AOI22_X1 port map( A1 => n107, A2 => regs(2534), B1 => n68, B2 => 
                           regs(2022), ZN => n1206);
   U1839 : NAND3_X1 port map( A1 => n1208, A2 => n1207, A3 => n1206, ZN => 
                           curr_proc_regs(486));
   U1840 : NAND2_X1 port map( A1 => regs(1511), A2 => n83, ZN => n1211);
   U1841 : AOI22_X1 port map( A1 => n52, A2 => regs(999), B1 => n39, B2 => 
                           regs(487), ZN => n1210);
   U1842 : AOI22_X1 port map( A1 => n108, A2 => regs(2535), B1 => n68, B2 => 
                           regs(2023), ZN => n1209);
   U1843 : NAND3_X1 port map( A1 => n1211, A2 => n1210, A3 => n1209, ZN => 
                           curr_proc_regs(487));
   U1844 : NAND2_X1 port map( A1 => regs(1000), A2 => n63, ZN => n1214);
   U1845 : AOI22_X1 port map( A1 => n86, A2 => regs(1512), B1 => n39, B2 => 
                           regs(488), ZN => n1213);
   U1846 : AOI22_X1 port map( A1 => n109, A2 => regs(2536), B1 => n68, B2 => 
                           regs(2024), ZN => n1212);
   U1847 : NAND3_X1 port map( A1 => n1214, A2 => n1213, A3 => n1212, ZN => 
                           curr_proc_regs(488));
   U1848 : NAND2_X1 port map( A1 => regs(1513), A2 => n86, ZN => n1217);
   U1849 : AOI22_X1 port map( A1 => n53, A2 => regs(1001), B1 => n39, B2 => 
                           regs(489), ZN => n1216);
   U1850 : AOI22_X1 port map( A1 => n107, A2 => regs(2537), B1 => n68, B2 => 
                           regs(2025), ZN => n1215);
   U1851 : NAND3_X1 port map( A1 => n1217, A2 => n1216, A3 => n1215, ZN => 
                           curr_proc_regs(489));
   U1852 : INV_X1 port map( A => regs(560), ZN => n1445);
   U1853 : AOI22_X1 port map( A1 => n108, A2 => regs(2096), B1 => n68, B2 => 
                           regs(1584), ZN => n1219);
   U1854 : AOI22_X1 port map( A1 => n79, A2 => regs(1072), B1 => n39, B2 => 
                           regs(48), ZN => n1218);
   U1855 : OAI211_X1 port map( C1 => n67, C2 => n1445, A => n1219, B => n1218, 
                           ZN => curr_proc_regs(48));
   U1856 : NAND2_X1 port map( A1 => regs(1002), A2 => n5, ZN => n1222);
   U1857 : AOI22_X1 port map( A1 => n79, A2 => regs(1514), B1 => n38, B2 => 
                           regs(490), ZN => n1221);
   U1858 : AOI22_X1 port map( A1 => n109, A2 => regs(2538), B1 => n68, B2 => 
                           regs(2026), ZN => n1220);
   U1859 : NAND3_X1 port map( A1 => n1222, A2 => n1221, A3 => n1220, ZN => 
                           curr_proc_regs(490));
   U1860 : NAND2_X1 port map( A1 => regs(1003), A2 => n63, ZN => n1225);
   U1861 : AOI22_X1 port map( A1 => n79, A2 => regs(1515), B1 => n38, B2 => 
                           regs(491), ZN => n1224);
   U1862 : AOI22_X1 port map( A1 => n109, A2 => regs(2539), B1 => n68, B2 => 
                           regs(2027), ZN => n1223);
   U1863 : NAND3_X1 port map( A1 => n1225, A2 => n1224, A3 => n1223, ZN => 
                           curr_proc_regs(491));
   U1864 : NAND2_X1 port map( A1 => regs(1516), A2 => n97, ZN => n1228);
   U1865 : AOI22_X1 port map( A1 => n54, A2 => regs(1004), B1 => n38, B2 => 
                           regs(492), ZN => n1227);
   U1866 : AOI22_X1 port map( A1 => n109, A2 => regs(2540), B1 => n72, B2 => 
                           regs(2028), ZN => n1226);
   U1867 : NAND3_X1 port map( A1 => n1228, A2 => n1227, A3 => n1226, ZN => 
                           curr_proc_regs(492));
   U1868 : NAND2_X1 port map( A1 => regs(1517), A2 => n93, ZN => n1231);
   U1869 : AOI22_X1 port map( A1 => n62, A2 => regs(1005), B1 => n38, B2 => 
                           regs(493), ZN => n1230);
   U1870 : AOI22_X1 port map( A1 => n109, A2 => regs(2541), B1 => n75, B2 => 
                           regs(2029), ZN => n1229);
   U1871 : NAND3_X1 port map( A1 => n1231, A2 => n1230, A3 => n1229, ZN => 
                           curr_proc_regs(493));
   U1872 : NAND2_X1 port map( A1 => regs(1518), A2 => n89, ZN => n1234);
   U1873 : AOI22_X1 port map( A1 => n56, A2 => regs(1006), B1 => n38, B2 => 
                           regs(494), ZN => n1233);
   U1874 : AOI22_X1 port map( A1 => n109, A2 => regs(2542), B1 => n68, B2 => 
                           regs(2030), ZN => n1232);
   U1875 : NAND3_X1 port map( A1 => n1234, A2 => n1233, A3 => n1232, ZN => 
                           curr_proc_regs(494));
   U1876 : NAND2_X1 port map( A1 => regs(1519), A2 => n83, ZN => n1237);
   U1877 : AOI22_X1 port map( A1 => n62, A2 => regs(1007), B1 => n38, B2 => 
                           regs(495), ZN => n1236);
   U1878 : AOI22_X1 port map( A1 => n109, A2 => regs(2543), B1 => n68, B2 => 
                           regs(2031), ZN => n1235);
   U1879 : NAND3_X1 port map( A1 => n1237, A2 => n1236, A3 => n1235, ZN => 
                           curr_proc_regs(495));
   U1880 : NAND2_X1 port map( A1 => regs(1008), A2 => n63, ZN => n1240);
   U1881 : AOI22_X1 port map( A1 => n79, A2 => regs(1520), B1 => n38, B2 => 
                           regs(496), ZN => n1239);
   U1882 : AOI22_X1 port map( A1 => n109, A2 => regs(2544), B1 => n68, B2 => 
                           regs(2032), ZN => n1238);
   U1883 : NAND3_X1 port map( A1 => n1240, A2 => n1239, A3 => n1238, ZN => 
                           curr_proc_regs(496));
   U1884 : NAND2_X1 port map( A1 => regs(1009), A2 => n63, ZN => n1243);
   U1885 : AOI22_X1 port map( A1 => n79, A2 => regs(1521), B1 => n40, B2 => 
                           regs(497), ZN => n1242);
   U1886 : AOI22_X1 port map( A1 => n109, A2 => regs(2545), B1 => n3, B2 => 
                           regs(2033), ZN => n1241);
   U1887 : NAND3_X1 port map( A1 => n1243, A2 => n1242, A3 => n1241, ZN => 
                           curr_proc_regs(497));
   U1888 : NAND2_X1 port map( A1 => regs(1010), A2 => n5, ZN => n1246);
   U1889 : AOI22_X1 port map( A1 => n79, A2 => regs(1522), B1 => n40, B2 => 
                           regs(498), ZN => n1245);
   U1890 : AOI22_X1 port map( A1 => n109, A2 => regs(2546), B1 => n12, B2 => 
                           regs(2034), ZN => n1244);
   U1891 : NAND3_X1 port map( A1 => n1246, A2 => n1245, A3 => n1244, ZN => 
                           curr_proc_regs(498));
   U1892 : NAND2_X1 port map( A1 => regs(1523), A2 => n96, ZN => n1249);
   U1893 : AOI22_X1 port map( A1 => n58, A2 => regs(1011), B1 => n40, B2 => 
                           regs(499), ZN => n1248);
   U1894 : AOI22_X1 port map( A1 => n109, A2 => regs(2547), B1 => n68, B2 => 
                           regs(2035), ZN => n1247);
   U1895 : NAND3_X1 port map( A1 => n1249, A2 => n1248, A3 => n1247, ZN => 
                           curr_proc_regs(499));
   U1896 : INV_X1 port map( A => regs(1073), ZN => n1448);
   U1897 : AOI22_X1 port map( A1 => n109, A2 => regs(2097), B1 => n2195, B2 => 
                           regs(1585), ZN => n1251);
   U1898 : AOI22_X1 port map( A1 => n60, A2 => regs(561), B1 => n40, B2 => 
                           regs(49), ZN => n1250);
   U1899 : OAI211_X1 port map( C1 => n2199, C2 => n1448, A => n1251, B => n1250
                           , ZN => curr_proc_regs(49));
   U1900 : INV_X1 port map( A => regs(1028), ZN => n1306);
   U1901 : AOI22_X1 port map( A1 => n109, A2 => regs(2052), B1 => n71, B2 => 
                           regs(1540), ZN => n1253);
   U1902 : AOI22_X1 port map( A1 => n49, A2 => regs(516), B1 => n39, B2 => 
                           regs(4), ZN => n1252);
   U1903 : OAI211_X1 port map( C1 => n99, C2 => n1306, A => n1253, B => n1252, 
                           ZN => curr_proc_regs(4));
   U1904 : NAND2_X1 port map( A1 => regs(1012), A2 => n5, ZN => n1256);
   U1905 : AOI22_X1 port map( A1 => n79, A2 => regs(1524), B1 => n39, B2 => 
                           regs(500), ZN => n1255);
   U1906 : AOI22_X1 port map( A1 => n108, A2 => regs(2548), B1 => n68, B2 => 
                           regs(2036), ZN => n1254);
   U1907 : NAND3_X1 port map( A1 => n1256, A2 => n1255, A3 => n1254, ZN => 
                           curr_proc_regs(500));
   U1908 : NAND2_X1 port map( A1 => regs(1525), A2 => n85, ZN => n1259);
   U1909 : AOI22_X1 port map( A1 => n51, A2 => regs(1013), B1 => n39, B2 => 
                           regs(501), ZN => n1258);
   U1910 : AOI22_X1 port map( A1 => n108, A2 => regs(2549), B1 => n73, B2 => 
                           regs(2037), ZN => n1257);
   U1911 : NAND3_X1 port map( A1 => n1259, A2 => n1258, A3 => n1257, ZN => 
                           curr_proc_regs(501));
   U1912 : NAND2_X1 port map( A1 => regs(1526), A2 => n81, ZN => n1262);
   U1913 : AOI22_X1 port map( A1 => n48, A2 => regs(1014), B1 => n39, B2 => 
                           regs(502), ZN => n1261);
   U1914 : AOI22_X1 port map( A1 => n108, A2 => regs(2550), B1 => n73, B2 => 
                           regs(2038), ZN => n1260);
   U1915 : NAND3_X1 port map( A1 => n1262, A2 => n1261, A3 => n1260, ZN => 
                           curr_proc_regs(502));
   U1916 : NAND2_X1 port map( A1 => regs(1527), A2 => n87, ZN => n1265);
   U1917 : AOI22_X1 port map( A1 => n48, A2 => regs(1015), B1 => n39, B2 => 
                           regs(503), ZN => n1264);
   U1918 : AOI22_X1 port map( A1 => n108, A2 => regs(2551), B1 => n16, B2 => 
                           regs(2039), ZN => n1263);
   U1919 : NAND3_X1 port map( A1 => n1265, A2 => n1264, A3 => n1263, ZN => 
                           curr_proc_regs(503));
   U1920 : NAND2_X1 port map( A1 => regs(1528), A2 => n14, ZN => n1268);
   U1921 : AOI22_X1 port map( A1 => n48, A2 => regs(1016), B1 => n39, B2 => 
                           regs(504), ZN => n1267);
   U1922 : AOI22_X1 port map( A1 => n108, A2 => regs(2552), B1 => n16, B2 => 
                           regs(2040), ZN => n1266);
   U1923 : NAND3_X1 port map( A1 => n1268, A2 => n1267, A3 => n1266, ZN => 
                           curr_proc_regs(504));
   U1924 : NAND2_X1 port map( A1 => regs(1017), A2 => n5, ZN => n1271);
   U1925 : AOI22_X1 port map( A1 => n79, A2 => regs(1529), B1 => n39, B2 => 
                           regs(505), ZN => n1270);
   U1926 : AOI22_X1 port map( A1 => n108, A2 => regs(2553), B1 => n16, B2 => 
                           regs(2041), ZN => n1269);
   U1927 : NAND3_X1 port map( A1 => n1271, A2 => n1270, A3 => n1269, ZN => 
                           curr_proc_regs(505));
   U1928 : NAND2_X1 port map( A1 => regs(1018), A2 => n5, ZN => n1274);
   U1929 : AOI22_X1 port map( A1 => n79, A2 => regs(1530), B1 => n41, B2 => 
                           regs(506), ZN => n1273);
   U1930 : AOI22_X1 port map( A1 => n108, A2 => regs(2554), B1 => n2195, B2 => 
                           regs(2042), ZN => n1272);
   U1931 : NAND3_X1 port map( A1 => n1274, A2 => n1273, A3 => n1272, ZN => 
                           curr_proc_regs(506));
   U1932 : NAND2_X1 port map( A1 => regs(1531), A2 => n14, ZN => n1277);
   U1933 : AOI22_X1 port map( A1 => n10, A2 => regs(1019), B1 => n41, B2 => 
                           regs(507), ZN => n1276);
   U1934 : AOI22_X1 port map( A1 => n108, A2 => regs(2555), B1 => n3, B2 => 
                           regs(2043), ZN => n1275);
   U1935 : NAND3_X1 port map( A1 => n1277, A2 => n1276, A3 => n1275, ZN => 
                           curr_proc_regs(507));
   U1936 : NAND2_X1 port map( A1 => regs(1020), A2 => n5, ZN => n1280);
   U1937 : AOI22_X1 port map( A1 => n79, A2 => regs(1532), B1 => n41, B2 => 
                           regs(508), ZN => n1279);
   U1938 : AOI22_X1 port map( A1 => n108, A2 => regs(2556), B1 => n2195, B2 => 
                           regs(2044), ZN => n1278);
   U1939 : NAND3_X1 port map( A1 => n1280, A2 => n1279, A3 => n1278, ZN => 
                           curr_proc_regs(508));
   U1940 : NAND2_X1 port map( A1 => regs(1021), A2 => n5, ZN => n1283);
   U1941 : AOI22_X1 port map( A1 => n79, A2 => regs(1533), B1 => n41, B2 => 
                           regs(509), ZN => n1282);
   U1942 : AOI22_X1 port map( A1 => n108, A2 => regs(2557), B1 => n71, B2 => 
                           regs(2045), ZN => n1281);
   U1943 : NAND3_X1 port map( A1 => n1283, A2 => n1282, A3 => n1281, ZN => 
                           curr_proc_regs(509));
   U1944 : INV_X1 port map( A => regs(562), ZN => n1451);
   U1945 : AOI22_X1 port map( A1 => n108, A2 => regs(2098), B1 => n68, B2 => 
                           regs(1586), ZN => n1285);
   U1946 : AOI22_X1 port map( A1 => n90, A2 => regs(1074), B1 => n40, B2 => 
                           regs(50), ZN => n1284);
   U1947 : OAI211_X1 port map( C1 => n6, C2 => n1451, A => n1285, B => n1284, 
                           ZN => curr_proc_regs(50));
   U1948 : NAND2_X1 port map( A1 => regs(1022), A2 => n62, ZN => n1288);
   U1949 : AOI22_X1 port map( A1 => n90, A2 => regs(1534), B1 => n40, B2 => 
                           regs(510), ZN => n1287);
   U1950 : AOI22_X1 port map( A1 => n107, A2 => regs(2558), B1 => n73, B2 => 
                           regs(2046), ZN => n1286);
   U1951 : NAND3_X1 port map( A1 => n1288, A2 => n1287, A3 => n1286, ZN => 
                           curr_proc_regs(510));
   U1952 : NAND2_X1 port map( A1 => regs(1535), A2 => n14, ZN => n1291);
   U1953 : AOI22_X1 port map( A1 => n62, A2 => regs(1023), B1 => n40, B2 => 
                           regs(511), ZN => n1290);
   U1954 : AOI22_X1 port map( A1 => n107, A2 => regs(2559), B1 => n71, B2 => 
                           regs(2047), ZN => n1289);
   U1955 : NAND3_X1 port map( A1 => n1291, A2 => n1290, A3 => n1289, ZN => 
                           curr_proc_regs(511));
   U1956 : AOI22_X1 port map( A1 => n107, A2 => regs(0), B1 => n16, B2 => 
                           regs(2048), ZN => n1293);
   U1957 : AOI22_X1 port map( A1 => n58, A2 => regs(1024), B1 => n98, B2 => 
                           regs(1536), ZN => n1292);
   U1958 : OAI211_X1 port map( C1 => n1294, C2 => n21, A => n1293, B => n1292, 
                           ZN => curr_proc_regs(512));
   U1959 : AOI22_X1 port map( A1 => n107, A2 => regs(1), B1 => n16, B2 => 
                           regs(2049), ZN => n1296);
   U1960 : AOI22_X1 port map( A1 => n60, A2 => regs(1025), B1 => n98, B2 => 
                           regs(1537), ZN => n1295);
   U1961 : OAI211_X1 port map( C1 => n21, C2 => n1297, A => n1296, B => n1295, 
                           ZN => curr_proc_regs(513));
   U1962 : AOI22_X1 port map( A1 => n107, A2 => regs(2), B1 => n2195, B2 => 
                           regs(2050), ZN => n1299);
   U1963 : AOI22_X1 port map( A1 => n10, A2 => regs(1026), B1 => n98, B2 => 
                           regs(1538), ZN => n1298);
   U1964 : OAI211_X1 port map( C1 => n21, C2 => n1300, A => n1299, B => n1298, 
                           ZN => curr_proc_regs(514));
   U1965 : AOI22_X1 port map( A1 => n107, A2 => regs(3), B1 => n3, B2 => 
                           regs(2051), ZN => n1302);
   U1966 : AOI22_X1 port map( A1 => n52, A2 => regs(1027), B1 => n98, B2 => 
                           regs(1539), ZN => n1301);
   U1967 : OAI211_X1 port map( C1 => n21, C2 => n1303, A => n1302, B => n1301, 
                           ZN => curr_proc_regs(515));
   U1968 : AOI22_X1 port map( A1 => n107, A2 => regs(4), B1 => n73, B2 => 
                           regs(2052), ZN => n1305);
   U1969 : AOI22_X1 port map( A1 => n96, A2 => regs(1540), B1 => n40, B2 => 
                           regs(516), ZN => n1304);
   U1970 : OAI211_X1 port map( C1 => n64, C2 => n1306, A => n1305, B => n1304, 
                           ZN => curr_proc_regs(516));
   U1971 : INV_X1 port map( A => regs(1541), ZN => n1309);
   U1972 : AOI22_X1 port map( A1 => n107, A2 => regs(5), B1 => n16, B2 => 
                           regs(2053), ZN => n1308);
   U1973 : AOI22_X1 port map( A1 => n10, A2 => regs(1029), B1 => n40, B2 => 
                           regs(517), ZN => n1307);
   U1974 : OAI211_X1 port map( C1 => n15, C2 => n1309, A => n1308, B => n1307, 
                           ZN => curr_proc_regs(517));
   U1975 : INV_X1 port map( A => regs(1030), ZN => n1892);
   U1976 : AOI22_X1 port map( A1 => n107, A2 => regs(6), B1 => n16, B2 => 
                           regs(2054), ZN => n1311);
   U1977 : AOI22_X1 port map( A1 => n92, A2 => regs(1542), B1 => n40, B2 => 
                           regs(518), ZN => n1310);
   U1978 : OAI211_X1 port map( C1 => n67, C2 => n1892, A => n1311, B => n1310, 
                           ZN => curr_proc_regs(518));
   U1979 : INV_X1 port map( A => regs(1031), ZN => n2130);
   U1980 : AOI22_X1 port map( A1 => n107, A2 => regs(7), B1 => n78, B2 => 
                           regs(2055), ZN => n1313);
   U1981 : AOI22_X1 port map( A1 => n79, A2 => regs(1543), B1 => n40, B2 => 
                           regs(519), ZN => n1312);
   U1982 : OAI211_X1 port map( C1 => n64, C2 => n2130, A => n1313, B => n1312, 
                           ZN => curr_proc_regs(519));
   U1983 : INV_X1 port map( A => regs(563), ZN => n1454);
   U1984 : AOI22_X1 port map( A1 => n107, A2 => regs(2099), B1 => n3, B2 => 
                           regs(1587), ZN => n1315);
   U1985 : AOI22_X1 port map( A1 => n96, A2 => regs(1075), B1 => n7, B2 => 
                           regs(51), ZN => n1314);
   U1986 : OAI211_X1 port map( C1 => n64, C2 => n1454, A => n1315, B => n1314, 
                           ZN => curr_proc_regs(51));
   U1987 : INV_X1 port map( A => regs(1032), ZN => n2163);
   U1988 : AOI22_X1 port map( A1 => n106, A2 => regs(8), B1 => n3, B2 => 
                           regs(2056), ZN => n1317);
   U1989 : AOI22_X1 port map( A1 => n82, A2 => regs(1544), B1 => n25, B2 => 
                           regs(520), ZN => n1316);
   U1990 : OAI211_X1 port map( C1 => n2185, C2 => n2163, A => n1317, B => n1316
                           , ZN => curr_proc_regs(520));
   U1991 : INV_X1 port map( A => regs(1545), ZN => n1320);
   U1992 : AOI22_X1 port map( A1 => n104, A2 => regs(9), B1 => n13, B2 => 
                           regs(2057), ZN => n1319);
   U1993 : AOI22_X1 port map( A1 => n48, A2 => regs(1033), B1 => n31, B2 => 
                           regs(521), ZN => n1318);
   U1994 : OAI211_X1 port map( C1 => n99, C2 => n1320, A => n1319, B => n1318, 
                           ZN => curr_proc_regs(521));
   U1995 : AOI22_X1 port map( A1 => n105, A2 => regs(10), B1 => n3, B2 => 
                           regs(2058), ZN => n1322);
   U1996 : AOI22_X1 port map( A1 => n10, A2 => regs(1034), B1 => n98, B2 => 
                           regs(1546), ZN => n1321);
   U1997 : OAI211_X1 port map( C1 => n21, C2 => n1323, A => n1322, B => n1321, 
                           ZN => curr_proc_regs(522));
   U1998 : AOI22_X1 port map( A1 => n105, A2 => regs(11), B1 => n71, B2 => 
                           regs(2059), ZN => n1325);
   U1999 : AOI22_X1 port map( A1 => n10, A2 => regs(1035), B1 => n98, B2 => 
                           regs(1547), ZN => n1324);
   U2000 : OAI211_X1 port map( C1 => n21, C2 => n1326, A => n1325, B => n1324, 
                           ZN => curr_proc_regs(523));
   U2001 : AOI22_X1 port map( A1 => n104, A2 => regs(12), B1 => n68, B2 => 
                           regs(2060), ZN => n1328);
   U2002 : AOI22_X1 port map( A1 => n61, A2 => regs(1036), B1 => n98, B2 => 
                           regs(1548), ZN => n1327);
   U2003 : OAI211_X1 port map( C1 => n21, C2 => n1329, A => n1328, B => n1327, 
                           ZN => curr_proc_regs(524));
   U2004 : AOI22_X1 port map( A1 => n106, A2 => regs(13), B1 => n73, B2 => 
                           regs(2061), ZN => n1331);
   U2005 : AOI22_X1 port map( A1 => n56, A2 => regs(1037), B1 => n98, B2 => 
                           regs(1549), ZN => n1330);
   U2006 : OAI211_X1 port map( C1 => n21, C2 => n1332, A => n1331, B => n1330, 
                           ZN => curr_proc_regs(525));
   U2007 : AOI22_X1 port map( A1 => n104, A2 => regs(14), B1 => n68, B2 => 
                           regs(2062), ZN => n1334);
   U2008 : AOI22_X1 port map( A1 => n92, A2 => regs(1550), B1 => n31, B2 => 
                           regs(526), ZN => n1333);
   U2009 : OAI211_X1 port map( C1 => n1, C2 => n1335, A => n1334, B => n1333, 
                           ZN => curr_proc_regs(526));
   U2010 : AOI22_X1 port map( A1 => n105, A2 => regs(15), B1 => n72, B2 => 
                           regs(2063), ZN => n1337);
   U2011 : AOI22_X1 port map( A1 => n79, A2 => regs(1551), B1 => n41, B2 => 
                           regs(527), ZN => n1336);
   U2012 : OAI211_X1 port map( C1 => n6, C2 => n1338, A => n1337, B => n1336, 
                           ZN => curr_proc_regs(527));
   U2013 : AOI22_X1 port map( A1 => n106, A2 => regs(16), B1 => n73, B2 => 
                           regs(2064), ZN => n1340);
   U2014 : AOI22_X1 port map( A1 => n82, A2 => regs(1552), B1 => n41, B2 => 
                           regs(528), ZN => n1339);
   U2015 : OAI211_X1 port map( C1 => n67, C2 => n1341, A => n1340, B => n1339, 
                           ZN => curr_proc_regs(528));
   U2016 : AOI22_X1 port map( A1 => n105, A2 => regs(17), B1 => n3, B2 => 
                           regs(2065), ZN => n1343);
   U2017 : AOI22_X1 port map( A1 => n83, A2 => regs(1553), B1 => n41, B2 => 
                           regs(529), ZN => n1342);
   U2018 : OAI211_X1 port map( C1 => n64, C2 => n1344, A => n1343, B => n1342, 
                           ZN => curr_proc_regs(529));
   U2019 : INV_X1 port map( A => regs(1076), ZN => n1457);
   U2020 : AOI22_X1 port map( A1 => n106, A2 => regs(2100), B1 => n16, B2 => 
                           regs(1588), ZN => n1346);
   U2021 : AOI22_X1 port map( A1 => n56, A2 => regs(564), B1 => n41, B2 => 
                           regs(52), ZN => n1345);
   U2022 : OAI211_X1 port map( C1 => n2199, C2 => n1457, A => n1346, B => n1345
                           , ZN => curr_proc_regs(52));
   U2023 : AOI22_X1 port map( A1 => n106, A2 => regs(18), B1 => n16, B2 => 
                           regs(2066), ZN => n1348);
   U2024 : AOI22_X1 port map( A1 => n80, A2 => regs(1554), B1 => n41, B2 => 
                           regs(530), ZN => n1347);
   U2025 : OAI211_X1 port map( C1 => n2185, C2 => n1349, A => n1348, B => n1347
                           , ZN => curr_proc_regs(530));
   U2026 : AOI22_X1 port map( A1 => n106, A2 => regs(19), B1 => n2195, B2 => 
                           regs(2067), ZN => n1351);
   U2027 : AOI22_X1 port map( A1 => n56, A2 => regs(1043), B1 => n83, B2 => 
                           regs(1555), ZN => n1350);
   U2028 : OAI211_X1 port map( C1 => n21, C2 => n1352, A => n1351, B => n1350, 
                           ZN => curr_proc_regs(531));
   U2029 : AOI22_X1 port map( A1 => n106, A2 => regs(20), B1 => n3, B2 => 
                           regs(2068), ZN => n1354);
   U2030 : AOI22_X1 port map( A1 => n81, A2 => regs(1556), B1 => n41, B2 => 
                           regs(532), ZN => n1353);
   U2031 : OAI211_X1 port map( C1 => n67, C2 => n1355, A => n1354, B => n1353, 
                           ZN => curr_proc_regs(532));
   U2032 : AOI22_X1 port map( A1 => n106, A2 => regs(21), B1 => n3, B2 => 
                           regs(2069), ZN => n1357);
   U2033 : AOI22_X1 port map( A1 => n56, A2 => regs(1045), B1 => n82, B2 => 
                           regs(1557), ZN => n1356);
   U2034 : OAI211_X1 port map( C1 => n21, C2 => n1358, A => n1357, B => n1356, 
                           ZN => curr_proc_regs(533));
   U2035 : AOI22_X1 port map( A1 => n106, A2 => regs(22), B1 => n12, B2 => 
                           regs(2070), ZN => n1360);
   U2036 : AOI22_X1 port map( A1 => n56, A2 => regs(1046), B1 => n85, B2 => 
                           regs(1558), ZN => n1359);
   U2037 : OAI211_X1 port map( C1 => n21, C2 => n1361, A => n1360, B => n1359, 
                           ZN => curr_proc_regs(534));
   U2038 : AOI22_X1 port map( A1 => n106, A2 => regs(23), B1 => n3, B2 => 
                           regs(2071), ZN => n1363);
   U2039 : AOI22_X1 port map( A1 => n94, A2 => regs(1559), B1 => n41, B2 => 
                           regs(535), ZN => n1362);
   U2040 : OAI211_X1 port map( C1 => n67, C2 => n1364, A => n1363, B => n1362, 
                           ZN => curr_proc_regs(535));
   U2041 : AOI22_X1 port map( A1 => n106, A2 => regs(24), B1 => n68, B2 => 
                           regs(2072), ZN => n1366);
   U2042 : AOI22_X1 port map( A1 => n56, A2 => regs(1048), B1 => n84, B2 => 
                           regs(1560), ZN => n1365);
   U2043 : OAI211_X1 port map( C1 => n21, C2 => n1367, A => n1366, B => n1365, 
                           ZN => curr_proc_regs(536));
   U2044 : AOI22_X1 port map( A1 => n106, A2 => regs(25), B1 => n73, B2 => 
                           regs(2073), ZN => n1369);
   U2045 : AOI22_X1 port map( A1 => n84, A2 => regs(1561), B1 => n23, B2 => 
                           regs(537), ZN => n1368);
   U2046 : OAI211_X1 port map( C1 => n67, C2 => n1370, A => n1369, B => n1368, 
                           ZN => curr_proc_regs(537));
   U2047 : AOI22_X1 port map( A1 => n106, A2 => regs(26), B1 => n68, B2 => 
                           regs(2074), ZN => n1372);
   U2048 : AOI22_X1 port map( A1 => n85, A2 => regs(1562), B1 => n23, B2 => 
                           regs(538), ZN => n1371);
   U2049 : OAI211_X1 port map( C1 => n67, C2 => n1373, A => n1372, B => n1371, 
                           ZN => curr_proc_regs(538));
   U2050 : AOI22_X1 port map( A1 => n106, A2 => regs(27), B1 => n68, B2 => 
                           regs(2075), ZN => n1375);
   U2051 : AOI22_X1 port map( A1 => n86, A2 => regs(1563), B1 => n23, B2 => 
                           regs(539), ZN => n1374);
   U2052 : OAI211_X1 port map( C1 => n67, C2 => n1376, A => n1375, B => n1374, 
                           ZN => curr_proc_regs(539));
   U2053 : INV_X1 port map( A => regs(565), ZN => n1460);
   U2054 : AOI22_X1 port map( A1 => n104, A2 => regs(2101), B1 => n73, B2 => 
                           regs(1589), ZN => n1378);
   U2055 : AOI22_X1 port map( A1 => n87, A2 => regs(1077), B1 => n23, B2 => 
                           regs(53), ZN => n1377);
   U2056 : OAI211_X1 port map( C1 => n67, C2 => n1460, A => n1378, B => n1377, 
                           ZN => curr_proc_regs(53));
   U2057 : AOI22_X1 port map( A1 => n106, A2 => regs(28), B1 => n73, B2 => 
                           regs(2076), ZN => n1380);
   U2058 : AOI22_X1 port map( A1 => n50, A2 => regs(1052), B1 => n86, B2 => 
                           regs(1564), ZN => n1379);
   U2059 : OAI211_X1 port map( C1 => n21, C2 => n1381, A => n1380, B => n1379, 
                           ZN => curr_proc_regs(540));
   U2060 : AOI22_X1 port map( A1 => n104, A2 => regs(29), B1 => n68, B2 => 
                           regs(2077), ZN => n1383);
   U2061 : AOI22_X1 port map( A1 => n88, A2 => regs(1565), B1 => n23, B2 => 
                           regs(541), ZN => n1382);
   U2062 : OAI211_X1 port map( C1 => n67, C2 => n1384, A => n1383, B => n1382, 
                           ZN => curr_proc_regs(541));
   U2063 : AOI22_X1 port map( A1 => n105, A2 => regs(30), B1 => n73, B2 => 
                           regs(2078), ZN => n1386);
   U2064 : AOI22_X1 port map( A1 => n88, A2 => regs(1566), B1 => n23, B2 => 
                           regs(542), ZN => n1385);
   U2065 : OAI211_X1 port map( C1 => n66, C2 => n1387, A => n1386, B => n1385, 
                           ZN => curr_proc_regs(542));
   U2066 : AOI22_X1 port map( A1 => n105, A2 => regs(31), B1 => n71, B2 => 
                           regs(2079), ZN => n1389);
   U2067 : AOI22_X1 port map( A1 => n53, A2 => regs(1055), B1 => n96, B2 => 
                           regs(1567), ZN => n1388);
   U2068 : OAI211_X1 port map( C1 => n21, C2 => n1390, A => n1389, B => n1388, 
                           ZN => curr_proc_regs(543));
   U2069 : AOI22_X1 port map( A1 => n106, A2 => regs(32), B1 => n16, B2 => 
                           regs(2080), ZN => n1392);
   U2070 : AOI22_X1 port map( A1 => n10, A2 => regs(1056), B1 => n98, B2 => 
                           regs(1568), ZN => n1391);
   U2071 : OAI211_X1 port map( C1 => n21, C2 => n1393, A => n1392, B => n1391, 
                           ZN => curr_proc_regs(544));
   U2072 : AOI22_X1 port map( A1 => n104, A2 => regs(33), B1 => n16, B2 => 
                           regs(2081), ZN => n1395);
   U2073 : AOI22_X1 port map( A1 => n96, A2 => regs(1569), B1 => n23, B2 => 
                           regs(545), ZN => n1394);
   U2074 : OAI211_X1 port map( C1 => n2185, C2 => n1396, A => n1395, B => n1394
                           , ZN => curr_proc_regs(545));
   U2075 : AOI22_X1 port map( A1 => n105, A2 => regs(34), B1 => n73, B2 => 
                           regs(2082), ZN => n1398);
   U2076 : AOI22_X1 port map( A1 => n10, A2 => regs(1058), B1 => n80, B2 => 
                           regs(1570), ZN => n1397);
   U2077 : OAI211_X1 port map( C1 => n22, C2 => n1399, A => n1398, B => n1397, 
                           ZN => curr_proc_regs(546));
   U2078 : AOI22_X1 port map( A1 => n106, A2 => regs(35), B1 => n16, B2 => 
                           regs(2083), ZN => n1401);
   U2079 : AOI22_X1 port map( A1 => n95, A2 => regs(1571), B1 => n23, B2 => 
                           regs(547), ZN => n1400);
   U2080 : OAI211_X1 port map( C1 => n66, C2 => n1402, A => n1401, B => n1400, 
                           ZN => curr_proc_regs(547));
   U2081 : AOI22_X1 port map( A1 => n106, A2 => regs(36), B1 => n16, B2 => 
                           regs(2084), ZN => n1404);
   U2082 : AOI22_X1 port map( A1 => n90, A2 => regs(1572), B1 => n23, B2 => 
                           regs(548), ZN => n1403);
   U2083 : OAI211_X1 port map( C1 => n2185, C2 => n1405, A => n1404, B => n1403
                           , ZN => curr_proc_regs(548));
   U2084 : AOI22_X1 port map( A1 => n104, A2 => regs(37), B1 => n77, B2 => 
                           regs(2085), ZN => n1407);
   U2085 : AOI22_X1 port map( A1 => n10, A2 => regs(1061), B1 => n87, B2 => 
                           regs(1573), ZN => n1406);
   U2086 : OAI211_X1 port map( C1 => n2112, C2 => n1408, A => n1407, B => n1406
                           , ZN => curr_proc_regs(549));
   U2087 : INV_X1 port map( A => regs(1078), ZN => n1463);
   U2088 : AOI22_X1 port map( A1 => n104, A2 => regs(2102), B1 => n3, B2 => 
                           regs(1590), ZN => n1410);
   U2089 : AOI22_X1 port map( A1 => n57, A2 => regs(566), B1 => n23, B2 => 
                           regs(54), ZN => n1409);
   U2090 : OAI211_X1 port map( C1 => n99, C2 => n1463, A => n1410, B => n1409, 
                           ZN => curr_proc_regs(54));
   U2091 : AOI22_X1 port map( A1 => n105, A2 => regs(38), B1 => n3, B2 => 
                           regs(2086), ZN => n1412);
   U2092 : AOI22_X1 port map( A1 => n57, A2 => regs(1062), B1 => n85, B2 => 
                           regs(1574), ZN => n1411);
   U2093 : OAI211_X1 port map( C1 => n2112, C2 => n1413, A => n1412, B => n1411
                           , ZN => curr_proc_regs(550));
   U2094 : AOI22_X1 port map( A1 => n106, A2 => regs(39), B1 => n68, B2 => 
                           regs(2087), ZN => n1415);
   U2095 : AOI22_X1 port map( A1 => n57, A2 => regs(1063), B1 => n84, B2 => 
                           regs(1575), ZN => n1414);
   U2096 : OAI211_X1 port map( C1 => n2112, C2 => n1416, A => n1415, B => n1414
                           , ZN => curr_proc_regs(551));
   U2097 : AOI22_X1 port map( A1 => n104, A2 => regs(40), B1 => n73, B2 => 
                           regs(2088), ZN => n1418);
   U2098 : AOI22_X1 port map( A1 => n57, A2 => regs(1064), B1 => n97, B2 => 
                           regs(1576), ZN => n1417);
   U2099 : OAI211_X1 port map( C1 => n2112, C2 => n1419, A => n1418, B => n1417
                           , ZN => curr_proc_regs(552));
   U2100 : AOI22_X1 port map( A1 => n105, A2 => regs(41), B1 => n9, B2 => 
                           regs(2089), ZN => n1421);
   U2101 : AOI22_X1 port map( A1 => n92, A2 => regs(1577), B1 => n23, B2 => 
                           regs(553), ZN => n1420);
   U2102 : OAI211_X1 port map( C1 => n2185, C2 => n1422, A => n1421, B => n1420
                           , ZN => curr_proc_regs(553));
   U2103 : AOI22_X1 port map( A1 => n106, A2 => regs(42), B1 => n73, B2 => 
                           regs(2090), ZN => n1424);
   U2104 : AOI22_X1 port map( A1 => n94, A2 => regs(1578), B1 => n24, B2 => 
                           regs(554), ZN => n1423);
   U2105 : OAI211_X1 port map( C1 => n2185, C2 => n1425, A => n1424, B => n1423
                           , ZN => curr_proc_regs(554));
   U2106 : AOI22_X1 port map( A1 => n104, A2 => regs(43), B1 => n71, B2 => 
                           regs(2091), ZN => n1427);
   U2107 : AOI22_X1 port map( A1 => n95, A2 => regs(1579), B1 => n24, B2 => 
                           regs(555), ZN => n1426);
   U2108 : OAI211_X1 port map( C1 => n66, C2 => n1428, A => n1427, B => n1426, 
                           ZN => curr_proc_regs(555));
   U2109 : AOI22_X1 port map( A1 => n105, A2 => regs(44), B1 => n11, B2 => 
                           regs(2092), ZN => n1430);
   U2110 : AOI22_X1 port map( A1 => n57, A2 => regs(1068), B1 => n82, B2 => 
                           regs(1580), ZN => n1429);
   U2111 : OAI211_X1 port map( C1 => n2112, C2 => n1431, A => n1430, B => n1429
                           , ZN => curr_proc_regs(556));
   U2112 : AOI22_X1 port map( A1 => n106, A2 => regs(45), B1 => n11, B2 => 
                           regs(2093), ZN => n1433);
   U2113 : AOI22_X1 port map( A1 => n57, A2 => regs(1069), B1 => n83, B2 => 
                           regs(1581), ZN => n1432);
   U2114 : OAI211_X1 port map( C1 => n21, C2 => n1434, A => n1433, B => n1432, 
                           ZN => curr_proc_regs(557));
   U2115 : AOI22_X1 port map( A1 => n104, A2 => regs(46), B1 => n78, B2 => 
                           regs(2094), ZN => n1436);
   U2116 : AOI22_X1 port map( A1 => n56, A2 => regs(1070), B1 => n79, B2 => 
                           regs(1582), ZN => n1435);
   U2117 : OAI211_X1 port map( C1 => n21, C2 => n1437, A => n1436, B => n1435, 
                           ZN => curr_proc_regs(558));
   U2118 : AOI22_X1 port map( A1 => n105, A2 => regs(47), B1 => n11, B2 => 
                           regs(2095), ZN => n1439);
   U2119 : AOI22_X1 port map( A1 => n56, A2 => regs(1071), B1 => n80, B2 => 
                           regs(1583), ZN => n1438);
   U2120 : OAI211_X1 port map( C1 => n21, C2 => n1440, A => n1439, B => n1438, 
                           ZN => curr_proc_regs(559));
   U2121 : INV_X1 port map( A => regs(1079), ZN => n1466);
   U2122 : AOI22_X1 port map( A1 => n105, A2 => regs(2103), B1 => n11, B2 => 
                           regs(1591), ZN => n1442);
   U2123 : AOI22_X1 port map( A1 => n56, A2 => regs(567), B1 => n24, B2 => 
                           regs(55), ZN => n1441);
   U2124 : OAI211_X1 port map( C1 => n102, C2 => n1466, A => n1442, B => n1441,
                           ZN => curr_proc_regs(55));
   U2125 : AOI22_X1 port map( A1 => n105, A2 => regs(48), B1 => n3, B2 => 
                           regs(2096), ZN => n1444);
   U2126 : AOI22_X1 port map( A1 => n56, A2 => regs(1072), B1 => n81, B2 => 
                           regs(1584), ZN => n1443);
   U2127 : OAI211_X1 port map( C1 => n21, C2 => n1445, A => n1444, B => n1443, 
                           ZN => curr_proc_regs(560));
   U2128 : AOI22_X1 port map( A1 => n105, A2 => regs(49), B1 => n78, B2 => 
                           regs(2097), ZN => n1447);
   U2129 : AOI22_X1 port map( A1 => n90, A2 => regs(1585), B1 => n24, B2 => 
                           regs(561), ZN => n1446);
   U2130 : OAI211_X1 port map( C1 => n64, C2 => n1448, A => n1447, B => n1446, 
                           ZN => curr_proc_regs(561));
   U2131 : AOI22_X1 port map( A1 => n105, A2 => regs(50), B1 => n11, B2 => 
                           regs(2098), ZN => n1450);
   U2132 : AOI22_X1 port map( A1 => n56, A2 => regs(1074), B1 => n83, B2 => 
                           regs(1586), ZN => n1449);
   U2133 : OAI211_X1 port map( C1 => n21, C2 => n1451, A => n1450, B => n1449, 
                           ZN => curr_proc_regs(562));
   U2134 : AOI22_X1 port map( A1 => n105, A2 => regs(51), B1 => n11, B2 => 
                           regs(2099), ZN => n1453);
   U2135 : AOI22_X1 port map( A1 => n58, A2 => regs(1075), B1 => n79, B2 => 
                           regs(1587), ZN => n1452);
   U2136 : OAI211_X1 port map( C1 => n21, C2 => n1454, A => n1453, B => n1452, 
                           ZN => curr_proc_regs(563));
   U2137 : AOI22_X1 port map( A1 => n105, A2 => regs(52), B1 => n3, B2 => 
                           regs(2100), ZN => n1456);
   U2138 : AOI22_X1 port map( A1 => n92, A2 => regs(1588), B1 => n24, B2 => 
                           regs(564), ZN => n1455);
   U2139 : OAI211_X1 port map( C1 => n66, C2 => n1457, A => n1456, B => n1455, 
                           ZN => curr_proc_regs(564));
   U2140 : AOI22_X1 port map( A1 => n105, A2 => regs(53), B1 => n78, B2 => 
                           regs(2101), ZN => n1459);
   U2141 : AOI22_X1 port map( A1 => n58, A2 => regs(1077), B1 => n81, B2 => 
                           regs(1589), ZN => n1458);
   U2142 : OAI211_X1 port map( C1 => n21, C2 => n1460, A => n1459, B => n1458, 
                           ZN => curr_proc_regs(565));
   U2143 : AOI22_X1 port map( A1 => n105, A2 => regs(54), B1 => n3, B2 => 
                           regs(2102), ZN => n1462);
   U2144 : AOI22_X1 port map( A1 => n94, A2 => regs(1590), B1 => n24, B2 => 
                           regs(566), ZN => n1461);
   U2145 : OAI211_X1 port map( C1 => n66, C2 => n1463, A => n1462, B => n1461, 
                           ZN => curr_proc_regs(566));
   U2146 : AOI22_X1 port map( A1 => n105, A2 => regs(55), B1 => n78, B2 => 
                           regs(2103), ZN => n1465);
   U2147 : AOI22_X1 port map( A1 => n95, A2 => regs(1591), B1 => n24, B2 => 
                           regs(567), ZN => n1464);
   U2148 : OAI211_X1 port map( C1 => n66, C2 => n1466, A => n1465, B => n1464, 
                           ZN => curr_proc_regs(567));
   U2149 : INV_X1 port map( A => regs(1592), ZN => n1469);
   U2150 : AOI22_X1 port map( A1 => n105, A2 => regs(56), B1 => n11, B2 => 
                           regs(2104), ZN => n1468);
   U2151 : AOI22_X1 port map( A1 => n58, A2 => regs(1080), B1 => n24, B2 => 
                           regs(568), ZN => n1467);
   U2152 : OAI211_X1 port map( C1 => n15, C2 => n1469, A => n1468, B => n1467, 
                           ZN => curr_proc_regs(568));
   U2153 : INV_X1 port map( A => regs(1593), ZN => n1472);
   U2154 : AOI22_X1 port map( A1 => n105, A2 => regs(57), B1 => n11, B2 => 
                           regs(2105), ZN => n1471);
   U2155 : AOI22_X1 port map( A1 => n58, A2 => regs(1081), B1 => n24, B2 => 
                           regs(569), ZN => n1470);
   U2156 : OAI211_X1 port map( C1 => n2199, C2 => n1472, A => n1471, B => n1470
                           , ZN => curr_proc_regs(569));
   U2157 : INV_X1 port map( A => regs(1080), ZN => n1475);
   U2158 : AOI22_X1 port map( A1 => n104, A2 => regs(2104), B1 => n11, B2 => 
                           regs(1592), ZN => n1474);
   U2159 : AOI22_X1 port map( A1 => n58, A2 => regs(568), B1 => n24, B2 => 
                           regs(56), ZN => n1473);
   U2160 : OAI211_X1 port map( C1 => n99, C2 => n1475, A => n1474, B => n1473, 
                           ZN => curr_proc_regs(56));
   U2161 : INV_X1 port map( A => regs(1594), ZN => n1478);
   U2162 : AOI22_X1 port map( A1 => n104, A2 => regs(58), B1 => n16, B2 => 
                           regs(2106), ZN => n1477);
   U2163 : AOI22_X1 port map( A1 => n58, A2 => regs(1082), B1 => n24, B2 => 
                           regs(570), ZN => n1476);
   U2164 : OAI211_X1 port map( C1 => n102, C2 => n1478, A => n1477, B => n1476,
                           ZN => curr_proc_regs(570));
   U2165 : INV_X1 port map( A => regs(1595), ZN => n1481);
   U2166 : AOI22_X1 port map( A1 => n104, A2 => regs(59), B1 => n78, B2 => 
                           regs(2107), ZN => n1480);
   U2167 : AOI22_X1 port map( A1 => n57, A2 => regs(1083), B1 => n31, B2 => 
                           regs(571), ZN => n1479);
   U2168 : OAI211_X1 port map( C1 => n15, C2 => n1481, A => n1480, B => n1479, 
                           ZN => curr_proc_regs(571));
   U2169 : INV_X1 port map( A => regs(1084), ZN => n1593);
   U2170 : AOI22_X1 port map( A1 => n104, A2 => regs(60), B1 => n11, B2 => 
                           regs(2108), ZN => n1483);
   U2171 : AOI22_X1 port map( A1 => n90, A2 => regs(1596), B1 => n29, B2 => 
                           regs(572), ZN => n1482);
   U2172 : OAI211_X1 port map( C1 => n2185, C2 => n1593, A => n1483, B => n1482
                           , ZN => curr_proc_regs(572));
   U2173 : INV_X1 port map( A => regs(1597), ZN => n1486);
   U2174 : AOI22_X1 port map( A1 => n104, A2 => regs(61), B1 => n11, B2 => 
                           regs(2109), ZN => n1485);
   U2175 : AOI22_X1 port map( A1 => n57, A2 => regs(1085), B1 => n38, B2 => 
                           regs(573), ZN => n1484);
   U2176 : OAI211_X1 port map( C1 => n15, C2 => n1486, A => n1485, B => n1484, 
                           ZN => curr_proc_regs(573));
   U2177 : INV_X1 port map( A => regs(1598), ZN => n1489);
   U2178 : AOI22_X1 port map( A1 => n104, A2 => regs(62), B1 => n11, B2 => 
                           regs(2110), ZN => n1488);
   U2179 : AOI22_X1 port map( A1 => n57, A2 => regs(1086), B1 => n41, B2 => 
                           regs(574), ZN => n1487);
   U2180 : OAI211_X1 port map( C1 => n100, C2 => n1489, A => n1488, B => n1487,
                           ZN => curr_proc_regs(574));
   U2181 : INV_X1 port map( A => regs(1599), ZN => n1492);
   U2182 : AOI22_X1 port map( A1 => n104, A2 => regs(63), B1 => n16, B2 => 
                           regs(2111), ZN => n1491);
   U2183 : AOI22_X1 port map( A1 => n57, A2 => regs(1087), B1 => n2, B2 => 
                           regs(575), ZN => n1490);
   U2184 : OAI211_X1 port map( C1 => n100, C2 => n1492, A => n1491, B => n1490,
                           ZN => curr_proc_regs(575));
   U2185 : INV_X1 port map( A => regs(1088), ZN => n1724);
   U2186 : AOI22_X1 port map( A1 => n104, A2 => regs(64), B1 => n11, B2 => 
                           regs(2112), ZN => n1494);
   U2187 : AOI22_X1 port map( A1 => n92, A2 => regs(1600), B1 => n2, B2 => 
                           regs(576), ZN => n1493);
   U2188 : OAI211_X1 port map( C1 => n66, C2 => n1724, A => n1494, B => n1493, 
                           ZN => curr_proc_regs(576));
   U2189 : INV_X1 port map( A => regs(1601), ZN => n1497);
   U2190 : AOI22_X1 port map( A1 => n104, A2 => regs(65), B1 => n11, B2 => 
                           regs(2113), ZN => n1496);
   U2191 : AOI22_X1 port map( A1 => n57, A2 => regs(1089), B1 => n7, B2 => 
                           regs(577), ZN => n1495);
   U2192 : OAI211_X1 port map( C1 => n100, C2 => n1497, A => n1496, B => n1495,
                           ZN => curr_proc_regs(577));
   U2193 : INV_X1 port map( A => regs(1090), ZN => n1790);
   U2194 : AOI22_X1 port map( A1 => n104, A2 => regs(66), B1 => n11, B2 => 
                           regs(2114), ZN => n1499);
   U2195 : AOI22_X1 port map( A1 => n79, A2 => regs(1602), B1 => n7, B2 => 
                           regs(578), ZN => n1498);
   U2196 : OAI211_X1 port map( C1 => n66, C2 => n1790, A => n1499, B => n1498, 
                           ZN => curr_proc_regs(578));
   U2197 : INV_X1 port map( A => regs(1603), ZN => n1502);
   U2198 : AOI22_X1 port map( A1 => n104, A2 => regs(67), B1 => n11, B2 => 
                           regs(2115), ZN => n1501);
   U2199 : AOI22_X1 port map( A1 => n59, A2 => regs(1091), B1 => n25, B2 => 
                           regs(579), ZN => n1500);
   U2200 : OAI211_X1 port map( C1 => n100, C2 => n1502, A => n1501, B => n1500,
                           ZN => curr_proc_regs(579));
   U2201 : INV_X1 port map( A => regs(569), ZN => n1505);
   U2202 : AOI22_X1 port map( A1 => n19, A2 => regs(2105), B1 => n11, B2 => 
                           regs(1593), ZN => n1504);
   U2203 : AOI22_X1 port map( A1 => n89, A2 => regs(1081), B1 => n31, B2 => 
                           regs(57), ZN => n1503);
   U2204 : OAI211_X1 port map( C1 => n2185, C2 => n1505, A => n1504, B => n1503
                           , ZN => curr_proc_regs(57));
   U2205 : INV_X1 port map( A => regs(1604), ZN => n1508);
   U2206 : AOI22_X1 port map( A1 => n19, A2 => regs(68), B1 => n11, B2 => 
                           regs(2116), ZN => n1507);
   U2207 : AOI22_X1 port map( A1 => n59, A2 => regs(1092), B1 => n29, B2 => 
                           regs(580), ZN => n1506);
   U2208 : OAI211_X1 port map( C1 => n100, C2 => n1508, A => n1507, B => n1506,
                           ZN => curr_proc_regs(580));
   U2209 : INV_X1 port map( A => regs(1605), ZN => n1511);
   U2210 : AOI22_X1 port map( A1 => n19, A2 => regs(69), B1 => n11, B2 => 
                           regs(2117), ZN => n1510);
   U2211 : AOI22_X1 port map( A1 => n59, A2 => regs(1093), B1 => n25, B2 => 
                           regs(581), ZN => n1509);
   U2212 : OAI211_X1 port map( C1 => n100, C2 => n1511, A => n1510, B => n1509,
                           ZN => curr_proc_regs(581));
   U2213 : INV_X1 port map( A => regs(1094), ZN => n1925);
   U2214 : AOI22_X1 port map( A1 => n19, A2 => regs(70), B1 => n11, B2 => 
                           regs(2118), ZN => n1513);
   U2215 : AOI22_X1 port map( A1 => n89, A2 => regs(1606), B1 => n25, B2 => 
                           regs(582), ZN => n1512);
   U2216 : OAI211_X1 port map( C1 => n2185, C2 => n1925, A => n1513, B => n1512
                           , ZN => curr_proc_regs(582));
   U2217 : INV_X1 port map( A => regs(1607), ZN => n1516);
   U2218 : AOI22_X1 port map( A1 => n19, A2 => regs(71), B1 => n11, B2 => 
                           regs(2119), ZN => n1515);
   U2219 : AOI22_X1 port map( A1 => n59, A2 => regs(1095), B1 => n25, B2 => 
                           regs(583), ZN => n1514);
   U2220 : OAI211_X1 port map( C1 => n100, C2 => n1516, A => n1515, B => n1514,
                           ZN => curr_proc_regs(583));
   U2221 : INV_X1 port map( A => regs(1096), ZN => n1991);
   U2222 : AOI22_X1 port map( A1 => n19, A2 => regs(72), B1 => n11, B2 => 
                           regs(2120), ZN => n1518);
   U2223 : AOI22_X1 port map( A1 => n89, A2 => regs(1608), B1 => n25, B2 => 
                           regs(584), ZN => n1517);
   U2224 : OAI211_X1 port map( C1 => n66, C2 => n1991, A => n1518, B => n1517, 
                           ZN => curr_proc_regs(584));
   U2225 : INV_X1 port map( A => regs(1097), ZN => n2024);
   U2226 : AOI22_X1 port map( A1 => n19, A2 => regs(73), B1 => n11, B2 => 
                           regs(2121), ZN => n1520);
   U2227 : AOI22_X1 port map( A1 => n89, A2 => regs(1609), B1 => n25, B2 => 
                           regs(585), ZN => n1519);
   U2228 : OAI211_X1 port map( C1 => n66, C2 => n2024, A => n1520, B => n1519, 
                           ZN => curr_proc_regs(585));
   U2229 : INV_X1 port map( A => regs(1098), ZN => n2057);
   U2230 : AOI22_X1 port map( A1 => n19, A2 => regs(74), B1 => n11, B2 => 
                           regs(2122), ZN => n1522);
   U2231 : AOI22_X1 port map( A1 => n89, A2 => regs(1610), B1 => n25, B2 => 
                           regs(586), ZN => n1521);
   U2232 : OAI211_X1 port map( C1 => n2185, C2 => n2057, A => n1522, B => n1521
                           , ZN => curr_proc_regs(586));
   U2233 : INV_X1 port map( A => regs(1611), ZN => n1525);
   U2234 : AOI22_X1 port map( A1 => n19, A2 => regs(75), B1 => n78, B2 => 
                           regs(2123), ZN => n1524);
   U2235 : AOI22_X1 port map( A1 => n59, A2 => regs(1099), B1 => n25, B2 => 
                           regs(587), ZN => n1523);
   U2236 : OAI211_X1 port map( C1 => n99, C2 => n1525, A => n1524, B => n1523, 
                           ZN => curr_proc_regs(587));
   U2237 : INV_X1 port map( A => regs(1100), ZN => n2118);
   U2238 : AOI22_X1 port map( A1 => n19, A2 => regs(76), B1 => n68, B2 => 
                           regs(2124), ZN => n1527);
   U2239 : AOI22_X1 port map( A1 => n89, A2 => regs(1612), B1 => n25, B2 => 
                           regs(588), ZN => n1526);
   U2240 : OAI211_X1 port map( C1 => n66, C2 => n2118, A => n1527, B => n1526, 
                           ZN => curr_proc_regs(588));
   U2241 : INV_X1 port map( A => regs(1613), ZN => n1530);
   U2242 : AOI22_X1 port map( A1 => n19, A2 => regs(77), B1 => n78, B2 => 
                           regs(2125), ZN => n1529);
   U2243 : AOI22_X1 port map( A1 => n59, A2 => regs(1101), B1 => n25, B2 => 
                           regs(589), ZN => n1528);
   U2244 : OAI211_X1 port map( C1 => n2199, C2 => n1530, A => n1529, B => n1528
                           , ZN => curr_proc_regs(589));
   U2245 : INV_X1 port map( A => regs(570), ZN => n1533);
   U2246 : AOI22_X1 port map( A1 => n19, A2 => regs(2106), B1 => n73, B2 => 
                           regs(1594), ZN => n1532);
   U2247 : AOI22_X1 port map( A1 => n89, A2 => regs(1082), B1 => n25, B2 => 
                           regs(58), ZN => n1531);
   U2248 : OAI211_X1 port map( C1 => n66, C2 => n1533, A => n1532, B => n1531, 
                           ZN => curr_proc_regs(58));
   U2249 : INV_X1 port map( A => regs(1102), ZN => n2124);
   U2250 : AOI22_X1 port map( A1 => n19, A2 => regs(78), B1 => n11, B2 => 
                           regs(2126), ZN => n1535);
   U2251 : AOI22_X1 port map( A1 => n89, A2 => regs(1614), B1 => n25, B2 => 
                           regs(590), ZN => n1534);
   U2252 : OAI211_X1 port map( C1 => n66, C2 => n2124, A => n1535, B => n1534, 
                           ZN => curr_proc_regs(590));
   U2253 : INV_X1 port map( A => regs(1103), ZN => n2127);
   U2254 : AOI22_X1 port map( A1 => n19, A2 => regs(79), B1 => n11, B2 => 
                           regs(2127), ZN => n1537);
   U2255 : AOI22_X1 port map( A1 => n88, A2 => regs(1615), B1 => n26, B2 => 
                           regs(591), ZN => n1536);
   U2256 : OAI211_X1 port map( C1 => n66, C2 => n2127, A => n1537, B => n1536, 
                           ZN => curr_proc_regs(591));
   U2257 : INV_X1 port map( A => regs(1104), ZN => n2133);
   U2258 : AOI22_X1 port map( A1 => n19, A2 => regs(80), B1 => n78, B2 => 
                           regs(2128), ZN => n1539);
   U2259 : AOI22_X1 port map( A1 => n88, A2 => regs(1616), B1 => n26, B2 => 
                           regs(592), ZN => n1538);
   U2260 : OAI211_X1 port map( C1 => n66, C2 => n2133, A => n1539, B => n1538, 
                           ZN => curr_proc_regs(592));
   U2261 : INV_X1 port map( A => regs(1105), ZN => n2136);
   U2262 : AOI22_X1 port map( A1 => n19, A2 => regs(81), B1 => n3, B2 => 
                           regs(2129), ZN => n1541);
   U2263 : AOI22_X1 port map( A1 => n88, A2 => regs(1617), B1 => n26, B2 => 
                           regs(593), ZN => n1540);
   U2264 : OAI211_X1 port map( C1 => n66, C2 => n2136, A => n1541, B => n1540, 
                           ZN => curr_proc_regs(593));
   U2265 : INV_X1 port map( A => regs(1618), ZN => n1544);
   U2266 : AOI22_X1 port map( A1 => n19, A2 => regs(82), B1 => n78, B2 => 
                           regs(2130), ZN => n1543);
   U2267 : AOI22_X1 port map( A1 => n59, A2 => regs(1106), B1 => n26, B2 => 
                           regs(594), ZN => n1542);
   U2268 : OAI211_X1 port map( C1 => n99, C2 => n1544, A => n1543, B => n1542, 
                           ZN => curr_proc_regs(594));
   U2269 : INV_X1 port map( A => regs(1619), ZN => n1547);
   U2270 : AOI22_X1 port map( A1 => n19, A2 => regs(83), B1 => n11, B2 => 
                           regs(2131), ZN => n1546);
   U2271 : AOI22_X1 port map( A1 => n58, A2 => regs(1107), B1 => n26, B2 => 
                           regs(595), ZN => n1545);
   U2272 : OAI211_X1 port map( C1 => n99, C2 => n1547, A => n1546, B => n1545, 
                           ZN => curr_proc_regs(595));
   U2273 : INV_X1 port map( A => regs(1620), ZN => n1550);
   U2274 : AOI22_X1 port map( A1 => n19, A2 => regs(84), B1 => n11, B2 => 
                           regs(2132), ZN => n1549);
   U2275 : AOI22_X1 port map( A1 => n58, A2 => regs(1108), B1 => n26, B2 => 
                           regs(596), ZN => n1548);
   U2276 : OAI211_X1 port map( C1 => n101, C2 => n1550, A => n1549, B => n1548,
                           ZN => curr_proc_regs(596));
   U2277 : INV_X1 port map( A => regs(1621), ZN => n1553);
   U2278 : AOI22_X1 port map( A1 => n19, A2 => regs(85), B1 => n11, B2 => 
                           regs(2133), ZN => n1552);
   U2279 : AOI22_X1 port map( A1 => n58, A2 => regs(1109), B1 => n26, B2 => 
                           regs(597), ZN => n1551);
   U2280 : OAI211_X1 port map( C1 => n15, C2 => n1553, A => n1552, B => n1551, 
                           ZN => curr_proc_regs(597));
   U2281 : INV_X1 port map( A => regs(1110), ZN => n2151);
   U2282 : AOI22_X1 port map( A1 => n19, A2 => regs(86), B1 => n3, B2 => 
                           regs(2134), ZN => n1555);
   U2283 : AOI22_X1 port map( A1 => n88, A2 => regs(1622), B1 => n26, B2 => 
                           regs(598), ZN => n1554);
   U2284 : OAI211_X1 port map( C1 => n66, C2 => n2151, A => n1555, B => n1554, 
                           ZN => curr_proc_regs(598));
   U2285 : INV_X1 port map( A => regs(1111), ZN => n2154);
   U2286 : AOI22_X1 port map( A1 => n19, A2 => regs(87), B1 => n78, B2 => 
                           regs(2135), ZN => n1557);
   U2287 : AOI22_X1 port map( A1 => n88, A2 => regs(1623), B1 => n26, B2 => 
                           regs(599), ZN => n1556);
   U2288 : OAI211_X1 port map( C1 => n66, C2 => n2154, A => n1557, B => n1556, 
                           ZN => curr_proc_regs(599));
   U2289 : INV_X1 port map( A => regs(571), ZN => n1560);
   U2290 : AOI22_X1 port map( A1 => n4, A2 => regs(2107), B1 => n78, B2 => 
                           regs(1595), ZN => n1559);
   U2291 : AOI22_X1 port map( A1 => n88, A2 => regs(1083), B1 => n26, B2 => 
                           regs(59), ZN => n1558);
   U2292 : OAI211_X1 port map( C1 => n67, C2 => n1560, A => n1559, B => n1558, 
                           ZN => curr_proc_regs(59));
   U2293 : INV_X1 port map( A => regs(517), ZN => n1563);
   U2294 : AOI22_X1 port map( A1 => n4, A2 => regs(2053), B1 => n11, B2 => 
                           regs(1541), ZN => n1562);
   U2295 : AOI22_X1 port map( A1 => n88, A2 => regs(1029), B1 => n26, B2 => 
                           regs(5), ZN => n1561);
   U2296 : OAI211_X1 port map( C1 => n65, C2 => n1563, A => n1562, B => n1561, 
                           ZN => curr_proc_regs(5));
   U2297 : INV_X1 port map( A => regs(1112), ZN => n2157);
   U2298 : AOI22_X1 port map( A1 => n4, A2 => regs(88), B1 => n11, B2 => 
                           regs(2136), ZN => n1565);
   U2299 : AOI22_X1 port map( A1 => n88, A2 => regs(1624), B1 => n27, B2 => 
                           regs(600), ZN => n1564);
   U2300 : OAI211_X1 port map( C1 => n65, C2 => n2157, A => n1565, B => n1564, 
                           ZN => curr_proc_regs(600));
   U2301 : INV_X1 port map( A => regs(1625), ZN => n1568);
   U2302 : AOI22_X1 port map( A1 => n4, A2 => regs(89), B1 => n11, B2 => 
                           regs(2137), ZN => n1567);
   U2303 : AOI22_X1 port map( A1 => n51, A2 => regs(1113), B1 => n27, B2 => 
                           regs(601), ZN => n1566);
   U2304 : OAI211_X1 port map( C1 => n99, C2 => n1568, A => n1567, B => n1566, 
                           ZN => curr_proc_regs(601));
   U2305 : INV_X1 port map( A => regs(1626), ZN => n1571);
   U2306 : AOI22_X1 port map( A1 => n4, A2 => regs(90), B1 => n11, B2 => 
                           regs(2138), ZN => n1570);
   U2307 : AOI22_X1 port map( A1 => n8, A2 => regs(1114), B1 => n27, B2 => 
                           regs(602), ZN => n1569);
   U2308 : OAI211_X1 port map( C1 => n102, C2 => n1571, A => n1570, B => n1569,
                           ZN => curr_proc_regs(602));
   U2309 : INV_X1 port map( A => regs(1627), ZN => n1574);
   U2310 : AOI22_X1 port map( A1 => n4, A2 => regs(91), B1 => n78, B2 => 
                           regs(2139), ZN => n1573);
   U2311 : AOI22_X1 port map( A1 => n10, A2 => regs(1115), B1 => n27, B2 => 
                           regs(603), ZN => n1572);
   U2312 : OAI211_X1 port map( C1 => n100, C2 => n1574, A => n1573, B => n1572,
                           ZN => curr_proc_regs(603));
   U2313 : INV_X1 port map( A => regs(1116), ZN => n2172);
   U2314 : AOI22_X1 port map( A1 => n4, A2 => regs(92), B1 => n78, B2 => 
                           regs(2140), ZN => n1576);
   U2315 : AOI22_X1 port map( A1 => n88, A2 => regs(1628), B1 => n27, B2 => 
                           regs(604), ZN => n1575);
   U2316 : OAI211_X1 port map( C1 => n65, C2 => n2172, A => n1576, B => n1575, 
                           ZN => curr_proc_regs(604));
   U2317 : INV_X1 port map( A => regs(1629), ZN => n1579);
   U2318 : AOI22_X1 port map( A1 => n4, A2 => regs(93), B1 => n3, B2 => 
                           regs(2141), ZN => n1578);
   U2319 : AOI22_X1 port map( A1 => n8, A2 => regs(1117), B1 => n27, B2 => 
                           regs(605), ZN => n1577);
   U2320 : OAI211_X1 port map( C1 => n101, C2 => n1579, A => n1578, B => n1577,
                           ZN => curr_proc_regs(605));
   U2321 : INV_X1 port map( A => regs(1630), ZN => n1582);
   U2322 : AOI22_X1 port map( A1 => n4, A2 => regs(94), B1 => n78, B2 => 
                           regs(2142), ZN => n1581);
   U2323 : AOI22_X1 port map( A1 => n8, A2 => regs(1118), B1 => n27, B2 => 
                           regs(606), ZN => n1580);
   U2324 : OAI211_X1 port map( C1 => n100, C2 => n1582, A => n1581, B => n1580,
                           ZN => curr_proc_regs(606));
   U2325 : INV_X1 port map( A => regs(1119), ZN => n2181);
   U2326 : AOI22_X1 port map( A1 => n4, A2 => regs(95), B1 => n78, B2 => 
                           regs(2143), ZN => n1584);
   U2327 : AOI22_X1 port map( A1 => n88, A2 => regs(1631), B1 => n27, B2 => 
                           regs(607), ZN => n1583);
   U2328 : OAI211_X1 port map( C1 => n65, C2 => n2181, A => n1584, B => n1583, 
                           ZN => curr_proc_regs(607));
   U2329 : INV_X1 port map( A => regs(1632), ZN => n1587);
   U2330 : AOI22_X1 port map( A1 => n4, A2 => regs(96), B1 => n78, B2 => 
                           regs(2144), ZN => n1586);
   U2331 : AOI22_X1 port map( A1 => n8, A2 => regs(1120), B1 => n27, B2 => 
                           regs(608), ZN => n1585);
   U2332 : OAI211_X1 port map( C1 => n102, C2 => n1587, A => n1586, B => n1585,
                           ZN => curr_proc_regs(608));
   U2333 : INV_X1 port map( A => regs(1633), ZN => n1590);
   U2334 : AOI22_X1 port map( A1 => n103, A2 => regs(97), B1 => n78, B2 => 
                           regs(2145), ZN => n1589);
   U2335 : AOI22_X1 port map( A1 => n8, A2 => regs(1121), B1 => n27, B2 => 
                           regs(609), ZN => n1588);
   U2336 : OAI211_X1 port map( C1 => n100, C2 => n1590, A => n1589, B => n1588,
                           ZN => curr_proc_regs(609));
   U2337 : AOI22_X1 port map( A1 => n103, A2 => regs(2108), B1 => n78, B2 => 
                           regs(1596), ZN => n1592);
   U2338 : AOI22_X1 port map( A1 => n8, A2 => regs(572), B1 => n27, B2 => 
                           regs(60), ZN => n1591);
   U2339 : OAI211_X1 port map( C1 => n100, C2 => n1593, A => n1592, B => n1591,
                           ZN => curr_proc_regs(60));
   U2340 : INV_X1 port map( A => regs(1634), ZN => n1596);
   U2341 : AOI22_X1 port map( A1 => n103, A2 => regs(98), B1 => n11, B2 => 
                           regs(2146), ZN => n1595);
   U2342 : AOI22_X1 port map( A1 => n59, A2 => regs(1122), B1 => n28, B2 => 
                           regs(610), ZN => n1594);
   U2343 : OAI211_X1 port map( C1 => n15, C2 => n1596, A => n1595, B => n1594, 
                           ZN => curr_proc_regs(610));
   U2344 : INV_X1 port map( A => regs(1123), ZN => n2194);
   U2345 : AOI22_X1 port map( A1 => n103, A2 => regs(99), B1 => n11, B2 => 
                           regs(2147), ZN => n1598);
   U2346 : AOI22_X1 port map( A1 => n88, A2 => regs(1635), B1 => n28, B2 => 
                           regs(611), ZN => n1597);
   U2347 : OAI211_X1 port map( C1 => n65, C2 => n2194, A => n1598, B => n1597, 
                           ZN => curr_proc_regs(611));
   U2348 : AOI22_X1 port map( A1 => n103, A2 => regs(100), B1 => n78, B2 => 
                           regs(2148), ZN => n1600);
   U2349 : AOI22_X1 port map( A1 => n87, A2 => regs(1636), B1 => n28, B2 => 
                           regs(612), ZN => n1599);
   U2350 : OAI211_X1 port map( C1 => n65, C2 => n1601, A => n1600, B => n1599, 
                           ZN => curr_proc_regs(612));
   U2351 : AOI22_X1 port map( A1 => n103, A2 => regs(101), B1 => n78, B2 => 
                           regs(2149), ZN => n1603);
   U2352 : AOI22_X1 port map( A1 => n8, A2 => regs(1125), B1 => n98, B2 => 
                           regs(1637), ZN => n1602);
   U2353 : OAI211_X1 port map( C1 => n21, C2 => n1604, A => n1603, B => n1602, 
                           ZN => curr_proc_regs(613));
   U2354 : AOI22_X1 port map( A1 => n103, A2 => regs(102), B1 => n78, B2 => 
                           regs(2150), ZN => n1606);
   U2355 : AOI22_X1 port map( A1 => n8, A2 => regs(1126), B1 => n98, B2 => 
                           regs(1638), ZN => n1605);
   U2356 : OAI211_X1 port map( C1 => n21, C2 => n1607, A => n1606, B => n1605, 
                           ZN => curr_proc_regs(614));
   U2357 : AOI22_X1 port map( A1 => n103, A2 => regs(103), B1 => n9, B2 => 
                           regs(2151), ZN => n1609);
   U2358 : AOI22_X1 port map( A1 => n57, A2 => regs(1127), B1 => n98, B2 => 
                           regs(1639), ZN => n1608);
   U2359 : OAI211_X1 port map( C1 => n21, C2 => n1610, A => n1609, B => n1608, 
                           ZN => curr_proc_regs(615));
   U2360 : AOI22_X1 port map( A1 => n103, A2 => regs(104), B1 => n9, B2 => 
                           regs(2152), ZN => n1612);
   U2361 : AOI22_X1 port map( A1 => n8, A2 => regs(1128), B1 => n88, B2 => 
                           regs(1640), ZN => n1611);
   U2362 : OAI211_X1 port map( C1 => n21, C2 => n1613, A => n1612, B => n1611, 
                           ZN => curr_proc_regs(616));
   U2363 : AOI22_X1 port map( A1 => n106, A2 => regs(105), B1 => n9, B2 => 
                           regs(2153), ZN => n1615);
   U2364 : AOI22_X1 port map( A1 => n8, A2 => regs(1129), B1 => n86, B2 => 
                           regs(1641), ZN => n1614);
   U2365 : OAI211_X1 port map( C1 => n2112, C2 => n1616, A => n1615, B => n1614
                           , ZN => curr_proc_regs(617));
   U2366 : AOI22_X1 port map( A1 => n113, A2 => regs(106), B1 => n9, B2 => 
                           regs(2154), ZN => n1618);
   U2367 : AOI22_X1 port map( A1 => n8, A2 => regs(1130), B1 => n84, B2 => 
                           regs(1642), ZN => n1617);
   U2368 : OAI211_X1 port map( C1 => n21, C2 => n1619, A => n1618, B => n1617, 
                           ZN => curr_proc_regs(618));
   U2369 : AOI22_X1 port map( A1 => n113, A2 => regs(107), B1 => n9, B2 => 
                           regs(2155), ZN => n1621);
   U2370 : AOI22_X1 port map( A1 => n87, A2 => regs(1643), B1 => n28, B2 => 
                           regs(619), ZN => n1620);
   U2371 : OAI211_X1 port map( C1 => n65, C2 => n1622, A => n1621, B => n1620, 
                           ZN => curr_proc_regs(619));
   U2372 : INV_X1 port map( A => regs(1085), ZN => n1625);
   U2373 : AOI22_X1 port map( A1 => n113, A2 => regs(2109), B1 => n9, B2 => 
                           regs(1597), ZN => n1624);
   U2374 : AOI22_X1 port map( A1 => n8, A2 => regs(573), B1 => n28, B2 => 
                           regs(61), ZN => n1623);
   U2375 : OAI211_X1 port map( C1 => n15, C2 => n1625, A => n1624, B => n1623, 
                           ZN => curr_proc_regs(61));
   U2376 : AOI22_X1 port map( A1 => n113, A2 => regs(108), B1 => n9, B2 => 
                           regs(2156), ZN => n1627);
   U2377 : AOI22_X1 port map( A1 => n8, A2 => regs(1132), B1 => n85, B2 => 
                           regs(1644), ZN => n1626);
   U2378 : OAI211_X1 port map( C1 => n21, C2 => n1628, A => n1627, B => n1626, 
                           ZN => curr_proc_regs(620));
   U2379 : AOI22_X1 port map( A1 => n113, A2 => regs(109), B1 => n9, B2 => 
                           regs(2157), ZN => n1630);
   U2380 : AOI22_X1 port map( A1 => n87, A2 => regs(1645), B1 => n28, B2 => 
                           regs(621), ZN => n1629);
   U2381 : OAI211_X1 port map( C1 => n1, C2 => n1631, A => n1630, B => n1629, 
                           ZN => curr_proc_regs(621));
   U2382 : AOI22_X1 port map( A1 => n113, A2 => regs(110), B1 => n9, B2 => 
                           regs(2158), ZN => n1633);
   U2383 : AOI22_X1 port map( A1 => n8, A2 => regs(1134), B1 => n82, B2 => 
                           regs(1646), ZN => n1632);
   U2384 : OAI211_X1 port map( C1 => n21, C2 => n1634, A => n1633, B => n1632, 
                           ZN => curr_proc_regs(622));
   U2385 : AOI22_X1 port map( A1 => n113, A2 => regs(111), B1 => n9, B2 => 
                           regs(2159), ZN => n1636);
   U2386 : AOI22_X1 port map( A1 => n8, A2 => regs(1135), B1 => n83, B2 => 
                           regs(1647), ZN => n1635);
   U2387 : OAI211_X1 port map( C1 => n21, C2 => n1637, A => n1636, B => n1635, 
                           ZN => curr_proc_regs(623));
   U2388 : AOI22_X1 port map( A1 => n113, A2 => regs(112), B1 => n9, B2 => 
                           regs(2160), ZN => n1639);
   U2389 : AOI22_X1 port map( A1 => n8, A2 => regs(1136), B1 => n97, B2 => 
                           regs(1648), ZN => n1638);
   U2390 : OAI211_X1 port map( C1 => n21, C2 => n1640, A => n1639, B => n1638, 
                           ZN => curr_proc_regs(624));
   U2391 : AOI22_X1 port map( A1 => n113, A2 => regs(113), B1 => n9, B2 => 
                           regs(2161), ZN => n1642);
   U2392 : AOI22_X1 port map( A1 => n8, A2 => regs(1137), B1 => n79, B2 => 
                           regs(1649), ZN => n1641);
   U2393 : OAI211_X1 port map( C1 => n21, C2 => n1643, A => n1642, B => n1641, 
                           ZN => curr_proc_regs(625));
   U2394 : AOI22_X1 port map( A1 => n113, A2 => regs(114), B1 => n77, B2 => 
                           regs(2162), ZN => n1645);
   U2395 : AOI22_X1 port map( A1 => n8, A2 => regs(1138), B1 => n98, B2 => 
                           regs(1650), ZN => n1644);
   U2396 : OAI211_X1 port map( C1 => n21, C2 => n1646, A => n1645, B => n1644, 
                           ZN => curr_proc_regs(626));
   U2397 : AOI22_X1 port map( A1 => n113, A2 => regs(115), B1 => n9, B2 => 
                           regs(2163), ZN => n1648);
   U2398 : AOI22_X1 port map( A1 => n8, A2 => regs(1139), B1 => n82, B2 => 
                           regs(1651), ZN => n1647);
   U2399 : OAI211_X1 port map( C1 => n21, C2 => n1649, A => n1648, B => n1647, 
                           ZN => curr_proc_regs(627));
   U2400 : AOI22_X1 port map( A1 => n116, A2 => regs(116), B1 => n9, B2 => 
                           regs(2164), ZN => n1651);
   U2401 : AOI22_X1 port map( A1 => n8, A2 => regs(1140), B1 => n88, B2 => 
                           regs(1652), ZN => n1650);
   U2402 : OAI211_X1 port map( C1 => n21, C2 => n1652, A => n1651, B => n1650, 
                           ZN => curr_proc_regs(628));
   U2403 : AOI22_X1 port map( A1 => n111, A2 => regs(117), B1 => n77, B2 => 
                           regs(2165), ZN => n1654);
   U2404 : AOI22_X1 port map( A1 => n8, A2 => regs(1141), B1 => n86, B2 => 
                           regs(1653), ZN => n1653);
   U2405 : OAI211_X1 port map( C1 => n21, C2 => n1655, A => n1654, B => n1653, 
                           ZN => curr_proc_regs(629));
   U2406 : INV_X1 port map( A => regs(1086), ZN => n1658);
   U2407 : AOI22_X1 port map( A1 => n112, A2 => regs(2110), B1 => n9, B2 => 
                           regs(1598), ZN => n1657);
   U2408 : AOI22_X1 port map( A1 => n53, A2 => regs(574), B1 => n28, B2 => 
                           regs(62), ZN => n1656);
   U2409 : OAI211_X1 port map( C1 => n15, C2 => n1658, A => n1657, B => n1656, 
                           ZN => curr_proc_regs(62));
   U2410 : AOI22_X1 port map( A1 => n112, A2 => regs(118), B1 => n9, B2 => 
                           regs(2166), ZN => n1660);
   U2411 : AOI22_X1 port map( A1 => n53, A2 => regs(1142), B1 => n81, B2 => 
                           regs(1654), ZN => n1659);
   U2412 : OAI211_X1 port map( C1 => n21, C2 => n1661, A => n1660, B => n1659, 
                           ZN => curr_proc_regs(630));
   U2413 : AOI22_X1 port map( A1 => n111, A2 => regs(119), B1 => n77, B2 => 
                           regs(2167), ZN => n1663);
   U2414 : AOI22_X1 port map( A1 => n87, A2 => regs(1655), B1 => n28, B2 => 
                           regs(631), ZN => n1662);
   U2415 : OAI211_X1 port map( C1 => n46, C2 => n1664, A => n1663, B => n1662, 
                           ZN => curr_proc_regs(631));
   U2416 : AOI22_X1 port map( A1 => n116, A2 => regs(120), B1 => n9, B2 => 
                           regs(2168), ZN => n1666);
   U2417 : AOI22_X1 port map( A1 => n87, A2 => regs(1656), B1 => n28, B2 => 
                           regs(632), ZN => n1665);
   U2418 : OAI211_X1 port map( C1 => n65, C2 => n1667, A => n1666, B => n1665, 
                           ZN => curr_proc_regs(632));
   U2419 : AOI22_X1 port map( A1 => n111, A2 => regs(121), B1 => n9, B2 => 
                           regs(2169), ZN => n1669);
   U2420 : AOI22_X1 port map( A1 => n53, A2 => regs(1145), B1 => n86, B2 => 
                           regs(1657), ZN => n1668);
   U2421 : OAI211_X1 port map( C1 => n21, C2 => n1670, A => n1669, B => n1668, 
                           ZN => curr_proc_regs(633));
   U2422 : AOI22_X1 port map( A1 => n112, A2 => regs(122), B1 => n77, B2 => 
                           regs(2170), ZN => n1672);
   U2423 : AOI22_X1 port map( A1 => n87, A2 => regs(1658), B1 => n28, B2 => 
                           regs(634), ZN => n1671);
   U2424 : OAI211_X1 port map( C1 => n66, C2 => n1673, A => n1672, B => n1671, 
                           ZN => curr_proc_regs(634));
   U2425 : AOI22_X1 port map( A1 => n116, A2 => regs(123), B1 => n9, B2 => 
                           regs(2171), ZN => n1675);
   U2426 : AOI22_X1 port map( A1 => n8, A2 => regs(1147), B1 => n87, B2 => 
                           regs(1659), ZN => n1674);
   U2427 : OAI211_X1 port map( C1 => n21, C2 => n1676, A => n1675, B => n1674, 
                           ZN => curr_proc_regs(635));
   U2428 : AOI22_X1 port map( A1 => n112, A2 => regs(124), B1 => n9, B2 => 
                           regs(2172), ZN => n1678);
   U2429 : AOI22_X1 port map( A1 => n87, A2 => regs(1660), B1 => n28, B2 => 
                           regs(636), ZN => n1677);
   U2430 : OAI211_X1 port map( C1 => n6, C2 => n1679, A => n1678, B => n1677, 
                           ZN => curr_proc_regs(636));
   U2431 : AOI22_X1 port map( A1 => n116, A2 => regs(125), B1 => n9, B2 => 
                           regs(2173), ZN => n1681);
   U2432 : AOI22_X1 port map( A1 => n87, A2 => regs(1661), B1 => n7, B2 => 
                           regs(637), ZN => n1680);
   U2433 : OAI211_X1 port map( C1 => n64, C2 => n1682, A => n1681, B => n1680, 
                           ZN => curr_proc_regs(637));
   U2434 : AOI22_X1 port map( A1 => n111, A2 => regs(126), B1 => n9, B2 => 
                           regs(2174), ZN => n1684);
   U2435 : AOI22_X1 port map( A1 => n87, A2 => regs(1662), B1 => n7, B2 => 
                           regs(638), ZN => n1683);
   U2436 : OAI211_X1 port map( C1 => n64, C2 => n1685, A => n1684, B => n1683, 
                           ZN => curr_proc_regs(638));
   U2437 : AOI22_X1 port map( A1 => n116, A2 => regs(127), B1 => n9, B2 => 
                           regs(2175), ZN => n1687);
   U2438 : AOI22_X1 port map( A1 => n87, A2 => regs(1663), B1 => n7, B2 => 
                           regs(639), ZN => n1686);
   U2439 : OAI211_X1 port map( C1 => n66, C2 => n1688, A => n1687, B => n1686, 
                           ZN => curr_proc_regs(639));
   U2440 : INV_X1 port map( A => regs(1087), ZN => n1691);
   U2441 : AOI22_X1 port map( A1 => n111, A2 => regs(2111), B1 => n9, B2 => 
                           regs(1599), ZN => n1690);
   U2442 : AOI22_X1 port map( A1 => n8, A2 => regs(575), B1 => n7, B2 => 
                           regs(63), ZN => n1689);
   U2443 : OAI211_X1 port map( C1 => n15, C2 => n1691, A => n1690, B => n1689, 
                           ZN => curr_proc_regs(63));
   U2444 : AOI22_X1 port map( A1 => n112, A2 => regs(128), B1 => n9, B2 => 
                           regs(2176), ZN => n1693);
   U2445 : AOI22_X1 port map( A1 => n87, A2 => regs(1664), B1 => n7, B2 => 
                           regs(640), ZN => n1692);
   U2446 : OAI211_X1 port map( C1 => n6, C2 => n1694, A => n1693, B => n1692, 
                           ZN => curr_proc_regs(640));
   U2447 : AOI22_X1 port map( A1 => n112, A2 => regs(129), B1 => n9, B2 => 
                           regs(2177), ZN => n1696);
   U2448 : AOI22_X1 port map( A1 => n8, A2 => regs(1153), B1 => n88, B2 => 
                           regs(1665), ZN => n1695);
   U2449 : OAI211_X1 port map( C1 => n21, C2 => n1697, A => n1696, B => n1695, 
                           ZN => curr_proc_regs(641));
   U2450 : AOI22_X1 port map( A1 => n116, A2 => regs(130), B1 => n9, B2 => 
                           regs(2178), ZN => n1699);
   U2451 : AOI22_X1 port map( A1 => n86, A2 => regs(1666), B1 => n7, B2 => 
                           regs(642), ZN => n1698);
   U2452 : OAI211_X1 port map( C1 => n64, C2 => n1700, A => n1699, B => n1698, 
                           ZN => curr_proc_regs(642));
   U2453 : AOI22_X1 port map( A1 => n111, A2 => regs(131), B1 => n9, B2 => 
                           regs(2179), ZN => n1702);
   U2454 : AOI22_X1 port map( A1 => n86, A2 => regs(1667), B1 => n7, B2 => 
                           regs(643), ZN => n1701);
   U2455 : OAI211_X1 port map( C1 => n64, C2 => n1703, A => n1702, B => n1701, 
                           ZN => curr_proc_regs(643));
   U2456 : AOI22_X1 port map( A1 => n112, A2 => regs(132), B1 => n9, B2 => 
                           regs(2180), ZN => n1705);
   U2457 : AOI22_X1 port map( A1 => n86, A2 => regs(1668), B1 => n7, B2 => 
                           regs(644), ZN => n1704);
   U2458 : OAI211_X1 port map( C1 => n67, C2 => n1706, A => n1705, B => n1704, 
                           ZN => curr_proc_regs(644));
   U2459 : AOI22_X1 port map( A1 => n116, A2 => regs(133), B1 => n77, B2 => 
                           regs(2181), ZN => n1708);
   U2460 : AOI22_X1 port map( A1 => n86, A2 => regs(1669), B1 => n7, B2 => 
                           regs(645), ZN => n1707);
   U2461 : OAI211_X1 port map( C1 => n1, C2 => n1709, A => n1708, B => n1707, 
                           ZN => curr_proc_regs(645));
   U2462 : AOI22_X1 port map( A1 => n116, A2 => regs(134), B1 => n9, B2 => 
                           regs(2182), ZN => n1711);
   U2463 : AOI22_X1 port map( A1 => n86, A2 => regs(1670), B1 => n7, B2 => 
                           regs(646), ZN => n1710);
   U2464 : OAI211_X1 port map( C1 => n66, C2 => n1712, A => n1711, B => n1710, 
                           ZN => curr_proc_regs(646));
   U2465 : AOI22_X1 port map( A1 => n111, A2 => regs(135), B1 => n9, B2 => 
                           regs(2183), ZN => n1714);
   U2466 : AOI22_X1 port map( A1 => n8, A2 => regs(1159), B1 => n79, B2 => 
                           regs(1671), ZN => n1713);
   U2467 : OAI211_X1 port map( C1 => n21, C2 => n1715, A => n1714, B => n1713, 
                           ZN => curr_proc_regs(647));
   U2468 : AOI22_X1 port map( A1 => n111, A2 => regs(136), B1 => n9, B2 => 
                           regs(2184), ZN => n1717);
   U2469 : AOI22_X1 port map( A1 => n8, A2 => regs(1160), B1 => n84, B2 => 
                           regs(1672), ZN => n1716);
   U2470 : OAI211_X1 port map( C1 => n21, C2 => n1718, A => n1717, B => n1716, 
                           ZN => curr_proc_regs(648));
   U2471 : AOI22_X1 port map( A1 => n112, A2 => regs(137), B1 => n77, B2 => 
                           regs(2185), ZN => n1720);
   U2472 : AOI22_X1 port map( A1 => n86, A2 => regs(1673), B1 => n7, B2 => 
                           regs(649), ZN => n1719);
   U2473 : OAI211_X1 port map( C1 => n65, C2 => n1721, A => n1720, B => n1719, 
                           ZN => curr_proc_regs(649));
   U2474 : AOI22_X1 port map( A1 => n116, A2 => regs(2112), B1 => n9, B2 => 
                           regs(1600), ZN => n1723);
   U2475 : AOI22_X1 port map( A1 => n8, A2 => regs(576), B1 => n7, B2 => 
                           regs(64), ZN => n1722);
   U2476 : OAI211_X1 port map( C1 => n15, C2 => n1724, A => n1723, B => n1722, 
                           ZN => curr_proc_regs(64));
   U2477 : AOI22_X1 port map( A1 => n111, A2 => regs(138), B1 => n9, B2 => 
                           regs(2186), ZN => n1726);
   U2478 : AOI22_X1 port map( A1 => n8, A2 => regs(1162), B1 => n82, B2 => 
                           regs(1674), ZN => n1725);
   U2479 : OAI211_X1 port map( C1 => n22, C2 => n1727, A => n1726, B => n1725, 
                           ZN => curr_proc_regs(650));
   U2480 : AOI22_X1 port map( A1 => n112, A2 => regs(139), B1 => n9, B2 => 
                           regs(2187), ZN => n1729);
   U2481 : AOI22_X1 port map( A1 => n86, A2 => regs(1675), B1 => n7, B2 => 
                           regs(651), ZN => n1728);
   U2482 : OAI211_X1 port map( C1 => n65, C2 => n1730, A => n1729, B => n1728, 
                           ZN => curr_proc_regs(651));
   U2483 : AOI22_X1 port map( A1 => n116, A2 => regs(140), B1 => n77, B2 => 
                           regs(2188), ZN => n1732);
   U2484 : AOI22_X1 port map( A1 => n8, A2 => regs(1164), B1 => n83, B2 => 
                           regs(1676), ZN => n1731);
   U2485 : OAI211_X1 port map( C1 => n22, C2 => n1733, A => n1732, B => n1731, 
                           ZN => curr_proc_regs(652));
   U2486 : AOI22_X1 port map( A1 => n111, A2 => regs(141), B1 => n77, B2 => 
                           regs(2189), ZN => n1735);
   U2487 : AOI22_X1 port map( A1 => n86, A2 => regs(1677), B1 => n7, B2 => 
                           regs(653), ZN => n1734);
   U2488 : OAI211_X1 port map( C1 => n65, C2 => n1736, A => n1735, B => n1734, 
                           ZN => curr_proc_regs(653));
   U2489 : AOI22_X1 port map( A1 => n112, A2 => regs(142), B1 => n9, B2 => 
                           regs(2190), ZN => n1738);
   U2490 : AOI22_X1 port map( A1 => n55, A2 => regs(1166), B1 => n87, B2 => 
                           regs(1678), ZN => n1737);
   U2491 : OAI211_X1 port map( C1 => n22, C2 => n1739, A => n1738, B => n1737, 
                           ZN => curr_proc_regs(654));
   U2492 : AOI22_X1 port map( A1 => n116, A2 => regs(143), B1 => n9, B2 => 
                           regs(2191), ZN => n1741);
   U2493 : AOI22_X1 port map( A1 => n86, A2 => regs(1679), B1 => n7, B2 => 
                           regs(655), ZN => n1740);
   U2494 : OAI211_X1 port map( C1 => n65, C2 => n1742, A => n1741, B => n1740, 
                           ZN => curr_proc_regs(655));
   U2495 : AOI22_X1 port map( A1 => n111, A2 => regs(144), B1 => n9, B2 => 
                           regs(2192), ZN => n1744);
   U2496 : AOI22_X1 port map( A1 => n86, A2 => regs(1680), B1 => n7, B2 => 
                           regs(656), ZN => n1743);
   U2497 : OAI211_X1 port map( C1 => n65, C2 => n1745, A => n1744, B => n1743, 
                           ZN => curr_proc_regs(656));
   U2498 : AOI22_X1 port map( A1 => n112, A2 => regs(145), B1 => n9, B2 => 
                           regs(2193), ZN => n1747);
   U2499 : AOI22_X1 port map( A1 => n55, A2 => regs(1169), B1 => n98, B2 => 
                           regs(1681), ZN => n1746);
   U2500 : OAI211_X1 port map( C1 => n22, C2 => n1748, A => n1747, B => n1746, 
                           ZN => curr_proc_regs(657));
   U2501 : AOI22_X1 port map( A1 => n112, A2 => regs(146), B1 => n9, B2 => 
                           regs(2194), ZN => n1750);
   U2502 : AOI22_X1 port map( A1 => n86, A2 => regs(1682), B1 => n7, B2 => 
                           regs(658), ZN => n1749);
   U2503 : OAI211_X1 port map( C1 => n65, C2 => n1751, A => n1750, B => n1749, 
                           ZN => curr_proc_regs(658));
   U2504 : AOI22_X1 port map( A1 => n112, A2 => regs(147), B1 => n77, B2 => 
                           regs(2195), ZN => n1753);
   U2505 : AOI22_X1 port map( A1 => n85, A2 => regs(1683), B1 => n7, B2 => 
                           regs(659), ZN => n1752);
   U2506 : OAI211_X1 port map( C1 => n65, C2 => n1754, A => n1753, B => n1752, 
                           ZN => curr_proc_regs(659));
   U2507 : INV_X1 port map( A => regs(577), ZN => n1757);
   U2508 : AOI22_X1 port map( A1 => n112, A2 => regs(2113), B1 => n77, B2 => 
                           regs(1601), ZN => n1756);
   U2509 : AOI22_X1 port map( A1 => n85, A2 => regs(1089), B1 => n7, B2 => 
                           regs(65), ZN => n1755);
   U2510 : OAI211_X1 port map( C1 => n66, C2 => n1757, A => n1756, B => n1755, 
                           ZN => curr_proc_regs(65));
   U2511 : AOI22_X1 port map( A1 => n112, A2 => regs(148), B1 => n9, B2 => 
                           regs(2196), ZN => n1759);
   U2512 : AOI22_X1 port map( A1 => n55, A2 => regs(1172), B1 => n85, B2 => 
                           regs(1684), ZN => n1758);
   U2513 : OAI211_X1 port map( C1 => n22, C2 => n1760, A => n1759, B => n1758, 
                           ZN => curr_proc_regs(660));
   U2514 : AOI22_X1 port map( A1 => n112, A2 => regs(149), B1 => n9, B2 => 
                           regs(2197), ZN => n1762);
   U2515 : AOI22_X1 port map( A1 => n85, A2 => regs(1685), B1 => n7, B2 => 
                           regs(661), ZN => n1761);
   U2516 : OAI211_X1 port map( C1 => n65, C2 => n1763, A => n1762, B => n1761, 
                           ZN => curr_proc_regs(661));
   U2517 : AOI22_X1 port map( A1 => n112, A2 => regs(150), B1 => n77, B2 => 
                           regs(2198), ZN => n1765);
   U2518 : AOI22_X1 port map( A1 => n85, A2 => regs(1686), B1 => n7, B2 => 
                           regs(662), ZN => n1764);
   U2519 : OAI211_X1 port map( C1 => n46, C2 => n1766, A => n1765, B => n1764, 
                           ZN => curr_proc_regs(662));
   U2520 : AOI22_X1 port map( A1 => n112, A2 => regs(151), B1 => n77, B2 => 
                           regs(2199), ZN => n1768);
   U2521 : AOI22_X1 port map( A1 => n85, A2 => regs(1687), B1 => n7, B2 => 
                           regs(663), ZN => n1767);
   U2522 : OAI211_X1 port map( C1 => n1, C2 => n1769, A => n1768, B => n1767, 
                           ZN => curr_proc_regs(663));
   U2523 : AOI22_X1 port map( A1 => n112, A2 => regs(152), B1 => n77, B2 => 
                           regs(2200), ZN => n1771);
   U2524 : AOI22_X1 port map( A1 => n55, A2 => regs(1176), B1 => n85, B2 => 
                           regs(1688), ZN => n1770);
   U2525 : OAI211_X1 port map( C1 => n22, C2 => n1772, A => n1771, B => n1770, 
                           ZN => curr_proc_regs(664));
   U2526 : AOI22_X1 port map( A1 => n112, A2 => regs(153), B1 => n9, B2 => 
                           regs(2201), ZN => n1774);
   U2527 : AOI22_X1 port map( A1 => n55, A2 => regs(1177), B1 => n79, B2 => 
                           regs(1689), ZN => n1773);
   U2528 : OAI211_X1 port map( C1 => n2112, C2 => n1775, A => n1774, B => n1773
                           , ZN => curr_proc_regs(665));
   U2529 : AOI22_X1 port map( A1 => n112, A2 => regs(154), B1 => n77, B2 => 
                           regs(2202), ZN => n1777);
   U2530 : AOI22_X1 port map( A1 => n55, A2 => regs(1178), B1 => n80, B2 => 
                           regs(1690), ZN => n1776);
   U2531 : OAI211_X1 port map( C1 => n22, C2 => n1778, A => n1777, B => n1776, 
                           ZN => curr_proc_regs(666));
   U2532 : AOI22_X1 port map( A1 => n112, A2 => regs(155), B1 => n77, B2 => 
                           regs(2203), ZN => n1780);
   U2533 : AOI22_X1 port map( A1 => n55, A2 => regs(1179), B1 => n81, B2 => 
                           regs(1691), ZN => n1779);
   U2534 : OAI211_X1 port map( C1 => n21, C2 => n1781, A => n1780, B => n1779, 
                           ZN => curr_proc_regs(667));
   U2535 : AOI22_X1 port map( A1 => n111, A2 => regs(156), B1 => n77, B2 => 
                           regs(2204), ZN => n1783);
   U2536 : AOI22_X1 port map( A1 => n55, A2 => regs(1180), B1 => n86, B2 => 
                           regs(1692), ZN => n1782);
   U2537 : OAI211_X1 port map( C1 => n2112, C2 => n1784, A => n1783, B => n1782
                           , ZN => curr_proc_regs(668));
   U2538 : AOI22_X1 port map( A1 => n111, A2 => regs(157), B1 => n77, B2 => 
                           regs(2205), ZN => n1786);
   U2539 : AOI22_X1 port map( A1 => n55, A2 => regs(1181), B1 => n87, B2 => 
                           regs(1693), ZN => n1785);
   U2540 : OAI211_X1 port map( C1 => n22, C2 => n1787, A => n1786, B => n1785, 
                           ZN => curr_proc_regs(669));
   U2541 : AOI22_X1 port map( A1 => n111, A2 => regs(2114), B1 => n9, B2 => 
                           regs(1602), ZN => n1789);
   U2542 : AOI22_X1 port map( A1 => n55, A2 => regs(578), B1 => n23, B2 => 
                           regs(66), ZN => n1788);
   U2543 : OAI211_X1 port map( C1 => n15, C2 => n1790, A => n1789, B => n1788, 
                           ZN => curr_proc_regs(66));
   U2544 : AOI22_X1 port map( A1 => n111, A2 => regs(158), B1 => n9, B2 => 
                           regs(2206), ZN => n1792);
   U2545 : AOI22_X1 port map( A1 => n85, A2 => regs(1694), B1 => n23, B2 => 
                           regs(670), ZN => n1791);
   U2546 : OAI211_X1 port map( C1 => n67, C2 => n1793, A => n1792, B => n1791, 
                           ZN => curr_proc_regs(670));
   U2547 : AOI22_X1 port map( A1 => n111, A2 => regs(159), B1 => n77, B2 => 
                           regs(2207), ZN => n1795);
   U2548 : AOI22_X1 port map( A1 => n85, A2 => regs(1695), B1 => n24, B2 => 
                           regs(671), ZN => n1794);
   U2549 : OAI211_X1 port map( C1 => n64, C2 => n1796, A => n1795, B => n1794, 
                           ZN => curr_proc_regs(671));
   U2550 : AOI22_X1 port map( A1 => n111, A2 => regs(160), B1 => n77, B2 => 
                           regs(2208), ZN => n1798);
   U2551 : AOI22_X1 port map( A1 => n85, A2 => regs(1696), B1 => n45, B2 => 
                           regs(672), ZN => n1797);
   U2552 : OAI211_X1 port map( C1 => n6, C2 => n1799, A => n1798, B => n1797, 
                           ZN => curr_proc_regs(672));
   U2553 : AOI22_X1 port map( A1 => n111, A2 => regs(161), B1 => n77, B2 => 
                           regs(2209), ZN => n1801);
   U2554 : AOI22_X1 port map( A1 => n51, A2 => regs(1185), B1 => n88, B2 => 
                           regs(1697), ZN => n1800);
   U2555 : OAI211_X1 port map( C1 => n21, C2 => n1802, A => n1801, B => n1800, 
                           ZN => curr_proc_regs(673));
   U2556 : AOI22_X1 port map( A1 => n111, A2 => regs(162), B1 => n77, B2 => 
                           regs(2210), ZN => n1804);
   U2557 : AOI22_X1 port map( A1 => n85, A2 => regs(1698), B1 => n42, B2 => 
                           regs(674), ZN => n1803);
   U2558 : OAI211_X1 port map( C1 => n6, C2 => n1805, A => n1804, B => n1803, 
                           ZN => curr_proc_regs(674));
   U2559 : AOI22_X1 port map( A1 => n111, A2 => regs(163), B1 => n3, B2 => 
                           regs(2211), ZN => n1807);
   U2560 : AOI22_X1 port map( A1 => n85, A2 => regs(1699), B1 => n42, B2 => 
                           regs(675), ZN => n1806);
   U2561 : OAI211_X1 port map( C1 => n6, C2 => n1808, A => n1807, B => n1806, 
                           ZN => curr_proc_regs(675));
   U2562 : AOI22_X1 port map( A1 => n111, A2 => regs(164), B1 => n3, B2 => 
                           regs(2212), ZN => n1810);
   U2563 : AOI22_X1 port map( A1 => n48, A2 => regs(1188), B1 => n86, B2 => 
                           regs(1700), ZN => n1809);
   U2564 : OAI211_X1 port map( C1 => n2112, C2 => n1811, A => n1810, B => n1809
                           , ZN => curr_proc_regs(676));
   U2565 : AOI22_X1 port map( A1 => n111, A2 => regs(165), B1 => n71, B2 => 
                           regs(2213), ZN => n1813);
   U2566 : AOI22_X1 port map( A1 => n85, A2 => regs(1701), B1 => n39, B2 => 
                           regs(677), ZN => n1812);
   U2567 : OAI211_X1 port map( C1 => n6, C2 => n1814, A => n1813, B => n1812, 
                           ZN => curr_proc_regs(677));
   U2568 : AOI22_X1 port map( A1 => n116, A2 => regs(166), B1 => n68, B2 => 
                           regs(2214), ZN => n1816);
   U2569 : AOI22_X1 port map( A1 => n48, A2 => regs(1190), B1 => n80, B2 => 
                           regs(1702), ZN => n1815);
   U2570 : OAI211_X1 port map( C1 => n22, C2 => n1817, A => n1816, B => n1815, 
                           ZN => curr_proc_regs(678));
   U2571 : AOI22_X1 port map( A1 => n116, A2 => regs(167), B1 => n73, B2 => 
                           regs(2215), ZN => n1819);
   U2572 : AOI22_X1 port map( A1 => n51, A2 => regs(1191), B1 => n98, B2 => 
                           regs(1703), ZN => n1818);
   U2573 : OAI211_X1 port map( C1 => n22, C2 => n1820, A => n1819, B => n1818, 
                           ZN => curr_proc_regs(679));
   U2574 : INV_X1 port map( A => regs(579), ZN => n1823);
   U2575 : AOI22_X1 port map( A1 => n116, A2 => regs(2115), B1 => n16, B2 => 
                           regs(1603), ZN => n1822);
   U2576 : AOI22_X1 port map( A1 => n84, A2 => regs(1091), B1 => n24, B2 => 
                           regs(67), ZN => n1821);
   U2577 : OAI211_X1 port map( C1 => n6, C2 => n1823, A => n1822, B => n1821, 
                           ZN => curr_proc_regs(67));
   U2578 : AOI22_X1 port map( A1 => n116, A2 => regs(168), B1 => n76, B2 => 
                           regs(2216), ZN => n1825);
   U2579 : AOI22_X1 port map( A1 => n50, A2 => regs(1192), B1 => n84, B2 => 
                           regs(1704), ZN => n1824);
   U2580 : OAI211_X1 port map( C1 => n22, C2 => n1826, A => n1825, B => n1824, 
                           ZN => curr_proc_regs(680));
   U2581 : AOI22_X1 port map( A1 => n116, A2 => regs(169), B1 => n76, B2 => 
                           regs(2217), ZN => n1828);
   U2582 : AOI22_X1 port map( A1 => n84, A2 => regs(1705), B1 => n23, B2 => 
                           regs(681), ZN => n1827);
   U2583 : OAI211_X1 port map( C1 => n6, C2 => n1829, A => n1828, B => n1827, 
                           ZN => curr_proc_regs(681));
   U2584 : AOI22_X1 port map( A1 => n116, A2 => regs(170), B1 => n76, B2 => 
                           regs(2218), ZN => n1831);
   U2585 : AOI22_X1 port map( A1 => n84, A2 => regs(1706), B1 => n39, B2 => 
                           regs(682), ZN => n1830);
   U2586 : OAI211_X1 port map( C1 => n6, C2 => n1832, A => n1831, B => n1830, 
                           ZN => curr_proc_regs(682));
   U2587 : AOI22_X1 port map( A1 => n116, A2 => regs(171), B1 => n76, B2 => 
                           regs(2219), ZN => n1834);
   U2588 : AOI22_X1 port map( A1 => n84, A2 => regs(1707), B1 => n23, B2 => 
                           regs(683), ZN => n1833);
   U2589 : OAI211_X1 port map( C1 => n6, C2 => n1835, A => n1834, B => n1833, 
                           ZN => curr_proc_regs(683));
   U2590 : AOI22_X1 port map( A1 => n116, A2 => regs(172), B1 => n76, B2 => 
                           regs(2220), ZN => n1837);
   U2591 : AOI22_X1 port map( A1 => n84, A2 => regs(1708), B1 => n2, B2 => 
                           regs(684), ZN => n1836);
   U2592 : OAI211_X1 port map( C1 => n64, C2 => n1838, A => n1837, B => n1836, 
                           ZN => curr_proc_regs(684));
   U2593 : AOI22_X1 port map( A1 => n116, A2 => regs(173), B1 => n76, B2 => 
                           regs(2221), ZN => n1840);
   U2594 : AOI22_X1 port map( A1 => n84, A2 => regs(1709), B1 => n2, B2 => 
                           regs(685), ZN => n1839);
   U2595 : OAI211_X1 port map( C1 => n47, C2 => n1841, A => n1840, B => n1839, 
                           ZN => curr_proc_regs(685));
   U2596 : AOI22_X1 port map( A1 => n116, A2 => regs(174), B1 => n76, B2 => 
                           regs(2222), ZN => n1843);
   U2597 : AOI22_X1 port map( A1 => n49, A2 => regs(1198), B1 => n97, B2 => 
                           regs(1710), ZN => n1842);
   U2598 : OAI211_X1 port map( C1 => n22, C2 => n1844, A => n1843, B => n1842, 
                           ZN => curr_proc_regs(686));
   U2599 : AOI22_X1 port map( A1 => n116, A2 => regs(175), B1 => n3, B2 => 
                           regs(2223), ZN => n1846);
   U2600 : AOI22_X1 port map( A1 => n56, A2 => regs(1199), B1 => n14, B2 => 
                           regs(1711), ZN => n1845);
   U2601 : OAI211_X1 port map( C1 => n22, C2 => n1847, A => n1846, B => n1845, 
                           ZN => curr_proc_regs(687));
   U2602 : AOI22_X1 port map( A1 => n4, A2 => regs(176), B1 => n76, B2 => 
                           regs(2224), ZN => n1849);
   U2603 : AOI22_X1 port map( A1 => n84, A2 => regs(1712), B1 => n2, B2 => 
                           regs(688), ZN => n1848);
   U2604 : OAI211_X1 port map( C1 => n46, C2 => n1850, A => n1849, B => n1848, 
                           ZN => curr_proc_regs(688));
   U2605 : AOI22_X1 port map( A1 => n116, A2 => regs(177), B1 => n76, B2 => 
                           regs(2225), ZN => n1852);
   U2606 : AOI22_X1 port map( A1 => n61, A2 => regs(1201), B1 => n14, B2 => 
                           regs(1713), ZN => n1851);
   U2607 : OAI211_X1 port map( C1 => n22, C2 => n1853, A => n1852, B => n1851, 
                           ZN => curr_proc_regs(689));
   U2608 : INV_X1 port map( A => regs(580), ZN => n1856);
   U2609 : AOI22_X1 port map( A1 => n116, A2 => regs(2116), B1 => n3, B2 => 
                           regs(1604), ZN => n1855);
   U2610 : AOI22_X1 port map( A1 => n84, A2 => regs(1092), B1 => n2, B2 => 
                           regs(68), ZN => n1854);
   U2611 : OAI211_X1 port map( C1 => n46, C2 => n1856, A => n1855, B => n1854, 
                           ZN => curr_proc_regs(68));
   U2612 : AOI22_X1 port map( A1 => n116, A2 => regs(178), B1 => n76, B2 => 
                           regs(2226), ZN => n1858);
   U2613 : AOI22_X1 port map( A1 => n84, A2 => regs(1714), B1 => n2, B2 => 
                           regs(690), ZN => n1857);
   U2614 : OAI211_X1 port map( C1 => n67, C2 => n1859, A => n1858, B => n1857, 
                           ZN => curr_proc_regs(690));
   U2615 : AOI22_X1 port map( A1 => n116, A2 => regs(179), B1 => n76, B2 => 
                           regs(2227), ZN => n1861);
   U2616 : AOI22_X1 port map( A1 => n59, A2 => regs(1203), B1 => n14, B2 => 
                           regs(1715), ZN => n1860);
   U2617 : OAI211_X1 port map( C1 => n22, C2 => n1862, A => n1861, B => n1860, 
                           ZN => curr_proc_regs(691));
   U2618 : AOI22_X1 port map( A1 => n4, A2 => regs(180), B1 => n77, B2 => 
                           regs(2228), ZN => n1864);
   U2619 : AOI22_X1 port map( A1 => n55, A2 => regs(1204), B1 => n14, B2 => 
                           regs(1716), ZN => n1863);
   U2620 : OAI211_X1 port map( C1 => n22, C2 => n1865, A => n1864, B => n1863, 
                           ZN => curr_proc_regs(692));
   U2621 : AOI22_X1 port map( A1 => n116, A2 => regs(181), B1 => n76, B2 => 
                           regs(2229), ZN => n1867);
   U2622 : AOI22_X1 port map( A1 => n54, A2 => regs(1205), B1 => n97, B2 => 
                           regs(1717), ZN => n1866);
   U2623 : OAI211_X1 port map( C1 => n22, C2 => n1868, A => n1867, B => n1866, 
                           ZN => curr_proc_regs(693));
   U2624 : AOI22_X1 port map( A1 => n116, A2 => regs(182), B1 => n76, B2 => 
                           regs(2230), ZN => n1870);
   U2625 : AOI22_X1 port map( A1 => n55, A2 => regs(1206), B1 => n14, B2 => 
                           regs(1718), ZN => n1869);
   U2626 : OAI211_X1 port map( C1 => n22, C2 => n1871, A => n1870, B => n1869, 
                           ZN => curr_proc_regs(694));
   U2627 : AOI22_X1 port map( A1 => n4, A2 => regs(183), B1 => n76, B2 => 
                           regs(2231), ZN => n1873);
   U2628 : AOI22_X1 port map( A1 => n59, A2 => regs(1207), B1 => n97, B2 => 
                           regs(1719), ZN => n1872);
   U2629 : OAI211_X1 port map( C1 => n22, C2 => n1874, A => n1873, B => n1872, 
                           ZN => curr_proc_regs(695));
   U2630 : AOI22_X1 port map( A1 => n116, A2 => regs(184), B1 => n76, B2 => 
                           regs(2232), ZN => n1876);
   U2631 : AOI22_X1 port map( A1 => n56, A2 => regs(1208), B1 => n14, B2 => 
                           regs(1720), ZN => n1875);
   U2632 : OAI211_X1 port map( C1 => n22, C2 => n1877, A => n1876, B => n1875, 
                           ZN => curr_proc_regs(696));
   U2633 : AOI22_X1 port map( A1 => n4, A2 => regs(185), B1 => n76, B2 => 
                           regs(2233), ZN => n1879);
   U2634 : AOI22_X1 port map( A1 => n49, A2 => regs(1209), B1 => n14, B2 => 
                           regs(1721), ZN => n1878);
   U2635 : OAI211_X1 port map( C1 => n22, C2 => n1880, A => n1879, B => n1878, 
                           ZN => curr_proc_regs(697));
   U2636 : AOI22_X1 port map( A1 => n4, A2 => regs(186), B1 => n76, B2 => 
                           regs(2234), ZN => n1882);
   U2637 : AOI22_X1 port map( A1 => n84, A2 => regs(1722), B1 => n2, B2 => 
                           regs(698), ZN => n1881);
   U2638 : OAI211_X1 port map( C1 => n64, C2 => n1883, A => n1882, B => n1881, 
                           ZN => curr_proc_regs(698));
   U2639 : AOI22_X1 port map( A1 => n4, A2 => regs(187), B1 => n76, B2 => 
                           regs(2235), ZN => n1885);
   U2640 : AOI22_X1 port map( A1 => n89, A2 => regs(1723), B1 => n2, B2 => 
                           regs(699), ZN => n1884);
   U2641 : OAI211_X1 port map( C1 => n46, C2 => n1886, A => n1885, B => n1884, 
                           ZN => curr_proc_regs(699));
   U2642 : INV_X1 port map( A => regs(581), ZN => n1889);
   U2643 : AOI22_X1 port map( A1 => n4, A2 => regs(2117), B1 => n76, B2 => 
                           regs(1605), ZN => n1888);
   U2644 : AOI22_X1 port map( A1 => n90, A2 => regs(1093), B1 => n2, B2 => 
                           regs(69), ZN => n1887);
   U2645 : OAI211_X1 port map( C1 => n6, C2 => n1889, A => n1888, B => n1887, 
                           ZN => curr_proc_regs(69));
   U2646 : AOI22_X1 port map( A1 => n4, A2 => regs(2054), B1 => n76, B2 => 
                           regs(1542), ZN => n1891);
   U2647 : AOI22_X1 port map( A1 => n50, A2 => regs(518), B1 => n2, B2 => 
                           regs(6), ZN => n1890);
   U2648 : OAI211_X1 port map( C1 => n15, C2 => n1892, A => n1891, B => n1890, 
                           ZN => curr_proc_regs(6));
   U2649 : AOI22_X1 port map( A1 => n4, A2 => regs(188), B1 => n76, B2 => 
                           regs(2236), ZN => n1894);
   U2650 : AOI22_X1 port map( A1 => n51, A2 => regs(1212), B1 => n97, B2 => 
                           regs(1724), ZN => n1893);
   U2651 : OAI211_X1 port map( C1 => n22, C2 => n1895, A => n1894, B => n1893, 
                           ZN => curr_proc_regs(700));
   U2652 : AOI22_X1 port map( A1 => n4, A2 => regs(189), B1 => n76, B2 => 
                           regs(2237), ZN => n1897);
   U2653 : AOI22_X1 port map( A1 => n48, A2 => regs(1213), B1 => n97, B2 => 
                           regs(1725), ZN => n1896);
   U2654 : OAI211_X1 port map( C1 => n22, C2 => n1898, A => n1897, B => n1896, 
                           ZN => curr_proc_regs(701));
   U2655 : AOI22_X1 port map( A1 => n4, A2 => regs(190), B1 => n76, B2 => 
                           regs(2238), ZN => n1900);
   U2656 : AOI22_X1 port map( A1 => n53, A2 => regs(1214), B1 => n97, B2 => 
                           regs(1726), ZN => n1899);
   U2657 : OAI211_X1 port map( C1 => n22, C2 => n1901, A => n1900, B => n1899, 
                           ZN => curr_proc_regs(702));
   U2658 : AOI22_X1 port map( A1 => n4, A2 => regs(191), B1 => n76, B2 => 
                           regs(2239), ZN => n1903);
   U2659 : AOI22_X1 port map( A1 => n52, A2 => regs(1215), B1 => n97, B2 => 
                           regs(1727), ZN => n1902);
   U2660 : OAI211_X1 port map( C1 => n22, C2 => n1904, A => n1903, B => n1902, 
                           ZN => curr_proc_regs(703));
   U2661 : AOI22_X1 port map( A1 => n4, A2 => regs(192), B1 => n76, B2 => 
                           regs(2240), ZN => n1906);
   U2662 : AOI22_X1 port map( A1 => n92, A2 => regs(1728), B1 => n2, B2 => 
                           regs(704), ZN => n1905);
   U2663 : OAI211_X1 port map( C1 => n6, C2 => n1907, A => n1906, B => n1905, 
                           ZN => curr_proc_regs(704));
   U2664 : AOI22_X1 port map( A1 => n4, A2 => regs(193), B1 => n68, B2 => 
                           regs(2241), ZN => n1909);
   U2665 : AOI22_X1 port map( A1 => n94, A2 => regs(1729), B1 => n2, B2 => 
                           regs(705), ZN => n1908);
   U2666 : OAI211_X1 port map( C1 => n6, C2 => n1910, A => n1909, B => n1908, 
                           ZN => curr_proc_regs(705));
   U2667 : AOI22_X1 port map( A1 => n116, A2 => regs(194), B1 => n73, B2 => 
                           regs(2242), ZN => n1912);
   U2668 : AOI22_X1 port map( A1 => n80, A2 => regs(1730), B1 => n2, B2 => 
                           regs(706), ZN => n1911);
   U2669 : OAI211_X1 port map( C1 => n6, C2 => n1913, A => n1912, B => n1911, 
                           ZN => curr_proc_regs(706));
   U2670 : AOI22_X1 port map( A1 => n4, A2 => regs(195), B1 => n76, B2 => 
                           regs(2243), ZN => n1915);
   U2671 : AOI22_X1 port map( A1 => n95, A2 => regs(1731), B1 => n2, B2 => 
                           regs(707), ZN => n1914);
   U2672 : OAI211_X1 port map( C1 => n6, C2 => n1916, A => n1915, B => n1914, 
                           ZN => curr_proc_regs(707));
   U2673 : AOI22_X1 port map( A1 => n116, A2 => regs(196), B1 => n76, B2 => 
                           regs(2244), ZN => n1918);
   U2674 : AOI22_X1 port map( A1 => n54, A2 => regs(1220), B1 => n97, B2 => 
                           regs(1732), ZN => n1917);
   U2675 : OAI211_X1 port map( C1 => n22, C2 => n1919, A => n1918, B => n1917, 
                           ZN => curr_proc_regs(708));
   U2676 : AOI22_X1 port map( A1 => n116, A2 => regs(197), B1 => n76, B2 => 
                           regs(2245), ZN => n1921);
   U2677 : AOI22_X1 port map( A1 => n90, A2 => regs(1733), B1 => n2, B2 => 
                           regs(709), ZN => n1920);
   U2678 : OAI211_X1 port map( C1 => n6, C2 => n1922, A => n1921, B => n1920, 
                           ZN => curr_proc_regs(709));
   U2679 : AOI22_X1 port map( A1 => n116, A2 => regs(2118), B1 => n16, B2 => 
                           regs(1606), ZN => n1924);
   U2680 : AOI22_X1 port map( A1 => n55, A2 => regs(582), B1 => n2, B2 => 
                           regs(70), ZN => n1923);
   U2681 : OAI211_X1 port map( C1 => n100, C2 => n1925, A => n1924, B => n1923,
                           ZN => curr_proc_regs(70));
   U2682 : AOI22_X1 port map( A1 => n4, A2 => regs(198), B1 => n76, B2 => 
                           regs(2246), ZN => n1927);
   U2683 : AOI22_X1 port map( A1 => n92, A2 => regs(1734), B1 => n2, B2 => 
                           regs(710), ZN => n1926);
   U2684 : OAI211_X1 port map( C1 => n6, C2 => n1928, A => n1927, B => n1926, 
                           ZN => curr_proc_regs(710));
   U2685 : AOI22_X1 port map( A1 => n116, A2 => regs(199), B1 => n76, B2 => 
                           regs(2247), ZN => n1930);
   U2686 : AOI22_X1 port map( A1 => n60, A2 => regs(1223), B1 => n14, B2 => 
                           regs(1735), ZN => n1929);
   U2687 : OAI211_X1 port map( C1 => n22, C2 => n1931, A => n1930, B => n1929, 
                           ZN => curr_proc_regs(711));
   U2688 : AOI22_X1 port map( A1 => n116, A2 => regs(200), B1 => n76, B2 => 
                           regs(2248), ZN => n1933);
   U2689 : AOI22_X1 port map( A1 => n94, A2 => regs(1736), B1 => n2, B2 => 
                           regs(712), ZN => n1932);
   U2690 : OAI211_X1 port map( C1 => n46, C2 => n1934, A => n1933, B => n1932, 
                           ZN => curr_proc_regs(712));
   U2691 : AOI22_X1 port map( A1 => n4, A2 => regs(201), B1 => n16, B2 => 
                           regs(2249), ZN => n1936);
   U2692 : AOI22_X1 port map( A1 => n97, A2 => regs(1737), B1 => n2, B2 => 
                           regs(713), ZN => n1935);
   U2693 : OAI211_X1 port map( C1 => n67, C2 => n1937, A => n1936, B => n1935, 
                           ZN => curr_proc_regs(713));
   U2694 : AOI22_X1 port map( A1 => n4, A2 => regs(202), B1 => n76, B2 => 
                           regs(2250), ZN => n1939);
   U2695 : AOI22_X1 port map( A1 => n63, A2 => regs(1226), B1 => n97, B2 => 
                           regs(1738), ZN => n1938);
   U2696 : OAI211_X1 port map( C1 => n22, C2 => n1940, A => n1939, B => n1938, 
                           ZN => curr_proc_regs(714));
   U2697 : AOI22_X1 port map( A1 => n116, A2 => regs(203), B1 => n3, B2 => 
                           regs(2251), ZN => n1942);
   U2698 : AOI22_X1 port map( A1 => n10, A2 => regs(1227), B1 => n97, B2 => 
                           regs(1739), ZN => n1941);
   U2699 : OAI211_X1 port map( C1 => n22, C2 => n1943, A => n1942, B => n1941, 
                           ZN => curr_proc_regs(715));
   U2700 : AOI22_X1 port map( A1 => n116, A2 => regs(204), B1 => n73, B2 => 
                           regs(2252), ZN => n1945);
   U2701 : AOI22_X1 port map( A1 => n98, A2 => regs(1740), B1 => n2, B2 => 
                           regs(716), ZN => n1944);
   U2702 : OAI211_X1 port map( C1 => n46, C2 => n1946, A => n1945, B => n1944, 
                           ZN => curr_proc_regs(716));
   U2703 : AOI22_X1 port map( A1 => n116, A2 => regs(205), B1 => n76, B2 => 
                           regs(2253), ZN => n1948);
   U2704 : AOI22_X1 port map( A1 => n98, A2 => regs(1741), B1 => n2, B2 => 
                           regs(717), ZN => n1947);
   U2705 : OAI211_X1 port map( C1 => n64, C2 => n1949, A => n1948, B => n1947, 
                           ZN => curr_proc_regs(717));
   U2706 : AOI22_X1 port map( A1 => n4, A2 => regs(206), B1 => n76, B2 => 
                           regs(2254), ZN => n1951);
   U2707 : AOI22_X1 port map( A1 => n10, A2 => regs(1230), B1 => n97, B2 => 
                           regs(1742), ZN => n1950);
   U2708 : OAI211_X1 port map( C1 => n22, C2 => n1952, A => n1951, B => n1950, 
                           ZN => curr_proc_regs(718));
   U2709 : AOI22_X1 port map( A1 => n116, A2 => regs(207), B1 => n76, B2 => 
                           regs(2255), ZN => n1954);
   U2710 : AOI22_X1 port map( A1 => n10, A2 => regs(1231), B1 => n14, B2 => 
                           regs(1743), ZN => n1953);
   U2711 : OAI211_X1 port map( C1 => n22, C2 => n1955, A => n1954, B => n1953, 
                           ZN => curr_proc_regs(719));
   U2712 : INV_X1 port map( A => regs(583), ZN => n1958);
   U2713 : AOI22_X1 port map( A1 => n116, A2 => regs(2119), B1 => n76, B2 => 
                           regs(1607), ZN => n1957);
   U2714 : AOI22_X1 port map( A1 => n92, A2 => regs(1095), B1 => n2, B2 => 
                           regs(71), ZN => n1956);
   U2715 : OAI211_X1 port map( C1 => n46, C2 => n1958, A => n1957, B => n1956, 
                           ZN => curr_proc_regs(71));
   U2716 : AOI22_X1 port map( A1 => n4, A2 => regs(208), B1 => n71, B2 => 
                           regs(2256), ZN => n1960);
   U2717 : AOI22_X1 port map( A1 => n80, A2 => regs(1744), B1 => n2, B2 => 
                           regs(720), ZN => n1959);
   U2718 : OAI211_X1 port map( C1 => n6, C2 => n1961, A => n1960, B => n1959, 
                           ZN => curr_proc_regs(720));
   U2719 : AOI22_X1 port map( A1 => n116, A2 => regs(209), B1 => n76, B2 => 
                           regs(2257), ZN => n1963);
   U2720 : AOI22_X1 port map( A1 => n87, A2 => regs(1745), B1 => n44, B2 => 
                           regs(721), ZN => n1962);
   U2721 : OAI211_X1 port map( C1 => n67, C2 => n1964, A => n1963, B => n1962, 
                           ZN => curr_proc_regs(721));
   U2722 : AOI22_X1 port map( A1 => n116, A2 => regs(210), B1 => n76, B2 => 
                           regs(2258), ZN => n1966);
   U2723 : AOI22_X1 port map( A1 => n95, A2 => regs(1746), B1 => n29, B2 => 
                           regs(722), ZN => n1965);
   U2724 : OAI211_X1 port map( C1 => n46, C2 => n1967, A => n1966, B => n1965, 
                           ZN => curr_proc_regs(722));
   U2725 : AOI22_X1 port map( A1 => n4, A2 => regs(211), B1 => n76, B2 => 
                           regs(2259), ZN => n1969);
   U2726 : AOI22_X1 port map( A1 => n96, A2 => regs(1747), B1 => n42, B2 => 
                           regs(723), ZN => n1968);
   U2727 : OAI211_X1 port map( C1 => n46, C2 => n1970, A => n1969, B => n1968, 
                           ZN => curr_proc_regs(723));
   U2728 : AOI22_X1 port map( A1 => n116, A2 => regs(212), B1 => n76, B2 => 
                           regs(2260), ZN => n1972);
   U2729 : AOI22_X1 port map( A1 => n58, A2 => regs(1236), B1 => n97, B2 => 
                           regs(1748), ZN => n1971);
   U2730 : OAI211_X1 port map( C1 => n22, C2 => n1973, A => n1972, B => n1971, 
                           ZN => curr_proc_regs(724));
   U2731 : AOI22_X1 port map( A1 => n116, A2 => regs(213), B1 => n76, B2 => 
                           regs(2261), ZN => n1975);
   U2732 : AOI22_X1 port map( A1 => n94, A2 => regs(1749), B1 => n39, B2 => 
                           regs(725), ZN => n1974);
   U2733 : OAI211_X1 port map( C1 => n46, C2 => n1976, A => n1975, B => n1974, 
                           ZN => curr_proc_regs(725));
   U2734 : AOI22_X1 port map( A1 => n116, A2 => regs(214), B1 => n76, B2 => 
                           regs(2262), ZN => n1978);
   U2735 : AOI22_X1 port map( A1 => n88, A2 => regs(1750), B1 => n42, B2 => 
                           regs(726), ZN => n1977);
   U2736 : OAI211_X1 port map( C1 => n46, C2 => n1979, A => n1978, B => n1977, 
                           ZN => curr_proc_regs(726));
   U2737 : AOI22_X1 port map( A1 => n116, A2 => regs(215), B1 => n76, B2 => 
                           regs(2263), ZN => n1981);
   U2738 : AOI22_X1 port map( A1 => n80, A2 => regs(1751), B1 => n24, B2 => 
                           regs(727), ZN => n1980);
   U2739 : OAI211_X1 port map( C1 => n46, C2 => n1982, A => n1981, B => n1980, 
                           ZN => curr_proc_regs(727));
   U2740 : AOI22_X1 port map( A1 => n116, A2 => regs(216), B1 => n76, B2 => 
                           regs(2264), ZN => n1984);
   U2741 : AOI22_X1 port map( A1 => n82, A2 => regs(1752), B1 => n23, B2 => 
                           regs(728), ZN => n1983);
   U2742 : OAI211_X1 port map( C1 => n1, C2 => n1985, A => n1984, B => n1983, 
                           ZN => curr_proc_regs(728));
   U2743 : AOI22_X1 port map( A1 => n116, A2 => regs(217), B1 => n3, B2 => 
                           regs(2265), ZN => n1987);
   U2744 : AOI22_X1 port map( A1 => n83, A2 => regs(1753), B1 => n39, B2 => 
                           regs(729), ZN => n1986);
   U2745 : OAI211_X1 port map( C1 => n46, C2 => n1988, A => n1987, B => n1986, 
                           ZN => curr_proc_regs(729));
   U2746 : AOI22_X1 port map( A1 => n116, A2 => regs(2120), B1 => n76, B2 => 
                           regs(1608), ZN => n1990);
   U2747 : AOI22_X1 port map( A1 => n54, A2 => regs(584), B1 => n36, B2 => 
                           regs(72), ZN => n1989);
   U2748 : OAI211_X1 port map( C1 => n101, C2 => n1991, A => n1990, B => n1989,
                           ZN => curr_proc_regs(72));
   U2749 : AOI22_X1 port map( A1 => n116, A2 => regs(218), B1 => n76, B2 => 
                           regs(2266), ZN => n1993);
   U2750 : AOI22_X1 port map( A1 => n83, A2 => regs(1754), B1 => n43, B2 => 
                           regs(730), ZN => n1992);
   U2751 : OAI211_X1 port map( C1 => n46, C2 => n1994, A => n1993, B => n1992, 
                           ZN => curr_proc_regs(730));
   U2752 : AOI22_X1 port map( A1 => n116, A2 => regs(219), B1 => n76, B2 => 
                           regs(2267), ZN => n1996);
   U2753 : AOI22_X1 port map( A1 => n62, A2 => regs(1243), B1 => n14, B2 => 
                           regs(1755), ZN => n1995);
   U2754 : OAI211_X1 port map( C1 => n22, C2 => n1997, A => n1996, B => n1995, 
                           ZN => curr_proc_regs(731));
   U2755 : AOI22_X1 port map( A1 => n116, A2 => regs(220), B1 => n76, B2 => 
                           regs(2268), ZN => n1999);
   U2756 : AOI22_X1 port map( A1 => n58, A2 => regs(1244), B1 => n14, B2 => 
                           regs(1756), ZN => n1998);
   U2757 : OAI211_X1 port map( C1 => n22, C2 => n2000, A => n1999, B => n1998, 
                           ZN => curr_proc_regs(732));
   U2758 : AOI22_X1 port map( A1 => n116, A2 => regs(221), B1 => n76, B2 => 
                           regs(2269), ZN => n2002);
   U2759 : AOI22_X1 port map( A1 => n83, A2 => regs(1757), B1 => n31, B2 => 
                           regs(733), ZN => n2001);
   U2760 : OAI211_X1 port map( C1 => n2185, C2 => n2003, A => n2002, B => n2001
                           , ZN => curr_proc_regs(733));
   U2761 : AOI22_X1 port map( A1 => n116, A2 => regs(222), B1 => n13, B2 => 
                           regs(2270), ZN => n2005);
   U2762 : AOI22_X1 port map( A1 => n60, A2 => regs(1246), B1 => n97, B2 => 
                           regs(1758), ZN => n2004);
   U2763 : OAI211_X1 port map( C1 => n22, C2 => n2006, A => n2005, B => n2004, 
                           ZN => curr_proc_regs(734));
   U2764 : AOI22_X1 port map( A1 => n116, A2 => regs(223), B1 => n69, B2 => 
                           regs(2271), ZN => n2008);
   U2765 : AOI22_X1 port map( A1 => n62, A2 => regs(1247), B1 => n14, B2 => 
                           regs(1759), ZN => n2007);
   U2766 : OAI211_X1 port map( C1 => n22, C2 => n2009, A => n2008, B => n2007, 
                           ZN => curr_proc_regs(735));
   U2767 : AOI22_X1 port map( A1 => n116, A2 => regs(224), B1 => n13, B2 => 
                           regs(2272), ZN => n2011);
   U2768 : AOI22_X1 port map( A1 => n83, A2 => regs(1760), B1 => n29, B2 => 
                           regs(736), ZN => n2010);
   U2769 : OAI211_X1 port map( C1 => n67, C2 => n2012, A => n2011, B => n2010, 
                           ZN => curr_proc_regs(736));
   U2770 : AOI22_X1 port map( A1 => n116, A2 => regs(225), B1 => n13, B2 => 
                           regs(2273), ZN => n2014);
   U2771 : AOI22_X1 port map( A1 => n83, A2 => regs(1761), B1 => n29, B2 => 
                           regs(737), ZN => n2013);
   U2772 : OAI211_X1 port map( C1 => n46, C2 => n2015, A => n2014, B => n2013, 
                           ZN => curr_proc_regs(737));
   U2773 : AOI22_X1 port map( A1 => n116, A2 => regs(226), B1 => n16, B2 => 
                           regs(2274), ZN => n2017);
   U2774 : AOI22_X1 port map( A1 => n58, A2 => regs(1250), B1 => n97, B2 => 
                           regs(1762), ZN => n2016);
   U2775 : OAI211_X1 port map( C1 => n2112, C2 => n2018, A => n2017, B => n2016
                           , ZN => curr_proc_regs(738));
   U2776 : AOI22_X1 port map( A1 => n116, A2 => regs(227), B1 => n16, B2 => 
                           regs(2275), ZN => n2020);
   U2777 : AOI22_X1 port map( A1 => n83, A2 => regs(1763), B1 => n29, B2 => 
                           regs(739), ZN => n2019);
   U2778 : OAI211_X1 port map( C1 => n46, C2 => n2021, A => n2020, B => n2019, 
                           ZN => curr_proc_regs(739));
   U2779 : AOI22_X1 port map( A1 => n116, A2 => regs(2121), B1 => n13, B2 => 
                           regs(1609), ZN => n2023);
   U2780 : AOI22_X1 port map( A1 => n62, A2 => regs(585), B1 => n29, B2 => 
                           regs(73), ZN => n2022);
   U2781 : OAI211_X1 port map( C1 => n100, C2 => n2024, A => n2023, B => n2022,
                           ZN => curr_proc_regs(73));
   U2782 : AOI22_X1 port map( A1 => n116, A2 => regs(228), B1 => n73, B2 => 
                           regs(2276), ZN => n2026);
   U2783 : AOI22_X1 port map( A1 => n83, A2 => regs(1764), B1 => n29, B2 => 
                           regs(740), ZN => n2025);
   U2784 : OAI211_X1 port map( C1 => n46, C2 => n2027, A => n2026, B => n2025, 
                           ZN => curr_proc_regs(740));
   U2785 : AOI22_X1 port map( A1 => n116, A2 => regs(229), B1 => n13, B2 => 
                           regs(2277), ZN => n2029);
   U2786 : AOI22_X1 port map( A1 => n83, A2 => regs(1765), B1 => n29, B2 => 
                           regs(741), ZN => n2028);
   U2787 : OAI211_X1 port map( C1 => n64, C2 => n2030, A => n2029, B => n2028, 
                           ZN => curr_proc_regs(741));
   U2788 : AOI22_X1 port map( A1 => n116, A2 => regs(230), B1 => n13, B2 => 
                           regs(2278), ZN => n2032);
   U2789 : AOI22_X1 port map( A1 => n83, A2 => regs(1766), B1 => n29, B2 => 
                           regs(742), ZN => n2031);
   U2790 : OAI211_X1 port map( C1 => n46, C2 => n2033, A => n2032, B => n2031, 
                           ZN => curr_proc_regs(742));
   U2791 : AOI22_X1 port map( A1 => n116, A2 => regs(231), B1 => n68, B2 => 
                           regs(2279), ZN => n2035);
   U2792 : AOI22_X1 port map( A1 => n83, A2 => regs(1767), B1 => n29, B2 => 
                           regs(743), ZN => n2034);
   U2793 : OAI211_X1 port map( C1 => n64, C2 => n2036, A => n2035, B => n2034, 
                           ZN => curr_proc_regs(743));
   U2794 : AOI22_X1 port map( A1 => n116, A2 => regs(232), B1 => n13, B2 => 
                           regs(2280), ZN => n2038);
   U2795 : AOI22_X1 port map( A1 => n83, A2 => regs(1768), B1 => n29, B2 => 
                           regs(744), ZN => n2037);
   U2796 : OAI211_X1 port map( C1 => n67, C2 => n2039, A => n2038, B => n2037, 
                           ZN => curr_proc_regs(744));
   U2797 : AOI22_X1 port map( A1 => n116, A2 => regs(233), B1 => n13, B2 => 
                           regs(2281), ZN => n2041);
   U2798 : AOI22_X1 port map( A1 => n83, A2 => regs(1769), B1 => n29, B2 => 
                           regs(745), ZN => n2040);
   U2799 : OAI211_X1 port map( C1 => n46, C2 => n2042, A => n2041, B => n2040, 
                           ZN => curr_proc_regs(745));
   U2800 : AOI22_X1 port map( A1 => n116, A2 => regs(234), B1 => n16, B2 => 
                           regs(2282), ZN => n2044);
   U2801 : AOI22_X1 port map( A1 => n79, A2 => regs(1770), B1 => n29, B2 => 
                           regs(746), ZN => n2043);
   U2802 : OAI211_X1 port map( C1 => n46, C2 => n2045, A => n2044, B => n2043, 
                           ZN => curr_proc_regs(746));
   U2803 : AOI22_X1 port map( A1 => n116, A2 => regs(235), B1 => n70, B2 => 
                           regs(2283), ZN => n2047);
   U2804 : AOI22_X1 port map( A1 => n55, A2 => regs(1259), B1 => n14, B2 => 
                           regs(1771), ZN => n2046);
   U2805 : OAI211_X1 port map( C1 => n21, C2 => n2048, A => n2047, B => n2046, 
                           ZN => curr_proc_regs(747));
   U2806 : AOI22_X1 port map( A1 => n110, A2 => regs(236), B1 => n13, B2 => 
                           regs(2284), ZN => n2050);
   U2807 : AOI22_X1 port map( A1 => n62, A2 => regs(1260), B1 => n14, B2 => 
                           regs(1772), ZN => n2049);
   U2808 : OAI211_X1 port map( C1 => n22, C2 => n2051, A => n2050, B => n2049, 
                           ZN => curr_proc_regs(748));
   U2809 : AOI22_X1 port map( A1 => n110, A2 => regs(237), B1 => n3, B2 => 
                           regs(2285), ZN => n2053);
   U2810 : AOI22_X1 port map( A1 => n80, A2 => regs(1773), B1 => n30, B2 => 
                           regs(749), ZN => n2052);
   U2811 : OAI211_X1 port map( C1 => n1, C2 => n2054, A => n2053, B => n2052, 
                           ZN => curr_proc_regs(749));
   U2812 : AOI22_X1 port map( A1 => n116, A2 => regs(2122), B1 => n3, B2 => 
                           regs(1610), ZN => n2056);
   U2813 : AOI22_X1 port map( A1 => n58, A2 => regs(586), B1 => n30, B2 => 
                           regs(74), ZN => n2055);
   U2814 : OAI211_X1 port map( C1 => n100, C2 => n2057, A => n2056, B => n2055,
                           ZN => curr_proc_regs(74));
   U2815 : AOI22_X1 port map( A1 => n110, A2 => regs(238), B1 => n9, B2 => 
                           regs(2286), ZN => n2059);
   U2816 : AOI22_X1 port map( A1 => n60, A2 => regs(1262), B1 => n14, B2 => 
                           regs(1774), ZN => n2058);
   U2817 : OAI211_X1 port map( C1 => n22, C2 => n2060, A => n2059, B => n2058, 
                           ZN => curr_proc_regs(750));
   U2818 : AOI22_X1 port map( A1 => n116, A2 => regs(239), B1 => n13, B2 => 
                           regs(2287), ZN => n2062);
   U2819 : AOI22_X1 port map( A1 => n58, A2 => regs(1263), B1 => n14, B2 => 
                           regs(1775), ZN => n2061);
   U2820 : OAI211_X1 port map( C1 => n22, C2 => n2063, A => n2062, B => n2061, 
                           ZN => curr_proc_regs(751));
   U2821 : AOI22_X1 port map( A1 => n110, A2 => regs(240), B1 => n73, B2 => 
                           regs(2288), ZN => n2065);
   U2822 : AOI22_X1 port map( A1 => n81, A2 => regs(1776), B1 => n30, B2 => 
                           regs(752), ZN => n2064);
   U2823 : OAI211_X1 port map( C1 => n46, C2 => n2066, A => n2065, B => n2064, 
                           ZN => curr_proc_regs(752));
   U2824 : AOI22_X1 port map( A1 => n103, A2 => regs(241), B1 => n71, B2 => 
                           regs(2289), ZN => n2068);
   U2825 : AOI22_X1 port map( A1 => n60, A2 => regs(1265), B1 => n14, B2 => 
                           regs(1777), ZN => n2067);
   U2826 : OAI211_X1 port map( C1 => n21, C2 => n2069, A => n2068, B => n2067, 
                           ZN => curr_proc_regs(753));
   U2827 : AOI22_X1 port map( A1 => n110, A2 => regs(242), B1 => n3, B2 => 
                           regs(2290), ZN => n2071);
   U2828 : AOI22_X1 port map( A1 => n90, A2 => regs(1778), B1 => n30, B2 => 
                           regs(754), ZN => n2070);
   U2829 : OAI211_X1 port map( C1 => n1, C2 => n2072, A => n2071, B => n2070, 
                           ZN => curr_proc_regs(754));
   U2830 : AOI22_X1 port map( A1 => win(4), A2 => regs(243), B1 => n3, B2 => 
                           regs(2291), ZN => n2074);
   U2831 : AOI22_X1 port map( A1 => n10, A2 => regs(1267), B1 => n14, B2 => 
                           regs(1779), ZN => n2073);
   U2832 : OAI211_X1 port map( C1 => n2112, C2 => n2075, A => n2074, B => n2073
                           , ZN => curr_proc_regs(755));
   U2833 : AOI22_X1 port map( A1 => n116, A2 => regs(244), B1 => n3, B2 => 
                           regs(2292), ZN => n2077);
   U2834 : AOI22_X1 port map( A1 => n10, A2 => regs(1268), B1 => n97, B2 => 
                           regs(1780), ZN => n2076);
   U2835 : OAI211_X1 port map( C1 => n22, C2 => n2078, A => n2077, B => n2076, 
                           ZN => curr_proc_regs(756));
   U2836 : AOI22_X1 port map( A1 => n116, A2 => regs(245), B1 => n3, B2 => 
                           regs(2293), ZN => n2080);
   U2837 : AOI22_X1 port map( A1 => n84, A2 => regs(1781), B1 => n30, B2 => 
                           regs(757), ZN => n2079);
   U2838 : OAI211_X1 port map( C1 => n1, C2 => n2081, A => n2080, B => n2079, 
                           ZN => curr_proc_regs(757));
   U2839 : AOI22_X1 port map( A1 => n116, A2 => regs(246), B1 => n71, B2 => 
                           regs(2294), ZN => n2083);
   U2840 : AOI22_X1 port map( A1 => n85, A2 => regs(1782), B1 => n30, B2 => 
                           regs(758), ZN => n2082);
   U2841 : OAI211_X1 port map( C1 => n1, C2 => n2084, A => n2083, B => n2082, 
                           ZN => curr_proc_regs(758));
   U2842 : AOI22_X1 port map( A1 => n110, A2 => regs(247), B1 => n68, B2 => 
                           regs(2295), ZN => n2086);
   U2843 : AOI22_X1 port map( A1 => n58, A2 => regs(1271), B1 => n97, B2 => 
                           regs(1783), ZN => n2085);
   U2844 : OAI211_X1 port map( C1 => n22, C2 => n2087, A => n2086, B => n2085, 
                           ZN => curr_proc_regs(759));
   U2845 : INV_X1 port map( A => regs(1099), ZN => n2090);
   U2846 : AOI22_X1 port map( A1 => n110, A2 => regs(2123), B1 => n73, B2 => 
                           regs(1611), ZN => n2089);
   U2847 : AOI22_X1 port map( A1 => n10, A2 => regs(587), B1 => n30, B2 => 
                           regs(75), ZN => n2088);
   U2848 : OAI211_X1 port map( C1 => n100, C2 => n2090, A => n2089, B => n2088,
                           ZN => curr_proc_regs(75));
   U2849 : AOI22_X1 port map( A1 => n116, A2 => regs(248), B1 => n16, B2 => 
                           regs(2296), ZN => n2092);
   U2850 : AOI22_X1 port map( A1 => n8, A2 => regs(1272), B1 => n14, B2 => 
                           regs(1784), ZN => n2091);
   U2851 : OAI211_X1 port map( C1 => n22, C2 => n2093, A => n2092, B => n2091, 
                           ZN => curr_proc_regs(760));
   U2852 : AOI22_X1 port map( A1 => n116, A2 => regs(249), B1 => n16, B2 => 
                           regs(2297), ZN => n2095);
   U2853 : AOI22_X1 port map( A1 => n10, A2 => regs(1273), B1 => n97, B2 => 
                           regs(1785), ZN => n2094);
   U2854 : OAI211_X1 port map( C1 => n2112, C2 => n2096, A => n2095, B => n2094
                           , ZN => curr_proc_regs(761));
   U2855 : AOI22_X1 port map( A1 => n110, A2 => regs(250), B1 => n78, B2 => 
                           regs(2298), ZN => n2098);
   U2856 : AOI22_X1 port map( A1 => n60, A2 => regs(1274), B1 => n14, B2 => 
                           regs(1786), ZN => n2097);
   U2857 : OAI211_X1 port map( C1 => n22, C2 => n2099, A => n2098, B => n2097, 
                           ZN => curr_proc_regs(762));
   U2858 : AOI22_X1 port map( A1 => n110, A2 => regs(251), B1 => n3, B2 => 
                           regs(2299), ZN => n2101);
   U2859 : AOI22_X1 port map( A1 => n86, A2 => regs(1787), B1 => n30, B2 => 
                           regs(763), ZN => n2100);
   U2860 : OAI211_X1 port map( C1 => n1, C2 => n2102, A => n2101, B => n2100, 
                           ZN => curr_proc_regs(763));
   U2861 : AOI22_X1 port map( A1 => n116, A2 => regs(252), B1 => n73, B2 => 
                           regs(2300), ZN => n2104);
   U2862 : AOI22_X1 port map( A1 => n87, A2 => regs(1788), B1 => n30, B2 => 
                           regs(764), ZN => n2103);
   U2863 : OAI211_X1 port map( C1 => n1, C2 => n2105, A => n2104, B => n2103, 
                           ZN => curr_proc_regs(764));
   U2864 : AOI22_X1 port map( A1 => n116, A2 => regs(253), B1 => n13, B2 => 
                           regs(2301), ZN => n2107);
   U2865 : AOI22_X1 port map( A1 => n57, A2 => regs(1277), B1 => n97, B2 => 
                           regs(1789), ZN => n2106);
   U2866 : OAI211_X1 port map( C1 => n22, C2 => n2108, A => n2107, B => n2106, 
                           ZN => curr_proc_regs(765));
   U2867 : AOI22_X1 port map( A1 => n116, A2 => regs(254), B1 => n71, B2 => 
                           regs(2302), ZN => n2110);
   U2868 : AOI22_X1 port map( A1 => n59, A2 => regs(1278), B1 => n97, B2 => 
                           regs(1790), ZN => n2109);
   U2869 : OAI211_X1 port map( C1 => n22, C2 => n2111, A => n2110, B => n2109, 
                           ZN => curr_proc_regs(766));
   U2870 : AOI22_X1 port map( A1 => n110, A2 => regs(255), B1 => n68, B2 => 
                           regs(2303), ZN => n2114);
   U2871 : AOI22_X1 port map( A1 => n88, A2 => regs(1791), B1 => n30, B2 => 
                           regs(767), ZN => n2113);
   U2872 : OAI211_X1 port map( C1 => n1, C2 => n2115, A => n2114, B => n2113, 
                           ZN => curr_proc_regs(767));
   U2873 : AOI22_X1 port map( A1 => n106, A2 => regs(2124), B1 => n13, B2 => 
                           regs(1612), ZN => n2117);
   U2874 : AOI22_X1 port map( A1 => n62, A2 => regs(588), B1 => n30, B2 => 
                           regs(76), ZN => n2116);
   U2875 : OAI211_X1 port map( C1 => n100, C2 => n2118, A => n2117, B => n2116,
                           ZN => curr_proc_regs(76));
   U2876 : INV_X1 port map( A => regs(589), ZN => n2121);
   U2877 : AOI22_X1 port map( A1 => n116, A2 => regs(2125), B1 => n13, B2 => 
                           regs(1613), ZN => n2120);
   U2878 : AOI22_X1 port map( A1 => n96, A2 => regs(1101), B1 => n31, B2 => 
                           regs(77), ZN => n2119);
   U2879 : OAI211_X1 port map( C1 => n1, C2 => n2121, A => n2120, B => n2119, 
                           ZN => curr_proc_regs(77));
   U2880 : AOI22_X1 port map( A1 => n110, A2 => regs(2126), B1 => n73, B2 => 
                           regs(1614), ZN => n2123);
   U2881 : AOI22_X1 port map( A1 => n58, A2 => regs(590), B1 => n31, B2 => 
                           regs(78), ZN => n2122);
   U2882 : OAI211_X1 port map( C1 => n100, C2 => n2124, A => n2123, B => n2122,
                           ZN => curr_proc_regs(78));
   U2883 : AOI22_X1 port map( A1 => n112, A2 => regs(2127), B1 => n16, B2 => 
                           regs(1615), ZN => n2126);
   U2884 : AOI22_X1 port map( A1 => n60, A2 => regs(591), B1 => n31, B2 => 
                           regs(79), ZN => n2125);
   U2885 : OAI211_X1 port map( C1 => n100, C2 => n2127, A => n2126, B => n2125,
                           ZN => curr_proc_regs(79));
   U2886 : AOI22_X1 port map( A1 => n116, A2 => regs(2055), B1 => n13, B2 => 
                           regs(1543), ZN => n2129);
   U2887 : AOI22_X1 port map( A1 => n62, A2 => regs(519), B1 => n31, B2 => 
                           regs(7), ZN => n2128);
   U2888 : OAI211_X1 port map( C1 => n100, C2 => n2130, A => n2129, B => n2128,
                           ZN => curr_proc_regs(7));
   U2889 : AOI22_X1 port map( A1 => n110, A2 => regs(2128), B1 => n13, B2 => 
                           regs(1616), ZN => n2132);
   U2890 : AOI22_X1 port map( A1 => n10, A2 => regs(592), B1 => n31, B2 => 
                           regs(80), ZN => n2131);
   U2891 : OAI211_X1 port map( C1 => n102, C2 => n2133, A => n2132, B => n2131,
                           ZN => curr_proc_regs(80));
   U2892 : AOI22_X1 port map( A1 => n111, A2 => regs(2129), B1 => n13, B2 => 
                           regs(1617), ZN => n2135);
   U2893 : AOI22_X1 port map( A1 => n58, A2 => regs(593), B1 => n31, B2 => 
                           regs(81), ZN => n2134);
   U2894 : OAI211_X1 port map( C1 => n100, C2 => n2136, A => n2135, B => n2134,
                           ZN => curr_proc_regs(81));
   U2895 : INV_X1 port map( A => regs(1106), ZN => n2139);
   U2896 : AOI22_X1 port map( A1 => n116, A2 => regs(2130), B1 => n3, B2 => 
                           regs(1618), ZN => n2138);
   U2897 : AOI22_X1 port map( A1 => n59, A2 => regs(594), B1 => n31, B2 => 
                           regs(82), ZN => n2137);
   U2898 : OAI211_X1 port map( C1 => n100, C2 => n2139, A => n2138, B => n2137,
                           ZN => curr_proc_regs(82));
   U2899 : INV_X1 port map( A => regs(1107), ZN => n2142);
   U2900 : AOI22_X1 port map( A1 => n110, A2 => regs(2131), B1 => n13, B2 => 
                           regs(1619), ZN => n2141);
   U2901 : AOI22_X1 port map( A1 => n60, A2 => regs(595), B1 => n31, B2 => 
                           regs(83), ZN => n2140);
   U2902 : OAI211_X1 port map( C1 => n101, C2 => n2142, A => n2141, B => n2140,
                           ZN => curr_proc_regs(83));
   U2903 : INV_X1 port map( A => regs(1108), ZN => n2145);
   U2904 : AOI22_X1 port map( A1 => n110, A2 => regs(2132), B1 => n13, B2 => 
                           regs(1620), ZN => n2144);
   U2905 : AOI22_X1 port map( A1 => n60, A2 => regs(596), B1 => n31, B2 => 
                           regs(84), ZN => n2143);
   U2906 : OAI211_X1 port map( C1 => n100, C2 => n2145, A => n2144, B => n2143,
                           ZN => curr_proc_regs(84));
   U2907 : INV_X1 port map( A => regs(597), ZN => n2148);
   U2908 : AOI22_X1 port map( A1 => n110, A2 => regs(2133), B1 => n13, B2 => 
                           regs(1621), ZN => n2147);
   U2909 : AOI22_X1 port map( A1 => n92, A2 => regs(1109), B1 => n31, B2 => 
                           regs(85), ZN => n2146);
   U2910 : OAI211_X1 port map( C1 => n46, C2 => n2148, A => n2147, B => n2146, 
                           ZN => curr_proc_regs(85));
   U2911 : AOI22_X1 port map( A1 => n110, A2 => regs(2134), B1 => n13, B2 => 
                           regs(1622), ZN => n2150);
   U2912 : AOI22_X1 port map( A1 => n59, A2 => regs(598), B1 => n31, B2 => 
                           regs(86), ZN => n2149);
   U2913 : OAI211_X1 port map( C1 => n100, C2 => n2151, A => n2150, B => n2149,
                           ZN => curr_proc_regs(86));
   U2914 : AOI22_X1 port map( A1 => n110, A2 => regs(2135), B1 => n3, B2 => 
                           regs(1623), ZN => n2153);
   U2915 : AOI22_X1 port map( A1 => n60, A2 => regs(599), B1 => n32, B2 => 
                           regs(87), ZN => n2152);
   U2916 : OAI211_X1 port map( C1 => n100, C2 => n2154, A => n2153, B => n2152,
                           ZN => curr_proc_regs(87));
   U2917 : AOI22_X1 port map( A1 => n110, A2 => regs(2136), B1 => n13, B2 => 
                           regs(1624), ZN => n2156);
   U2918 : AOI22_X1 port map( A1 => n60, A2 => regs(600), B1 => n32, B2 => 
                           regs(88), ZN => n2155);
   U2919 : OAI211_X1 port map( C1 => n102, C2 => n2157, A => n2156, B => n2155,
                           ZN => curr_proc_regs(88));
   U2920 : INV_X1 port map( A => regs(1113), ZN => n2160);
   U2921 : AOI22_X1 port map( A1 => n110, A2 => regs(2137), B1 => n13, B2 => 
                           regs(1625), ZN => n2159);
   U2922 : AOI22_X1 port map( A1 => n60, A2 => regs(601), B1 => n32, B2 => 
                           regs(89), ZN => n2158);
   U2923 : OAI211_X1 port map( C1 => n100, C2 => n2160, A => n2159, B => n2158,
                           ZN => curr_proc_regs(89));
   U2924 : AOI22_X1 port map( A1 => n110, A2 => regs(2056), B1 => n3, B2 => 
                           regs(1544), ZN => n2162);
   U2925 : AOI22_X1 port map( A1 => n59, A2 => regs(520), B1 => n32, B2 => 
                           regs(8), ZN => n2161);
   U2926 : OAI211_X1 port map( C1 => n100, C2 => n2163, A => n2162, B => n2161,
                           ZN => curr_proc_regs(8));
   U2927 : INV_X1 port map( A => regs(602), ZN => n2166);
   U2928 : AOI22_X1 port map( A1 => n110, A2 => regs(2138), B1 => n13, B2 => 
                           regs(1626), ZN => n2165);
   U2929 : AOI22_X1 port map( A1 => n82, A2 => regs(1114), B1 => n32, B2 => 
                           regs(90), ZN => n2164);
   U2930 : OAI211_X1 port map( C1 => n67, C2 => n2166, A => n2165, B => n2164, 
                           ZN => curr_proc_regs(90));
   U2931 : INV_X1 port map( A => regs(603), ZN => n2169);
   U2932 : AOI22_X1 port map( A1 => n110, A2 => regs(2139), B1 => n13, B2 => 
                           regs(1627), ZN => n2168);
   U2933 : AOI22_X1 port map( A1 => n84, A2 => regs(1115), B1 => n32, B2 => 
                           regs(91), ZN => n2167);
   U2934 : OAI211_X1 port map( C1 => n46, C2 => n2169, A => n2168, B => n2167, 
                           ZN => curr_proc_regs(91));
   U2935 : AOI22_X1 port map( A1 => n110, A2 => regs(2140), B1 => n11, B2 => 
                           regs(1628), ZN => n2171);
   U2936 : AOI22_X1 port map( A1 => n60, A2 => regs(604), B1 => n32, B2 => 
                           regs(92), ZN => n2170);
   U2937 : OAI211_X1 port map( C1 => n102, C2 => n2172, A => n2171, B => n2170,
                           ZN => curr_proc_regs(92));
   U2938 : INV_X1 port map( A => regs(1117), ZN => n2175);
   U2939 : AOI22_X1 port map( A1 => n110, A2 => regs(2141), B1 => n13, B2 => 
                           regs(1629), ZN => n2174);
   U2940 : AOI22_X1 port map( A1 => n59, A2 => regs(605), B1 => n32, B2 => 
                           regs(93), ZN => n2173);
   U2941 : OAI211_X1 port map( C1 => n100, C2 => n2175, A => n2174, B => n2173,
                           ZN => curr_proc_regs(93));
   U2942 : INV_X1 port map( A => regs(1118), ZN => n2178);
   U2943 : AOI22_X1 port map( A1 => n114, A2 => regs(2142), B1 => n73, B2 => 
                           regs(1630), ZN => n2177);
   U2944 : AOI22_X1 port map( A1 => n61, A2 => regs(606), B1 => n32, B2 => 
                           regs(94), ZN => n2176);
   U2945 : OAI211_X1 port map( C1 => n100, C2 => n2178, A => n2177, B => n2176,
                           ZN => curr_proc_regs(94));
   U2946 : AOI22_X1 port map( A1 => n113, A2 => regs(2143), B1 => n13, B2 => 
                           regs(1631), ZN => n2180);
   U2947 : AOI22_X1 port map( A1 => n61, A2 => regs(607), B1 => n32, B2 => 
                           regs(95), ZN => n2179);
   U2948 : OAI211_X1 port map( C1 => n100, C2 => n2181, A => n2180, B => n2179,
                           ZN => curr_proc_regs(95));
   U2949 : INV_X1 port map( A => regs(608), ZN => n2184);
   U2950 : AOI22_X1 port map( A1 => n107, A2 => regs(2144), B1 => n71, B2 => 
                           regs(1632), ZN => n2183);
   U2951 : AOI22_X1 port map( A1 => n95, A2 => regs(1120), B1 => n32, B2 => 
                           regs(96), ZN => n2182);
   U2952 : OAI211_X1 port map( C1 => n6, C2 => n2184, A => n2183, B => n2182, 
                           ZN => curr_proc_regs(96));
   U2953 : INV_X1 port map( A => regs(1121), ZN => n2188);
   U2954 : AOI22_X1 port map( A1 => n108, A2 => regs(2145), B1 => n68, B2 => 
                           regs(1633), ZN => n2187);
   U2955 : AOI22_X1 port map( A1 => n61, A2 => regs(609), B1 => n33, B2 => 
                           regs(97), ZN => n2186);
   U2956 : OAI211_X1 port map( C1 => n102, C2 => n2188, A => n2187, B => n2186,
                           ZN => curr_proc_regs(97));
   U2957 : INV_X1 port map( A => regs(1122), ZN => n2191);
   U2958 : AOI22_X1 port map( A1 => n4, A2 => regs(2146), B1 => n16, B2 => 
                           regs(1634), ZN => n2190);
   U2959 : AOI22_X1 port map( A1 => n60, A2 => regs(610), B1 => n33, B2 => 
                           regs(98), ZN => n2189);
   U2960 : OAI211_X1 port map( C1 => n100, C2 => n2191, A => n2190, B => n2189,
                           ZN => curr_proc_regs(98));
   U2961 : AOI22_X1 port map( A1 => n103, A2 => regs(2147), B1 => n16, B2 => 
                           regs(1635), ZN => n2193);
   U2962 : AOI22_X1 port map( A1 => n61, A2 => regs(611), B1 => n33, B2 => 
                           regs(99), ZN => n2192);
   U2963 : OAI211_X1 port map( C1 => n100, C2 => n2194, A => n2193, B => n2192,
                           ZN => curr_proc_regs(99));
   U2964 : INV_X1 port map( A => regs(1033), ZN => n2198);
   U2965 : AOI22_X1 port map( A1 => n105, A2 => regs(2057), B1 => n74, B2 => 
                           regs(1545), ZN => n2197);
   U2966 : AOI22_X1 port map( A1 => n5, A2 => regs(521), B1 => n33, B2 => 
                           regs(9), ZN => n2196);
   U2967 : OAI211_X1 port map( C1 => n100, C2 => n2198, A => n2197, B => n2196,
                           ZN => curr_proc_regs(9));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32.all;

entity mux_N32_M5_1 is

   port( S : in std_logic_vector (4 downto 0);  Q : in std_logic_vector (1023 
         downto 0);  Y : out std_logic_vector (31 downto 0));

end mux_N32_M5_1;

architecture SYN_behav of mux_N32_M5_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n546, n547, 
      n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, 
      n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, 
      n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, 
      n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, 
      n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, 
      n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, 
      n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, 
      n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, 
      n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, 
      n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, 
      n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, 
      n680, n681, n682, n683, n684, n685, n686, n687, n688 : std_logic;

begin
   
   U2 : AOI22_X1 port map( A1 => n674, A2 => Q(499), B1 => n673, B2 => Q(563), 
                           ZN => n1);
   U3 : AOI22_X1 port map( A1 => n676, A2 => Q(659), B1 => n675, B2 => Q(467), 
                           ZN => n2);
   U4 : AOI22_X1 port map( A1 => n678, A2 => Q(371), B1 => n677, B2 => Q(307), 
                           ZN => n3);
   U5 : AOI22_X1 port map( A1 => n680, A2 => Q(403), B1 => n679, B2 => Q(275), 
                           ZN => n4);
   U6 : NAND4_X1 port map( A1 => n1, A2 => n2, A3 => n3, A4 => n4, ZN => n5);
   U7 : AOI22_X1 port map( A1 => n682, A2 => Q(339), B1 => n681, B2 => Q(435), 
                           ZN => n6);
   U8 : AOI22_X1 port map( A1 => n684, A2 => Q(243), B1 => n683, B2 => Q(147), 
                           ZN => n7);
   U9 : AOI22_X1 port map( A1 => n686, A2 => Q(83), B1 => n685, B2 => Q(179), 
                           ZN => n8);
   U10 : AOI22_X1 port map( A1 => n688, A2 => Q(211), B1 => n687, B2 => Q(51), 
                           ZN => n9);
   U11 : NAND4_X1 port map( A1 => n6, A2 => n7, A3 => n8, A4 => n9, ZN => n10);
   U12 : AOI22_X1 port map( A1 => n657, A2 => Q(1011), B1 => n656, B2 => Q(947)
                           , ZN => n11);
   U13 : AOI22_X1 port map( A1 => n659, A2 => Q(979), B1 => n658, B2 => Q(915),
                           ZN => n12);
   U14 : AOI222_X1 port map( A1 => n661, A2 => Q(819), B1 => n662, B2 => Q(115)
                           , C1 => n660, C2 => Q(755), ZN => n13);
   U15 : NAND3_X1 port map( A1 => n11, A2 => n12, A3 => n13, ZN => n14);
   U16 : AOI22_X1 port map( A1 => n664, A2 => Q(851), B1 => n663, B2 => Q(723),
                           ZN => n15);
   U17 : AOI22_X1 port map( A1 => n666, A2 => Q(787), B1 => n665, B2 => Q(883),
                           ZN => n16);
   U18 : NAND4_X1 port map( A1 => n614, A2 => n615, A3 => n15, A4 => n16, ZN =>
                           n17);
   U19 : OR4_X1 port map( A1 => n5, A2 => n10, A3 => n14, A4 => n17, ZN => 
                           Y(19));
   U20 : AOI22_X1 port map( A1 => n674, A2 => Q(509), B1 => n673, B2 => Q(573),
                           ZN => n18);
   U21 : AOI22_X1 port map( A1 => n676, A2 => Q(669), B1 => n675, B2 => Q(477),
                           ZN => n19);
   U22 : AOI22_X1 port map( A1 => n678, A2 => Q(381), B1 => n677, B2 => Q(317),
                           ZN => n20);
   U23 : AOI22_X1 port map( A1 => n680, A2 => Q(413), B1 => n679, B2 => Q(285),
                           ZN => n21);
   U24 : NAND4_X1 port map( A1 => n18, A2 => n19, A3 => n20, A4 => n21, ZN => 
                           n22);
   U25 : AOI22_X1 port map( A1 => n682, A2 => Q(349), B1 => n681, B2 => Q(445),
                           ZN => n23);
   U26 : AOI22_X1 port map( A1 => n684, A2 => Q(253), B1 => n683, B2 => Q(157),
                           ZN => n24);
   U27 : AOI22_X1 port map( A1 => n686, A2 => Q(93), B1 => n685, B2 => Q(189), 
                           ZN => n25);
   U28 : AOI22_X1 port map( A1 => n688, A2 => Q(221), B1 => n687, B2 => Q(61), 
                           ZN => n26);
   U29 : NAND4_X1 port map( A1 => n23, A2 => n24, A3 => n25, A4 => n26, ZN => 
                           n27);
   U30 : AOI22_X1 port map( A1 => n657, A2 => Q(1021), B1 => n656, B2 => Q(957)
                           , ZN => n28);
   U31 : AOI22_X1 port map( A1 => n659, A2 => Q(989), B1 => n658, B2 => Q(925),
                           ZN => n29);
   U32 : AOI222_X1 port map( A1 => n661, A2 => Q(829), B1 => n662, B2 => Q(125)
                           , C1 => n660, C2 => Q(765), ZN => n30);
   U33 : NAND3_X1 port map( A1 => n28, A2 => n29, A3 => n30, ZN => n31);
   U34 : AOI22_X1 port map( A1 => n664, A2 => Q(861), B1 => n663, B2 => Q(733),
                           ZN => n32);
   U35 : AOI22_X1 port map( A1 => n666, A2 => Q(797), B1 => n665, B2 => Q(893),
                           ZN => n33);
   U36 : NAND4_X1 port map( A1 => n636, A2 => n637, A3 => n32, A4 => n33, ZN =>
                           n34);
   U37 : OR4_X1 port map( A1 => n22, A2 => n27, A3 => n31, A4 => n34, ZN => 
                           Y(29));
   U38 : AOI22_X1 port map( A1 => n674, A2 => Q(497), B1 => n673, B2 => Q(561),
                           ZN => n35);
   U39 : AOI22_X1 port map( A1 => n676, A2 => Q(657), B1 => n675, B2 => Q(465),
                           ZN => n36);
   U40 : AOI22_X1 port map( A1 => n678, A2 => Q(369), B1 => n677, B2 => Q(305),
                           ZN => n37);
   U41 : AOI22_X1 port map( A1 => n680, A2 => Q(401), B1 => n679, B2 => Q(273),
                           ZN => n38);
   U42 : NAND4_X1 port map( A1 => n35, A2 => n36, A3 => n37, A4 => n38, ZN => 
                           n39);
   U43 : AOI22_X1 port map( A1 => n682, A2 => Q(337), B1 => n681, B2 => Q(433),
                           ZN => n40);
   U44 : AOI22_X1 port map( A1 => n684, A2 => Q(241), B1 => n683, B2 => Q(145),
                           ZN => n41);
   U45 : AOI22_X1 port map( A1 => n686, A2 => Q(81), B1 => n685, B2 => Q(177), 
                           ZN => n42);
   U46 : AOI22_X1 port map( A1 => n688, A2 => Q(209), B1 => n687, B2 => Q(49), 
                           ZN => n43);
   U47 : NAND4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n44);
   U48 : AOI22_X1 port map( A1 => n657, A2 => Q(1009), B1 => n656, B2 => Q(945)
                           , ZN => n45);
   U49 : AOI22_X1 port map( A1 => n659, A2 => Q(977), B1 => n658, B2 => Q(913),
                           ZN => n46);
   U50 : AOI222_X1 port map( A1 => n661, A2 => Q(817), B1 => n662, B2 => Q(113)
                           , C1 => n660, C2 => Q(753), ZN => n47);
   U51 : NAND3_X1 port map( A1 => n45, A2 => n46, A3 => n47, ZN => n48);
   U52 : AOI22_X1 port map( A1 => n664, A2 => Q(849), B1 => n663, B2 => Q(721),
                           ZN => n49);
   U53 : AOI22_X1 port map( A1 => n666, A2 => Q(785), B1 => n665, B2 => Q(881),
                           ZN => n50);
   U54 : NAND4_X1 port map( A1 => n610, A2 => n611, A3 => n49, A4 => n50, ZN =>
                           n51);
   U55 : OR4_X1 port map( A1 => n39, A2 => n44, A3 => n48, A4 => n51, ZN => 
                           Y(17));
   U56 : AOI22_X1 port map( A1 => n674, A2 => Q(498), B1 => n673, B2 => Q(562),
                           ZN => n52);
   U57 : AOI22_X1 port map( A1 => n676, A2 => Q(658), B1 => n675, B2 => Q(466),
                           ZN => n53);
   U58 : AOI22_X1 port map( A1 => n678, A2 => Q(370), B1 => n677, B2 => Q(306),
                           ZN => n54);
   U59 : AOI22_X1 port map( A1 => n680, A2 => Q(402), B1 => n679, B2 => Q(274),
                           ZN => n55);
   U60 : NAND4_X1 port map( A1 => n52, A2 => n53, A3 => n54, A4 => n55, ZN => 
                           n56);
   U61 : AOI22_X1 port map( A1 => n682, A2 => Q(338), B1 => n681, B2 => Q(434),
                           ZN => n57);
   U62 : AOI22_X1 port map( A1 => n684, A2 => Q(242), B1 => n683, B2 => Q(146),
                           ZN => n58);
   U63 : AOI22_X1 port map( A1 => n686, A2 => Q(82), B1 => n685, B2 => Q(178), 
                           ZN => n59);
   U64 : AOI22_X1 port map( A1 => n688, A2 => Q(210), B1 => n687, B2 => Q(50), 
                           ZN => n60);
   U65 : NAND4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           n61);
   U66 : AOI22_X1 port map( A1 => n657, A2 => Q(1010), B1 => n656, B2 => Q(946)
                           , ZN => n62);
   U67 : AOI22_X1 port map( A1 => n659, A2 => Q(978), B1 => n658, B2 => Q(914),
                           ZN => n63);
   U68 : AOI222_X1 port map( A1 => n661, A2 => Q(818), B1 => n662, B2 => Q(114)
                           , C1 => n660, C2 => Q(754), ZN => n64);
   U69 : NAND3_X1 port map( A1 => n62, A2 => n63, A3 => n64, ZN => n65);
   U70 : AOI22_X1 port map( A1 => n664, A2 => Q(850), B1 => n663, B2 => Q(722),
                           ZN => n66);
   U71 : AOI22_X1 port map( A1 => n666, A2 => Q(786), B1 => n665, B2 => Q(882),
                           ZN => n67);
   U72 : NAND4_X1 port map( A1 => n612, A2 => n613, A3 => n66, A4 => n67, ZN =>
                           n68);
   U73 : OR4_X1 port map( A1 => n56, A2 => n61, A3 => n65, A4 => n68, ZN => 
                           Y(18));
   U74 : AOI22_X1 port map( A1 => n674, A2 => Q(495), B1 => n673, B2 => Q(559),
                           ZN => n69);
   U75 : AOI22_X1 port map( A1 => n676, A2 => Q(655), B1 => n675, B2 => Q(463),
                           ZN => n70);
   U76 : AOI22_X1 port map( A1 => n678, A2 => Q(367), B1 => n677, B2 => Q(303),
                           ZN => n71);
   U77 : AOI22_X1 port map( A1 => n680, A2 => Q(399), B1 => n679, B2 => Q(271),
                           ZN => n72);
   U78 : NAND4_X1 port map( A1 => n69, A2 => n70, A3 => n71, A4 => n72, ZN => 
                           n73);
   U79 : AOI22_X1 port map( A1 => n682, A2 => Q(335), B1 => n681, B2 => Q(431),
                           ZN => n74);
   U80 : AOI22_X1 port map( A1 => n684, A2 => Q(239), B1 => n683, B2 => Q(143),
                           ZN => n75);
   U81 : AOI22_X1 port map( A1 => n686, A2 => Q(79), B1 => n685, B2 => Q(175), 
                           ZN => n76);
   U82 : AOI22_X1 port map( A1 => n688, A2 => Q(207), B1 => n687, B2 => Q(47), 
                           ZN => n77);
   U83 : NAND4_X1 port map( A1 => n74, A2 => n75, A3 => n76, A4 => n77, ZN => 
                           n78);
   U84 : AOI22_X1 port map( A1 => n657, A2 => Q(1007), B1 => n656, B2 => Q(943)
                           , ZN => n79);
   U85 : AOI22_X1 port map( A1 => n659, A2 => Q(975), B1 => n658, B2 => Q(911),
                           ZN => n80);
   U86 : AOI222_X1 port map( A1 => n661, A2 => Q(815), B1 => n662, B2 => Q(111)
                           , C1 => n660, C2 => Q(751), ZN => n81);
   U87 : NAND3_X1 port map( A1 => n79, A2 => n80, A3 => n81, ZN => n82);
   U88 : AOI22_X1 port map( A1 => n664, A2 => Q(847), B1 => n663, B2 => Q(719),
                           ZN => n83);
   U89 : AOI22_X1 port map( A1 => n666, A2 => Q(783), B1 => n665, B2 => Q(879),
                           ZN => n84);
   U90 : NAND4_X1 port map( A1 => n606, A2 => n607, A3 => n83, A4 => n84, ZN =>
                           n85);
   U91 : OR4_X1 port map( A1 => n73, A2 => n78, A3 => n82, A4 => n85, ZN => 
                           Y(15));
   U92 : AOI22_X1 port map( A1 => n674, A2 => Q(496), B1 => n673, B2 => Q(560),
                           ZN => n86);
   U93 : AOI22_X1 port map( A1 => n676, A2 => Q(656), B1 => n675, B2 => Q(464),
                           ZN => n87);
   U94 : AOI22_X1 port map( A1 => n678, A2 => Q(368), B1 => n677, B2 => Q(304),
                           ZN => n88);
   U95 : AOI22_X1 port map( A1 => n680, A2 => Q(400), B1 => n679, B2 => Q(272),
                           ZN => n89);
   U96 : NAND4_X1 port map( A1 => n86, A2 => n87, A3 => n88, A4 => n89, ZN => 
                           n90);
   U97 : AOI22_X1 port map( A1 => n682, A2 => Q(336), B1 => n681, B2 => Q(432),
                           ZN => n91);
   U98 : AOI22_X1 port map( A1 => n684, A2 => Q(240), B1 => n683, B2 => Q(144),
                           ZN => n92);
   U99 : AOI22_X1 port map( A1 => n686, A2 => Q(80), B1 => n685, B2 => Q(176), 
                           ZN => n93);
   U100 : AOI22_X1 port map( A1 => n688, A2 => Q(208), B1 => n687, B2 => Q(48),
                           ZN => n94);
   U101 : NAND4_X1 port map( A1 => n91, A2 => n92, A3 => n93, A4 => n94, ZN => 
                           n95);
   U102 : AOI22_X1 port map( A1 => n657, A2 => Q(1008), B1 => n656, B2 => 
                           Q(944), ZN => n96);
   U103 : AOI22_X1 port map( A1 => n659, A2 => Q(976), B1 => n658, B2 => Q(912)
                           , ZN => n97);
   U104 : AOI222_X1 port map( A1 => n661, A2 => Q(816), B1 => n662, B2 => 
                           Q(112), C1 => n660, C2 => Q(752), ZN => n98);
   U105 : NAND3_X1 port map( A1 => n96, A2 => n97, A3 => n98, ZN => n99);
   U106 : AOI22_X1 port map( A1 => n664, A2 => Q(848), B1 => n663, B2 => Q(720)
                           , ZN => n100);
   U107 : AOI22_X1 port map( A1 => n666, A2 => Q(784), B1 => n665, B2 => Q(880)
                           , ZN => n101);
   U108 : NAND4_X1 port map( A1 => n608, A2 => n609, A3 => n100, A4 => n101, ZN
                           => n102);
   U109 : OR4_X1 port map( A1 => n90, A2 => n95, A3 => n99, A4 => n102, ZN => 
                           Y(16));
   U110 : AOI22_X1 port map( A1 => n674, A2 => Q(493), B1 => n673, B2 => Q(557)
                           , ZN => n103);
   U111 : AOI22_X1 port map( A1 => n676, A2 => Q(653), B1 => n675, B2 => Q(461)
                           , ZN => n104);
   U112 : AOI22_X1 port map( A1 => n678, A2 => Q(365), B1 => n677, B2 => Q(301)
                           , ZN => n105);
   U113 : AOI22_X1 port map( A1 => n680, A2 => Q(397), B1 => n679, B2 => Q(269)
                           , ZN => n106);
   U114 : NAND4_X1 port map( A1 => n103, A2 => n104, A3 => n105, A4 => n106, ZN
                           => n107);
   U115 : AOI22_X1 port map( A1 => n682, A2 => Q(333), B1 => n681, B2 => Q(429)
                           , ZN => n108);
   U116 : AOI22_X1 port map( A1 => n684, A2 => Q(237), B1 => n683, B2 => Q(141)
                           , ZN => n109);
   U117 : AOI22_X1 port map( A1 => n686, A2 => Q(77), B1 => n685, B2 => Q(173),
                           ZN => n110);
   U118 : AOI22_X1 port map( A1 => n688, A2 => Q(205), B1 => n687, B2 => Q(45),
                           ZN => n111);
   U119 : NAND4_X1 port map( A1 => n108, A2 => n109, A3 => n110, A4 => n111, ZN
                           => n112);
   U120 : AOI22_X1 port map( A1 => n657, A2 => Q(1005), B1 => n656, B2 => 
                           Q(941), ZN => n113);
   U121 : AOI22_X1 port map( A1 => n659, A2 => Q(973), B1 => n658, B2 => Q(909)
                           , ZN => n114);
   U122 : AOI222_X1 port map( A1 => n661, A2 => Q(813), B1 => n662, B2 => 
                           Q(109), C1 => n660, C2 => Q(749), ZN => n115);
   U123 : NAND3_X1 port map( A1 => n113, A2 => n114, A3 => n115, ZN => n116);
   U124 : AOI22_X1 port map( A1 => n664, A2 => Q(845), B1 => n663, B2 => Q(717)
                           , ZN => n117);
   U125 : AOI22_X1 port map( A1 => n666, A2 => Q(781), B1 => n665, B2 => Q(877)
                           , ZN => n118);
   U126 : NAND4_X1 port map( A1 => n602, A2 => n603, A3 => n117, A4 => n118, ZN
                           => n119);
   U127 : OR4_X1 port map( A1 => n107, A2 => n112, A3 => n116, A4 => n119, ZN 
                           => Y(13));
   U128 : AOI22_X1 port map( A1 => n674, A2 => Q(494), B1 => n673, B2 => Q(558)
                           , ZN => n120);
   U129 : AOI22_X1 port map( A1 => n676, A2 => Q(654), B1 => n675, B2 => Q(462)
                           , ZN => n121);
   U130 : AOI22_X1 port map( A1 => n678, A2 => Q(366), B1 => n677, B2 => Q(302)
                           , ZN => n122);
   U131 : AOI22_X1 port map( A1 => n680, A2 => Q(398), B1 => n679, B2 => Q(270)
                           , ZN => n123);
   U132 : NAND4_X1 port map( A1 => n120, A2 => n121, A3 => n122, A4 => n123, ZN
                           => n124);
   U133 : AOI22_X1 port map( A1 => n682, A2 => Q(334), B1 => n681, B2 => Q(430)
                           , ZN => n125);
   U134 : AOI22_X1 port map( A1 => n684, A2 => Q(238), B1 => n683, B2 => Q(142)
                           , ZN => n126);
   U135 : AOI22_X1 port map( A1 => n686, A2 => Q(78), B1 => n685, B2 => Q(174),
                           ZN => n127);
   U136 : AOI22_X1 port map( A1 => n688, A2 => Q(206), B1 => n687, B2 => Q(46),
                           ZN => n128);
   U137 : NAND4_X1 port map( A1 => n125, A2 => n126, A3 => n127, A4 => n128, ZN
                           => n129);
   U138 : AOI22_X1 port map( A1 => n657, A2 => Q(1006), B1 => n656, B2 => 
                           Q(942), ZN => n130);
   U139 : AOI22_X1 port map( A1 => n659, A2 => Q(974), B1 => n658, B2 => Q(910)
                           , ZN => n131);
   U140 : AOI222_X1 port map( A1 => n661, A2 => Q(814), B1 => n662, B2 => 
                           Q(110), C1 => n660, C2 => Q(750), ZN => n132);
   U141 : NAND3_X1 port map( A1 => n130, A2 => n131, A3 => n132, ZN => n133);
   U142 : AOI22_X1 port map( A1 => n664, A2 => Q(846), B1 => n663, B2 => Q(718)
                           , ZN => n134);
   U143 : AOI22_X1 port map( A1 => n666, A2 => Q(782), B1 => n665, B2 => Q(878)
                           , ZN => n135);
   U144 : NAND4_X1 port map( A1 => n604, A2 => n605, A3 => n134, A4 => n135, ZN
                           => n136);
   U145 : OR4_X1 port map( A1 => n124, A2 => n129, A3 => n133, A4 => n136, ZN 
                           => Y(14));
   U146 : AOI22_X1 port map( A1 => n562, A2 => Q(510), B1 => n561, B2 => Q(574)
                           , ZN => n137);
   U147 : AOI22_X1 port map( A1 => n564, A2 => Q(670), B1 => n563, B2 => Q(478)
                           , ZN => n138);
   U148 : AOI22_X1 port map( A1 => n566, A2 => Q(382), B1 => n565, B2 => Q(318)
                           , ZN => n139);
   U149 : AOI22_X1 port map( A1 => n568, A2 => Q(414), B1 => n567, B2 => Q(286)
                           , ZN => n140);
   U150 : NAND4_X1 port map( A1 => n137, A2 => n138, A3 => n139, A4 => n140, ZN
                           => n141);
   U151 : AOI22_X1 port map( A1 => n570, A2 => Q(350), B1 => n569, B2 => Q(446)
                           , ZN => n142);
   U152 : AOI22_X1 port map( A1 => n572, A2 => Q(254), B1 => n571, B2 => Q(158)
                           , ZN => n143);
   U153 : AOI22_X1 port map( A1 => n574, A2 => Q(94), B1 => n573, B2 => Q(190),
                           ZN => n144);
   U154 : AOI22_X1 port map( A1 => n576, A2 => Q(222), B1 => n575, B2 => Q(62),
                           ZN => n145);
   U155 : NAND4_X1 port map( A1 => n142, A2 => n143, A3 => n144, A4 => n145, ZN
                           => n146);
   U156 : AOI22_X1 port map( A1 => n547, A2 => Q(1022), B1 => n546, B2 => 
                           Q(958), ZN => n147);
   U157 : AOI22_X1 port map( A1 => n549, A2 => Q(990), B1 => n548, B2 => Q(926)
                           , ZN => n148);
   U158 : AOI222_X1 port map( A1 => n551, A2 => Q(830), B1 => n552, B2 => 
                           Q(126), C1 => n550, C2 => Q(766), ZN => n149);
   U159 : NAND3_X1 port map( A1 => n147, A2 => n148, A3 => n149, ZN => n150);
   U160 : AOI22_X1 port map( A1 => n554, A2 => Q(862), B1 => n553, B2 => Q(734)
                           , ZN => n151);
   U161 : AOI22_X1 port map( A1 => n556, A2 => Q(798), B1 => n555, B2 => Q(894)
                           , ZN => n152);
   U162 : NAND4_X1 port map( A1 => n640, A2 => n641, A3 => n151, A4 => n152, ZN
                           => n153);
   U163 : OR4_X1 port map( A1 => n141, A2 => n146, A3 => n150, A4 => n153, ZN 
                           => Y(30));
   U164 : AOI22_X1 port map( A1 => n562, A2 => Q(508), B1 => n561, B2 => Q(572)
                           , ZN => n154);
   U165 : AOI22_X1 port map( A1 => n564, A2 => Q(668), B1 => n563, B2 => Q(476)
                           , ZN => n155);
   U166 : AOI22_X1 port map( A1 => n566, A2 => Q(380), B1 => n565, B2 => Q(316)
                           , ZN => n156);
   U167 : AOI22_X1 port map( A1 => n568, A2 => Q(412), B1 => n567, B2 => Q(284)
                           , ZN => n157);
   U168 : NAND4_X1 port map( A1 => n154, A2 => n155, A3 => n156, A4 => n157, ZN
                           => n158);
   U169 : AOI22_X1 port map( A1 => n570, A2 => Q(348), B1 => n569, B2 => Q(444)
                           , ZN => n159);
   U170 : AOI22_X1 port map( A1 => n572, A2 => Q(252), B1 => n571, B2 => Q(156)
                           , ZN => n160);
   U171 : AOI22_X1 port map( A1 => n574, A2 => Q(92), B1 => n573, B2 => Q(188),
                           ZN => n161);
   U172 : AOI22_X1 port map( A1 => n576, A2 => Q(220), B1 => n575, B2 => Q(60),
                           ZN => n162);
   U173 : NAND4_X1 port map( A1 => n159, A2 => n160, A3 => n161, A4 => n162, ZN
                           => n163);
   U174 : AOI22_X1 port map( A1 => n547, A2 => Q(1020), B1 => n546, B2 => 
                           Q(956), ZN => n164);
   U175 : AOI22_X1 port map( A1 => n549, A2 => Q(988), B1 => n548, B2 => Q(924)
                           , ZN => n165);
   U176 : AOI222_X1 port map( A1 => n551, A2 => Q(828), B1 => n552, B2 => 
                           Q(124), C1 => n550, C2 => Q(764), ZN => n166);
   U177 : NAND3_X1 port map( A1 => n164, A2 => n165, A3 => n166, ZN => n167);
   U178 : AOI22_X1 port map( A1 => n554, A2 => Q(860), B1 => n553, B2 => Q(732)
                           , ZN => n168);
   U179 : AOI22_X1 port map( A1 => n556, A2 => Q(796), B1 => n555, B2 => Q(892)
                           , ZN => n169);
   U180 : NAND4_X1 port map( A1 => n634, A2 => n635, A3 => n168, A4 => n169, ZN
                           => n170);
   U181 : OR4_X1 port map( A1 => n158, A2 => n163, A3 => n167, A4 => n170, ZN 
                           => Y(28));
   U182 : AOI22_X1 port map( A1 => n562, A2 => Q(507), B1 => n561, B2 => Q(571)
                           , ZN => n171);
   U183 : AOI22_X1 port map( A1 => n564, A2 => Q(667), B1 => n563, B2 => Q(475)
                           , ZN => n172);
   U184 : AOI22_X1 port map( A1 => n566, A2 => Q(379), B1 => n565, B2 => Q(315)
                           , ZN => n173);
   U185 : AOI22_X1 port map( A1 => n568, A2 => Q(411), B1 => n567, B2 => Q(283)
                           , ZN => n174);
   U186 : NAND4_X1 port map( A1 => n171, A2 => n172, A3 => n173, A4 => n174, ZN
                           => n175);
   U187 : AOI22_X1 port map( A1 => n570, A2 => Q(347), B1 => n569, B2 => Q(443)
                           , ZN => n176);
   U188 : AOI22_X1 port map( A1 => n572, A2 => Q(251), B1 => n571, B2 => Q(155)
                           , ZN => n177);
   U189 : AOI22_X1 port map( A1 => n574, A2 => Q(91), B1 => n573, B2 => Q(187),
                           ZN => n178);
   U190 : AOI22_X1 port map( A1 => n576, A2 => Q(219), B1 => n575, B2 => Q(59),
                           ZN => n179);
   U191 : NAND4_X1 port map( A1 => n176, A2 => n177, A3 => n178, A4 => n179, ZN
                           => n180);
   U192 : AOI22_X1 port map( A1 => n547, A2 => Q(1019), B1 => n546, B2 => 
                           Q(955), ZN => n181);
   U193 : AOI22_X1 port map( A1 => n549, A2 => Q(987), B1 => n548, B2 => Q(923)
                           , ZN => n182);
   U194 : AOI222_X1 port map( A1 => n551, A2 => Q(827), B1 => n552, B2 => 
                           Q(123), C1 => n550, C2 => Q(763), ZN => n183);
   U195 : NAND3_X1 port map( A1 => n181, A2 => n182, A3 => n183, ZN => n184);
   U196 : AOI22_X1 port map( A1 => n554, A2 => Q(859), B1 => n553, B2 => Q(731)
                           , ZN => n185);
   U197 : AOI22_X1 port map( A1 => n556, A2 => Q(795), B1 => n555, B2 => Q(891)
                           , ZN => n186);
   U198 : NAND4_X1 port map( A1 => n632, A2 => n633, A3 => n185, A4 => n186, ZN
                           => n187);
   U199 : OR4_X1 port map( A1 => n175, A2 => n180, A3 => n184, A4 => n187, ZN 
                           => Y(27));
   U200 : AOI22_X1 port map( A1 => n562, A2 => Q(506), B1 => n561, B2 => Q(570)
                           , ZN => n188);
   U201 : AOI22_X1 port map( A1 => n564, A2 => Q(666), B1 => n563, B2 => Q(474)
                           , ZN => n189);
   U202 : AOI22_X1 port map( A1 => n566, A2 => Q(378), B1 => n565, B2 => Q(314)
                           , ZN => n190);
   U203 : AOI22_X1 port map( A1 => n568, A2 => Q(410), B1 => n567, B2 => Q(282)
                           , ZN => n191);
   U204 : NAND4_X1 port map( A1 => n188, A2 => n189, A3 => n190, A4 => n191, ZN
                           => n192);
   U205 : AOI22_X1 port map( A1 => n570, A2 => Q(346), B1 => n569, B2 => Q(442)
                           , ZN => n193);
   U206 : AOI22_X1 port map( A1 => n572, A2 => Q(250), B1 => n571, B2 => Q(154)
                           , ZN => n194);
   U207 : AOI22_X1 port map( A1 => n574, A2 => Q(90), B1 => n573, B2 => Q(186),
                           ZN => n195);
   U208 : AOI22_X1 port map( A1 => n576, A2 => Q(218), B1 => n575, B2 => Q(58),
                           ZN => n196);
   U209 : NAND4_X1 port map( A1 => n193, A2 => n194, A3 => n195, A4 => n196, ZN
                           => n197);
   U210 : AOI22_X1 port map( A1 => n547, A2 => Q(1018), B1 => n546, B2 => 
                           Q(954), ZN => n198);
   U211 : AOI22_X1 port map( A1 => n549, A2 => Q(986), B1 => n548, B2 => Q(922)
                           , ZN => n199);
   U212 : AOI222_X1 port map( A1 => n551, A2 => Q(826), B1 => n552, B2 => 
                           Q(122), C1 => n550, C2 => Q(762), ZN => n200);
   U213 : NAND3_X1 port map( A1 => n198, A2 => n199, A3 => n200, ZN => n201);
   U214 : AOI22_X1 port map( A1 => n554, A2 => Q(858), B1 => n553, B2 => Q(730)
                           , ZN => n202);
   U215 : AOI22_X1 port map( A1 => n556, A2 => Q(794), B1 => n555, B2 => Q(890)
                           , ZN => n203);
   U216 : NAND4_X1 port map( A1 => n630, A2 => n631, A3 => n202, A4 => n203, ZN
                           => n204);
   U217 : OR4_X1 port map( A1 => n192, A2 => n197, A3 => n201, A4 => n204, ZN 
                           => Y(26));
   U218 : AOI22_X1 port map( A1 => n562, A2 => Q(505), B1 => n561, B2 => Q(569)
                           , ZN => n205);
   U219 : AOI22_X1 port map( A1 => n564, A2 => Q(665), B1 => n563, B2 => Q(473)
                           , ZN => n206);
   U220 : AOI22_X1 port map( A1 => n566, A2 => Q(377), B1 => n565, B2 => Q(313)
                           , ZN => n207);
   U221 : AOI22_X1 port map( A1 => n568, A2 => Q(409), B1 => n567, B2 => Q(281)
                           , ZN => n208);
   U222 : NAND4_X1 port map( A1 => n205, A2 => n206, A3 => n207, A4 => n208, ZN
                           => n209);
   U223 : AOI22_X1 port map( A1 => n570, A2 => Q(345), B1 => n569, B2 => Q(441)
                           , ZN => n210);
   U224 : AOI22_X1 port map( A1 => n572, A2 => Q(249), B1 => n571, B2 => Q(153)
                           , ZN => n211);
   U225 : AOI22_X1 port map( A1 => n574, A2 => Q(89), B1 => n573, B2 => Q(185),
                           ZN => n212);
   U226 : AOI22_X1 port map( A1 => n576, A2 => Q(217), B1 => n575, B2 => Q(57),
                           ZN => n213);
   U227 : NAND4_X1 port map( A1 => n210, A2 => n211, A3 => n212, A4 => n213, ZN
                           => n214);
   U228 : AOI22_X1 port map( A1 => n547, A2 => Q(1017), B1 => n546, B2 => 
                           Q(953), ZN => n215);
   U229 : AOI22_X1 port map( A1 => n549, A2 => Q(985), B1 => n548, B2 => Q(921)
                           , ZN => n216);
   U230 : AOI222_X1 port map( A1 => n551, A2 => Q(825), B1 => n552, B2 => 
                           Q(121), C1 => n550, C2 => Q(761), ZN => n217);
   U231 : NAND3_X1 port map( A1 => n215, A2 => n216, A3 => n217, ZN => n218);
   U232 : AOI22_X1 port map( A1 => n554, A2 => Q(857), B1 => n553, B2 => Q(729)
                           , ZN => n219);
   U233 : AOI22_X1 port map( A1 => n556, A2 => Q(793), B1 => n555, B2 => Q(889)
                           , ZN => n220);
   U234 : NAND4_X1 port map( A1 => n628, A2 => n629, A3 => n219, A4 => n220, ZN
                           => n221);
   U235 : OR4_X1 port map( A1 => n209, A2 => n214, A3 => n218, A4 => n221, ZN 
                           => Y(25));
   U236 : AOI22_X1 port map( A1 => n562, A2 => Q(504), B1 => n561, B2 => Q(568)
                           , ZN => n222);
   U237 : AOI22_X1 port map( A1 => n564, A2 => Q(664), B1 => n563, B2 => Q(472)
                           , ZN => n223);
   U238 : AOI22_X1 port map( A1 => n566, A2 => Q(376), B1 => n565, B2 => Q(312)
                           , ZN => n224);
   U239 : AOI22_X1 port map( A1 => n568, A2 => Q(408), B1 => n567, B2 => Q(280)
                           , ZN => n225);
   U240 : NAND4_X1 port map( A1 => n222, A2 => n223, A3 => n224, A4 => n225, ZN
                           => n226);
   U241 : AOI22_X1 port map( A1 => n570, A2 => Q(344), B1 => n569, B2 => Q(440)
                           , ZN => n227);
   U242 : AOI22_X1 port map( A1 => n572, A2 => Q(248), B1 => n571, B2 => Q(152)
                           , ZN => n228);
   U243 : AOI22_X1 port map( A1 => n574, A2 => Q(88), B1 => n573, B2 => Q(184),
                           ZN => n229);
   U244 : AOI22_X1 port map( A1 => n576, A2 => Q(216), B1 => n575, B2 => Q(56),
                           ZN => n230);
   U245 : NAND4_X1 port map( A1 => n227, A2 => n228, A3 => n229, A4 => n230, ZN
                           => n231);
   U246 : AOI22_X1 port map( A1 => n547, A2 => Q(1016), B1 => n546, B2 => 
                           Q(952), ZN => n232);
   U247 : AOI22_X1 port map( A1 => n549, A2 => Q(984), B1 => n548, B2 => Q(920)
                           , ZN => n233);
   U248 : AOI222_X1 port map( A1 => n551, A2 => Q(824), B1 => n552, B2 => 
                           Q(120), C1 => n550, C2 => Q(760), ZN => n234);
   U249 : NAND3_X1 port map( A1 => n232, A2 => n233, A3 => n234, ZN => n235);
   U250 : AOI22_X1 port map( A1 => n554, A2 => Q(856), B1 => n553, B2 => Q(728)
                           , ZN => n236);
   U251 : AOI22_X1 port map( A1 => n556, A2 => Q(792), B1 => n555, B2 => Q(888)
                           , ZN => n237);
   U252 : NAND4_X1 port map( A1 => n626, A2 => n627, A3 => n236, A4 => n237, ZN
                           => n238);
   U253 : OR4_X1 port map( A1 => n226, A2 => n231, A3 => n235, A4 => n238, ZN 
                           => Y(24));
   U254 : AOI22_X1 port map( A1 => n562, A2 => Q(503), B1 => n561, B2 => Q(567)
                           , ZN => n239);
   U255 : AOI22_X1 port map( A1 => n564, A2 => Q(663), B1 => n563, B2 => Q(471)
                           , ZN => n240);
   U256 : AOI22_X1 port map( A1 => n566, A2 => Q(375), B1 => n565, B2 => Q(311)
                           , ZN => n241);
   U257 : AOI22_X1 port map( A1 => n568, A2 => Q(407), B1 => n567, B2 => Q(279)
                           , ZN => n242);
   U258 : NAND4_X1 port map( A1 => n239, A2 => n240, A3 => n241, A4 => n242, ZN
                           => n243);
   U259 : AOI22_X1 port map( A1 => n570, A2 => Q(343), B1 => n569, B2 => Q(439)
                           , ZN => n244);
   U260 : AOI22_X1 port map( A1 => n572, A2 => Q(247), B1 => n571, B2 => Q(151)
                           , ZN => n245);
   U261 : AOI22_X1 port map( A1 => n574, A2 => Q(87), B1 => n573, B2 => Q(183),
                           ZN => n246);
   U262 : AOI22_X1 port map( A1 => n576, A2 => Q(215), B1 => n575, B2 => Q(55),
                           ZN => n247);
   U263 : NAND4_X1 port map( A1 => n244, A2 => n245, A3 => n246, A4 => n247, ZN
                           => n248);
   U264 : AOI22_X1 port map( A1 => n547, A2 => Q(1015), B1 => n546, B2 => 
                           Q(951), ZN => n249);
   U265 : AOI22_X1 port map( A1 => n549, A2 => Q(983), B1 => n548, B2 => Q(919)
                           , ZN => n250);
   U266 : AOI222_X1 port map( A1 => n551, A2 => Q(823), B1 => n552, B2 => 
                           Q(119), C1 => n550, C2 => Q(759), ZN => n251);
   U267 : NAND3_X1 port map( A1 => n249, A2 => n250, A3 => n251, ZN => n252);
   U268 : AOI22_X1 port map( A1 => n554, A2 => Q(855), B1 => n553, B2 => Q(727)
                           , ZN => n253);
   U269 : AOI22_X1 port map( A1 => n556, A2 => Q(791), B1 => n555, B2 => Q(887)
                           , ZN => n254);
   U270 : NAND4_X1 port map( A1 => n624, A2 => n625, A3 => n253, A4 => n254, ZN
                           => n255);
   U271 : OR4_X1 port map( A1 => n243, A2 => n248, A3 => n252, A4 => n255, ZN 
                           => Y(23));
   U272 : AOI22_X1 port map( A1 => n562, A2 => Q(502), B1 => n561, B2 => Q(566)
                           , ZN => n256);
   U273 : AOI22_X1 port map( A1 => n564, A2 => Q(662), B1 => n563, B2 => Q(470)
                           , ZN => n257);
   U274 : AOI22_X1 port map( A1 => n566, A2 => Q(374), B1 => n565, B2 => Q(310)
                           , ZN => n258);
   U275 : AOI22_X1 port map( A1 => n568, A2 => Q(406), B1 => n567, B2 => Q(278)
                           , ZN => n259);
   U276 : NAND4_X1 port map( A1 => n256, A2 => n257, A3 => n258, A4 => n259, ZN
                           => n260);
   U277 : AOI22_X1 port map( A1 => n570, A2 => Q(342), B1 => n569, B2 => Q(438)
                           , ZN => n261);
   U278 : AOI22_X1 port map( A1 => n572, A2 => Q(246), B1 => n571, B2 => Q(150)
                           , ZN => n262);
   U279 : AOI22_X1 port map( A1 => n574, A2 => Q(86), B1 => n573, B2 => Q(182),
                           ZN => n263);
   U280 : AOI22_X1 port map( A1 => n576, A2 => Q(214), B1 => n575, B2 => Q(54),
                           ZN => n264);
   U281 : NAND4_X1 port map( A1 => n261, A2 => n262, A3 => n263, A4 => n264, ZN
                           => n265);
   U282 : AOI22_X1 port map( A1 => n547, A2 => Q(1014), B1 => n546, B2 => 
                           Q(950), ZN => n266);
   U283 : AOI22_X1 port map( A1 => n549, A2 => Q(982), B1 => n548, B2 => Q(918)
                           , ZN => n267);
   U284 : AOI222_X1 port map( A1 => n551, A2 => Q(822), B1 => n552, B2 => 
                           Q(118), C1 => n550, C2 => Q(758), ZN => n268);
   U285 : NAND3_X1 port map( A1 => n266, A2 => n267, A3 => n268, ZN => n269);
   U286 : AOI22_X1 port map( A1 => n554, A2 => Q(854), B1 => n553, B2 => Q(726)
                           , ZN => n270);
   U287 : AOI22_X1 port map( A1 => n556, A2 => Q(790), B1 => n555, B2 => Q(886)
                           , ZN => n271);
   U288 : NAND4_X1 port map( A1 => n622, A2 => n623, A3 => n270, A4 => n271, ZN
                           => n272);
   U289 : OR4_X1 port map( A1 => n260, A2 => n265, A3 => n269, A4 => n272, ZN 
                           => Y(22));
   U290 : AOI22_X1 port map( A1 => n562, A2 => Q(501), B1 => n561, B2 => Q(565)
                           , ZN => n273);
   U291 : AOI22_X1 port map( A1 => n564, A2 => Q(661), B1 => n563, B2 => Q(469)
                           , ZN => n274);
   U292 : AOI22_X1 port map( A1 => n566, A2 => Q(373), B1 => n565, B2 => Q(309)
                           , ZN => n275);
   U293 : AOI22_X1 port map( A1 => n568, A2 => Q(405), B1 => n567, B2 => Q(277)
                           , ZN => n276);
   U294 : NAND4_X1 port map( A1 => n273, A2 => n274, A3 => n275, A4 => n276, ZN
                           => n277);
   U295 : AOI22_X1 port map( A1 => n570, A2 => Q(341), B1 => n569, B2 => Q(437)
                           , ZN => n278);
   U296 : AOI22_X1 port map( A1 => n572, A2 => Q(245), B1 => n571, B2 => Q(149)
                           , ZN => n279);
   U297 : AOI22_X1 port map( A1 => n574, A2 => Q(85), B1 => n573, B2 => Q(181),
                           ZN => n280);
   U298 : AOI22_X1 port map( A1 => n576, A2 => Q(213), B1 => n575, B2 => Q(53),
                           ZN => n281);
   U299 : NAND4_X1 port map( A1 => n278, A2 => n279, A3 => n280, A4 => n281, ZN
                           => n282);
   U300 : AOI22_X1 port map( A1 => n547, A2 => Q(1013), B1 => n546, B2 => 
                           Q(949), ZN => n283);
   U301 : AOI22_X1 port map( A1 => n549, A2 => Q(981), B1 => n548, B2 => Q(917)
                           , ZN => n284);
   U302 : AOI222_X1 port map( A1 => n551, A2 => Q(821), B1 => n552, B2 => 
                           Q(117), C1 => n550, C2 => Q(757), ZN => n285);
   U303 : NAND3_X1 port map( A1 => n283, A2 => n284, A3 => n285, ZN => n286);
   U304 : AOI22_X1 port map( A1 => n554, A2 => Q(853), B1 => n553, B2 => Q(725)
                           , ZN => n287);
   U305 : AOI22_X1 port map( A1 => n556, A2 => Q(789), B1 => n555, B2 => Q(885)
                           , ZN => n288);
   U306 : NAND4_X1 port map( A1 => n620, A2 => n621, A3 => n287, A4 => n288, ZN
                           => n289);
   U307 : OR4_X1 port map( A1 => n277, A2 => n282, A3 => n286, A4 => n289, ZN 
                           => Y(21));
   U308 : AOI22_X1 port map( A1 => n562, A2 => Q(500), B1 => n561, B2 => Q(564)
                           , ZN => n290);
   U309 : AOI22_X1 port map( A1 => n564, A2 => Q(660), B1 => n563, B2 => Q(468)
                           , ZN => n291);
   U310 : AOI22_X1 port map( A1 => n566, A2 => Q(372), B1 => n565, B2 => Q(308)
                           , ZN => n292);
   U311 : AOI22_X1 port map( A1 => n568, A2 => Q(404), B1 => n567, B2 => Q(276)
                           , ZN => n293);
   U312 : NAND4_X1 port map( A1 => n290, A2 => n291, A3 => n292, A4 => n293, ZN
                           => n294);
   U313 : AOI22_X1 port map( A1 => n570, A2 => Q(340), B1 => n569, B2 => Q(436)
                           , ZN => n295);
   U314 : AOI22_X1 port map( A1 => n572, A2 => Q(244), B1 => n571, B2 => Q(148)
                           , ZN => n296);
   U315 : AOI22_X1 port map( A1 => n574, A2 => Q(84), B1 => n573, B2 => Q(180),
                           ZN => n297);
   U316 : AOI22_X1 port map( A1 => n576, A2 => Q(212), B1 => n575, B2 => Q(52),
                           ZN => n298);
   U317 : NAND4_X1 port map( A1 => n295, A2 => n296, A3 => n297, A4 => n298, ZN
                           => n299);
   U318 : AOI22_X1 port map( A1 => n547, A2 => Q(1012), B1 => n546, B2 => 
                           Q(948), ZN => n300);
   U319 : AOI22_X1 port map( A1 => n549, A2 => Q(980), B1 => n548, B2 => Q(916)
                           , ZN => n301);
   U320 : AOI222_X1 port map( A1 => n551, A2 => Q(820), B1 => n552, B2 => 
                           Q(116), C1 => n550, C2 => Q(756), ZN => n302);
   U321 : NAND3_X1 port map( A1 => n300, A2 => n301, A3 => n302, ZN => n303);
   U322 : AOI22_X1 port map( A1 => n554, A2 => Q(852), B1 => n553, B2 => Q(724)
                           , ZN => n304);
   U323 : AOI22_X1 port map( A1 => n556, A2 => Q(788), B1 => n555, B2 => Q(884)
                           , ZN => n305);
   U324 : NAND4_X1 port map( A1 => n618, A2 => n619, A3 => n304, A4 => n305, ZN
                           => n306);
   U325 : OR4_X1 port map( A1 => n294, A2 => n299, A3 => n303, A4 => n306, ZN 
                           => Y(20));
   U326 : AOI22_X1 port map( A1 => n674, A2 => Q(491), B1 => n673, B2 => Q(555)
                           , ZN => n307);
   U327 : AOI22_X1 port map( A1 => n676, A2 => Q(651), B1 => n675, B2 => Q(459)
                           , ZN => n308);
   U328 : AOI22_X1 port map( A1 => n678, A2 => Q(363), B1 => n677, B2 => Q(299)
                           , ZN => n309);
   U329 : AOI22_X1 port map( A1 => n680, A2 => Q(395), B1 => n679, B2 => Q(267)
                           , ZN => n310);
   U330 : NAND4_X1 port map( A1 => n307, A2 => n308, A3 => n309, A4 => n310, ZN
                           => n311);
   U331 : AOI22_X1 port map( A1 => n682, A2 => Q(331), B1 => n681, B2 => Q(427)
                           , ZN => n312);
   U332 : AOI22_X1 port map( A1 => n684, A2 => Q(235), B1 => n683, B2 => Q(139)
                           , ZN => n313);
   U333 : AOI22_X1 port map( A1 => n686, A2 => Q(75), B1 => n685, B2 => Q(171),
                           ZN => n314);
   U334 : AOI22_X1 port map( A1 => n688, A2 => Q(203), B1 => n687, B2 => Q(43),
                           ZN => n315);
   U335 : NAND4_X1 port map( A1 => n312, A2 => n313, A3 => n314, A4 => n315, ZN
                           => n316);
   U336 : AOI22_X1 port map( A1 => n657, A2 => Q(1003), B1 => n656, B2 => 
                           Q(939), ZN => n317);
   U337 : AOI22_X1 port map( A1 => n659, A2 => Q(971), B1 => n658, B2 => Q(907)
                           , ZN => n318);
   U338 : AOI222_X1 port map( A1 => n661, A2 => Q(811), B1 => n662, B2 => 
                           Q(107), C1 => n660, C2 => Q(747), ZN => n319);
   U339 : NAND3_X1 port map( A1 => n317, A2 => n318, A3 => n319, ZN => n320);
   U340 : AOI22_X1 port map( A1 => n664, A2 => Q(843), B1 => n663, B2 => Q(715)
                           , ZN => n321);
   U341 : AOI22_X1 port map( A1 => n666, A2 => Q(779), B1 => n665, B2 => Q(875)
                           , ZN => n322);
   U342 : NAND4_X1 port map( A1 => n598, A2 => n599, A3 => n321, A4 => n322, ZN
                           => n323);
   U343 : OR4_X1 port map( A1 => n311, A2 => n316, A3 => n320, A4 => n323, ZN 
                           => Y(11));
   U344 : AOI22_X1 port map( A1 => n562, A2 => Q(490), B1 => n561, B2 => Q(554)
                           , ZN => n324);
   U345 : AOI22_X1 port map( A1 => n564, A2 => Q(650), B1 => n563, B2 => Q(458)
                           , ZN => n325);
   U346 : AOI22_X1 port map( A1 => n566, A2 => Q(362), B1 => n565, B2 => Q(298)
                           , ZN => n326);
   U347 : AOI22_X1 port map( A1 => n568, A2 => Q(394), B1 => n567, B2 => Q(266)
                           , ZN => n327);
   U348 : NAND4_X1 port map( A1 => n324, A2 => n325, A3 => n326, A4 => n327, ZN
                           => n328);
   U349 : AOI22_X1 port map( A1 => n570, A2 => Q(330), B1 => n569, B2 => Q(426)
                           , ZN => n329);
   U350 : AOI22_X1 port map( A1 => n572, A2 => Q(234), B1 => n571, B2 => Q(138)
                           , ZN => n330);
   U351 : AOI22_X1 port map( A1 => n574, A2 => Q(74), B1 => n573, B2 => Q(170),
                           ZN => n331);
   U352 : AOI22_X1 port map( A1 => n576, A2 => Q(202), B1 => n575, B2 => Q(42),
                           ZN => n332);
   U353 : NAND4_X1 port map( A1 => n329, A2 => n330, A3 => n331, A4 => n332, ZN
                           => n333);
   U354 : AOI22_X1 port map( A1 => n547, A2 => Q(1002), B1 => n546, B2 => 
                           Q(938), ZN => n334);
   U355 : AOI22_X1 port map( A1 => n549, A2 => Q(970), B1 => n548, B2 => Q(906)
                           , ZN => n335);
   U356 : AOI222_X1 port map( A1 => n551, A2 => Q(810), B1 => n552, B2 => 
                           Q(106), C1 => n550, C2 => Q(746), ZN => n336);
   U357 : NAND3_X1 port map( A1 => n334, A2 => n335, A3 => n336, ZN => n337);
   U358 : AOI22_X1 port map( A1 => n554, A2 => Q(842), B1 => n553, B2 => Q(714)
                           , ZN => n338);
   U359 : AOI22_X1 port map( A1 => n556, A2 => Q(778), B1 => n555, B2 => Q(874)
                           , ZN => n339);
   U360 : NAND4_X1 port map( A1 => n596, A2 => n597, A3 => n338, A4 => n339, ZN
                           => n340);
   U361 : OR4_X1 port map( A1 => n328, A2 => n333, A3 => n337, A4 => n340, ZN 
                           => Y(10));
   U362 : AOI22_X1 port map( A1 => n562, A2 => Q(489), B1 => n561, B2 => Q(553)
                           , ZN => n341);
   U363 : AOI22_X1 port map( A1 => n564, A2 => Q(649), B1 => n563, B2 => Q(457)
                           , ZN => n342);
   U364 : AOI22_X1 port map( A1 => n566, A2 => Q(361), B1 => n565, B2 => Q(297)
                           , ZN => n343);
   U365 : AOI22_X1 port map( A1 => n568, A2 => Q(393), B1 => n567, B2 => Q(265)
                           , ZN => n344);
   U366 : NAND4_X1 port map( A1 => n341, A2 => n342, A3 => n343, A4 => n344, ZN
                           => n345);
   U367 : AOI22_X1 port map( A1 => n570, A2 => Q(329), B1 => n569, B2 => Q(425)
                           , ZN => n346);
   U368 : AOI22_X1 port map( A1 => n572, A2 => Q(233), B1 => n571, B2 => Q(137)
                           , ZN => n347);
   U369 : AOI22_X1 port map( A1 => n574, A2 => Q(73), B1 => n573, B2 => Q(169),
                           ZN => n348);
   U370 : AOI22_X1 port map( A1 => n576, A2 => Q(201), B1 => n575, B2 => Q(41),
                           ZN => n349);
   U371 : NAND4_X1 port map( A1 => n346, A2 => n347, A3 => n348, A4 => n349, ZN
                           => n350);
   U372 : AOI22_X1 port map( A1 => n547, A2 => Q(1001), B1 => n546, B2 => 
                           Q(937), ZN => n351);
   U373 : AOI22_X1 port map( A1 => n549, A2 => Q(969), B1 => n548, B2 => Q(905)
                           , ZN => n352);
   U374 : AOI222_X1 port map( A1 => n551, A2 => Q(809), B1 => n552, B2 => 
                           Q(105), C1 => n550, C2 => Q(745), ZN => n353);
   U375 : NAND3_X1 port map( A1 => n351, A2 => n352, A3 => n353, ZN => n354);
   U376 : AOI22_X1 port map( A1 => n554, A2 => Q(841), B1 => n553, B2 => Q(713)
                           , ZN => n355);
   U377 : AOI22_X1 port map( A1 => n556, A2 => Q(777), B1 => n555, B2 => Q(873)
                           , ZN => n356);
   U378 : NAND4_X1 port map( A1 => n671, A2 => n672, A3 => n355, A4 => n356, ZN
                           => n357);
   U379 : OR4_X1 port map( A1 => n345, A2 => n350, A3 => n354, A4 => n357, ZN 
                           => Y(9));
   U380 : AOI22_X1 port map( A1 => n562, A2 => Q(488), B1 => n561, B2 => Q(552)
                           , ZN => n358);
   U381 : AOI22_X1 port map( A1 => n564, A2 => Q(648), B1 => n563, B2 => Q(456)
                           , ZN => n359);
   U382 : AOI22_X1 port map( A1 => n566, A2 => Q(360), B1 => n565, B2 => Q(296)
                           , ZN => n360);
   U383 : AOI22_X1 port map( A1 => n568, A2 => Q(392), B1 => n567, B2 => Q(264)
                           , ZN => n361);
   U384 : NAND4_X1 port map( A1 => n358, A2 => n359, A3 => n360, A4 => n361, ZN
                           => n362);
   U385 : AOI22_X1 port map( A1 => n570, A2 => Q(328), B1 => n569, B2 => Q(424)
                           , ZN => n363);
   U386 : AOI22_X1 port map( A1 => n572, A2 => Q(232), B1 => n571, B2 => Q(136)
                           , ZN => n364);
   U387 : AOI22_X1 port map( A1 => n574, A2 => Q(72), B1 => n573, B2 => Q(168),
                           ZN => n365);
   U388 : AOI22_X1 port map( A1 => n576, A2 => Q(200), B1 => n575, B2 => Q(40),
                           ZN => n366);
   U389 : NAND4_X1 port map( A1 => n363, A2 => n364, A3 => n365, A4 => n366, ZN
                           => n367);
   U390 : AOI22_X1 port map( A1 => n547, A2 => Q(1000), B1 => n546, B2 => 
                           Q(936), ZN => n368);
   U391 : AOI22_X1 port map( A1 => n549, A2 => Q(968), B1 => n548, B2 => Q(904)
                           , ZN => n369);
   U392 : AOI222_X1 port map( A1 => n551, A2 => Q(808), B1 => n552, B2 => 
                           Q(104), C1 => n550, C2 => Q(744), ZN => n370);
   U393 : NAND3_X1 port map( A1 => n368, A2 => n369, A3 => n370, ZN => n371);
   U394 : AOI22_X1 port map( A1 => n554, A2 => Q(840), B1 => n553, B2 => Q(712)
                           , ZN => n372);
   U395 : AOI22_X1 port map( A1 => n556, A2 => Q(776), B1 => n555, B2 => Q(872)
                           , ZN => n373);
   U396 : NAND4_X1 port map( A1 => n654, A2 => n655, A3 => n372, A4 => n373, ZN
                           => n374);
   U397 : OR4_X1 port map( A1 => n362, A2 => n367, A3 => n371, A4 => n374, ZN 
                           => Y(8));
   U398 : AOI22_X1 port map( A1 => n562, A2 => Q(487), B1 => n561, B2 => Q(551)
                           , ZN => n375);
   U399 : AOI22_X1 port map( A1 => n564, A2 => Q(647), B1 => n563, B2 => Q(455)
                           , ZN => n376);
   U400 : AOI22_X1 port map( A1 => n566, A2 => Q(359), B1 => n565, B2 => Q(295)
                           , ZN => n377);
   U401 : AOI22_X1 port map( A1 => n568, A2 => Q(391), B1 => n567, B2 => Q(263)
                           , ZN => n378);
   U402 : NAND4_X1 port map( A1 => n375, A2 => n376, A3 => n377, A4 => n378, ZN
                           => n379);
   U403 : AOI22_X1 port map( A1 => n570, A2 => Q(327), B1 => n569, B2 => Q(423)
                           , ZN => n380);
   U404 : AOI22_X1 port map( A1 => n572, A2 => Q(231), B1 => n571, B2 => Q(135)
                           , ZN => n381);
   U405 : AOI22_X1 port map( A1 => n574, A2 => Q(71), B1 => n573, B2 => Q(167),
                           ZN => n382);
   U406 : AOI22_X1 port map( A1 => n576, A2 => Q(199), B1 => n575, B2 => Q(39),
                           ZN => n383);
   U407 : NAND4_X1 port map( A1 => n380, A2 => n381, A3 => n382, A4 => n383, ZN
                           => n384);
   U408 : AOI22_X1 port map( A1 => n547, A2 => Q(999), B1 => n546, B2 => Q(935)
                           , ZN => n385);
   U409 : AOI22_X1 port map( A1 => n549, A2 => Q(967), B1 => n548, B2 => Q(903)
                           , ZN => n386);
   U410 : AOI222_X1 port map( A1 => n551, A2 => Q(807), B1 => n552, B2 => 
                           Q(103), C1 => n550, C2 => Q(743), ZN => n387);
   U411 : NAND3_X1 port map( A1 => n385, A2 => n386, A3 => n387, ZN => n388);
   U412 : AOI22_X1 port map( A1 => n554, A2 => Q(839), B1 => n553, B2 => Q(711)
                           , ZN => n389);
   U413 : AOI22_X1 port map( A1 => n556, A2 => Q(775), B1 => n555, B2 => Q(871)
                           , ZN => n390);
   U414 : NAND4_X1 port map( A1 => n652, A2 => n653, A3 => n389, A4 => n390, ZN
                           => n391);
   U415 : OR4_X1 port map( A1 => n379, A2 => n384, A3 => n388, A4 => n391, ZN 
                           => Y(7));
   U416 : AOI22_X1 port map( A1 => n562, A2 => Q(486), B1 => n561, B2 => Q(550)
                           , ZN => n392);
   U417 : AOI22_X1 port map( A1 => n564, A2 => Q(646), B1 => n563, B2 => Q(454)
                           , ZN => n393);
   U418 : AOI22_X1 port map( A1 => n566, A2 => Q(358), B1 => n565, B2 => Q(294)
                           , ZN => n394);
   U419 : AOI22_X1 port map( A1 => n568, A2 => Q(390), B1 => n567, B2 => Q(262)
                           , ZN => n395);
   U420 : NAND4_X1 port map( A1 => n392, A2 => n393, A3 => n394, A4 => n395, ZN
                           => n396);
   U421 : AOI22_X1 port map( A1 => n570, A2 => Q(326), B1 => n569, B2 => Q(422)
                           , ZN => n397);
   U422 : AOI22_X1 port map( A1 => n572, A2 => Q(230), B1 => n571, B2 => Q(134)
                           , ZN => n398);
   U423 : AOI22_X1 port map( A1 => n574, A2 => Q(70), B1 => n573, B2 => Q(166),
                           ZN => n399);
   U424 : AOI22_X1 port map( A1 => n576, A2 => Q(198), B1 => n575, B2 => Q(38),
                           ZN => n400);
   U425 : NAND4_X1 port map( A1 => n397, A2 => n398, A3 => n399, A4 => n400, ZN
                           => n401);
   U426 : AOI22_X1 port map( A1 => n547, A2 => Q(998), B1 => n546, B2 => Q(934)
                           , ZN => n402);
   U427 : AOI22_X1 port map( A1 => n549, A2 => Q(966), B1 => n548, B2 => Q(902)
                           , ZN => n403);
   U428 : AOI222_X1 port map( A1 => n551, A2 => Q(806), B1 => n552, B2 => 
                           Q(102), C1 => n550, C2 => Q(742), ZN => n404);
   U429 : NAND3_X1 port map( A1 => n402, A2 => n403, A3 => n404, ZN => n405);
   U430 : AOI22_X1 port map( A1 => n554, A2 => Q(838), B1 => n553, B2 => Q(710)
                           , ZN => n406);
   U431 : AOI22_X1 port map( A1 => n556, A2 => Q(774), B1 => n555, B2 => Q(870)
                           , ZN => n407);
   U432 : NAND4_X1 port map( A1 => n650, A2 => n651, A3 => n406, A4 => n407, ZN
                           => n408);
   U433 : OR4_X1 port map( A1 => n396, A2 => n401, A3 => n405, A4 => n408, ZN 
                           => Y(6));
   U434 : AOI22_X1 port map( A1 => n562, A2 => Q(485), B1 => n561, B2 => Q(549)
                           , ZN => n409);
   U435 : AOI22_X1 port map( A1 => n564, A2 => Q(645), B1 => n563, B2 => Q(453)
                           , ZN => n410);
   U436 : AOI22_X1 port map( A1 => n566, A2 => Q(357), B1 => n565, B2 => Q(293)
                           , ZN => n411);
   U437 : AOI22_X1 port map( A1 => n568, A2 => Q(389), B1 => n567, B2 => Q(261)
                           , ZN => n412);
   U438 : NAND4_X1 port map( A1 => n409, A2 => n410, A3 => n411, A4 => n412, ZN
                           => n413);
   U439 : AOI22_X1 port map( A1 => n570, A2 => Q(325), B1 => n569, B2 => Q(421)
                           , ZN => n414);
   U440 : AOI22_X1 port map( A1 => n572, A2 => Q(229), B1 => n571, B2 => Q(133)
                           , ZN => n415);
   U441 : AOI22_X1 port map( A1 => n574, A2 => Q(69), B1 => n573, B2 => Q(165),
                           ZN => n416);
   U442 : AOI22_X1 port map( A1 => n576, A2 => Q(197), B1 => n575, B2 => Q(37),
                           ZN => n417);
   U443 : NAND4_X1 port map( A1 => n414, A2 => n415, A3 => n416, A4 => n417, ZN
                           => n418);
   U444 : AOI22_X1 port map( A1 => n547, A2 => Q(997), B1 => n546, B2 => Q(933)
                           , ZN => n419);
   U445 : AOI22_X1 port map( A1 => n549, A2 => Q(965), B1 => n548, B2 => Q(901)
                           , ZN => n420);
   U446 : AOI222_X1 port map( A1 => n551, A2 => Q(805), B1 => n552, B2 => 
                           Q(101), C1 => n550, C2 => Q(741), ZN => n421);
   U447 : NAND3_X1 port map( A1 => n419, A2 => n420, A3 => n421, ZN => n422);
   U448 : AOI22_X1 port map( A1 => n554, A2 => Q(837), B1 => n553, B2 => Q(709)
                           , ZN => n423);
   U449 : AOI22_X1 port map( A1 => n556, A2 => Q(773), B1 => n555, B2 => Q(869)
                           , ZN => n424);
   U450 : NAND4_X1 port map( A1 => n648, A2 => n649, A3 => n423, A4 => n424, ZN
                           => n425);
   U451 : OR4_X1 port map( A1 => n413, A2 => n418, A3 => n422, A4 => n425, ZN 
                           => Y(5));
   U452 : AOI22_X1 port map( A1 => n562, A2 => Q(484), B1 => n561, B2 => Q(548)
                           , ZN => n426);
   U453 : AOI22_X1 port map( A1 => n564, A2 => Q(644), B1 => n563, B2 => Q(452)
                           , ZN => n427);
   U454 : AOI22_X1 port map( A1 => n566, A2 => Q(356), B1 => n565, B2 => Q(292)
                           , ZN => n428);
   U455 : AOI22_X1 port map( A1 => n568, A2 => Q(388), B1 => n567, B2 => Q(260)
                           , ZN => n429);
   U456 : NAND4_X1 port map( A1 => n426, A2 => n427, A3 => n428, A4 => n429, ZN
                           => n430);
   U457 : AOI22_X1 port map( A1 => n570, A2 => Q(324), B1 => n569, B2 => Q(420)
                           , ZN => n431);
   U458 : AOI22_X1 port map( A1 => n572, A2 => Q(228), B1 => n571, B2 => Q(132)
                           , ZN => n432);
   U459 : AOI22_X1 port map( A1 => n574, A2 => Q(68), B1 => n573, B2 => Q(164),
                           ZN => n433);
   U460 : AOI22_X1 port map( A1 => n576, A2 => Q(196), B1 => n575, B2 => Q(36),
                           ZN => n434);
   U461 : NAND4_X1 port map( A1 => n431, A2 => n432, A3 => n433, A4 => n434, ZN
                           => n435);
   U462 : AOI22_X1 port map( A1 => n547, A2 => Q(996), B1 => n546, B2 => Q(932)
                           , ZN => n436);
   U463 : AOI22_X1 port map( A1 => n549, A2 => Q(964), B1 => n548, B2 => Q(900)
                           , ZN => n437);
   U464 : AOI222_X1 port map( A1 => n551, A2 => Q(804), B1 => n552, B2 => 
                           Q(100), C1 => n550, C2 => Q(740), ZN => n438);
   U465 : NAND3_X1 port map( A1 => n436, A2 => n437, A3 => n438, ZN => n439);
   U466 : AOI22_X1 port map( A1 => n554, A2 => Q(836), B1 => n553, B2 => Q(708)
                           , ZN => n440);
   U467 : AOI22_X1 port map( A1 => n556, A2 => Q(772), B1 => n555, B2 => Q(868)
                           , ZN => n441);
   U468 : NAND4_X1 port map( A1 => n646, A2 => n647, A3 => n440, A4 => n441, ZN
                           => n442);
   U469 : OR4_X1 port map( A1 => n430, A2 => n435, A3 => n439, A4 => n442, ZN 
                           => Y(4));
   U470 : AOI22_X1 port map( A1 => n562, A2 => Q(483), B1 => n561, B2 => Q(547)
                           , ZN => n443);
   U471 : AOI22_X1 port map( A1 => n564, A2 => Q(643), B1 => n563, B2 => Q(451)
                           , ZN => n444);
   U472 : AOI22_X1 port map( A1 => n566, A2 => Q(355), B1 => n565, B2 => Q(291)
                           , ZN => n445);
   U473 : AOI22_X1 port map( A1 => n568, A2 => Q(387), B1 => n567, B2 => Q(259)
                           , ZN => n446);
   U474 : NAND4_X1 port map( A1 => n443, A2 => n444, A3 => n445, A4 => n446, ZN
                           => n447);
   U475 : AOI22_X1 port map( A1 => n570, A2 => Q(323), B1 => n569, B2 => Q(419)
                           , ZN => n448);
   U476 : AOI22_X1 port map( A1 => n572, A2 => Q(227), B1 => n571, B2 => Q(131)
                           , ZN => n449);
   U477 : AOI22_X1 port map( A1 => n574, A2 => Q(67), B1 => n573, B2 => Q(163),
                           ZN => n450);
   U478 : AOI22_X1 port map( A1 => n576, A2 => Q(195), B1 => n575, B2 => Q(35),
                           ZN => n451);
   U479 : NAND4_X1 port map( A1 => n448, A2 => n449, A3 => n450, A4 => n451, ZN
                           => n452);
   U480 : AOI22_X1 port map( A1 => n547, A2 => Q(995), B1 => n546, B2 => Q(931)
                           , ZN => n453);
   U481 : AOI22_X1 port map( A1 => n549, A2 => Q(963), B1 => n548, B2 => Q(899)
                           , ZN => n454);
   U482 : AOI222_X1 port map( A1 => n551, A2 => Q(803), B1 => n552, B2 => Q(99)
                           , C1 => n550, C2 => Q(739), ZN => n455);
   U483 : NAND3_X1 port map( A1 => n453, A2 => n454, A3 => n455, ZN => n456);
   U484 : AOI22_X1 port map( A1 => n554, A2 => Q(835), B1 => n553, B2 => Q(707)
                           , ZN => n457);
   U485 : AOI22_X1 port map( A1 => n556, A2 => Q(771), B1 => n555, B2 => Q(867)
                           , ZN => n458);
   U486 : NAND4_X1 port map( A1 => n644, A2 => n645, A3 => n457, A4 => n458, ZN
                           => n459);
   U487 : OR4_X1 port map( A1 => n447, A2 => n452, A3 => n456, A4 => n459, ZN 
                           => Y(3));
   U488 : AOI22_X1 port map( A1 => n562, A2 => Q(482), B1 => n561, B2 => Q(546)
                           , ZN => n460);
   U489 : AOI22_X1 port map( A1 => n564, A2 => Q(642), B1 => n563, B2 => Q(450)
                           , ZN => n461);
   U490 : AOI22_X1 port map( A1 => n566, A2 => Q(354), B1 => n565, B2 => Q(290)
                           , ZN => n462);
   U491 : AOI22_X1 port map( A1 => n568, A2 => Q(386), B1 => n567, B2 => Q(258)
                           , ZN => n463);
   U492 : NAND4_X1 port map( A1 => n460, A2 => n461, A3 => n462, A4 => n463, ZN
                           => n464);
   U493 : AOI22_X1 port map( A1 => n570, A2 => Q(322), B1 => n569, B2 => Q(418)
                           , ZN => n465);
   U494 : AOI22_X1 port map( A1 => n572, A2 => Q(226), B1 => n571, B2 => Q(130)
                           , ZN => n466);
   U495 : AOI22_X1 port map( A1 => n574, A2 => Q(66), B1 => n573, B2 => Q(162),
                           ZN => n467);
   U496 : AOI22_X1 port map( A1 => n576, A2 => Q(194), B1 => n575, B2 => Q(34),
                           ZN => n468);
   U497 : NAND4_X1 port map( A1 => n465, A2 => n466, A3 => n467, A4 => n468, ZN
                           => n469);
   U498 : AOI22_X1 port map( A1 => n547, A2 => Q(994), B1 => n546, B2 => Q(930)
                           , ZN => n470);
   U499 : AOI22_X1 port map( A1 => n549, A2 => Q(962), B1 => n548, B2 => Q(898)
                           , ZN => n471);
   U500 : AOI222_X1 port map( A1 => n551, A2 => Q(802), B1 => n552, B2 => Q(98)
                           , C1 => n550, C2 => Q(738), ZN => n472);
   U501 : NAND3_X1 port map( A1 => n470, A2 => n471, A3 => n472, ZN => n473);
   U502 : AOI22_X1 port map( A1 => n554, A2 => Q(834), B1 => n553, B2 => Q(706)
                           , ZN => n474);
   U503 : AOI22_X1 port map( A1 => n556, A2 => Q(770), B1 => n555, B2 => Q(866)
                           , ZN => n475);
   U504 : NAND4_X1 port map( A1 => n638, A2 => n639, A3 => n474, A4 => n475, ZN
                           => n476);
   U505 : OR4_X1 port map( A1 => n464, A2 => n469, A3 => n473, A4 => n476, ZN 
                           => Y(2));
   U506 : AOI22_X1 port map( A1 => n562, A2 => Q(481), B1 => n561, B2 => Q(545)
                           , ZN => n477);
   U507 : AOI22_X1 port map( A1 => n564, A2 => Q(641), B1 => n563, B2 => Q(449)
                           , ZN => n478);
   U508 : AOI22_X1 port map( A1 => n566, A2 => Q(353), B1 => n565, B2 => Q(289)
                           , ZN => n479);
   U509 : AOI22_X1 port map( A1 => n568, A2 => Q(385), B1 => n567, B2 => Q(257)
                           , ZN => n480);
   U510 : NAND4_X1 port map( A1 => n477, A2 => n478, A3 => n479, A4 => n480, ZN
                           => n481);
   U511 : AOI22_X1 port map( A1 => n570, A2 => Q(321), B1 => n569, B2 => Q(417)
                           , ZN => n482);
   U512 : AOI22_X1 port map( A1 => n572, A2 => Q(225), B1 => n571, B2 => Q(129)
                           , ZN => n483);
   U513 : AOI22_X1 port map( A1 => n574, A2 => Q(65), B1 => n573, B2 => Q(161),
                           ZN => n484);
   U514 : AOI22_X1 port map( A1 => n576, A2 => Q(193), B1 => n575, B2 => Q(33),
                           ZN => n485);
   U515 : NAND4_X1 port map( A1 => n482, A2 => n483, A3 => n484, A4 => n485, ZN
                           => n486);
   U516 : AOI22_X1 port map( A1 => n547, A2 => Q(993), B1 => n546, B2 => Q(929)
                           , ZN => n487);
   U517 : AOI22_X1 port map( A1 => n549, A2 => Q(961), B1 => n548, B2 => Q(897)
                           , ZN => n488);
   U518 : AOI222_X1 port map( A1 => n551, A2 => Q(801), B1 => n552, B2 => Q(97)
                           , C1 => n550, C2 => Q(737), ZN => n489);
   U519 : NAND3_X1 port map( A1 => n487, A2 => n488, A3 => n489, ZN => n490);
   U520 : AOI22_X1 port map( A1 => n554, A2 => Q(833), B1 => n553, B2 => Q(705)
                           , ZN => n491);
   U521 : AOI22_X1 port map( A1 => n556, A2 => Q(769), B1 => n555, B2 => Q(865)
                           , ZN => n492);
   U522 : NAND4_X1 port map( A1 => n616, A2 => n617, A3 => n491, A4 => n492, ZN
                           => n493);
   U523 : OR4_X1 port map( A1 => n481, A2 => n486, A3 => n490, A4 => n493, ZN 
                           => Y(1));
   U524 : AOI22_X1 port map( A1 => n562, A2 => Q(480), B1 => n561, B2 => Q(544)
                           , ZN => n494);
   U525 : AOI22_X1 port map( A1 => n564, A2 => Q(640), B1 => n563, B2 => Q(448)
                           , ZN => n495);
   U526 : AOI22_X1 port map( A1 => n566, A2 => Q(352), B1 => n565, B2 => Q(288)
                           , ZN => n496);
   U527 : AOI22_X1 port map( A1 => n568, A2 => Q(384), B1 => n567, B2 => Q(256)
                           , ZN => n497);
   U528 : NAND4_X1 port map( A1 => n494, A2 => n495, A3 => n496, A4 => n497, ZN
                           => n498);
   U529 : AOI22_X1 port map( A1 => n570, A2 => Q(320), B1 => n569, B2 => Q(416)
                           , ZN => n499);
   U530 : AOI22_X1 port map( A1 => n572, A2 => Q(224), B1 => n571, B2 => Q(128)
                           , ZN => n500);
   U531 : AOI22_X1 port map( A1 => n574, A2 => Q(64), B1 => n573, B2 => Q(160),
                           ZN => n501);
   U532 : AOI22_X1 port map( A1 => n576, A2 => Q(192), B1 => n575, B2 => Q(32),
                           ZN => n502);
   U533 : NAND4_X1 port map( A1 => n499, A2 => n500, A3 => n501, A4 => n502, ZN
                           => n503);
   U534 : AOI22_X1 port map( A1 => n547, A2 => Q(992), B1 => n546, B2 => Q(928)
                           , ZN => n504);
   U535 : AOI22_X1 port map( A1 => n549, A2 => Q(960), B1 => n548, B2 => Q(896)
                           , ZN => n505);
   U536 : AOI222_X1 port map( A1 => n551, A2 => Q(800), B1 => n552, B2 => Q(96)
                           , C1 => n550, C2 => Q(736), ZN => n506);
   U537 : NAND3_X1 port map( A1 => n504, A2 => n505, A3 => n506, ZN => n507);
   U538 : AOI22_X1 port map( A1 => n554, A2 => Q(832), B1 => n553, B2 => Q(704)
                           , ZN => n508);
   U539 : AOI22_X1 port map( A1 => n556, A2 => Q(768), B1 => n555, B2 => Q(864)
                           , ZN => n509);
   U540 : NAND4_X1 port map( A1 => n581, A2 => n582, A3 => n508, A4 => n509, ZN
                           => n510);
   U541 : OR4_X1 port map( A1 => n498, A2 => n503, A3 => n507, A4 => n510, ZN 
                           => Y(0));
   U542 : AOI22_X1 port map( A1 => n674, A2 => Q(492), B1 => n673, B2 => Q(556)
                           , ZN => n511);
   U543 : AOI22_X1 port map( A1 => n676, A2 => Q(652), B1 => n675, B2 => Q(460)
                           , ZN => n512);
   U544 : AOI22_X1 port map( A1 => n678, A2 => Q(364), B1 => n677, B2 => Q(300)
                           , ZN => n513);
   U545 : AOI22_X1 port map( A1 => n680, A2 => Q(396), B1 => n679, B2 => Q(268)
                           , ZN => n514);
   U546 : NAND4_X1 port map( A1 => n511, A2 => n512, A3 => n513, A4 => n514, ZN
                           => n515);
   U547 : AOI22_X1 port map( A1 => n682, A2 => Q(332), B1 => n681, B2 => Q(428)
                           , ZN => n516);
   U548 : AOI22_X1 port map( A1 => n684, A2 => Q(236), B1 => n683, B2 => Q(140)
                           , ZN => n517);
   U549 : AOI22_X1 port map( A1 => n686, A2 => Q(76), B1 => n685, B2 => Q(172),
                           ZN => n518);
   U550 : AOI22_X1 port map( A1 => n688, A2 => Q(204), B1 => n687, B2 => Q(44),
                           ZN => n519);
   U551 : NAND4_X1 port map( A1 => n516, A2 => n517, A3 => n518, A4 => n519, ZN
                           => n520);
   U552 : AOI22_X1 port map( A1 => n657, A2 => Q(1004), B1 => n656, B2 => 
                           Q(940), ZN => n521);
   U553 : AOI22_X1 port map( A1 => n659, A2 => Q(972), B1 => n658, B2 => Q(908)
                           , ZN => n522);
   U554 : AOI222_X1 port map( A1 => n661, A2 => Q(812), B1 => n662, B2 => 
                           Q(108), C1 => n660, C2 => Q(748), ZN => n523);
   U555 : NAND3_X1 port map( A1 => n521, A2 => n522, A3 => n523, ZN => n524);
   U556 : AOI22_X1 port map( A1 => n664, A2 => Q(844), B1 => n663, B2 => Q(716)
                           , ZN => n525);
   U557 : AOI22_X1 port map( A1 => n666, A2 => Q(780), B1 => n665, B2 => Q(876)
                           , ZN => n526);
   U558 : NAND4_X1 port map( A1 => n600, A2 => n601, A3 => n525, A4 => n526, ZN
                           => n527);
   U559 : OR4_X1 port map( A1 => n515, A2 => n520, A3 => n524, A4 => n527, ZN 
                           => Y(12));
   U560 : AOI22_X1 port map( A1 => n562, A2 => Q(511), B1 => n561, B2 => Q(575)
                           , ZN => n528);
   U561 : AOI22_X1 port map( A1 => n564, A2 => Q(671), B1 => n563, B2 => Q(479)
                           , ZN => n529);
   U562 : AOI22_X1 port map( A1 => n566, A2 => Q(383), B1 => n565, B2 => Q(319)
                           , ZN => n530);
   U563 : AOI22_X1 port map( A1 => n568, A2 => Q(415), B1 => n567, B2 => Q(287)
                           , ZN => n531);
   U564 : NAND4_X1 port map( A1 => n528, A2 => n529, A3 => n530, A4 => n531, ZN
                           => n532);
   U565 : AOI22_X1 port map( A1 => n570, A2 => Q(351), B1 => n569, B2 => Q(447)
                           , ZN => n533);
   U566 : AOI22_X1 port map( A1 => n572, A2 => Q(255), B1 => n571, B2 => Q(159)
                           , ZN => n534);
   U567 : AOI22_X1 port map( A1 => n574, A2 => Q(95), B1 => n573, B2 => Q(191),
                           ZN => n535);
   U568 : AOI22_X1 port map( A1 => n576, A2 => Q(223), B1 => n575, B2 => Q(63),
                           ZN => n536);
   U569 : NAND4_X1 port map( A1 => n533, A2 => n534, A3 => n535, A4 => n536, ZN
                           => n537);
   U570 : AOI22_X1 port map( A1 => n547, A2 => Q(1023), B1 => n546, B2 => 
                           Q(959), ZN => n538);
   U571 : AOI22_X1 port map( A1 => n549, A2 => Q(991), B1 => n548, B2 => Q(927)
                           , ZN => n539);
   U572 : AOI222_X1 port map( A1 => n551, A2 => Q(831), B1 => n552, B2 => 
                           Q(127), C1 => n550, C2 => Q(767), ZN => n540);
   U573 : NAND3_X1 port map( A1 => n538, A2 => n539, A3 => n540, ZN => n541);
   U574 : AOI22_X1 port map( A1 => n554, A2 => Q(863), B1 => n553, B2 => Q(735)
                           , ZN => n542);
   U575 : AOI22_X1 port map( A1 => n556, A2 => Q(799), B1 => n555, B2 => Q(895)
                           , ZN => n543);
   U576 : NAND4_X1 port map( A1 => n642, A2 => n643, A3 => n542, A4 => n543, ZN
                           => n544);
   U577 : OR4_X1 port map( A1 => n532, A2 => n537, A3 => n541, A4 => n544, ZN 
                           => Y(31));
   U578 : BUF_X1 port map( A => n687, Z => n575);
   U579 : BUF_X1 port map( A => n688, Z => n576);
   U580 : BUF_X1 port map( A => n685, Z => n573);
   U581 : BUF_X1 port map( A => n686, Z => n574);
   U582 : BUF_X1 port map( A => n683, Z => n571);
   U583 : BUF_X1 port map( A => n684, Z => n572);
   U584 : BUF_X1 port map( A => n681, Z => n569);
   U585 : BUF_X1 port map( A => n682, Z => n570);
   U586 : BUF_X1 port map( A => n679, Z => n567);
   U587 : BUF_X1 port map( A => n680, Z => n568);
   U588 : BUF_X1 port map( A => n677, Z => n565);
   U589 : BUF_X1 port map( A => n678, Z => n566);
   U590 : BUF_X1 port map( A => n675, Z => n563);
   U591 : BUF_X1 port map( A => n676, Z => n564);
   U592 : BUF_X1 port map( A => n673, Z => n561);
   U593 : BUF_X1 port map( A => n674, Z => n562);
   U594 : BUF_X1 port map( A => n669, Z => n559);
   U595 : BUF_X1 port map( A => n670, Z => n560);
   U596 : BUF_X1 port map( A => n667, Z => n557);
   U597 : BUF_X1 port map( A => n668, Z => n558);
   U598 : BUF_X1 port map( A => n665, Z => n555);
   U599 : BUF_X1 port map( A => n666, Z => n556);
   U600 : BUF_X1 port map( A => n663, Z => n553);
   U601 : BUF_X1 port map( A => n664, Z => n554);
   U602 : BUF_X1 port map( A => n662, Z => n552);
   U603 : BUF_X1 port map( A => n660, Z => n550);
   U604 : BUF_X1 port map( A => n661, Z => n551);
   U605 : BUF_X1 port map( A => n658, Z => n548);
   U606 : BUF_X1 port map( A => n659, Z => n549);
   U607 : BUF_X1 port map( A => n656, Z => n546);
   U608 : OR2_X1 port map( A1 => n577, A2 => S(1), ZN => n591);
   U609 : BUF_X1 port map( A => n657, Z => n547);
   U610 : NAND2_X1 port map( A1 => S(1), A2 => S(2), ZN => n593);
   U611 : NAND3_X1 port map( A1 => S(3), A2 => S(4), A3 => S(0), ZN => n580);
   U612 : NOR2_X1 port map( A1 => n593, A2 => n580, ZN => n657);
   U613 : INV_X1 port map( A => S(2), ZN => n577);
   U614 : NOR2_X1 port map( A1 => n580, A2 => n591, ZN => n656);
   U615 : INV_X1 port map( A => S(0), ZN => n578);
   U616 : NAND3_X1 port map( A1 => S(4), A2 => S(3), A3 => n578, ZN => n579);
   U617 : NOR2_X1 port map( A1 => n593, A2 => n579, ZN => n659);
   U618 : NOR2_X1 port map( A1 => n591, A2 => n579, ZN => n658);
   U619 : OR2_X1 port map( A1 => S(1), A2 => S(2), ZN => n594);
   U620 : NOR2_X1 port map( A1 => n580, A2 => n594, ZN => n661);
   U621 : INV_X1 port map( A => S(3), ZN => n588);
   U622 : NAND3_X1 port map( A1 => S(4), A2 => S(0), A3 => n588, ZN => n584);
   U623 : NOR2_X1 port map( A1 => n593, A2 => n584, ZN => n660);
   U624 : NAND2_X1 port map( A1 => S(1), A2 => n577, ZN => n590);
   U625 : INV_X1 port map( A => S(4), ZN => n583);
   U626 : NAND3_X1 port map( A1 => S(0), A2 => n588, A3 => n583, ZN => n595);
   U627 : NOR2_X1 port map( A1 => n590, A2 => n595, ZN => n662);
   U628 : NOR2_X1 port map( A1 => n590, A2 => n579, ZN => n664);
   U629 : NAND3_X1 port map( A1 => S(4), A2 => n588, A3 => n578, ZN => n585);
   U630 : NOR2_X1 port map( A1 => n593, A2 => n585, ZN => n663);
   U631 : NOR2_X1 port map( A1 => n579, A2 => n594, ZN => n666);
   U632 : NOR2_X1 port map( A1 => n590, A2 => n580, ZN => n665);
   U633 : NOR2_X1 port map( A1 => n591, A2 => n584, ZN => n668);
   U634 : NOR2_X1 port map( A1 => n590, A2 => n585, ZN => n667);
   U635 : AOI22_X1 port map( A1 => n558, A2 => Q(672), B1 => n557, B2 => Q(576)
                           , ZN => n582);
   U636 : NOR2_X1 port map( A1 => n594, A2 => n585, ZN => n670);
   U637 : NOR2_X1 port map( A1 => n590, A2 => n584, ZN => n669);
   U638 : AOI22_X1 port map( A1 => n560, A2 => Q(512), B1 => n559, B2 => Q(608)
                           , ZN => n581);
   U639 : NAND3_X1 port map( A1 => S(3), A2 => S(0), A3 => n583, ZN => n587);
   U640 : NOR2_X1 port map( A1 => n593, A2 => n587, ZN => n674);
   U641 : NOR2_X1 port map( A1 => n594, A2 => n584, ZN => n673);
   U642 : NOR2_X1 port map( A1 => n591, A2 => n585, ZN => n676);
   U643 : NOR2_X1 port map( A1 => S(4), A2 => S(0), ZN => n589);
   U644 : NAND2_X1 port map( A1 => S(3), A2 => n589, ZN => n586);
   U645 : NOR2_X1 port map( A1 => n593, A2 => n586, ZN => n675);
   U646 : NOR2_X1 port map( A1 => n590, A2 => n587, ZN => n678);
   U647 : NOR2_X1 port map( A1 => n594, A2 => n587, ZN => n677);
   U648 : NOR2_X1 port map( A1 => n591, A2 => n586, ZN => n680);
   U649 : NOR2_X1 port map( A1 => n594, A2 => n586, ZN => n679);
   U650 : NOR2_X1 port map( A1 => n590, A2 => n586, ZN => n682);
   U651 : NOR2_X1 port map( A1 => n591, A2 => n587, ZN => n681);
   U652 : NOR2_X1 port map( A1 => n595, A2 => n593, ZN => n684);
   U653 : NAND2_X1 port map( A1 => n589, A2 => n588, ZN => n592);
   U654 : NOR2_X1 port map( A1 => n591, A2 => n592, ZN => n683);
   U655 : NOR2_X1 port map( A1 => n590, A2 => n592, ZN => n686);
   U656 : NOR2_X1 port map( A1 => n595, A2 => n591, ZN => n685);
   U657 : NOR2_X1 port map( A1 => n593, A2 => n592, ZN => n688);
   U658 : NOR2_X1 port map( A1 => n595, A2 => n594, ZN => n687);
   U659 : AOI22_X1 port map( A1 => n558, A2 => Q(682), B1 => n557, B2 => Q(586)
                           , ZN => n597);
   U660 : AOI22_X1 port map( A1 => n560, A2 => Q(522), B1 => n559, B2 => Q(618)
                           , ZN => n596);
   U661 : AOI22_X1 port map( A1 => n668, A2 => Q(683), B1 => n667, B2 => Q(587)
                           , ZN => n599);
   U662 : AOI22_X1 port map( A1 => n670, A2 => Q(523), B1 => n669, B2 => Q(619)
                           , ZN => n598);
   U663 : AOI22_X1 port map( A1 => n668, A2 => Q(684), B1 => n667, B2 => Q(588)
                           , ZN => n601);
   U664 : AOI22_X1 port map( A1 => n670, A2 => Q(524), B1 => n669, B2 => Q(620)
                           , ZN => n600);
   U665 : AOI22_X1 port map( A1 => n668, A2 => Q(685), B1 => n667, B2 => Q(589)
                           , ZN => n603);
   U666 : AOI22_X1 port map( A1 => n670, A2 => Q(525), B1 => n669, B2 => Q(621)
                           , ZN => n602);
   U667 : AOI22_X1 port map( A1 => n668, A2 => Q(686), B1 => n667, B2 => Q(590)
                           , ZN => n605);
   U668 : AOI22_X1 port map( A1 => n670, A2 => Q(526), B1 => n669, B2 => Q(622)
                           , ZN => n604);
   U669 : AOI22_X1 port map( A1 => n668, A2 => Q(687), B1 => n667, B2 => Q(591)
                           , ZN => n607);
   U670 : AOI22_X1 port map( A1 => n670, A2 => Q(527), B1 => n669, B2 => Q(623)
                           , ZN => n606);
   U671 : AOI22_X1 port map( A1 => n668, A2 => Q(688), B1 => n667, B2 => Q(592)
                           , ZN => n609);
   U672 : AOI22_X1 port map( A1 => n670, A2 => Q(528), B1 => n669, B2 => Q(624)
                           , ZN => n608);
   U673 : AOI22_X1 port map( A1 => n668, A2 => Q(689), B1 => n667, B2 => Q(593)
                           , ZN => n611);
   U674 : AOI22_X1 port map( A1 => n670, A2 => Q(529), B1 => n669, B2 => Q(625)
                           , ZN => n610);
   U675 : AOI22_X1 port map( A1 => n668, A2 => Q(690), B1 => n667, B2 => Q(594)
                           , ZN => n613);
   U676 : AOI22_X1 port map( A1 => n670, A2 => Q(530), B1 => n669, B2 => Q(626)
                           , ZN => n612);
   U677 : AOI22_X1 port map( A1 => n668, A2 => Q(691), B1 => n667, B2 => Q(595)
                           , ZN => n615);
   U678 : AOI22_X1 port map( A1 => n670, A2 => Q(531), B1 => n669, B2 => Q(627)
                           , ZN => n614);
   U679 : AOI22_X1 port map( A1 => n558, A2 => Q(673), B1 => n557, B2 => Q(577)
                           , ZN => n617);
   U680 : AOI22_X1 port map( A1 => n560, A2 => Q(513), B1 => n559, B2 => Q(609)
                           , ZN => n616);
   U681 : AOI22_X1 port map( A1 => n558, A2 => Q(692), B1 => n557, B2 => Q(596)
                           , ZN => n619);
   U682 : AOI22_X1 port map( A1 => n560, A2 => Q(532), B1 => n559, B2 => Q(628)
                           , ZN => n618);
   U683 : AOI22_X1 port map( A1 => n558, A2 => Q(693), B1 => n557, B2 => Q(597)
                           , ZN => n621);
   U684 : AOI22_X1 port map( A1 => n560, A2 => Q(533), B1 => n559, B2 => Q(629)
                           , ZN => n620);
   U685 : AOI22_X1 port map( A1 => n558, A2 => Q(694), B1 => n557, B2 => Q(598)
                           , ZN => n623);
   U686 : AOI22_X1 port map( A1 => n560, A2 => Q(534), B1 => n559, B2 => Q(630)
                           , ZN => n622);
   U687 : AOI22_X1 port map( A1 => n558, A2 => Q(695), B1 => n557, B2 => Q(599)
                           , ZN => n625);
   U688 : AOI22_X1 port map( A1 => n560, A2 => Q(535), B1 => n559, B2 => Q(631)
                           , ZN => n624);
   U689 : AOI22_X1 port map( A1 => n558, A2 => Q(696), B1 => n557, B2 => Q(600)
                           , ZN => n627);
   U690 : AOI22_X1 port map( A1 => n560, A2 => Q(536), B1 => n559, B2 => Q(632)
                           , ZN => n626);
   U691 : AOI22_X1 port map( A1 => n558, A2 => Q(697), B1 => n557, B2 => Q(601)
                           , ZN => n629);
   U692 : AOI22_X1 port map( A1 => n560, A2 => Q(537), B1 => n559, B2 => Q(633)
                           , ZN => n628);
   U693 : AOI22_X1 port map( A1 => n558, A2 => Q(698), B1 => n557, B2 => Q(602)
                           , ZN => n631);
   U694 : AOI22_X1 port map( A1 => n560, A2 => Q(538), B1 => n559, B2 => Q(634)
                           , ZN => n630);
   U695 : AOI22_X1 port map( A1 => n558, A2 => Q(699), B1 => n557, B2 => Q(603)
                           , ZN => n633);
   U696 : AOI22_X1 port map( A1 => n560, A2 => Q(539), B1 => n559, B2 => Q(635)
                           , ZN => n632);
   U697 : AOI22_X1 port map( A1 => n558, A2 => Q(700), B1 => n557, B2 => Q(604)
                           , ZN => n635);
   U698 : AOI22_X1 port map( A1 => n560, A2 => Q(540), B1 => n559, B2 => Q(636)
                           , ZN => n634);
   U699 : AOI22_X1 port map( A1 => n668, A2 => Q(701), B1 => n667, B2 => Q(605)
                           , ZN => n637);
   U700 : AOI22_X1 port map( A1 => n670, A2 => Q(541), B1 => n669, B2 => Q(637)
                           , ZN => n636);
   U701 : AOI22_X1 port map( A1 => n558, A2 => Q(674), B1 => n557, B2 => Q(578)
                           , ZN => n639);
   U702 : AOI22_X1 port map( A1 => n560, A2 => Q(514), B1 => n559, B2 => Q(610)
                           , ZN => n638);
   U703 : AOI22_X1 port map( A1 => n558, A2 => Q(702), B1 => n557, B2 => Q(606)
                           , ZN => n641);
   U704 : AOI22_X1 port map( A1 => n560, A2 => Q(542), B1 => n559, B2 => Q(638)
                           , ZN => n640);
   U705 : AOI22_X1 port map( A1 => n558, A2 => Q(703), B1 => n557, B2 => Q(607)
                           , ZN => n643);
   U706 : AOI22_X1 port map( A1 => n560, A2 => Q(543), B1 => n559, B2 => Q(639)
                           , ZN => n642);
   U707 : AOI22_X1 port map( A1 => n558, A2 => Q(675), B1 => n557, B2 => Q(579)
                           , ZN => n645);
   U708 : AOI22_X1 port map( A1 => n560, A2 => Q(515), B1 => n559, B2 => Q(611)
                           , ZN => n644);
   U709 : AOI22_X1 port map( A1 => n558, A2 => Q(676), B1 => n557, B2 => Q(580)
                           , ZN => n647);
   U710 : AOI22_X1 port map( A1 => n560, A2 => Q(516), B1 => n559, B2 => Q(612)
                           , ZN => n646);
   U711 : AOI22_X1 port map( A1 => n558, A2 => Q(677), B1 => n557, B2 => Q(581)
                           , ZN => n649);
   U712 : AOI22_X1 port map( A1 => n560, A2 => Q(517), B1 => n559, B2 => Q(613)
                           , ZN => n648);
   U713 : AOI22_X1 port map( A1 => n558, A2 => Q(678), B1 => n557, B2 => Q(582)
                           , ZN => n651);
   U714 : AOI22_X1 port map( A1 => n560, A2 => Q(518), B1 => n559, B2 => Q(614)
                           , ZN => n650);
   U715 : AOI22_X1 port map( A1 => n558, A2 => Q(679), B1 => n557, B2 => Q(583)
                           , ZN => n653);
   U716 : AOI22_X1 port map( A1 => n560, A2 => Q(519), B1 => n559, B2 => Q(615)
                           , ZN => n652);
   U717 : AOI22_X1 port map( A1 => n558, A2 => Q(680), B1 => n557, B2 => Q(584)
                           , ZN => n655);
   U718 : AOI22_X1 port map( A1 => n560, A2 => Q(520), B1 => n559, B2 => Q(616)
                           , ZN => n654);
   U719 : AOI22_X1 port map( A1 => n558, A2 => Q(681), B1 => n557, B2 => Q(585)
                           , ZN => n672);
   U720 : AOI22_X1 port map( A1 => n560, A2 => Q(521), B1 => n559, B2 => Q(617)
                           , ZN => n671);

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32.all;

entity in_loc_selblock_NBIT_DATA32_N8_F5 is

   port( regs : in std_logic_vector (2559 downto 0);  win : in std_logic_vector
         (4 downto 0);  curr_proc_regs : out std_logic_vector (511 downto 0));

end in_loc_selblock_NBIT_DATA32_N8_F5;

architecture SYN_behav of in_loc_selblock_NBIT_DATA32_N8_F5 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X32
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, 
      n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, 
      n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, 
      n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, 
      n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, 
      n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, 
      n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, 
      n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, 
      n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, 
      n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, 
      n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, 
      n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, 
      n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, 
      n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, 
      n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, 
      n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, 
      n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, 
      n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, 
      n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, 
      n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, 
      n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, 
      n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, 
      n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, 
      n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, 
      n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, 
      n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, 
      n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, 
      n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, 
      n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, 
      n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, 
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, 
      n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, 
      n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, 
      n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, 
      n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, 
      n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, 
      n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, 
      n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, 
      n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, 
      n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, 
      n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, 
      n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, 
      n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, 
      n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, 
      n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, 
      n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, 
      n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, 
      n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, 
      n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, 
      n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, 
      n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, 
      n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, 
      n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, 
      n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, 
      n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, 
      n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, 
      n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, 
      n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, 
      n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, 
      n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, 
      n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, 
      n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, 
      n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, 
      n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591 : std_logic
      ;

begin
   
   U2 : CLKBUF_X3 port map( A => n20, Z => n7);
   U3 : BUF_X2 port map( A => n21, Z => n1);
   U4 : BUF_X2 port map( A => n6, Z => n2);
   U5 : BUF_X4 port map( A => n28, Z => n31);
   U6 : BUF_X4 port map( A => n37, Z => n36);
   U7 : CLKBUF_X2 port map( A => n39, Z => n9);
   U8 : BUF_X2 port map( A => n1588, Z => n39);
   U9 : CLKBUF_X3 port map( A => n1588, Z => n35);
   U10 : BUF_X4 port map( A => n1586, Z => n3);
   U11 : BUF_X4 port map( A => n38, Z => n4);
   U12 : NOR3_X2 port map( A1 => win(3), A2 => n12, A3 => n50, ZN => n1587);
   U13 : BUF_X2 port map( A => n40, Z => n5);
   U14 : BUF_X2 port map( A => n2, Z => n22);
   U15 : BUF_X2 port map( A => n2, Z => n18);
   U16 : BUF_X2 port map( A => n17, Z => n6);
   U17 : BUF_X2 port map( A => n3, Z => n30);
   U18 : BUF_X2 port map( A => n1585, Z => n19);
   U19 : BUF_X4 port map( A => n29, Z => n8);
   U20 : AND3_X2 port map( A1 => n49, A2 => win(0), A3 => n48, ZN => n1586);
   U21 : AND2_X2 port map( A1 => n49, A2 => win(1), ZN => n1585);
   U22 : BUF_X2 port map( A => n46, Z => n10);
   U23 : BUF_X2 port map( A => n44, Z => n11);
   U24 : BUF_X2 port map( A => n43, Z => n12);
   U25 : BUF_X2 port map( A => n5, Z => n13);
   U26 : BUF_X2 port map( A => n5, Z => n14);
   U27 : BUF_X2 port map( A => n45, Z => n15);
   U28 : BUF_X2 port map( A => n47, Z => n16);
   U29 : BUF_X2 port map( A => win(4), Z => n40);
   U30 : BUF_X32 port map( A => n1587, Z => n32);
   U31 : BUF_X1 port map( A => n40, Z => n41);
   U32 : BUF_X1 port map( A => n40, Z => n42);
   U33 : BUF_X1 port map( A => n8, Z => n26);
   U34 : BUF_X1 port map( A => n1588, Z => n33);
   U35 : BUF_X1 port map( A => n40, Z => n45);
   U36 : BUF_X1 port map( A => n18, Z => n24);
   U37 : BUF_X1 port map( A => n40, Z => n44);
   U38 : BUF_X1 port map( A => n30, Z => n25);
   U39 : BUF_X1 port map( A => n20, Z => n21);
   U40 : BUF_X1 port map( A => n40, Z => n47);
   U41 : BUF_X1 port map( A => n22, Z => n23);
   U42 : BUF_X1 port map( A => n7, Z => n17);
   U43 : BUF_X1 port map( A => n1585, Z => n20);
   U44 : BUF_X1 port map( A => n31, Z => n27);
   U45 : BUF_X1 port map( A => n1586, Z => n29);
   U46 : BUF_X1 port map( A => n1588, Z => n38);
   U47 : BUF_X1 port map( A => n40, Z => n46);
   U48 : NOR2_X1 port map( A1 => n14, A2 => n51, ZN => n1588);
   U49 : BUF_X1 port map( A => n40, Z => n43);
   U50 : BUF_X2 port map( A => n33, Z => n37);
   U51 : BUF_X2 port map( A => n1588, Z => n34);
   U52 : BUF_X2 port map( A => n29, Z => n28);
   U53 : NOR3_X1 port map( A1 => win(2), A2 => win(3), A3 => n12, ZN => n49);
   U54 : INV_X1 port map( A => win(1), ZN => n48);
   U55 : NAND2_X1 port map( A1 => regs(0), A2 => n1586, ZN => n54);
   U56 : INV_X1 port map( A => win(2), ZN => n50);
   U57 : AOI22_X1 port map( A1 => n7, A2 => regs(512), B1 => n32, B2 => 
                           regs(1024), ZN => n53);
   U58 : INV_X1 port map( A => win(3), ZN => n51);
   U59 : AOI22_X1 port map( A1 => n40, A2 => regs(2048), B1 => n34, B2 => 
                           regs(1536), ZN => n52);
   U60 : NAND3_X1 port map( A1 => n54, A2 => n53, A3 => n52, ZN => 
                           curr_proc_regs(0));
   U61 : NAND2_X1 port map( A1 => regs(612), A2 => n7, ZN => n57);
   U62 : AOI22_X1 port map( A1 => n32, A2 => regs(1124), B1 => n25, B2 => 
                           regs(100), ZN => n56);
   U63 : AOI22_X1 port map( A1 => n40, A2 => regs(2148), B1 => n4, B2 => 
                           regs(1636), ZN => n55);
   U64 : NAND3_X1 port map( A1 => n57, A2 => n56, A3 => n55, ZN => 
                           curr_proc_regs(100));
   U65 : NAND2_X1 port map( A1 => regs(613), A2 => n7, ZN => n60);
   U66 : AOI22_X1 port map( A1 => n32, A2 => regs(1125), B1 => n25, B2 => 
                           regs(101), ZN => n59);
   U67 : AOI22_X1 port map( A1 => n40, A2 => regs(2149), B1 => n36, B2 => 
                           regs(1637), ZN => n58);
   U68 : NAND3_X1 port map( A1 => n60, A2 => n59, A3 => n58, ZN => 
                           curr_proc_regs(101));
   U69 : NAND2_X1 port map( A1 => regs(614), A2 => n7, ZN => n63);
   U70 : AOI22_X1 port map( A1 => n32, A2 => regs(1126), B1 => n26, B2 => 
                           regs(102), ZN => n62);
   U71 : AOI22_X1 port map( A1 => n42, A2 => regs(2150), B1 => n9, B2 => 
                           regs(1638), ZN => n61);
   U72 : NAND3_X1 port map( A1 => n63, A2 => n62, A3 => n61, ZN => 
                           curr_proc_regs(102));
   U73 : NAND2_X1 port map( A1 => regs(615), A2 => n21, ZN => n66);
   U74 : AOI22_X1 port map( A1 => n32, A2 => regs(1127), B1 => n1586, B2 => 
                           regs(103), ZN => n65);
   U75 : AOI22_X1 port map( A1 => n41, A2 => regs(2151), B1 => n35, B2 => 
                           regs(1639), ZN => n64);
   U76 : NAND3_X1 port map( A1 => n66, A2 => n65, A3 => n64, ZN => 
                           curr_proc_regs(103));
   U77 : NAND2_X1 port map( A1 => regs(616), A2 => n7, ZN => n69);
   U78 : AOI22_X1 port map( A1 => n32, A2 => regs(1128), B1 => n1586, B2 => 
                           regs(104), ZN => n68);
   U79 : AOI22_X1 port map( A1 => n40, A2 => regs(2152), B1 => n9, B2 => 
                           regs(1640), ZN => n67);
   U80 : NAND3_X1 port map( A1 => n69, A2 => n68, A3 => n67, ZN => 
                           curr_proc_regs(104));
   U81 : NAND2_X1 port map( A1 => regs(617), A2 => n23, ZN => n72);
   U82 : AOI22_X1 port map( A1 => n32, A2 => regs(1129), B1 => n26, B2 => 
                           regs(105), ZN => n71);
   U83 : AOI22_X1 port map( A1 => n40, A2 => regs(2153), B1 => n4, B2 => 
                           regs(1641), ZN => n70);
   U84 : NAND3_X1 port map( A1 => n72, A2 => n71, A3 => n70, ZN => 
                           curr_proc_regs(105));
   U85 : NAND2_X1 port map( A1 => regs(618), A2 => n7, ZN => n75);
   U86 : AOI22_X1 port map( A1 => n32, A2 => regs(1130), B1 => n25, B2 => 
                           regs(106), ZN => n74);
   U87 : AOI22_X1 port map( A1 => n41, A2 => regs(2154), B1 => n9, B2 => 
                           regs(1642), ZN => n73);
   U88 : NAND3_X1 port map( A1 => n75, A2 => n74, A3 => n73, ZN => 
                           curr_proc_regs(106));
   U89 : NAND2_X1 port map( A1 => regs(619), A2 => n19, ZN => n78);
   U90 : AOI22_X1 port map( A1 => n32, A2 => regs(1131), B1 => n26, B2 => 
                           regs(107), ZN => n77);
   U91 : AOI22_X1 port map( A1 => n42, A2 => regs(2155), B1 => n36, B2 => 
                           regs(1643), ZN => n76);
   U92 : NAND3_X1 port map( A1 => n78, A2 => n77, A3 => n76, ZN => 
                           curr_proc_regs(107));
   U93 : NAND2_X1 port map( A1 => regs(620), A2 => n7, ZN => n81);
   U94 : AOI22_X1 port map( A1 => n32, A2 => regs(1132), B1 => n1586, B2 => 
                           regs(108), ZN => n80);
   U95 : AOI22_X1 port map( A1 => n42, A2 => regs(2156), B1 => n1588, B2 => 
                           regs(1644), ZN => n79);
   U96 : NAND3_X1 port map( A1 => n81, A2 => n80, A3 => n79, ZN => 
                           curr_proc_regs(108));
   U97 : NAND2_X1 port map( A1 => regs(621), A2 => n1585, ZN => n84);
   U98 : AOI22_X1 port map( A1 => n32, A2 => regs(1133), B1 => n28, B2 => 
                           regs(109), ZN => n83);
   U99 : AOI22_X1 port map( A1 => n41, A2 => regs(2157), B1 => n36, B2 => 
                           regs(1645), ZN => n82);
   U100 : NAND3_X1 port map( A1 => n84, A2 => n83, A3 => n82, ZN => 
                           curr_proc_regs(109));
   U101 : NAND2_X1 port map( A1 => regs(522), A2 => n6, ZN => n87);
   U102 : AOI22_X1 port map( A1 => n32, A2 => regs(1034), B1 => n8, B2 => 
                           regs(10), ZN => n86);
   U103 : AOI22_X1 port map( A1 => n42, A2 => regs(2058), B1 => n34, B2 => 
                           regs(1546), ZN => n85);
   U104 : NAND3_X1 port map( A1 => n87, A2 => n86, A3 => n85, ZN => 
                           curr_proc_regs(10));
   U105 : NAND2_X1 port map( A1 => regs(622), A2 => n22, ZN => n90);
   U106 : AOI22_X1 port map( A1 => n32, A2 => regs(1134), B1 => n28, B2 => 
                           regs(110), ZN => n89);
   U107 : AOI22_X1 port map( A1 => n40, A2 => regs(2158), B1 => n34, B2 => 
                           regs(1646), ZN => n88);
   U108 : NAND3_X1 port map( A1 => n90, A2 => n89, A3 => n88, ZN => 
                           curr_proc_regs(110));
   U109 : NAND2_X1 port map( A1 => regs(623), A2 => n1585, ZN => n93);
   U110 : AOI22_X1 port map( A1 => n32, A2 => regs(1135), B1 => n8, B2 => 
                           regs(111), ZN => n92);
   U111 : AOI22_X1 port map( A1 => n40, A2 => regs(2159), B1 => n34, B2 => 
                           regs(1647), ZN => n91);
   U112 : NAND3_X1 port map( A1 => n93, A2 => n92, A3 => n91, ZN => 
                           curr_proc_regs(111));
   U113 : NAND2_X1 port map( A1 => regs(624), A2 => n19, ZN => n96);
   U114 : AOI22_X1 port map( A1 => n32, A2 => regs(1136), B1 => n8, B2 => 
                           regs(112), ZN => n95);
   U115 : AOI22_X1 port map( A1 => n41, A2 => regs(2160), B1 => n34, B2 => 
                           regs(1648), ZN => n94);
   U116 : NAND3_X1 port map( A1 => n96, A2 => n95, A3 => n94, ZN => 
                           curr_proc_regs(112));
   U117 : NAND2_X1 port map( A1 => regs(625), A2 => n6, ZN => n99);
   U118 : AOI22_X1 port map( A1 => n32, A2 => regs(1137), B1 => n31, B2 => 
                           regs(113), ZN => n98);
   U119 : AOI22_X1 port map( A1 => n42, A2 => regs(2161), B1 => n34, B2 => 
                           regs(1649), ZN => n97);
   U120 : NAND3_X1 port map( A1 => n99, A2 => n98, A3 => n97, ZN => 
                           curr_proc_regs(113));
   U121 : NAND2_X1 port map( A1 => regs(626), A2 => n2, ZN => n102);
   U122 : AOI22_X1 port map( A1 => n32, A2 => regs(1138), B1 => n3, B2 => 
                           regs(114), ZN => n101);
   U123 : AOI22_X1 port map( A1 => n41, A2 => regs(2162), B1 => n34, B2 => 
                           regs(1650), ZN => n100);
   U124 : NAND3_X1 port map( A1 => n102, A2 => n101, A3 => n100, ZN => 
                           curr_proc_regs(114));
   U125 : NAND2_X1 port map( A1 => regs(627), A2 => n22, ZN => n105);
   U126 : AOI22_X1 port map( A1 => n32, A2 => regs(1139), B1 => n28, B2 => 
                           regs(115), ZN => n104);
   U127 : AOI22_X1 port map( A1 => n40, A2 => regs(2163), B1 => n34, B2 => 
                           regs(1651), ZN => n103);
   U128 : NAND3_X1 port map( A1 => n105, A2 => n104, A3 => n103, ZN => 
                           curr_proc_regs(115));
   U129 : NAND2_X1 port map( A1 => regs(628), A2 => n1585, ZN => n108);
   U130 : AOI22_X1 port map( A1 => n32, A2 => regs(1140), B1 => n1586, B2 => 
                           regs(116), ZN => n107);
   U131 : AOI22_X1 port map( A1 => n41, A2 => regs(2164), B1 => n34, B2 => 
                           regs(1652), ZN => n106);
   U132 : NAND3_X1 port map( A1 => n108, A2 => n107, A3 => n106, ZN => 
                           curr_proc_regs(116));
   U133 : NAND2_X1 port map( A1 => regs(629), A2 => n19, ZN => n111);
   U134 : AOI22_X1 port map( A1 => n32, A2 => regs(1141), B1 => n8, B2 => 
                           regs(117), ZN => n110);
   U135 : AOI22_X1 port map( A1 => n42, A2 => regs(2165), B1 => n34, B2 => 
                           regs(1653), ZN => n109);
   U136 : NAND3_X1 port map( A1 => n111, A2 => n110, A3 => n109, ZN => 
                           curr_proc_regs(117));
   U137 : NAND2_X1 port map( A1 => regs(630), A2 => n6, ZN => n114);
   U138 : AOI22_X1 port map( A1 => n32, A2 => regs(1142), B1 => n26, B2 => 
                           regs(118), ZN => n113);
   U139 : AOI22_X1 port map( A1 => n42, A2 => regs(2166), B1 => n34, B2 => 
                           regs(1654), ZN => n112);
   U140 : NAND3_X1 port map( A1 => n114, A2 => n113, A3 => n112, ZN => 
                           curr_proc_regs(118));
   U141 : NAND2_X1 port map( A1 => regs(631), A2 => n2, ZN => n117);
   U142 : AOI22_X1 port map( A1 => n32, A2 => regs(1143), B1 => n3, B2 => 
                           regs(119), ZN => n116);
   U143 : AOI22_X1 port map( A1 => n40, A2 => regs(2167), B1 => n34, B2 => 
                           regs(1655), ZN => n115);
   U144 : NAND3_X1 port map( A1 => n117, A2 => n116, A3 => n115, ZN => 
                           curr_proc_regs(119));
   U145 : NAND2_X1 port map( A1 => regs(523), A2 => n17, ZN => n120);
   U146 : AOI22_X1 port map( A1 => n32, A2 => regs(1035), B1 => n26, B2 => 
                           regs(11), ZN => n119);
   U147 : AOI22_X1 port map( A1 => n40, A2 => regs(2059), B1 => n9, B2 => 
                           regs(1547), ZN => n118);
   U148 : NAND3_X1 port map( A1 => n120, A2 => n119, A3 => n118, ZN => 
                           curr_proc_regs(11));
   U149 : NAND2_X1 port map( A1 => regs(632), A2 => n17, ZN => n123);
   U150 : AOI22_X1 port map( A1 => n32, A2 => regs(1144), B1 => n1586, B2 => 
                           regs(120), ZN => n122);
   U151 : AOI22_X1 port map( A1 => n41, A2 => regs(2168), B1 => n1588, B2 => 
                           regs(1656), ZN => n121);
   U152 : NAND3_X1 port map( A1 => n123, A2 => n122, A3 => n121, ZN => 
                           curr_proc_regs(120));
   U153 : NAND2_X1 port map( A1 => regs(633), A2 => n17, ZN => n126);
   U154 : AOI22_X1 port map( A1 => n32, A2 => regs(1145), B1 => n8, B2 => 
                           regs(121), ZN => n125);
   U155 : AOI22_X1 port map( A1 => n42, A2 => regs(2169), B1 => n4, B2 => 
                           regs(1657), ZN => n124);
   U156 : NAND3_X1 port map( A1 => n126, A2 => n125, A3 => n124, ZN => 
                           curr_proc_regs(121));
   U157 : NAND2_X1 port map( A1 => regs(634), A2 => n17, ZN => n129);
   U158 : AOI22_X1 port map( A1 => n32, A2 => regs(1146), B1 => n25, B2 => 
                           regs(122), ZN => n128);
   U159 : AOI22_X1 port map( A1 => n40, A2 => regs(2170), B1 => n9, B2 => 
                           regs(1658), ZN => n127);
   U160 : NAND3_X1 port map( A1 => n129, A2 => n128, A3 => n127, ZN => 
                           curr_proc_regs(122));
   U161 : NAND2_X1 port map( A1 => regs(635), A2 => n17, ZN => n132);
   U162 : AOI22_X1 port map( A1 => n32, A2 => regs(1147), B1 => n26, B2 => 
                           regs(123), ZN => n131);
   U163 : AOI22_X1 port map( A1 => n41, A2 => regs(2171), B1 => n34, B2 => 
                           regs(1659), ZN => n130);
   U164 : NAND3_X1 port map( A1 => n132, A2 => n131, A3 => n130, ZN => 
                           curr_proc_regs(123));
   U165 : NAND2_X1 port map( A1 => regs(636), A2 => n17, ZN => n135);
   U166 : AOI22_X1 port map( A1 => n32, A2 => regs(1148), B1 => n1586, B2 => 
                           regs(124), ZN => n134);
   U167 : AOI22_X1 port map( A1 => n42, A2 => regs(2172), B1 => n36, B2 => 
                           regs(1660), ZN => n133);
   U168 : NAND3_X1 port map( A1 => n135, A2 => n134, A3 => n133, ZN => 
                           curr_proc_regs(124));
   U169 : NAND2_X1 port map( A1 => regs(637), A2 => n17, ZN => n138);
   U170 : AOI22_X1 port map( A1 => n32, A2 => regs(1149), B1 => n3, B2 => 
                           regs(125), ZN => n137);
   U171 : AOI22_X1 port map( A1 => n40, A2 => regs(2173), B1 => n9, B2 => 
                           regs(1661), ZN => n136);
   U172 : NAND3_X1 port map( A1 => n138, A2 => n137, A3 => n136, ZN => 
                           curr_proc_regs(125));
   U173 : NAND2_X1 port map( A1 => regs(638), A2 => n17, ZN => n141);
   U174 : AOI22_X1 port map( A1 => n32, A2 => regs(1150), B1 => n25, B2 => 
                           regs(126), ZN => n140);
   U175 : AOI22_X1 port map( A1 => n41, A2 => regs(2174), B1 => n35, B2 => 
                           regs(1662), ZN => n139);
   U176 : NAND3_X1 port map( A1 => n141, A2 => n140, A3 => n139, ZN => 
                           curr_proc_regs(126));
   U177 : NAND2_X1 port map( A1 => regs(639), A2 => n17, ZN => n144);
   U178 : AOI22_X1 port map( A1 => n32, A2 => regs(1151), B1 => n26, B2 => 
                           regs(127), ZN => n143);
   U179 : AOI22_X1 port map( A1 => n42, A2 => regs(2175), B1 => n4, B2 => 
                           regs(1663), ZN => n142);
   U180 : NAND3_X1 port map( A1 => n144, A2 => n143, A3 => n142, ZN => 
                           curr_proc_regs(127));
   U181 : NAND2_X1 port map( A1 => regs(640), A2 => n17, ZN => n147);
   U182 : AOI22_X1 port map( A1 => n32, A2 => regs(1152), B1 => n1586, B2 => 
                           regs(128), ZN => n146);
   U183 : AOI22_X1 port map( A1 => n40, A2 => regs(2176), B1 => n9, B2 => 
                           regs(1664), ZN => n145);
   U184 : NAND3_X1 port map( A1 => n147, A2 => n146, A3 => n145, ZN => 
                           curr_proc_regs(128));
   U185 : NAND2_X1 port map( A1 => regs(641), A2 => n17, ZN => n150);
   U186 : AOI22_X1 port map( A1 => n32, A2 => regs(1153), B1 => n8, B2 => 
                           regs(129), ZN => n149);
   U187 : AOI22_X1 port map( A1 => n40, A2 => regs(2177), B1 => n35, B2 => 
                           regs(1665), ZN => n148);
   U188 : NAND3_X1 port map( A1 => n150, A2 => n149, A3 => n148, ZN => 
                           curr_proc_regs(129));
   U189 : NAND2_X1 port map( A1 => regs(524), A2 => n18, ZN => n153);
   U190 : AOI22_X1 port map( A1 => n32, A2 => regs(1036), B1 => n31, B2 => 
                           regs(12), ZN => n152);
   U191 : AOI22_X1 port map( A1 => n42, A2 => regs(2060), B1 => n35, B2 => 
                           regs(1548), ZN => n151);
   U192 : NAND3_X1 port map( A1 => n153, A2 => n152, A3 => n151, ZN => 
                           curr_proc_regs(12));
   U193 : NAND2_X1 port map( A1 => regs(642), A2 => n18, ZN => n156);
   U194 : AOI22_X1 port map( A1 => n32, A2 => regs(1154), B1 => n8, B2 => 
                           regs(130), ZN => n155);
   U195 : AOI22_X1 port map( A1 => n42, A2 => regs(2178), B1 => n35, B2 => 
                           regs(1666), ZN => n154);
   U196 : NAND3_X1 port map( A1 => n156, A2 => n155, A3 => n154, ZN => 
                           curr_proc_regs(130));
   U197 : NAND2_X1 port map( A1 => regs(643), A2 => n18, ZN => n159);
   U198 : AOI22_X1 port map( A1 => n32, A2 => regs(1155), B1 => n8, B2 => 
                           regs(131), ZN => n158);
   U199 : AOI22_X1 port map( A1 => n42, A2 => regs(2179), B1 => n35, B2 => 
                           regs(1667), ZN => n157);
   U200 : NAND3_X1 port map( A1 => n159, A2 => n158, A3 => n157, ZN => 
                           curr_proc_regs(131));
   U201 : NAND2_X1 port map( A1 => regs(644), A2 => n18, ZN => n162);
   U202 : AOI22_X1 port map( A1 => n32, A2 => regs(1156), B1 => n3, B2 => 
                           regs(132), ZN => n161);
   U203 : AOI22_X1 port map( A1 => n42, A2 => regs(2180), B1 => n35, B2 => 
                           regs(1668), ZN => n160);
   U204 : NAND3_X1 port map( A1 => n162, A2 => n161, A3 => n160, ZN => 
                           curr_proc_regs(132));
   U205 : NAND2_X1 port map( A1 => regs(645), A2 => n18, ZN => n165);
   U206 : AOI22_X1 port map( A1 => n32, A2 => regs(1157), B1 => n28, B2 => 
                           regs(133), ZN => n164);
   U207 : AOI22_X1 port map( A1 => n42, A2 => regs(2181), B1 => n35, B2 => 
                           regs(1669), ZN => n163);
   U208 : NAND3_X1 port map( A1 => n165, A2 => n164, A3 => n163, ZN => 
                           curr_proc_regs(133));
   U209 : NAND2_X1 port map( A1 => regs(646), A2 => n18, ZN => n168);
   U210 : AOI22_X1 port map( A1 => n32, A2 => regs(1158), B1 => n8, B2 => 
                           regs(134), ZN => n167);
   U211 : AOI22_X1 port map( A1 => n42, A2 => regs(2182), B1 => n35, B2 => 
                           regs(1670), ZN => n166);
   U212 : NAND3_X1 port map( A1 => n168, A2 => n167, A3 => n166, ZN => 
                           curr_proc_regs(134));
   U213 : NAND2_X1 port map( A1 => regs(647), A2 => n18, ZN => n171);
   U214 : AOI22_X1 port map( A1 => n32, A2 => regs(1159), B1 => n8, B2 => 
                           regs(135), ZN => n170);
   U215 : AOI22_X1 port map( A1 => n42, A2 => regs(2183), B1 => n35, B2 => 
                           regs(1671), ZN => n169);
   U216 : NAND3_X1 port map( A1 => n171, A2 => n170, A3 => n169, ZN => 
                           curr_proc_regs(135));
   U217 : NAND2_X1 port map( A1 => regs(648), A2 => n18, ZN => n174);
   U218 : AOI22_X1 port map( A1 => n32, A2 => regs(1160), B1 => n31, B2 => 
                           regs(136), ZN => n173);
   U219 : AOI22_X1 port map( A1 => n42, A2 => regs(2184), B1 => n35, B2 => 
                           regs(1672), ZN => n172);
   U220 : NAND3_X1 port map( A1 => n174, A2 => n173, A3 => n172, ZN => 
                           curr_proc_regs(136));
   U221 : NAND2_X1 port map( A1 => regs(649), A2 => n18, ZN => n177);
   U222 : AOI22_X1 port map( A1 => n32, A2 => regs(1161), B1 => n28, B2 => 
                           regs(137), ZN => n176);
   U223 : AOI22_X1 port map( A1 => n42, A2 => regs(2185), B1 => n35, B2 => 
                           regs(1673), ZN => n175);
   U224 : NAND3_X1 port map( A1 => n177, A2 => n176, A3 => n175, ZN => 
                           curr_proc_regs(137));
   U225 : NAND2_X1 port map( A1 => regs(650), A2 => n18, ZN => n180);
   U226 : AOI22_X1 port map( A1 => n32, A2 => regs(1162), B1 => n8, B2 => 
                           regs(138), ZN => n179);
   U227 : AOI22_X1 port map( A1 => n42, A2 => regs(2186), B1 => n35, B2 => 
                           regs(1674), ZN => n178);
   U228 : NAND3_X1 port map( A1 => n180, A2 => n179, A3 => n178, ZN => 
                           curr_proc_regs(138));
   U229 : NAND2_X1 port map( A1 => regs(651), A2 => n18, ZN => n183);
   U230 : AOI22_X1 port map( A1 => n32, A2 => regs(1163), B1 => n28, B2 => 
                           regs(139), ZN => n182);
   U231 : AOI22_X1 port map( A1 => n42, A2 => regs(2187), B1 => n35, B2 => 
                           regs(1675), ZN => n181);
   U232 : NAND3_X1 port map( A1 => n183, A2 => n182, A3 => n181, ZN => 
                           curr_proc_regs(139));
   U233 : NAND2_X1 port map( A1 => regs(525), A2 => n19, ZN => n186);
   U234 : AOI22_X1 port map( A1 => n32, A2 => regs(1037), B1 => n25, B2 => 
                           regs(13), ZN => n185);
   U235 : AOI22_X1 port map( A1 => n41, A2 => regs(2061), B1 => n36, B2 => 
                           regs(1549), ZN => n184);
   U236 : NAND3_X1 port map( A1 => n186, A2 => n185, A3 => n184, ZN => 
                           curr_proc_regs(13));
   U237 : NAND2_X1 port map( A1 => regs(652), A2 => n19, ZN => n189);
   U238 : AOI22_X1 port map( A1 => n32, A2 => regs(1164), B1 => n25, B2 => 
                           regs(140), ZN => n188);
   U239 : AOI22_X1 port map( A1 => n41, A2 => regs(2188), B1 => n4, B2 => 
                           regs(1676), ZN => n187);
   U240 : NAND3_X1 port map( A1 => n189, A2 => n188, A3 => n187, ZN => 
                           curr_proc_regs(140));
   U241 : NAND2_X1 port map( A1 => regs(653), A2 => n19, ZN => n192);
   U242 : AOI22_X1 port map( A1 => n32, A2 => regs(1165), B1 => n25, B2 => 
                           regs(141), ZN => n191);
   U243 : AOI22_X1 port map( A1 => n41, A2 => regs(2189), B1 => n36, B2 => 
                           regs(1677), ZN => n190);
   U244 : NAND3_X1 port map( A1 => n192, A2 => n191, A3 => n190, ZN => 
                           curr_proc_regs(141));
   U245 : NAND2_X1 port map( A1 => regs(654), A2 => n19, ZN => n195);
   U246 : AOI22_X1 port map( A1 => n32, A2 => regs(1166), B1 => n25, B2 => 
                           regs(142), ZN => n194);
   U247 : AOI22_X1 port map( A1 => n41, A2 => regs(2190), B1 => n4, B2 => 
                           regs(1678), ZN => n193);
   U248 : NAND3_X1 port map( A1 => n195, A2 => n194, A3 => n193, ZN => 
                           curr_proc_regs(142));
   U249 : NAND2_X1 port map( A1 => regs(655), A2 => n19, ZN => n198);
   U250 : AOI22_X1 port map( A1 => n32, A2 => regs(1167), B1 => n25, B2 => 
                           regs(143), ZN => n197);
   U251 : AOI22_X1 port map( A1 => n41, A2 => regs(2191), B1 => n36, B2 => 
                           regs(1679), ZN => n196);
   U252 : NAND3_X1 port map( A1 => n198, A2 => n197, A3 => n196, ZN => 
                           curr_proc_regs(143));
   U253 : NAND2_X1 port map( A1 => regs(656), A2 => n19, ZN => n201);
   U254 : AOI22_X1 port map( A1 => n32, A2 => regs(1168), B1 => n25, B2 => 
                           regs(144), ZN => n200);
   U255 : AOI22_X1 port map( A1 => n41, A2 => regs(2192), B1 => n4, B2 => 
                           regs(1680), ZN => n199);
   U256 : NAND3_X1 port map( A1 => n201, A2 => n200, A3 => n199, ZN => 
                           curr_proc_regs(144));
   U257 : NAND2_X1 port map( A1 => regs(657), A2 => n19, ZN => n204);
   U258 : AOI22_X1 port map( A1 => n32, A2 => regs(1169), B1 => n25, B2 => 
                           regs(145), ZN => n203);
   U259 : AOI22_X1 port map( A1 => n41, A2 => regs(2193), B1 => n36, B2 => 
                           regs(1681), ZN => n202);
   U260 : NAND3_X1 port map( A1 => n204, A2 => n203, A3 => n202, ZN => 
                           curr_proc_regs(145));
   U261 : NAND2_X1 port map( A1 => regs(658), A2 => n19, ZN => n207);
   U262 : AOI22_X1 port map( A1 => n32, A2 => regs(1170), B1 => n25, B2 => 
                           regs(146), ZN => n206);
   U263 : AOI22_X1 port map( A1 => n41, A2 => regs(2194), B1 => n4, B2 => 
                           regs(1682), ZN => n205);
   U264 : NAND3_X1 port map( A1 => n207, A2 => n206, A3 => n205, ZN => 
                           curr_proc_regs(146));
   U265 : NAND2_X1 port map( A1 => regs(659), A2 => n19, ZN => n210);
   U266 : AOI22_X1 port map( A1 => n32, A2 => regs(1171), B1 => n25, B2 => 
                           regs(147), ZN => n209);
   U267 : AOI22_X1 port map( A1 => n41, A2 => regs(2195), B1 => n36, B2 => 
                           regs(1683), ZN => n208);
   U268 : NAND3_X1 port map( A1 => n210, A2 => n209, A3 => n208, ZN => 
                           curr_proc_regs(147));
   U269 : NAND2_X1 port map( A1 => regs(660), A2 => n19, ZN => n213);
   U270 : AOI22_X1 port map( A1 => n32, A2 => regs(1172), B1 => n25, B2 => 
                           regs(148), ZN => n212);
   U271 : AOI22_X1 port map( A1 => n41, A2 => regs(2196), B1 => n4, B2 => 
                           regs(1684), ZN => n211);
   U272 : NAND3_X1 port map( A1 => n213, A2 => n212, A3 => n211, ZN => 
                           curr_proc_regs(148));
   U273 : NAND2_X1 port map( A1 => regs(661), A2 => n19, ZN => n216);
   U274 : AOI22_X1 port map( A1 => n32, A2 => regs(1173), B1 => n25, B2 => 
                           regs(149), ZN => n215);
   U275 : AOI22_X1 port map( A1 => n41, A2 => regs(2197), B1 => n36, B2 => 
                           regs(1685), ZN => n214);
   U276 : NAND3_X1 port map( A1 => n216, A2 => n215, A3 => n214, ZN => 
                           curr_proc_regs(149));
   U277 : NAND2_X1 port map( A1 => regs(526), A2 => n19, ZN => n219);
   U278 : AOI22_X1 port map( A1 => n32, A2 => regs(1038), B1 => n26, B2 => 
                           regs(14), ZN => n218);
   U279 : AOI22_X1 port map( A1 => n40, A2 => regs(2062), B1 => n9, B2 => 
                           regs(1550), ZN => n217);
   U280 : NAND3_X1 port map( A1 => n219, A2 => n218, A3 => n217, ZN => 
                           curr_proc_regs(14));
   U281 : NAND2_X1 port map( A1 => regs(662), A2 => n6, ZN => n222);
   U282 : AOI22_X1 port map( A1 => n32, A2 => regs(1174), B1 => n1586, B2 => 
                           regs(150), ZN => n221);
   U283 : AOI22_X1 port map( A1 => n40, A2 => regs(2198), B1 => n36, B2 => 
                           regs(1686), ZN => n220);
   U284 : NAND3_X1 port map( A1 => n222, A2 => n221, A3 => n220, ZN => 
                           curr_proc_regs(150));
   U285 : NAND2_X1 port map( A1 => regs(663), A2 => n2, ZN => n225);
   U286 : AOI22_X1 port map( A1 => n32, A2 => regs(1175), B1 => n3, B2 => 
                           regs(151), ZN => n224);
   U287 : AOI22_X1 port map( A1 => n40, A2 => regs(2199), B1 => n4, B2 => 
                           regs(1687), ZN => n223);
   U288 : NAND3_X1 port map( A1 => n225, A2 => n224, A3 => n223, ZN => 
                           curr_proc_regs(151));
   U289 : NAND2_X1 port map( A1 => regs(664), A2 => n22, ZN => n228);
   U290 : AOI22_X1 port map( A1 => n32, A2 => regs(1176), B1 => n1586, B2 => 
                           regs(152), ZN => n227);
   U291 : AOI22_X1 port map( A1 => n40, A2 => regs(2200), B1 => n9, B2 => 
                           regs(1688), ZN => n226);
   U292 : NAND3_X1 port map( A1 => n228, A2 => n227, A3 => n226, ZN => 
                           curr_proc_regs(152));
   U293 : NAND2_X1 port map( A1 => regs(665), A2 => n1585, ZN => n231);
   U294 : AOI22_X1 port map( A1 => n32, A2 => regs(1177), B1 => n28, B2 => 
                           regs(153), ZN => n230);
   U295 : AOI22_X1 port map( A1 => n41, A2 => regs(2201), B1 => n34, B2 => 
                           regs(1689), ZN => n229);
   U296 : NAND3_X1 port map( A1 => n231, A2 => n230, A3 => n229, ZN => 
                           curr_proc_regs(153));
   U297 : NAND2_X1 port map( A1 => regs(666), A2 => n19, ZN => n234);
   U298 : AOI22_X1 port map( A1 => n32, A2 => regs(1178), B1 => n25, B2 => 
                           regs(154), ZN => n233);
   U299 : AOI22_X1 port map( A1 => n42, A2 => regs(2202), B1 => n34, B2 => 
                           regs(1690), ZN => n232);
   U300 : NAND3_X1 port map( A1 => n234, A2 => n233, A3 => n232, ZN => 
                           curr_proc_regs(154));
   U301 : NAND2_X1 port map( A1 => regs(667), A2 => n6, ZN => n237);
   U302 : AOI22_X1 port map( A1 => n32, A2 => regs(1179), B1 => n26, B2 => 
                           regs(155), ZN => n236);
   U303 : AOI22_X1 port map( A1 => n40, A2 => regs(2203), B1 => n9, B2 => 
                           regs(1691), ZN => n235);
   U304 : NAND3_X1 port map( A1 => n237, A2 => n236, A3 => n235, ZN => 
                           curr_proc_regs(155));
   U305 : NAND2_X1 port map( A1 => regs(668), A2 => n2, ZN => n240);
   U306 : AOI22_X1 port map( A1 => n32, A2 => regs(1180), B1 => n1586, B2 => 
                           regs(156), ZN => n239);
   U307 : AOI22_X1 port map( A1 => n13, A2 => regs(2204), B1 => n36, B2 => 
                           regs(1692), ZN => n238);
   U308 : NAND3_X1 port map( A1 => n240, A2 => n239, A3 => n238, ZN => 
                           curr_proc_regs(156));
   U309 : NAND2_X1 port map( A1 => regs(669), A2 => n22, ZN => n243);
   U310 : AOI22_X1 port map( A1 => n32, A2 => regs(1181), B1 => n3, B2 => 
                           regs(157), ZN => n242);
   U311 : AOI22_X1 port map( A1 => n40, A2 => regs(2205), B1 => n9, B2 => 
                           regs(1693), ZN => n241);
   U312 : NAND3_X1 port map( A1 => n243, A2 => n242, A3 => n241, ZN => 
                           curr_proc_regs(157));
   U313 : NAND2_X1 port map( A1 => regs(670), A2 => n1585, ZN => n246);
   U314 : AOI22_X1 port map( A1 => n32, A2 => regs(1182), B1 => n28, B2 => 
                           regs(158), ZN => n245);
   U315 : AOI22_X1 port map( A1 => n40, A2 => regs(2206), B1 => n34, B2 => 
                           regs(1694), ZN => n244);
   U316 : NAND3_X1 port map( A1 => n246, A2 => n245, A3 => n244, ZN => 
                           curr_proc_regs(158));
   U317 : NAND2_X1 port map( A1 => regs(671), A2 => n19, ZN => n249);
   U318 : AOI22_X1 port map( A1 => n32, A2 => regs(1183), B1 => n1586, B2 => 
                           regs(159), ZN => n248);
   U319 : AOI22_X1 port map( A1 => n41, A2 => regs(2207), B1 => n4, B2 => 
                           regs(1695), ZN => n247);
   U320 : NAND3_X1 port map( A1 => n249, A2 => n248, A3 => n247, ZN => 
                           curr_proc_regs(159));
   U321 : NAND2_X1 port map( A1 => regs(527), A2 => n2, ZN => n252);
   U322 : AOI22_X1 port map( A1 => n32, A2 => regs(1039), B1 => n26, B2 => 
                           regs(15), ZN => n251);
   U323 : AOI22_X1 port map( A1 => n44, A2 => regs(2063), B1 => n9, B2 => 
                           regs(1551), ZN => n250);
   U324 : NAND3_X1 port map( A1 => n252, A2 => n251, A3 => n250, ZN => 
                           curr_proc_regs(15));
   U325 : NAND2_X1 port map( A1 => regs(672), A2 => n2, ZN => n255);
   U326 : AOI22_X1 port map( A1 => n32, A2 => regs(1184), B1 => n26, B2 => 
                           regs(160), ZN => n254);
   U327 : AOI22_X1 port map( A1 => n44, A2 => regs(2208), B1 => n9, B2 => 
                           regs(1696), ZN => n253);
   U328 : NAND3_X1 port map( A1 => n255, A2 => n254, A3 => n253, ZN => 
                           curr_proc_regs(160));
   U329 : NAND2_X1 port map( A1 => regs(673), A2 => n2, ZN => n258);
   U330 : AOI22_X1 port map( A1 => n32, A2 => regs(1185), B1 => n26, B2 => 
                           regs(161), ZN => n257);
   U331 : AOI22_X1 port map( A1 => n44, A2 => regs(2209), B1 => n9, B2 => 
                           regs(1697), ZN => n256);
   U332 : NAND3_X1 port map( A1 => n258, A2 => n257, A3 => n256, ZN => 
                           curr_proc_regs(161));
   U333 : NAND2_X1 port map( A1 => regs(674), A2 => n2, ZN => n261);
   U334 : AOI22_X1 port map( A1 => n32, A2 => regs(1186), B1 => n26, B2 => 
                           regs(162), ZN => n260);
   U335 : AOI22_X1 port map( A1 => n11, A2 => regs(2210), B1 => n9, B2 => 
                           regs(1698), ZN => n259);
   U336 : NAND3_X1 port map( A1 => n261, A2 => n260, A3 => n259, ZN => 
                           curr_proc_regs(162));
   U337 : NAND2_X1 port map( A1 => regs(675), A2 => n2, ZN => n264);
   U338 : AOI22_X1 port map( A1 => n32, A2 => regs(1187), B1 => n26, B2 => 
                           regs(163), ZN => n263);
   U339 : AOI22_X1 port map( A1 => n11, A2 => regs(2211), B1 => n9, B2 => 
                           regs(1699), ZN => n262);
   U340 : NAND3_X1 port map( A1 => n264, A2 => n263, A3 => n262, ZN => 
                           curr_proc_regs(163));
   U341 : NAND2_X1 port map( A1 => regs(676), A2 => n2, ZN => n267);
   U342 : AOI22_X1 port map( A1 => n32, A2 => regs(1188), B1 => n26, B2 => 
                           regs(164), ZN => n266);
   U343 : AOI22_X1 port map( A1 => n44, A2 => regs(2212), B1 => n9, B2 => 
                           regs(1700), ZN => n265);
   U344 : NAND3_X1 port map( A1 => n267, A2 => n266, A3 => n265, ZN => 
                           curr_proc_regs(164));
   U345 : NAND2_X1 port map( A1 => regs(677), A2 => n2, ZN => n270);
   U346 : AOI22_X1 port map( A1 => n32, A2 => regs(1189), B1 => n26, B2 => 
                           regs(165), ZN => n269);
   U347 : AOI22_X1 port map( A1 => n44, A2 => regs(2213), B1 => n9, B2 => 
                           regs(1701), ZN => n268);
   U348 : NAND3_X1 port map( A1 => n270, A2 => n269, A3 => n268, ZN => 
                           curr_proc_regs(165));
   U349 : NAND2_X1 port map( A1 => regs(678), A2 => n2, ZN => n273);
   U350 : AOI22_X1 port map( A1 => n32, A2 => regs(1190), B1 => n26, B2 => 
                           regs(166), ZN => n272);
   U351 : AOI22_X1 port map( A1 => n11, A2 => regs(2214), B1 => n9, B2 => 
                           regs(1702), ZN => n271);
   U352 : NAND3_X1 port map( A1 => n273, A2 => n272, A3 => n271, ZN => 
                           curr_proc_regs(166));
   U353 : NAND2_X1 port map( A1 => regs(679), A2 => n2, ZN => n276);
   U354 : AOI22_X1 port map( A1 => n32, A2 => regs(1191), B1 => n26, B2 => 
                           regs(167), ZN => n275);
   U355 : AOI22_X1 port map( A1 => n11, A2 => regs(2215), B1 => n9, B2 => 
                           regs(1703), ZN => n274);
   U356 : NAND3_X1 port map( A1 => n276, A2 => n275, A3 => n274, ZN => 
                           curr_proc_regs(167));
   U357 : NAND2_X1 port map( A1 => regs(680), A2 => n2, ZN => n279);
   U358 : AOI22_X1 port map( A1 => n32, A2 => regs(1192), B1 => n26, B2 => 
                           regs(168), ZN => n278);
   U359 : AOI22_X1 port map( A1 => n11, A2 => regs(2216), B1 => n9, B2 => 
                           regs(1704), ZN => n277);
   U360 : NAND3_X1 port map( A1 => n279, A2 => n278, A3 => n277, ZN => 
                           curr_proc_regs(168));
   U361 : NAND2_X1 port map( A1 => regs(681), A2 => n2, ZN => n282);
   U362 : AOI22_X1 port map( A1 => n32, A2 => regs(1193), B1 => n26, B2 => 
                           regs(169), ZN => n281);
   U363 : AOI22_X1 port map( A1 => n11, A2 => regs(2217), B1 => n9, B2 => 
                           regs(1705), ZN => n280);
   U364 : NAND3_X1 port map( A1 => n282, A2 => n281, A3 => n280, ZN => 
                           curr_proc_regs(169));
   U365 : NAND2_X1 port map( A1 => regs(528), A2 => n22, ZN => n285);
   U366 : AOI22_X1 port map( A1 => n32, A2 => regs(1040), B1 => n31, B2 => 
                           regs(16), ZN => n284);
   U367 : AOI22_X1 port map( A1 => n11, A2 => regs(2064), B1 => n35, B2 => 
                           regs(1552), ZN => n283);
   U368 : NAND3_X1 port map( A1 => n285, A2 => n284, A3 => n283, ZN => 
                           curr_proc_regs(16));
   U369 : NAND2_X1 port map( A1 => regs(682), A2 => n22, ZN => n288);
   U370 : AOI22_X1 port map( A1 => n32, A2 => regs(1194), B1 => n1586, B2 => 
                           regs(170), ZN => n287);
   U371 : AOI22_X1 port map( A1 => n44, A2 => regs(2218), B1 => n37, B2 => 
                           regs(1706), ZN => n286);
   U372 : NAND3_X1 port map( A1 => n288, A2 => n287, A3 => n286, ZN => 
                           curr_proc_regs(170));
   U373 : NAND2_X1 port map( A1 => regs(683), A2 => n22, ZN => n291);
   U374 : AOI22_X1 port map( A1 => n32, A2 => regs(1195), B1 => n1586, B2 => 
                           regs(171), ZN => n290);
   U375 : AOI22_X1 port map( A1 => n44, A2 => regs(2219), B1 => n34, B2 => 
                           regs(1707), ZN => n289);
   U376 : NAND3_X1 port map( A1 => n291, A2 => n290, A3 => n289, ZN => 
                           curr_proc_regs(171));
   U377 : NAND2_X1 port map( A1 => regs(684), A2 => n22, ZN => n294);
   U378 : AOI22_X1 port map( A1 => n32, A2 => regs(1196), B1 => n8, B2 => 
                           regs(172), ZN => n293);
   U379 : AOI22_X1 port map( A1 => n11, A2 => regs(2220), B1 => n35, B2 => 
                           regs(1708), ZN => n292);
   U380 : NAND3_X1 port map( A1 => n294, A2 => n293, A3 => n292, ZN => 
                           curr_proc_regs(172));
   U381 : NAND2_X1 port map( A1 => regs(685), A2 => n22, ZN => n297);
   U382 : AOI22_X1 port map( A1 => n32, A2 => regs(1197), B1 => n26, B2 => 
                           regs(173), ZN => n296);
   U383 : AOI22_X1 port map( A1 => n11, A2 => regs(2221), B1 => n37, B2 => 
                           regs(1709), ZN => n295);
   U384 : NAND3_X1 port map( A1 => n297, A2 => n296, A3 => n295, ZN => 
                           curr_proc_regs(173));
   U385 : NAND2_X1 port map( A1 => regs(686), A2 => n22, ZN => n300);
   U386 : AOI22_X1 port map( A1 => n32, A2 => regs(1198), B1 => n3, B2 => 
                           regs(174), ZN => n299);
   U387 : AOI22_X1 port map( A1 => n11, A2 => regs(2222), B1 => n34, B2 => 
                           regs(1710), ZN => n298);
   U388 : NAND3_X1 port map( A1 => n300, A2 => n299, A3 => n298, ZN => 
                           curr_proc_regs(174));
   U389 : NAND2_X1 port map( A1 => regs(687), A2 => n22, ZN => n303);
   U390 : AOI22_X1 port map( A1 => n32, A2 => regs(1199), B1 => n8, B2 => 
                           regs(175), ZN => n302);
   U391 : AOI22_X1 port map( A1 => n44, A2 => regs(2223), B1 => n35, B2 => 
                           regs(1711), ZN => n301);
   U392 : NAND3_X1 port map( A1 => n303, A2 => n302, A3 => n301, ZN => 
                           curr_proc_regs(175));
   U393 : NAND2_X1 port map( A1 => regs(688), A2 => n22, ZN => n306);
   U394 : AOI22_X1 port map( A1 => n32, A2 => regs(1200), B1 => n27, B2 => 
                           regs(176), ZN => n305);
   U395 : AOI22_X1 port map( A1 => n11, A2 => regs(2224), B1 => n37, B2 => 
                           regs(1712), ZN => n304);
   U396 : NAND3_X1 port map( A1 => n306, A2 => n305, A3 => n304, ZN => 
                           curr_proc_regs(176));
   U397 : NAND2_X1 port map( A1 => regs(689), A2 => n22, ZN => n309);
   U398 : AOI22_X1 port map( A1 => n32, A2 => regs(1201), B1 => n31, B2 => 
                           regs(177), ZN => n308);
   U399 : AOI22_X1 port map( A1 => n11, A2 => regs(2225), B1 => n34, B2 => 
                           regs(1713), ZN => n307);
   U400 : NAND3_X1 port map( A1 => n309, A2 => n308, A3 => n307, ZN => 
                           curr_proc_regs(177));
   U401 : NAND2_X1 port map( A1 => regs(690), A2 => n22, ZN => n312);
   U402 : AOI22_X1 port map( A1 => n32, A2 => regs(1202), B1 => n25, B2 => 
                           regs(178), ZN => n311);
   U403 : AOI22_X1 port map( A1 => n11, A2 => regs(2226), B1 => n35, B2 => 
                           regs(1714), ZN => n310);
   U404 : NAND3_X1 port map( A1 => n312, A2 => n311, A3 => n310, ZN => 
                           curr_proc_regs(178));
   U405 : NAND2_X1 port map( A1 => regs(691), A2 => n22, ZN => n315);
   U406 : AOI22_X1 port map( A1 => n32, A2 => regs(1203), B1 => n3, B2 => 
                           regs(179), ZN => n314);
   U407 : AOI22_X1 port map( A1 => n44, A2 => regs(2227), B1 => n37, B2 => 
                           regs(1715), ZN => n313);
   U408 : NAND3_X1 port map( A1 => n315, A2 => n314, A3 => n313, ZN => 
                           curr_proc_regs(179));
   U409 : NAND2_X1 port map( A1 => regs(529), A2 => n20, ZN => n318);
   U410 : AOI22_X1 port map( A1 => n32, A2 => regs(1041), B1 => n25, B2 => 
                           regs(17), ZN => n317);
   U411 : AOI22_X1 port map( A1 => n44, A2 => regs(2065), B1 => n37, B2 => 
                           regs(1553), ZN => n316);
   U412 : NAND3_X1 port map( A1 => n318, A2 => n317, A3 => n316, ZN => 
                           curr_proc_regs(17));
   U413 : NAND2_X1 port map( A1 => regs(692), A2 => n20, ZN => n321);
   U414 : AOI22_X1 port map( A1 => n32, A2 => regs(1204), B1 => n3, B2 => 
                           regs(180), ZN => n320);
   U415 : AOI22_X1 port map( A1 => n11, A2 => regs(2228), B1 => n34, B2 => 
                           regs(1716), ZN => n319);
   U416 : NAND3_X1 port map( A1 => n321, A2 => n320, A3 => n319, ZN => 
                           curr_proc_regs(180));
   U417 : NAND2_X1 port map( A1 => regs(693), A2 => n20, ZN => n324);
   U418 : AOI22_X1 port map( A1 => n32, A2 => regs(1205), B1 => n8, B2 => 
                           regs(181), ZN => n323);
   U419 : AOI22_X1 port map( A1 => n11, A2 => regs(2229), B1 => n9, B2 => 
                           regs(1717), ZN => n322);
   U420 : NAND3_X1 port map( A1 => n324, A2 => n323, A3 => n322, ZN => 
                           curr_proc_regs(181));
   U421 : NAND2_X1 port map( A1 => regs(694), A2 => n20, ZN => n327);
   U422 : AOI22_X1 port map( A1 => n32, A2 => regs(1206), B1 => n25, B2 => 
                           regs(182), ZN => n326);
   U423 : AOI22_X1 port map( A1 => n44, A2 => regs(2230), B1 => n37, B2 => 
                           regs(1718), ZN => n325);
   U424 : NAND3_X1 port map( A1 => n327, A2 => n326, A3 => n325, ZN => 
                           curr_proc_regs(182));
   U425 : NAND2_X1 port map( A1 => regs(695), A2 => n20, ZN => n330);
   U426 : AOI22_X1 port map( A1 => n32, A2 => regs(1207), B1 => n26, B2 => 
                           regs(183), ZN => n329);
   U427 : AOI22_X1 port map( A1 => n11, A2 => regs(2231), B1 => n4, B2 => 
                           regs(1719), ZN => n328);
   U428 : NAND3_X1 port map( A1 => n330, A2 => n329, A3 => n328, ZN => 
                           curr_proc_regs(183));
   U429 : NAND2_X1 port map( A1 => regs(696), A2 => n20, ZN => n333);
   U430 : AOI22_X1 port map( A1 => n32, A2 => regs(1208), B1 => n1586, B2 => 
                           regs(184), ZN => n332);
   U431 : AOI22_X1 port map( A1 => n11, A2 => regs(2232), B1 => n9, B2 => 
                           regs(1720), ZN => n331);
   U432 : NAND3_X1 port map( A1 => n333, A2 => n332, A3 => n331, ZN => 
                           curr_proc_regs(184));
   U433 : NAND2_X1 port map( A1 => regs(697), A2 => n20, ZN => n336);
   U434 : AOI22_X1 port map( A1 => n32, A2 => regs(1209), B1 => n3, B2 => 
                           regs(185), ZN => n335);
   U435 : AOI22_X1 port map( A1 => n44, A2 => regs(2233), B1 => n4, B2 => 
                           regs(1721), ZN => n334);
   U436 : NAND3_X1 port map( A1 => n336, A2 => n335, A3 => n334, ZN => 
                           curr_proc_regs(185));
   U437 : NAND2_X1 port map( A1 => regs(698), A2 => n20, ZN => n339);
   U438 : AOI22_X1 port map( A1 => n32, A2 => regs(1210), B1 => n31, B2 => 
                           regs(186), ZN => n338);
   U439 : AOI22_X1 port map( A1 => n11, A2 => regs(2234), B1 => n37, B2 => 
                           regs(1722), ZN => n337);
   U440 : NAND3_X1 port map( A1 => n339, A2 => n338, A3 => n337, ZN => 
                           curr_proc_regs(186));
   U441 : NAND2_X1 port map( A1 => regs(699), A2 => n20, ZN => n342);
   U442 : AOI22_X1 port map( A1 => n32, A2 => regs(1211), B1 => n8, B2 => 
                           regs(187), ZN => n341);
   U443 : AOI22_X1 port map( A1 => n11, A2 => regs(2235), B1 => n35, B2 => 
                           regs(1723), ZN => n340);
   U444 : NAND3_X1 port map( A1 => n342, A2 => n341, A3 => n340, ZN => 
                           curr_proc_regs(187));
   U445 : NAND2_X1 port map( A1 => regs(700), A2 => n20, ZN => n345);
   U446 : AOI22_X1 port map( A1 => n32, A2 => regs(1212), B1 => n25, B2 => 
                           regs(188), ZN => n344);
   U447 : AOI22_X1 port map( A1 => n44, A2 => regs(2236), B1 => n36, B2 => 
                           regs(1724), ZN => n343);
   U448 : NAND3_X1 port map( A1 => n345, A2 => n344, A3 => n343, ZN => 
                           curr_proc_regs(188));
   U449 : NAND2_X1 port map( A1 => regs(701), A2 => n20, ZN => n348);
   U450 : AOI22_X1 port map( A1 => n32, A2 => regs(1213), B1 => n29, B2 => 
                           regs(189), ZN => n347);
   U451 : AOI22_X1 port map( A1 => n11, A2 => regs(2237), B1 => n9, B2 => 
                           regs(1725), ZN => n346);
   U452 : NAND3_X1 port map( A1 => n348, A2 => n347, A3 => n346, ZN => 
                           curr_proc_regs(189));
   U453 : NAND2_X1 port map( A1 => regs(530), A2 => n21, ZN => n351);
   U454 : AOI22_X1 port map( A1 => n32, A2 => regs(1042), B1 => n1586, B2 => 
                           regs(18), ZN => n350);
   U455 : AOI22_X1 port map( A1 => n11, A2 => regs(2066), B1 => n34, B2 => 
                           regs(1554), ZN => n349);
   U456 : NAND3_X1 port map( A1 => n351, A2 => n350, A3 => n349, ZN => 
                           curr_proc_regs(18));
   U457 : NAND2_X1 port map( A1 => regs(702), A2 => n21, ZN => n354);
   U458 : AOI22_X1 port map( A1 => n32, A2 => regs(1214), B1 => n8, B2 => 
                           regs(190), ZN => n353);
   U459 : AOI22_X1 port map( A1 => n11, A2 => regs(2238), B1 => n35, B2 => 
                           regs(1726), ZN => n352);
   U460 : NAND3_X1 port map( A1 => n354, A2 => n353, A3 => n352, ZN => 
                           curr_proc_regs(190));
   U461 : NAND2_X1 port map( A1 => regs(703), A2 => n21, ZN => n357);
   U462 : AOI22_X1 port map( A1 => n32, A2 => regs(1215), B1 => n26, B2 => 
                           regs(191), ZN => n356);
   U463 : AOI22_X1 port map( A1 => n11, A2 => regs(2239), B1 => n34, B2 => 
                           regs(1727), ZN => n355);
   U464 : NAND3_X1 port map( A1 => n357, A2 => n356, A3 => n355, ZN => 
                           curr_proc_regs(191));
   U465 : NAND2_X1 port map( A1 => regs(704), A2 => n21, ZN => n360);
   U466 : AOI22_X1 port map( A1 => n32, A2 => regs(1216), B1 => n3, B2 => 
                           regs(192), ZN => n359);
   U467 : AOI22_X1 port map( A1 => n11, A2 => regs(2240), B1 => n34, B2 => 
                           regs(1728), ZN => n358);
   U468 : NAND3_X1 port map( A1 => n360, A2 => n359, A3 => n358, ZN => 
                           curr_proc_regs(192));
   U469 : NAND2_X1 port map( A1 => regs(705), A2 => n21, ZN => n363);
   U470 : AOI22_X1 port map( A1 => n32, A2 => regs(1217), B1 => n8, B2 => 
                           regs(193), ZN => n362);
   U471 : AOI22_X1 port map( A1 => n11, A2 => regs(2241), B1 => n35, B2 => 
                           regs(1729), ZN => n361);
   U472 : NAND3_X1 port map( A1 => n363, A2 => n362, A3 => n361, ZN => 
                           curr_proc_regs(193));
   U473 : NAND2_X1 port map( A1 => regs(706), A2 => n21, ZN => n366);
   U474 : AOI22_X1 port map( A1 => n32, A2 => regs(1218), B1 => n31, B2 => 
                           regs(194), ZN => n365);
   U475 : AOI22_X1 port map( A1 => n11, A2 => regs(2242), B1 => n35, B2 => 
                           regs(1730), ZN => n364);
   U476 : NAND3_X1 port map( A1 => n366, A2 => n365, A3 => n364, ZN => 
                           curr_proc_regs(194));
   U477 : NAND2_X1 port map( A1 => regs(707), A2 => n21, ZN => n369);
   U478 : AOI22_X1 port map( A1 => n32, A2 => regs(1219), B1 => n25, B2 => 
                           regs(195), ZN => n368);
   U479 : AOI22_X1 port map( A1 => n11, A2 => regs(2243), B1 => n34, B2 => 
                           regs(1731), ZN => n367);
   U480 : NAND3_X1 port map( A1 => n369, A2 => n368, A3 => n367, ZN => 
                           curr_proc_regs(195));
   U481 : NAND2_X1 port map( A1 => regs(708), A2 => n21, ZN => n372);
   U482 : AOI22_X1 port map( A1 => n32, A2 => regs(1220), B1 => n28, B2 => 
                           regs(196), ZN => n371);
   U483 : AOI22_X1 port map( A1 => n11, A2 => regs(2244), B1 => n35, B2 => 
                           regs(1732), ZN => n370);
   U484 : NAND3_X1 port map( A1 => n372, A2 => n371, A3 => n370, ZN => 
                           curr_proc_regs(196));
   U485 : NAND2_X1 port map( A1 => regs(709), A2 => n21, ZN => n375);
   U486 : AOI22_X1 port map( A1 => n32, A2 => regs(1221), B1 => n27, B2 => 
                           regs(197), ZN => n374);
   U487 : AOI22_X1 port map( A1 => n11, A2 => regs(2245), B1 => n37, B2 => 
                           regs(1733), ZN => n373);
   U488 : NAND3_X1 port map( A1 => n375, A2 => n374, A3 => n373, ZN => 
                           curr_proc_regs(197));
   U489 : NAND2_X1 port map( A1 => regs(710), A2 => n21, ZN => n378);
   U490 : AOI22_X1 port map( A1 => n32, A2 => regs(1222), B1 => n8, B2 => 
                           regs(198), ZN => n377);
   U491 : AOI22_X1 port map( A1 => n11, A2 => regs(2246), B1 => n34, B2 => 
                           regs(1734), ZN => n376);
   U492 : NAND3_X1 port map( A1 => n378, A2 => n377, A3 => n376, ZN => 
                           curr_proc_regs(198));
   U493 : NAND2_X1 port map( A1 => regs(711), A2 => n21, ZN => n381);
   U494 : AOI22_X1 port map( A1 => n32, A2 => regs(1223), B1 => n29, B2 => 
                           regs(199), ZN => n380);
   U495 : AOI22_X1 port map( A1 => n11, A2 => regs(2247), B1 => n35, B2 => 
                           regs(1735), ZN => n379);
   U496 : NAND3_X1 port map( A1 => n381, A2 => n380, A3 => n379, ZN => 
                           curr_proc_regs(199));
   U497 : NAND2_X1 port map( A1 => regs(531), A2 => n1, ZN => n384);
   U498 : AOI22_X1 port map( A1 => n32, A2 => regs(1043), B1 => n3, B2 => 
                           regs(19), ZN => n383);
   U499 : AOI22_X1 port map( A1 => n11, A2 => regs(2067), B1 => n4, B2 => 
                           regs(1555), ZN => n382);
   U500 : NAND3_X1 port map( A1 => n384, A2 => n383, A3 => n382, ZN => 
                           curr_proc_regs(19));
   U501 : NAND2_X1 port map( A1 => regs(513), A2 => n1, ZN => n387);
   U502 : AOI22_X1 port map( A1 => n32, A2 => regs(1025), B1 => n28, B2 => 
                           regs(1), ZN => n386);
   U503 : AOI22_X1 port map( A1 => n11, A2 => regs(2049), B1 => n1588, B2 => 
                           regs(1537), ZN => n385);
   U504 : NAND3_X1 port map( A1 => n387, A2 => n386, A3 => n385, ZN => 
                           curr_proc_regs(1));
   U505 : NAND2_X1 port map( A1 => regs(712), A2 => n1, ZN => n390);
   U506 : AOI22_X1 port map( A1 => n32, A2 => regs(1224), B1 => n25, B2 => 
                           regs(200), ZN => n389);
   U507 : AOI22_X1 port map( A1 => n11, A2 => regs(2248), B1 => n34, B2 => 
                           regs(1736), ZN => n388);
   U508 : NAND3_X1 port map( A1 => n390, A2 => n389, A3 => n388, ZN => 
                           curr_proc_regs(200));
   U509 : NAND2_X1 port map( A1 => regs(713), A2 => n1, ZN => n393);
   U510 : AOI22_X1 port map( A1 => n32, A2 => regs(1225), B1 => n8, B2 => 
                           regs(201), ZN => n392);
   U511 : AOI22_X1 port map( A1 => n11, A2 => regs(2249), B1 => n35, B2 => 
                           regs(1737), ZN => n391);
   U512 : NAND3_X1 port map( A1 => n393, A2 => n392, A3 => n391, ZN => 
                           curr_proc_regs(201));
   U513 : NAND2_X1 port map( A1 => regs(714), A2 => n1, ZN => n396);
   U514 : AOI22_X1 port map( A1 => n32, A2 => regs(1226), B1 => n29, B2 => 
                           regs(202), ZN => n395);
   U515 : AOI22_X1 port map( A1 => n11, A2 => regs(2250), B1 => n36, B2 => 
                           regs(1738), ZN => n394);
   U516 : NAND3_X1 port map( A1 => n396, A2 => n395, A3 => n394, ZN => 
                           curr_proc_regs(202));
   U517 : NAND2_X1 port map( A1 => regs(715), A2 => n1, ZN => n399);
   U518 : AOI22_X1 port map( A1 => n32, A2 => regs(1227), B1 => n31, B2 => 
                           regs(203), ZN => n398);
   U519 : AOI22_X1 port map( A1 => n11, A2 => regs(2251), B1 => n39, B2 => 
                           regs(1739), ZN => n397);
   U520 : NAND3_X1 port map( A1 => n399, A2 => n398, A3 => n397, ZN => 
                           curr_proc_regs(203));
   U521 : NAND2_X1 port map( A1 => regs(716), A2 => n1, ZN => n402);
   U522 : AOI22_X1 port map( A1 => n32, A2 => regs(1228), B1 => n28, B2 => 
                           regs(204), ZN => n401);
   U523 : AOI22_X1 port map( A1 => n11, A2 => regs(2252), B1 => n38, B2 => 
                           regs(1740), ZN => n400);
   U524 : NAND3_X1 port map( A1 => n402, A2 => n401, A3 => n400, ZN => 
                           curr_proc_regs(204));
   U525 : NAND2_X1 port map( A1 => regs(717), A2 => n1, ZN => n405);
   U526 : AOI22_X1 port map( A1 => n32, A2 => regs(1229), B1 => n29, B2 => 
                           regs(205), ZN => n404);
   U527 : AOI22_X1 port map( A1 => n11, A2 => regs(2253), B1 => n35, B2 => 
                           regs(1741), ZN => n403);
   U528 : NAND3_X1 port map( A1 => n405, A2 => n404, A3 => n403, ZN => 
                           curr_proc_regs(205));
   U529 : NAND2_X1 port map( A1 => regs(718), A2 => n1, ZN => n408);
   U530 : AOI22_X1 port map( A1 => n32, A2 => regs(1230), B1 => n8, B2 => 
                           regs(206), ZN => n407);
   U531 : AOI22_X1 port map( A1 => n11, A2 => regs(2254), B1 => n34, B2 => 
                           regs(1742), ZN => n406);
   U532 : NAND3_X1 port map( A1 => n408, A2 => n407, A3 => n406, ZN => 
                           curr_proc_regs(206));
   U533 : NAND2_X1 port map( A1 => regs(719), A2 => n1, ZN => n411);
   U534 : AOI22_X1 port map( A1 => n32, A2 => regs(1231), B1 => n31, B2 => 
                           regs(207), ZN => n410);
   U535 : AOI22_X1 port map( A1 => n11, A2 => regs(2255), B1 => n39, B2 => 
                           regs(1743), ZN => n409);
   U536 : NAND3_X1 port map( A1 => n411, A2 => n410, A3 => n409, ZN => 
                           curr_proc_regs(207));
   U537 : NAND2_X1 port map( A1 => regs(720), A2 => n1, ZN => n414);
   U538 : AOI22_X1 port map( A1 => n32, A2 => regs(1232), B1 => n8, B2 => 
                           regs(208), ZN => n413);
   U539 : AOI22_X1 port map( A1 => n11, A2 => regs(2256), B1 => n9, B2 => 
                           regs(1744), ZN => n412);
   U540 : NAND3_X1 port map( A1 => n414, A2 => n413, A3 => n412, ZN => 
                           curr_proc_regs(208));
   U541 : NAND2_X1 port map( A1 => regs(721), A2 => n7, ZN => n417);
   U542 : AOI22_X1 port map( A1 => n32, A2 => regs(1233), B1 => n31, B2 => 
                           regs(209), ZN => n416);
   U543 : AOI22_X1 port map( A1 => n44, A2 => regs(2257), B1 => n9, B2 => 
                           regs(1745), ZN => n415);
   U544 : NAND3_X1 port map( A1 => n417, A2 => n416, A3 => n415, ZN => 
                           curr_proc_regs(209));
   U545 : NAND2_X1 port map( A1 => regs(532), A2 => n7, ZN => n420);
   U546 : AOI22_X1 port map( A1 => n32, A2 => regs(1044), B1 => n31, B2 => 
                           regs(20), ZN => n419);
   U547 : AOI22_X1 port map( A1 => n44, A2 => regs(2068), B1 => n9, B2 => 
                           regs(1556), ZN => n418);
   U548 : NAND3_X1 port map( A1 => n420, A2 => n419, A3 => n418, ZN => 
                           curr_proc_regs(20));
   U549 : NAND2_X1 port map( A1 => regs(722), A2 => n7, ZN => n423);
   U550 : AOI22_X1 port map( A1 => n32, A2 => regs(1234), B1 => n31, B2 => 
                           regs(210), ZN => n422);
   U551 : AOI22_X1 port map( A1 => n44, A2 => regs(2258), B1 => n9, B2 => 
                           regs(1746), ZN => n421);
   U552 : NAND3_X1 port map( A1 => n423, A2 => n422, A3 => n421, ZN => 
                           curr_proc_regs(210));
   U553 : NAND2_X1 port map( A1 => regs(723), A2 => n7, ZN => n426);
   U554 : AOI22_X1 port map( A1 => n32, A2 => regs(1235), B1 => n31, B2 => 
                           regs(211), ZN => n425);
   U555 : AOI22_X1 port map( A1 => n44, A2 => regs(2259), B1 => n9, B2 => 
                           regs(1747), ZN => n424);
   U556 : NAND3_X1 port map( A1 => n426, A2 => n425, A3 => n424, ZN => 
                           curr_proc_regs(211));
   U557 : NAND2_X1 port map( A1 => regs(724), A2 => n7, ZN => n429);
   U558 : AOI22_X1 port map( A1 => n32, A2 => regs(1236), B1 => n31, B2 => 
                           regs(212), ZN => n428);
   U559 : AOI22_X1 port map( A1 => n11, A2 => regs(2260), B1 => n9, B2 => 
                           regs(1748), ZN => n427);
   U560 : NAND3_X1 port map( A1 => n429, A2 => n428, A3 => n427, ZN => 
                           curr_proc_regs(212));
   U561 : NAND2_X1 port map( A1 => regs(725), A2 => n7, ZN => n432);
   U562 : AOI22_X1 port map( A1 => n32, A2 => regs(1237), B1 => n31, B2 => 
                           regs(213), ZN => n431);
   U563 : AOI22_X1 port map( A1 => n11, A2 => regs(2261), B1 => n9, B2 => 
                           regs(1749), ZN => n430);
   U564 : NAND3_X1 port map( A1 => n432, A2 => n431, A3 => n430, ZN => 
                           curr_proc_regs(213));
   U565 : NAND2_X1 port map( A1 => regs(726), A2 => n7, ZN => n435);
   U566 : AOI22_X1 port map( A1 => n32, A2 => regs(1238), B1 => n31, B2 => 
                           regs(214), ZN => n434);
   U567 : AOI22_X1 port map( A1 => n40, A2 => regs(2262), B1 => n9, B2 => 
                           regs(1750), ZN => n433);
   U568 : NAND3_X1 port map( A1 => n435, A2 => n434, A3 => n433, ZN => 
                           curr_proc_regs(214));
   U569 : NAND2_X1 port map( A1 => regs(727), A2 => n7, ZN => n438);
   U570 : AOI22_X1 port map( A1 => n32, A2 => regs(1239), B1 => n31, B2 => 
                           regs(215), ZN => n437);
   U571 : AOI22_X1 port map( A1 => n43, A2 => regs(2263), B1 => n9, B2 => 
                           regs(1751), ZN => n436);
   U572 : NAND3_X1 port map( A1 => n438, A2 => n437, A3 => n436, ZN => 
                           curr_proc_regs(215));
   U573 : NAND2_X1 port map( A1 => regs(728), A2 => n7, ZN => n441);
   U574 : AOI22_X1 port map( A1 => n32, A2 => regs(1240), B1 => n31, B2 => 
                           regs(216), ZN => n440);
   U575 : AOI22_X1 port map( A1 => n12, A2 => regs(2264), B1 => n9, B2 => 
                           regs(1752), ZN => n439);
   U576 : NAND3_X1 port map( A1 => n441, A2 => n440, A3 => n439, ZN => 
                           curr_proc_regs(216));
   U577 : NAND2_X1 port map( A1 => regs(729), A2 => n7, ZN => n444);
   U578 : AOI22_X1 port map( A1 => n32, A2 => regs(1241), B1 => n31, B2 => 
                           regs(217), ZN => n443);
   U579 : AOI22_X1 port map( A1 => n43, A2 => regs(2265), B1 => n9, B2 => 
                           regs(1753), ZN => n442);
   U580 : NAND3_X1 port map( A1 => n444, A2 => n443, A3 => n442, ZN => 
                           curr_proc_regs(217));
   U581 : NAND2_X1 port map( A1 => regs(730), A2 => n7, ZN => n447);
   U582 : AOI22_X1 port map( A1 => n32, A2 => regs(1242), B1 => n31, B2 => 
                           regs(218), ZN => n446);
   U583 : AOI22_X1 port map( A1 => n43, A2 => regs(2266), B1 => n9, B2 => 
                           regs(1754), ZN => n445);
   U584 : NAND3_X1 port map( A1 => n447, A2 => n446, A3 => n445, ZN => 
                           curr_proc_regs(218));
   U585 : NAND2_X1 port map( A1 => regs(731), A2 => n1, ZN => n450);
   U586 : AOI22_X1 port map( A1 => n32, A2 => regs(1243), B1 => n27, B2 => 
                           regs(219), ZN => n449);
   U587 : AOI22_X1 port map( A1 => n12, A2 => regs(2267), B1 => n39, B2 => 
                           regs(1755), ZN => n448);
   U588 : NAND3_X1 port map( A1 => n450, A2 => n449, A3 => n448, ZN => 
                           curr_proc_regs(219));
   U589 : NAND2_X1 port map( A1 => regs(533), A2 => n23, ZN => n453);
   U590 : AOI22_X1 port map( A1 => n32, A2 => regs(1045), B1 => n31, B2 => 
                           regs(21), ZN => n452);
   U591 : AOI22_X1 port map( A1 => n43, A2 => regs(2069), B1 => n39, B2 => 
                           regs(1557), ZN => n451);
   U592 : NAND3_X1 port map( A1 => n453, A2 => n452, A3 => n451, ZN => 
                           curr_proc_regs(21));
   U593 : NAND2_X1 port map( A1 => regs(732), A2 => n17, ZN => n456);
   U594 : AOI22_X1 port map( A1 => n32, A2 => regs(1244), B1 => n31, B2 => 
                           regs(220), ZN => n455);
   U595 : AOI22_X1 port map( A1 => n12, A2 => regs(2268), B1 => n9, B2 => 
                           regs(1756), ZN => n454);
   U596 : NAND3_X1 port map( A1 => n456, A2 => n455, A3 => n454, ZN => 
                           curr_proc_regs(220));
   U597 : NAND2_X1 port map( A1 => regs(733), A2 => n22, ZN => n459);
   U598 : AOI22_X1 port map( A1 => n32, A2 => regs(1245), B1 => n27, B2 => 
                           regs(221), ZN => n458);
   U599 : AOI22_X1 port map( A1 => n12, A2 => regs(2269), B1 => n39, B2 => 
                           regs(1757), ZN => n457);
   U600 : NAND3_X1 port map( A1 => n459, A2 => n458, A3 => n457, ZN => 
                           curr_proc_regs(221));
   U601 : NAND2_X1 port map( A1 => regs(734), A2 => n7, ZN => n462);
   U602 : AOI22_X1 port map( A1 => n32, A2 => regs(1246), B1 => n31, B2 => 
                           regs(222), ZN => n461);
   U603 : AOI22_X1 port map( A1 => n43, A2 => regs(2270), B1 => n39, B2 => 
                           regs(1758), ZN => n460);
   U604 : NAND3_X1 port map( A1 => n462, A2 => n461, A3 => n460, ZN => 
                           curr_proc_regs(222));
   U605 : NAND2_X1 port map( A1 => regs(735), A2 => n1585, ZN => n465);
   U606 : AOI22_X1 port map( A1 => n32, A2 => regs(1247), B1 => n31, B2 => 
                           regs(223), ZN => n464);
   U607 : AOI22_X1 port map( A1 => n12, A2 => regs(2271), B1 => n9, B2 => 
                           regs(1759), ZN => n463);
   U608 : NAND3_X1 port map( A1 => n465, A2 => n464, A3 => n463, ZN => 
                           curr_proc_regs(223));
   U609 : NAND2_X1 port map( A1 => regs(736), A2 => n1585, ZN => n468);
   U610 : AOI22_X1 port map( A1 => n32, A2 => regs(1248), B1 => n27, B2 => 
                           regs(224), ZN => n467);
   U611 : AOI22_X1 port map( A1 => n12, A2 => regs(2272), B1 => n39, B2 => 
                           regs(1760), ZN => n466);
   U612 : NAND3_X1 port map( A1 => n468, A2 => n467, A3 => n466, ZN => 
                           curr_proc_regs(224));
   U613 : NAND2_X1 port map( A1 => regs(737), A2 => n6, ZN => n471);
   U614 : AOI22_X1 port map( A1 => n32, A2 => regs(1249), B1 => n31, B2 => 
                           regs(225), ZN => n470);
   U615 : AOI22_X1 port map( A1 => n12, A2 => regs(2273), B1 => n39, B2 => 
                           regs(1761), ZN => n469);
   U616 : NAND3_X1 port map( A1 => n471, A2 => n470, A3 => n469, ZN => 
                           curr_proc_regs(225));
   U617 : NAND2_X1 port map( A1 => regs(738), A2 => n1585, ZN => n474);
   U618 : AOI22_X1 port map( A1 => n32, A2 => regs(1250), B1 => n31, B2 => 
                           regs(226), ZN => n473);
   U619 : AOI22_X1 port map( A1 => n43, A2 => regs(2274), B1 => n9, B2 => 
                           regs(1762), ZN => n472);
   U620 : NAND3_X1 port map( A1 => n474, A2 => n473, A3 => n472, ZN => 
                           curr_proc_regs(226));
   U621 : NAND2_X1 port map( A1 => regs(739), A2 => n18, ZN => n477);
   U622 : AOI22_X1 port map( A1 => n32, A2 => regs(1251), B1 => n27, B2 => 
                           regs(227), ZN => n476);
   U623 : AOI22_X1 port map( A1 => n43, A2 => regs(2275), B1 => n39, B2 => 
                           regs(1763), ZN => n475);
   U624 : NAND3_X1 port map( A1 => n477, A2 => n476, A3 => n475, ZN => 
                           curr_proc_regs(227));
   U625 : NAND2_X1 port map( A1 => regs(740), A2 => n2, ZN => n480);
   U626 : AOI22_X1 port map( A1 => n32, A2 => regs(1252), B1 => n31, B2 => 
                           regs(228), ZN => n479);
   U627 : AOI22_X1 port map( A1 => n12, A2 => regs(2276), B1 => n39, B2 => 
                           regs(1764), ZN => n478);
   U628 : NAND3_X1 port map( A1 => n480, A2 => n479, A3 => n478, ZN => 
                           curr_proc_regs(228));
   U629 : NAND2_X1 port map( A1 => regs(741), A2 => n19, ZN => n483);
   U630 : AOI22_X1 port map( A1 => n32, A2 => regs(1253), B1 => n27, B2 => 
                           regs(229), ZN => n482);
   U631 : AOI22_X1 port map( A1 => n12, A2 => regs(2277), B1 => n39, B2 => 
                           regs(1765), ZN => n481);
   U632 : NAND3_X1 port map( A1 => n483, A2 => n482, A3 => n481, ZN => 
                           curr_proc_regs(229));
   U633 : NAND2_X1 port map( A1 => regs(534), A2 => n19, ZN => n486);
   U634 : AOI22_X1 port map( A1 => n32, A2 => regs(1046), B1 => n27, B2 => 
                           regs(22), ZN => n485);
   U635 : AOI22_X1 port map( A1 => n43, A2 => regs(2070), B1 => n39, B2 => 
                           regs(1558), ZN => n484);
   U636 : NAND3_X1 port map( A1 => n486, A2 => n485, A3 => n484, ZN => 
                           curr_proc_regs(22));
   U637 : NAND2_X1 port map( A1 => regs(742), A2 => n19, ZN => n489);
   U638 : AOI22_X1 port map( A1 => n32, A2 => regs(1254), B1 => n27, B2 => 
                           regs(230), ZN => n488);
   U639 : AOI22_X1 port map( A1 => n12, A2 => regs(2278), B1 => n39, B2 => 
                           regs(1766), ZN => n487);
   U640 : NAND3_X1 port map( A1 => n489, A2 => n488, A3 => n487, ZN => 
                           curr_proc_regs(230));
   U641 : NAND2_X1 port map( A1 => regs(743), A2 => n19, ZN => n492);
   U642 : AOI22_X1 port map( A1 => n32, A2 => regs(1255), B1 => n27, B2 => 
                           regs(231), ZN => n491);
   U643 : AOI22_X1 port map( A1 => n12, A2 => regs(2279), B1 => n39, B2 => 
                           regs(1767), ZN => n490);
   U644 : NAND3_X1 port map( A1 => n492, A2 => n491, A3 => n490, ZN => 
                           curr_proc_regs(231));
   U645 : NAND2_X1 port map( A1 => regs(744), A2 => n19, ZN => n495);
   U646 : AOI22_X1 port map( A1 => n32, A2 => regs(1256), B1 => n27, B2 => 
                           regs(232), ZN => n494);
   U647 : AOI22_X1 port map( A1 => n43, A2 => regs(2280), B1 => n39, B2 => 
                           regs(1768), ZN => n493);
   U648 : NAND3_X1 port map( A1 => n495, A2 => n494, A3 => n493, ZN => 
                           curr_proc_regs(232));
   U649 : NAND2_X1 port map( A1 => regs(745), A2 => n19, ZN => n498);
   U650 : AOI22_X1 port map( A1 => n32, A2 => regs(1257), B1 => n27, B2 => 
                           regs(233), ZN => n497);
   U651 : AOI22_X1 port map( A1 => n12, A2 => regs(2281), B1 => n39, B2 => 
                           regs(1769), ZN => n496);
   U652 : NAND3_X1 port map( A1 => n498, A2 => n497, A3 => n496, ZN => 
                           curr_proc_regs(233));
   U653 : NAND2_X1 port map( A1 => regs(746), A2 => n19, ZN => n501);
   U654 : AOI22_X1 port map( A1 => n32, A2 => regs(1258), B1 => n27, B2 => 
                           regs(234), ZN => n500);
   U655 : AOI22_X1 port map( A1 => n12, A2 => regs(2282), B1 => n39, B2 => 
                           regs(1770), ZN => n499);
   U656 : NAND3_X1 port map( A1 => n501, A2 => n500, A3 => n499, ZN => 
                           curr_proc_regs(234));
   U657 : NAND2_X1 port map( A1 => regs(747), A2 => n19, ZN => n504);
   U658 : AOI22_X1 port map( A1 => n32, A2 => regs(1259), B1 => n27, B2 => 
                           regs(235), ZN => n503);
   U659 : AOI22_X1 port map( A1 => n12, A2 => regs(2283), B1 => n39, B2 => 
                           regs(1771), ZN => n502);
   U660 : NAND3_X1 port map( A1 => n504, A2 => n503, A3 => n502, ZN => 
                           curr_proc_regs(235));
   U661 : NAND2_X1 port map( A1 => regs(748), A2 => n19, ZN => n507);
   U662 : AOI22_X1 port map( A1 => n32, A2 => regs(1260), B1 => n27, B2 => 
                           regs(236), ZN => n506);
   U663 : AOI22_X1 port map( A1 => n12, A2 => regs(2284), B1 => n39, B2 => 
                           regs(1772), ZN => n505);
   U664 : NAND3_X1 port map( A1 => n507, A2 => n506, A3 => n505, ZN => 
                           curr_proc_regs(236));
   U665 : NAND2_X1 port map( A1 => regs(749), A2 => n19, ZN => n510);
   U666 : AOI22_X1 port map( A1 => n32, A2 => regs(1261), B1 => n27, B2 => 
                           regs(237), ZN => n509);
   U667 : AOI22_X1 port map( A1 => n43, A2 => regs(2285), B1 => n39, B2 => 
                           regs(1773), ZN => n508);
   U668 : NAND3_X1 port map( A1 => n510, A2 => n509, A3 => n508, ZN => 
                           curr_proc_regs(237));
   U669 : NAND2_X1 port map( A1 => regs(750), A2 => n19, ZN => n513);
   U670 : AOI22_X1 port map( A1 => n32, A2 => regs(1262), B1 => n27, B2 => 
                           regs(238), ZN => n512);
   U671 : AOI22_X1 port map( A1 => n43, A2 => regs(2286), B1 => n39, B2 => 
                           regs(1774), ZN => n511);
   U672 : NAND3_X1 port map( A1 => n513, A2 => n512, A3 => n511, ZN => 
                           curr_proc_regs(238));
   U673 : NAND2_X1 port map( A1 => regs(751), A2 => n22, ZN => n516);
   U674 : AOI22_X1 port map( A1 => n32, A2 => regs(1263), B1 => n31, B2 => 
                           regs(239), ZN => n515);
   U675 : AOI22_X1 port map( A1 => n12, A2 => regs(2287), B1 => n39, B2 => 
                           regs(1775), ZN => n514);
   U676 : NAND3_X1 port map( A1 => n516, A2 => n515, A3 => n514, ZN => 
                           curr_proc_regs(239));
   U677 : NAND2_X1 port map( A1 => regs(535), A2 => n22, ZN => n519);
   U678 : AOI22_X1 port map( A1 => n32, A2 => regs(1047), B1 => n31, B2 => 
                           regs(23), ZN => n518);
   U679 : AOI22_X1 port map( A1 => n12, A2 => regs(2071), B1 => n9, B2 => 
                           regs(1559), ZN => n517);
   U680 : NAND3_X1 port map( A1 => n519, A2 => n518, A3 => n517, ZN => 
                           curr_proc_regs(23));
   U681 : NAND2_X1 port map( A1 => regs(752), A2 => n22, ZN => n522);
   U682 : AOI22_X1 port map( A1 => n32, A2 => regs(1264), B1 => n31, B2 => 
                           regs(240), ZN => n521);
   U683 : AOI22_X1 port map( A1 => n12, A2 => regs(2288), B1 => n9, B2 => 
                           regs(1776), ZN => n520);
   U684 : NAND3_X1 port map( A1 => n522, A2 => n521, A3 => n520, ZN => 
                           curr_proc_regs(240));
   U685 : NAND2_X1 port map( A1 => regs(753), A2 => n22, ZN => n525);
   U686 : AOI22_X1 port map( A1 => n32, A2 => regs(1265), B1 => n27, B2 => 
                           regs(241), ZN => n524);
   U687 : AOI22_X1 port map( A1 => n12, A2 => regs(2289), B1 => n39, B2 => 
                           regs(1777), ZN => n523);
   U688 : NAND3_X1 port map( A1 => n525, A2 => n524, A3 => n523, ZN => 
                           curr_proc_regs(241));
   U689 : NAND2_X1 port map( A1 => regs(754), A2 => n22, ZN => n528);
   U690 : AOI22_X1 port map( A1 => n32, A2 => regs(1266), B1 => n31, B2 => 
                           regs(242), ZN => n527);
   U691 : AOI22_X1 port map( A1 => n12, A2 => regs(2290), B1 => n39, B2 => 
                           regs(1778), ZN => n526);
   U692 : NAND3_X1 port map( A1 => n528, A2 => n527, A3 => n526, ZN => 
                           curr_proc_regs(242));
   U693 : NAND2_X1 port map( A1 => regs(755), A2 => n22, ZN => n531);
   U694 : AOI22_X1 port map( A1 => n32, A2 => regs(1267), B1 => n27, B2 => 
                           regs(243), ZN => n530);
   U695 : AOI22_X1 port map( A1 => n12, A2 => regs(2291), B1 => n39, B2 => 
                           regs(1779), ZN => n529);
   U696 : NAND3_X1 port map( A1 => n531, A2 => n530, A3 => n529, ZN => 
                           curr_proc_regs(243));
   U697 : NAND2_X1 port map( A1 => regs(756), A2 => n22, ZN => n534);
   U698 : AOI22_X1 port map( A1 => n32, A2 => regs(1268), B1 => n31, B2 => 
                           regs(244), ZN => n533);
   U699 : AOI22_X1 port map( A1 => n12, A2 => regs(2292), B1 => n9, B2 => 
                           regs(1780), ZN => n532);
   U700 : NAND3_X1 port map( A1 => n534, A2 => n533, A3 => n532, ZN => 
                           curr_proc_regs(244));
   U701 : NAND2_X1 port map( A1 => regs(757), A2 => n22, ZN => n537);
   U702 : AOI22_X1 port map( A1 => n32, A2 => regs(1269), B1 => n27, B2 => 
                           regs(245), ZN => n536);
   U703 : AOI22_X1 port map( A1 => n12, A2 => regs(2293), B1 => n39, B2 => 
                           regs(1781), ZN => n535);
   U704 : NAND3_X1 port map( A1 => n537, A2 => n536, A3 => n535, ZN => 
                           curr_proc_regs(245));
   U705 : NAND2_X1 port map( A1 => regs(758), A2 => n22, ZN => n540);
   U706 : AOI22_X1 port map( A1 => n32, A2 => regs(1270), B1 => n31, B2 => 
                           regs(246), ZN => n539);
   U707 : AOI22_X1 port map( A1 => n12, A2 => regs(2294), B1 => n39, B2 => 
                           regs(1782), ZN => n538);
   U708 : NAND3_X1 port map( A1 => n540, A2 => n539, A3 => n538, ZN => 
                           curr_proc_regs(246));
   U709 : NAND2_X1 port map( A1 => regs(759), A2 => n22, ZN => n543);
   U710 : AOI22_X1 port map( A1 => n32, A2 => regs(1271), B1 => n31, B2 => 
                           regs(247), ZN => n542);
   U711 : AOI22_X1 port map( A1 => n12, A2 => regs(2295), B1 => n39, B2 => 
                           regs(1783), ZN => n541);
   U712 : NAND3_X1 port map( A1 => n543, A2 => n542, A3 => n541, ZN => 
                           curr_proc_regs(247));
   U713 : NAND2_X1 port map( A1 => regs(760), A2 => n22, ZN => n546);
   U714 : AOI22_X1 port map( A1 => n32, A2 => regs(1272), B1 => n31, B2 => 
                           regs(248), ZN => n545);
   U715 : AOI22_X1 port map( A1 => n12, A2 => regs(2296), B1 => n9, B2 => 
                           regs(1784), ZN => n544);
   U716 : NAND3_X1 port map( A1 => n546, A2 => n545, A3 => n544, ZN => 
                           curr_proc_regs(248));
   U717 : NAND2_X1 port map( A1 => regs(761), A2 => n23, ZN => n549);
   U718 : AOI22_X1 port map( A1 => n32, A2 => regs(1273), B1 => n27, B2 => 
                           regs(249), ZN => n548);
   U719 : AOI22_X1 port map( A1 => n12, A2 => regs(2297), B1 => n39, B2 => 
                           regs(1785), ZN => n547);
   U720 : NAND3_X1 port map( A1 => n549, A2 => n548, A3 => n547, ZN => 
                           curr_proc_regs(249));
   U721 : NAND2_X1 port map( A1 => regs(536), A2 => n23, ZN => n552);
   U722 : AOI22_X1 port map( A1 => n32, A2 => regs(1048), B1 => n31, B2 => 
                           regs(24), ZN => n551);
   U723 : AOI22_X1 port map( A1 => n12, A2 => regs(2072), B1 => n9, B2 => 
                           regs(1560), ZN => n550);
   U724 : NAND3_X1 port map( A1 => n552, A2 => n551, A3 => n550, ZN => 
                           curr_proc_regs(24));
   U725 : NAND2_X1 port map( A1 => regs(762), A2 => n23, ZN => n555);
   U726 : AOI22_X1 port map( A1 => n32, A2 => regs(1274), B1 => n31, B2 => 
                           regs(250), ZN => n554);
   U727 : AOI22_X1 port map( A1 => n12, A2 => regs(2298), B1 => n9, B2 => 
                           regs(1786), ZN => n553);
   U728 : NAND3_X1 port map( A1 => n555, A2 => n554, A3 => n553, ZN => 
                           curr_proc_regs(250));
   U729 : NAND2_X1 port map( A1 => regs(763), A2 => n23, ZN => n558);
   U730 : AOI22_X1 port map( A1 => n32, A2 => regs(1275), B1 => n27, B2 => 
                           regs(251), ZN => n557);
   U731 : AOI22_X1 port map( A1 => n12, A2 => regs(2299), B1 => n39, B2 => 
                           regs(1787), ZN => n556);
   U732 : NAND3_X1 port map( A1 => n558, A2 => n557, A3 => n556, ZN => 
                           curr_proc_regs(251));
   U733 : NAND2_X1 port map( A1 => regs(764), A2 => n23, ZN => n561);
   U734 : AOI22_X1 port map( A1 => n32, A2 => regs(1276), B1 => n31, B2 => 
                           regs(252), ZN => n560);
   U735 : AOI22_X1 port map( A1 => n12, A2 => regs(2300), B1 => n39, B2 => 
                           regs(1788), ZN => n559);
   U736 : NAND3_X1 port map( A1 => n561, A2 => n560, A3 => n559, ZN => 
                           curr_proc_regs(252));
   U737 : NAND2_X1 port map( A1 => regs(765), A2 => n23, ZN => n564);
   U738 : AOI22_X1 port map( A1 => n32, A2 => regs(1277), B1 => n31, B2 => 
                           regs(253), ZN => n563);
   U739 : AOI22_X1 port map( A1 => n12, A2 => regs(2301), B1 => n39, B2 => 
                           regs(1789), ZN => n562);
   U740 : NAND3_X1 port map( A1 => n564, A2 => n563, A3 => n562, ZN => 
                           curr_proc_regs(253));
   U741 : NAND2_X1 port map( A1 => regs(766), A2 => n23, ZN => n567);
   U742 : AOI22_X1 port map( A1 => n32, A2 => regs(1278), B1 => n27, B2 => 
                           regs(254), ZN => n566);
   U743 : AOI22_X1 port map( A1 => n12, A2 => regs(2302), B1 => n39, B2 => 
                           regs(1790), ZN => n565);
   U744 : NAND3_X1 port map( A1 => n567, A2 => n566, A3 => n565, ZN => 
                           curr_proc_regs(254));
   U745 : NAND2_X1 port map( A1 => regs(767), A2 => n23, ZN => n570);
   U746 : AOI22_X1 port map( A1 => n32, A2 => regs(1279), B1 => n31, B2 => 
                           regs(255), ZN => n569);
   U747 : AOI22_X1 port map( A1 => n12, A2 => regs(2303), B1 => n9, B2 => 
                           regs(1791), ZN => n568);
   U748 : NAND3_X1 port map( A1 => n570, A2 => n569, A3 => n568, ZN => 
                           curr_proc_regs(255));
   U749 : NAND2_X1 port map( A1 => regs(768), A2 => n23, ZN => n573);
   U750 : AOI22_X1 port map( A1 => n32, A2 => regs(1280), B1 => n31, B2 => 
                           regs(256), ZN => n572);
   U751 : AOI22_X1 port map( A1 => n12, A2 => regs(2304), B1 => n39, B2 => 
                           regs(1792), ZN => n571);
   U752 : NAND3_X1 port map( A1 => n573, A2 => n572, A3 => n571, ZN => 
                           curr_proc_regs(256));
   U753 : NAND2_X1 port map( A1 => regs(769), A2 => n23, ZN => n576);
   U754 : AOI22_X1 port map( A1 => n32, A2 => regs(1281), B1 => n31, B2 => 
                           regs(257), ZN => n575);
   U755 : AOI22_X1 port map( A1 => n12, A2 => regs(2305), B1 => n39, B2 => 
                           regs(1793), ZN => n574);
   U756 : NAND3_X1 port map( A1 => n576, A2 => n575, A3 => n574, ZN => 
                           curr_proc_regs(257));
   U757 : NAND2_X1 port map( A1 => regs(770), A2 => n23, ZN => n579);
   U758 : AOI22_X1 port map( A1 => n32, A2 => regs(1282), B1 => n31, B2 => 
                           regs(258), ZN => n578);
   U759 : AOI22_X1 port map( A1 => n12, A2 => regs(2306), B1 => n39, B2 => 
                           regs(1794), ZN => n577);
   U760 : NAND3_X1 port map( A1 => n579, A2 => n578, A3 => n577, ZN => 
                           curr_proc_regs(258));
   U761 : NAND2_X1 port map( A1 => regs(771), A2 => n7, ZN => n582);
   U762 : AOI22_X1 port map( A1 => n32, A2 => regs(1283), B1 => n27, B2 => 
                           regs(259), ZN => n581);
   U763 : AOI22_X1 port map( A1 => n12, A2 => regs(2307), B1 => n39, B2 => 
                           regs(1795), ZN => n580);
   U764 : NAND3_X1 port map( A1 => n582, A2 => n581, A3 => n580, ZN => 
                           curr_proc_regs(259));
   U765 : NAND2_X1 port map( A1 => regs(537), A2 => n7, ZN => n585);
   U766 : AOI22_X1 port map( A1 => n32, A2 => regs(1049), B1 => n31, B2 => 
                           regs(25), ZN => n584);
   U767 : AOI22_X1 port map( A1 => n12, A2 => regs(2073), B1 => n39, B2 => 
                           regs(1561), ZN => n583);
   U768 : NAND3_X1 port map( A1 => n585, A2 => n584, A3 => n583, ZN => 
                           curr_proc_regs(25));
   U769 : NAND2_X1 port map( A1 => regs(772), A2 => n7, ZN => n588);
   U770 : AOI22_X1 port map( A1 => n32, A2 => regs(1284), B1 => n31, B2 => 
                           regs(260), ZN => n587);
   U771 : AOI22_X1 port map( A1 => n12, A2 => regs(2308), B1 => n39, B2 => 
                           regs(1796), ZN => n586);
   U772 : NAND3_X1 port map( A1 => n588, A2 => n587, A3 => n586, ZN => 
                           curr_proc_regs(260));
   U773 : NAND2_X1 port map( A1 => regs(773), A2 => n7, ZN => n591);
   U774 : AOI22_X1 port map( A1 => n32, A2 => regs(1285), B1 => n31, B2 => 
                           regs(261), ZN => n590);
   U775 : AOI22_X1 port map( A1 => n43, A2 => regs(2309), B1 => n39, B2 => 
                           regs(1797), ZN => n589);
   U776 : NAND3_X1 port map( A1 => n591, A2 => n590, A3 => n589, ZN => 
                           curr_proc_regs(261));
   U777 : NAND2_X1 port map( A1 => regs(774), A2 => n7, ZN => n594);
   U778 : AOI22_X1 port map( A1 => n32, A2 => regs(1286), B1 => n31, B2 => 
                           regs(262), ZN => n593);
   U779 : AOI22_X1 port map( A1 => n43, A2 => regs(2310), B1 => n39, B2 => 
                           regs(1798), ZN => n592);
   U780 : NAND3_X1 port map( A1 => n594, A2 => n593, A3 => n592, ZN => 
                           curr_proc_regs(262));
   U781 : NAND2_X1 port map( A1 => regs(775), A2 => n7, ZN => n597);
   U782 : AOI22_X1 port map( A1 => n32, A2 => regs(1287), B1 => n31, B2 => 
                           regs(263), ZN => n596);
   U783 : AOI22_X1 port map( A1 => n43, A2 => regs(2311), B1 => n9, B2 => 
                           regs(1799), ZN => n595);
   U784 : NAND3_X1 port map( A1 => n597, A2 => n596, A3 => n595, ZN => 
                           curr_proc_regs(263));
   U785 : NAND2_X1 port map( A1 => regs(776), A2 => n7, ZN => n600);
   U786 : AOI22_X1 port map( A1 => n32, A2 => regs(1288), B1 => n27, B2 => 
                           regs(264), ZN => n599);
   U787 : AOI22_X1 port map( A1 => n43, A2 => regs(2312), B1 => n39, B2 => 
                           regs(1800), ZN => n598);
   U788 : NAND3_X1 port map( A1 => n600, A2 => n599, A3 => n598, ZN => 
                           curr_proc_regs(264));
   U789 : NAND2_X1 port map( A1 => regs(777), A2 => n7, ZN => n603);
   U790 : AOI22_X1 port map( A1 => n32, A2 => regs(1289), B1 => n31, B2 => 
                           regs(265), ZN => n602);
   U791 : AOI22_X1 port map( A1 => n43, A2 => regs(2313), B1 => n39, B2 => 
                           regs(1801), ZN => n601);
   U792 : NAND3_X1 port map( A1 => n603, A2 => n602, A3 => n601, ZN => 
                           curr_proc_regs(265));
   U793 : NAND2_X1 port map( A1 => regs(778), A2 => n7, ZN => n606);
   U794 : AOI22_X1 port map( A1 => n32, A2 => regs(1290), B1 => n31, B2 => 
                           regs(266), ZN => n605);
   U795 : AOI22_X1 port map( A1 => n43, A2 => regs(2314), B1 => n39, B2 => 
                           regs(1802), ZN => n604);
   U796 : NAND3_X1 port map( A1 => n606, A2 => n605, A3 => n604, ZN => 
                           curr_proc_regs(266));
   U797 : NAND2_X1 port map( A1 => regs(779), A2 => n7, ZN => n609);
   U798 : AOI22_X1 port map( A1 => n32, A2 => regs(1291), B1 => n31, B2 => 
                           regs(267), ZN => n608);
   U799 : AOI22_X1 port map( A1 => n12, A2 => regs(2315), B1 => n39, B2 => 
                           regs(1803), ZN => n607);
   U800 : NAND3_X1 port map( A1 => n609, A2 => n608, A3 => n607, ZN => 
                           curr_proc_regs(267));
   U801 : NAND2_X1 port map( A1 => regs(780), A2 => n7, ZN => n612);
   U802 : AOI22_X1 port map( A1 => n32, A2 => regs(1292), B1 => n31, B2 => 
                           regs(268), ZN => n611);
   U803 : AOI22_X1 port map( A1 => n43, A2 => regs(2316), B1 => n39, B2 => 
                           regs(1804), ZN => n610);
   U804 : NAND3_X1 port map( A1 => n612, A2 => n611, A3 => n610, ZN => 
                           curr_proc_regs(268));
   U805 : NAND2_X1 port map( A1 => regs(781), A2 => n6, ZN => n615);
   U806 : AOI22_X1 port map( A1 => n32, A2 => regs(1293), B1 => n25, B2 => 
                           regs(269), ZN => n614);
   U807 : AOI22_X1 port map( A1 => n43, A2 => regs(2317), B1 => n1588, B2 => 
                           regs(1805), ZN => n613);
   U808 : NAND3_X1 port map( A1 => n615, A2 => n614, A3 => n613, ZN => 
                           curr_proc_regs(269));
   U809 : NAND2_X1 port map( A1 => regs(538), A2 => n6, ZN => n618);
   U810 : AOI22_X1 port map( A1 => n32, A2 => regs(1050), B1 => n1586, B2 => 
                           regs(26), ZN => n617);
   U811 : AOI22_X1 port map( A1 => n12, A2 => regs(2074), B1 => n1588, B2 => 
                           regs(1562), ZN => n616);
   U812 : NAND3_X1 port map( A1 => n618, A2 => n617, A3 => n616, ZN => 
                           curr_proc_regs(26));
   U813 : NAND2_X1 port map( A1 => regs(782), A2 => n6, ZN => n621);
   U814 : AOI22_X1 port map( A1 => n32, A2 => regs(1294), B1 => n1586, B2 => 
                           regs(270), ZN => n620);
   U815 : AOI22_X1 port map( A1 => n13, A2 => regs(2318), B1 => n1588, B2 => 
                           regs(1806), ZN => n619);
   U816 : NAND3_X1 port map( A1 => n621, A2 => n620, A3 => n619, ZN => 
                           curr_proc_regs(270));
   U817 : NAND2_X1 port map( A1 => regs(783), A2 => n6, ZN => n624);
   U818 : AOI22_X1 port map( A1 => n32, A2 => regs(1295), B1 => n1586, B2 => 
                           regs(271), ZN => n623);
   U819 : AOI22_X1 port map( A1 => n43, A2 => regs(2319), B1 => n34, B2 => 
                           regs(1807), ZN => n622);
   U820 : NAND3_X1 port map( A1 => n624, A2 => n623, A3 => n622, ZN => 
                           curr_proc_regs(271));
   U821 : NAND2_X1 port map( A1 => regs(784), A2 => n6, ZN => n627);
   U822 : AOI22_X1 port map( A1 => n32, A2 => regs(1296), B1 => n1586, B2 => 
                           regs(272), ZN => n626);
   U823 : AOI22_X1 port map( A1 => n13, A2 => regs(2320), B1 => n35, B2 => 
                           regs(1808), ZN => n625);
   U824 : NAND3_X1 port map( A1 => n627, A2 => n626, A3 => n625, ZN => 
                           curr_proc_regs(272));
   U825 : NAND2_X1 port map( A1 => regs(785), A2 => n6, ZN => n630);
   U826 : AOI22_X1 port map( A1 => n32, A2 => regs(1297), B1 => n1586, B2 => 
                           regs(273), ZN => n629);
   U827 : AOI22_X1 port map( A1 => n13, A2 => regs(2321), B1 => n34, B2 => 
                           regs(1809), ZN => n628);
   U828 : NAND3_X1 port map( A1 => n630, A2 => n629, A3 => n628, ZN => 
                           curr_proc_regs(273));
   U829 : NAND2_X1 port map( A1 => regs(786), A2 => n6, ZN => n633);
   U830 : AOI22_X1 port map( A1 => n32, A2 => regs(1298), B1 => n30, B2 => 
                           regs(274), ZN => n632);
   U831 : AOI22_X1 port map( A1 => n13, A2 => regs(2322), B1 => n36, B2 => 
                           regs(1810), ZN => n631);
   U832 : NAND3_X1 port map( A1 => n633, A2 => n632, A3 => n631, ZN => 
                           curr_proc_regs(274));
   U833 : NAND2_X1 port map( A1 => regs(787), A2 => n6, ZN => n636);
   U834 : AOI22_X1 port map( A1 => n32, A2 => regs(1299), B1 => n30, B2 => 
                           regs(275), ZN => n635);
   U835 : AOI22_X1 port map( A1 => n13, A2 => regs(2323), B1 => n36, B2 => 
                           regs(1811), ZN => n634);
   U836 : NAND3_X1 port map( A1 => n636, A2 => n635, A3 => n634, ZN => 
                           curr_proc_regs(275));
   U837 : NAND2_X1 port map( A1 => regs(788), A2 => n6, ZN => n639);
   U838 : AOI22_X1 port map( A1 => n32, A2 => regs(1300), B1 => n30, B2 => 
                           regs(276), ZN => n638);
   U839 : AOI22_X1 port map( A1 => n13, A2 => regs(2324), B1 => n36, B2 => 
                           regs(1812), ZN => n637);
   U840 : NAND3_X1 port map( A1 => n639, A2 => n638, A3 => n637, ZN => 
                           curr_proc_regs(276));
   U841 : NAND2_X1 port map( A1 => regs(789), A2 => n6, ZN => n642);
   U842 : AOI22_X1 port map( A1 => n32, A2 => regs(1301), B1 => n30, B2 => 
                           regs(277), ZN => n641);
   U843 : AOI22_X1 port map( A1 => n13, A2 => regs(2325), B1 => n36, B2 => 
                           regs(1813), ZN => n640);
   U844 : NAND3_X1 port map( A1 => n642, A2 => n641, A3 => n640, ZN => 
                           curr_proc_regs(277));
   U845 : NAND2_X1 port map( A1 => regs(790), A2 => n6, ZN => n645);
   U846 : AOI22_X1 port map( A1 => n32, A2 => regs(1302), B1 => n30, B2 => 
                           regs(278), ZN => n644);
   U847 : AOI22_X1 port map( A1 => n13, A2 => regs(2326), B1 => n36, B2 => 
                           regs(1814), ZN => n643);
   U848 : NAND3_X1 port map( A1 => n645, A2 => n644, A3 => n643, ZN => 
                           curr_proc_regs(278));
   U849 : NAND2_X1 port map( A1 => regs(791), A2 => n6, ZN => n648);
   U850 : AOI22_X1 port map( A1 => n32, A2 => regs(1303), B1 => n30, B2 => 
                           regs(279), ZN => n647);
   U851 : AOI22_X1 port map( A1 => n13, A2 => regs(2327), B1 => n36, B2 => 
                           regs(1815), ZN => n646);
   U852 : NAND3_X1 port map( A1 => n648, A2 => n647, A3 => n646, ZN => 
                           curr_proc_regs(279));
   U853 : NAND2_X1 port map( A1 => regs(539), A2 => n2, ZN => n651);
   U854 : AOI22_X1 port map( A1 => n32, A2 => regs(1051), B1 => n30, B2 => 
                           regs(27), ZN => n650);
   U855 : AOI22_X1 port map( A1 => n13, A2 => regs(2075), B1 => n36, B2 => 
                           regs(1563), ZN => n649);
   U856 : NAND3_X1 port map( A1 => n651, A2 => n650, A3 => n649, ZN => 
                           curr_proc_regs(27));
   U857 : NAND2_X1 port map( A1 => regs(792), A2 => n6, ZN => n654);
   U858 : AOI22_X1 port map( A1 => n32, A2 => regs(1304), B1 => n3, B2 => 
                           regs(280), ZN => n653);
   U859 : AOI22_X1 port map( A1 => n5, A2 => regs(2328), B1 => n37, B2 => 
                           regs(1816), ZN => n652);
   U860 : NAND3_X1 port map( A1 => n654, A2 => n653, A3 => n652, ZN => 
                           curr_proc_regs(280));
   U861 : NAND2_X1 port map( A1 => regs(793), A2 => n2, ZN => n657);
   U862 : AOI22_X1 port map( A1 => n32, A2 => regs(1305), B1 => n30, B2 => 
                           regs(281), ZN => n656);
   U863 : AOI22_X1 port map( A1 => n5, A2 => regs(2329), B1 => n36, B2 => 
                           regs(1817), ZN => n655);
   U864 : NAND3_X1 port map( A1 => n657, A2 => n656, A3 => n655, ZN => 
                           curr_proc_regs(281));
   U865 : NAND2_X1 port map( A1 => regs(794), A2 => n6, ZN => n660);
   U866 : AOI22_X1 port map( A1 => n32, A2 => regs(1306), B1 => n30, B2 => 
                           regs(282), ZN => n659);
   U867 : AOI22_X1 port map( A1 => n5, A2 => regs(2330), B1 => n36, B2 => 
                           regs(1818), ZN => n658);
   U868 : NAND3_X1 port map( A1 => n660, A2 => n659, A3 => n658, ZN => 
                           curr_proc_regs(282));
   U869 : NAND2_X1 port map( A1 => regs(795), A2 => n2, ZN => n663);
   U870 : AOI22_X1 port map( A1 => n32, A2 => regs(1307), B1 => n1586, B2 => 
                           regs(283), ZN => n662);
   U871 : AOI22_X1 port map( A1 => n13, A2 => regs(2331), B1 => n35, B2 => 
                           regs(1819), ZN => n661);
   U872 : NAND3_X1 port map( A1 => n663, A2 => n662, A3 => n661, ZN => 
                           curr_proc_regs(283));
   U873 : NAND2_X1 port map( A1 => regs(796), A2 => n6, ZN => n666);
   U874 : AOI22_X1 port map( A1 => n32, A2 => regs(1308), B1 => n30, B2 => 
                           regs(284), ZN => n665);
   U875 : AOI22_X1 port map( A1 => n13, A2 => regs(2332), B1 => n36, B2 => 
                           regs(1820), ZN => n664);
   U876 : NAND3_X1 port map( A1 => n666, A2 => n665, A3 => n664, ZN => 
                           curr_proc_regs(284));
   U877 : NAND2_X1 port map( A1 => regs(797), A2 => n2, ZN => n669);
   U878 : AOI22_X1 port map( A1 => n32, A2 => regs(1309), B1 => n30, B2 => 
                           regs(285), ZN => n668);
   U879 : AOI22_X1 port map( A1 => n5, A2 => regs(2333), B1 => n36, B2 => 
                           regs(1821), ZN => n667);
   U880 : NAND3_X1 port map( A1 => n669, A2 => n668, A3 => n667, ZN => 
                           curr_proc_regs(285));
   U881 : NAND2_X1 port map( A1 => regs(798), A2 => n6, ZN => n672);
   U882 : AOI22_X1 port map( A1 => n32, A2 => regs(1310), B1 => n3, B2 => 
                           regs(286), ZN => n671);
   U883 : AOI22_X1 port map( A1 => n5, A2 => regs(2334), B1 => n34, B2 => 
                           regs(1822), ZN => n670);
   U884 : NAND3_X1 port map( A1 => n672, A2 => n671, A3 => n670, ZN => 
                           curr_proc_regs(286));
   U885 : NAND2_X1 port map( A1 => regs(799), A2 => n2, ZN => n675);
   U886 : AOI22_X1 port map( A1 => n32, A2 => regs(1311), B1 => n30, B2 => 
                           regs(287), ZN => n674);
   U887 : AOI22_X1 port map( A1 => n13, A2 => regs(2335), B1 => n36, B2 => 
                           regs(1823), ZN => n673);
   U888 : NAND3_X1 port map( A1 => n675, A2 => n674, A3 => n673, ZN => 
                           curr_proc_regs(287));
   U889 : NAND2_X1 port map( A1 => regs(800), A2 => n6, ZN => n678);
   U890 : AOI22_X1 port map( A1 => n32, A2 => regs(1312), B1 => n30, B2 => 
                           regs(288), ZN => n677);
   U891 : AOI22_X1 port map( A1 => n13, A2 => regs(2336), B1 => n36, B2 => 
                           regs(1824), ZN => n676);
   U892 : NAND3_X1 port map( A1 => n678, A2 => n677, A3 => n676, ZN => 
                           curr_proc_regs(288));
   U893 : NAND2_X1 port map( A1 => regs(801), A2 => n17, ZN => n681);
   U894 : AOI22_X1 port map( A1 => n32, A2 => regs(1313), B1 => n30, B2 => 
                           regs(289), ZN => n680);
   U895 : AOI22_X1 port map( A1 => n13, A2 => regs(2337), B1 => n36, B2 => 
                           regs(1825), ZN => n679);
   U896 : NAND3_X1 port map( A1 => n681, A2 => n680, A3 => n679, ZN => 
                           curr_proc_regs(289));
   U897 : NAND2_X1 port map( A1 => regs(540), A2 => n22, ZN => n684);
   U898 : AOI22_X1 port map( A1 => n32, A2 => regs(1052), B1 => n30, B2 => 
                           regs(28), ZN => n683);
   U899 : AOI22_X1 port map( A1 => n13, A2 => regs(2076), B1 => n36, B2 => 
                           regs(1564), ZN => n682);
   U900 : NAND3_X1 port map( A1 => n684, A2 => n683, A3 => n682, ZN => 
                           curr_proc_regs(28));
   U901 : NAND2_X1 port map( A1 => regs(802), A2 => n7, ZN => n687);
   U902 : AOI22_X1 port map( A1 => n32, A2 => regs(1314), B1 => n30, B2 => 
                           regs(290), ZN => n686);
   U903 : AOI22_X1 port map( A1 => n13, A2 => regs(2338), B1 => n36, B2 => 
                           regs(1826), ZN => n685);
   U904 : NAND3_X1 port map( A1 => n687, A2 => n686, A3 => n685, ZN => 
                           curr_proc_regs(290));
   U905 : NAND2_X1 port map( A1 => regs(803), A2 => n22, ZN => n690);
   U906 : AOI22_X1 port map( A1 => n32, A2 => regs(1315), B1 => n30, B2 => 
                           regs(291), ZN => n689);
   U907 : AOI22_X1 port map( A1 => n5, A2 => regs(2339), B1 => n36, B2 => 
                           regs(1827), ZN => n688);
   U908 : NAND3_X1 port map( A1 => n690, A2 => n689, A3 => n688, ZN => 
                           curr_proc_regs(291));
   U909 : NAND2_X1 port map( A1 => regs(804), A2 => n6, ZN => n693);
   U910 : AOI22_X1 port map( A1 => n32, A2 => regs(1316), B1 => n30, B2 => 
                           regs(292), ZN => n692);
   U911 : AOI22_X1 port map( A1 => n5, A2 => regs(2340), B1 => n36, B2 => 
                           regs(1828), ZN => n691);
   U912 : NAND3_X1 port map( A1 => n693, A2 => n692, A3 => n691, ZN => 
                           curr_proc_regs(292));
   U913 : NAND2_X1 port map( A1 => regs(805), A2 => n22, ZN => n696);
   U914 : AOI22_X1 port map( A1 => n32, A2 => regs(1317), B1 => n30, B2 => 
                           regs(293), ZN => n695);
   U915 : AOI22_X1 port map( A1 => n13, A2 => regs(2341), B1 => n36, B2 => 
                           regs(1829), ZN => n694);
   U916 : NAND3_X1 port map( A1 => n696, A2 => n695, A3 => n694, ZN => 
                           curr_proc_regs(293));
   U917 : NAND2_X1 port map( A1 => regs(806), A2 => n18, ZN => n699);
   U918 : AOI22_X1 port map( A1 => n32, A2 => regs(1318), B1 => n30, B2 => 
                           regs(294), ZN => n698);
   U919 : AOI22_X1 port map( A1 => n13, A2 => regs(2342), B1 => n36, B2 => 
                           regs(1830), ZN => n697);
   U920 : NAND3_X1 port map( A1 => n699, A2 => n698, A3 => n697, ZN => 
                           curr_proc_regs(294));
   U921 : NAND2_X1 port map( A1 => regs(807), A2 => n22, ZN => n702);
   U922 : AOI22_X1 port map( A1 => n32, A2 => regs(1319), B1 => n30, B2 => 
                           regs(295), ZN => n701);
   U923 : AOI22_X1 port map( A1 => n13, A2 => regs(2343), B1 => n36, B2 => 
                           regs(1831), ZN => n700);
   U924 : NAND3_X1 port map( A1 => n702, A2 => n701, A3 => n700, ZN => 
                           curr_proc_regs(295));
   U925 : NAND2_X1 port map( A1 => regs(808), A2 => n2, ZN => n705);
   U926 : AOI22_X1 port map( A1 => n32, A2 => regs(1320), B1 => n30, B2 => 
                           regs(296), ZN => n704);
   U927 : AOI22_X1 port map( A1 => n5, A2 => regs(2344), B1 => n36, B2 => 
                           regs(1832), ZN => n703);
   U928 : NAND3_X1 port map( A1 => n705, A2 => n704, A3 => n703, ZN => 
                           curr_proc_regs(296));
   U929 : NAND2_X1 port map( A1 => regs(809), A2 => n22, ZN => n708);
   U930 : AOI22_X1 port map( A1 => n32, A2 => regs(1321), B1 => n30, B2 => 
                           regs(297), ZN => n707);
   U931 : AOI22_X1 port map( A1 => n13, A2 => regs(2345), B1 => n36, B2 => 
                           regs(1833), ZN => n706);
   U932 : NAND3_X1 port map( A1 => n708, A2 => n707, A3 => n706, ZN => 
                           curr_proc_regs(297));
   U933 : NAND2_X1 port map( A1 => regs(810), A2 => n22, ZN => n711);
   U934 : AOI22_X1 port map( A1 => n32, A2 => regs(1322), B1 => n30, B2 => 
                           regs(298), ZN => n710);
   U935 : AOI22_X1 port map( A1 => n13, A2 => regs(2346), B1 => n36, B2 => 
                           regs(1834), ZN => n709);
   U936 : NAND3_X1 port map( A1 => n711, A2 => n710, A3 => n709, ZN => 
                           curr_proc_regs(298));
   U937 : NAND2_X1 port map( A1 => regs(811), A2 => n7, ZN => n714);
   U938 : AOI22_X1 port map( A1 => n32, A2 => regs(1323), B1 => n30, B2 => 
                           regs(299), ZN => n713);
   U939 : AOI22_X1 port map( A1 => n13, A2 => regs(2347), B1 => n36, B2 => 
                           regs(1835), ZN => n712);
   U940 : NAND3_X1 port map( A1 => n714, A2 => n713, A3 => n712, ZN => 
                           curr_proc_regs(299));
   U941 : NAND2_X1 port map( A1 => regs(541), A2 => n7, ZN => n717);
   U942 : AOI22_X1 port map( A1 => n32, A2 => regs(1053), B1 => n8, B2 => 
                           regs(29), ZN => n716);
   U943 : AOI22_X1 port map( A1 => n5, A2 => regs(2077), B1 => n35, B2 => 
                           regs(1565), ZN => n715);
   U944 : NAND3_X1 port map( A1 => n717, A2 => n716, A3 => n715, ZN => 
                           curr_proc_regs(29));
   U945 : NAND2_X1 port map( A1 => regs(514), A2 => n7, ZN => n720);
   U946 : AOI22_X1 port map( A1 => n32, A2 => regs(1026), B1 => n1586, B2 => 
                           regs(2), ZN => n719);
   U947 : AOI22_X1 port map( A1 => n5, A2 => regs(2050), B1 => n4, B2 => 
                           regs(1538), ZN => n718);
   U948 : NAND3_X1 port map( A1 => n720, A2 => n719, A3 => n718, ZN => 
                           curr_proc_regs(2));
   U949 : NAND2_X1 port map( A1 => regs(812), A2 => n7, ZN => n723);
   U950 : AOI22_X1 port map( A1 => n32, A2 => regs(1324), B1 => n30, B2 => 
                           regs(300), ZN => n722);
   U951 : AOI22_X1 port map( A1 => n13, A2 => regs(2348), B1 => n36, B2 => 
                           regs(1836), ZN => n721);
   U952 : NAND3_X1 port map( A1 => n723, A2 => n722, A3 => n721, ZN => 
                           curr_proc_regs(300));
   U953 : NAND2_X1 port map( A1 => regs(813), A2 => n7, ZN => n726);
   U954 : AOI22_X1 port map( A1 => n32, A2 => regs(1325), B1 => n30, B2 => 
                           regs(301), ZN => n725);
   U955 : AOI22_X1 port map( A1 => n13, A2 => regs(2349), B1 => n36, B2 => 
                           regs(1837), ZN => n724);
   U956 : NAND3_X1 port map( A1 => n726, A2 => n725, A3 => n724, ZN => 
                           curr_proc_regs(301));
   U957 : NAND2_X1 port map( A1 => regs(814), A2 => n7, ZN => n729);
   U958 : AOI22_X1 port map( A1 => n32, A2 => regs(1326), B1 => n30, B2 => 
                           regs(302), ZN => n728);
   U959 : AOI22_X1 port map( A1 => n5, A2 => regs(2350), B1 => n36, B2 => 
                           regs(1838), ZN => n727);
   U960 : NAND3_X1 port map( A1 => n729, A2 => n728, A3 => n727, ZN => 
                           curr_proc_regs(302));
   U961 : NAND2_X1 port map( A1 => regs(815), A2 => n7, ZN => n732);
   U962 : AOI22_X1 port map( A1 => n32, A2 => regs(1327), B1 => n26, B2 => 
                           regs(303), ZN => n731);
   U963 : AOI22_X1 port map( A1 => n13, A2 => regs(2351), B1 => n4, B2 => 
                           regs(1839), ZN => n730);
   U964 : NAND3_X1 port map( A1 => n732, A2 => n731, A3 => n730, ZN => 
                           curr_proc_regs(303));
   U965 : NAND2_X1 port map( A1 => regs(816), A2 => n7, ZN => n735);
   U966 : AOI22_X1 port map( A1 => n32, A2 => regs(1328), B1 => n30, B2 => 
                           regs(304), ZN => n734);
   U967 : AOI22_X1 port map( A1 => n13, A2 => regs(2352), B1 => n36, B2 => 
                           regs(1840), ZN => n733);
   U968 : NAND3_X1 port map( A1 => n735, A2 => n734, A3 => n733, ZN => 
                           curr_proc_regs(304));
   U969 : NAND2_X1 port map( A1 => regs(817), A2 => n7, ZN => n738);
   U970 : AOI22_X1 port map( A1 => n32, A2 => regs(1329), B1 => n30, B2 => 
                           regs(305), ZN => n737);
   U971 : AOI22_X1 port map( A1 => n5, A2 => regs(2353), B1 => n36, B2 => 
                           regs(1841), ZN => n736);
   U972 : NAND3_X1 port map( A1 => n738, A2 => n737, A3 => n736, ZN => 
                           curr_proc_regs(305));
   U973 : NAND2_X1 port map( A1 => regs(818), A2 => n7, ZN => n741);
   U974 : AOI22_X1 port map( A1 => n32, A2 => regs(1330), B1 => n30, B2 => 
                           regs(306), ZN => n740);
   U975 : AOI22_X1 port map( A1 => n13, A2 => regs(2354), B1 => n36, B2 => 
                           regs(1842), ZN => n739);
   U976 : NAND3_X1 port map( A1 => n741, A2 => n740, A3 => n739, ZN => 
                           curr_proc_regs(306));
   U977 : NAND2_X1 port map( A1 => regs(819), A2 => n7, ZN => n744);
   U978 : AOI22_X1 port map( A1 => n32, A2 => regs(1331), B1 => n1586, B2 => 
                           regs(307), ZN => n743);
   U979 : AOI22_X1 port map( A1 => n13, A2 => regs(2355), B1 => n1588, B2 => 
                           regs(1843), ZN => n742);
   U980 : NAND3_X1 port map( A1 => n744, A2 => n743, A3 => n742, ZN => 
                           curr_proc_regs(307));
   U981 : NAND2_X1 port map( A1 => regs(820), A2 => n18, ZN => n747);
   U982 : AOI22_X1 port map( A1 => n32, A2 => regs(1332), B1 => n30, B2 => 
                           regs(308), ZN => n746);
   U983 : AOI22_X1 port map( A1 => n5, A2 => regs(2356), B1 => n36, B2 => 
                           regs(1844), ZN => n745);
   U984 : NAND3_X1 port map( A1 => n747, A2 => n746, A3 => n745, ZN => 
                           curr_proc_regs(308));
   U985 : NAND2_X1 port map( A1 => regs(821), A2 => n22, ZN => n750);
   U986 : AOI22_X1 port map( A1 => n32, A2 => regs(1333), B1 => n1586, B2 => 
                           regs(309), ZN => n749);
   U987 : AOI22_X1 port map( A1 => n13, A2 => regs(2357), B1 => n9, B2 => 
                           regs(1845), ZN => n748);
   U988 : NAND3_X1 port map( A1 => n750, A2 => n749, A3 => n748, ZN => 
                           curr_proc_regs(309));
   U989 : NAND2_X1 port map( A1 => regs(542), A2 => n1585, ZN => n753);
   U990 : AOI22_X1 port map( A1 => n32, A2 => regs(1054), B1 => n28, B2 => 
                           regs(30), ZN => n752);
   U991 : AOI22_X1 port map( A1 => n13, A2 => regs(2078), B1 => n34, B2 => 
                           regs(1566), ZN => n751);
   U992 : NAND3_X1 port map( A1 => n753, A2 => n752, A3 => n751, ZN => 
                           curr_proc_regs(30));
   U993 : NAND2_X1 port map( A1 => regs(822), A2 => n19, ZN => n756);
   U994 : AOI22_X1 port map( A1 => n32, A2 => regs(1334), B1 => n30, B2 => 
                           regs(310), ZN => n755);
   U995 : AOI22_X1 port map( A1 => n13, A2 => regs(2358), B1 => n36, B2 => 
                           regs(1846), ZN => n754);
   U996 : NAND3_X1 port map( A1 => n756, A2 => n755, A3 => n754, ZN => 
                           curr_proc_regs(310));
   U997 : NAND2_X1 port map( A1 => regs(823), A2 => n6, ZN => n759);
   U998 : AOI22_X1 port map( A1 => n32, A2 => regs(1335), B1 => n30, B2 => 
                           regs(311), ZN => n758);
   U999 : AOI22_X1 port map( A1 => n13, A2 => regs(2359), B1 => n36, B2 => 
                           regs(1847), ZN => n757);
   U1000 : NAND3_X1 port map( A1 => n759, A2 => n758, A3 => n757, ZN => 
                           curr_proc_regs(311));
   U1001 : NAND2_X1 port map( A1 => regs(824), A2 => n2, ZN => n762);
   U1002 : AOI22_X1 port map( A1 => n32, A2 => regs(1336), B1 => n30, B2 => 
                           regs(312), ZN => n761);
   U1003 : AOI22_X1 port map( A1 => n13, A2 => regs(2360), B1 => n36, B2 => 
                           regs(1848), ZN => n760);
   U1004 : NAND3_X1 port map( A1 => n762, A2 => n761, A3 => n760, ZN => 
                           curr_proc_regs(312));
   U1005 : NAND2_X1 port map( A1 => regs(825), A2 => n18, ZN => n765);
   U1006 : AOI22_X1 port map( A1 => n32, A2 => regs(1337), B1 => n30, B2 => 
                           regs(313), ZN => n764);
   U1007 : AOI22_X1 port map( A1 => n13, A2 => regs(2361), B1 => n36, B2 => 
                           regs(1849), ZN => n763);
   U1008 : NAND3_X1 port map( A1 => n765, A2 => n764, A3 => n763, ZN => 
                           curr_proc_regs(313));
   U1009 : NAND2_X1 port map( A1 => regs(826), A2 => n22, ZN => n768);
   U1010 : AOI22_X1 port map( A1 => n32, A2 => regs(1338), B1 => n31, B2 => 
                           regs(314), ZN => n767);
   U1011 : AOI22_X1 port map( A1 => n13, A2 => regs(2362), B1 => n35, B2 => 
                           regs(1850), ZN => n766);
   U1012 : NAND3_X1 port map( A1 => n768, A2 => n767, A3 => n766, ZN => 
                           curr_proc_regs(314));
   U1013 : NAND2_X1 port map( A1 => regs(827), A2 => n1585, ZN => n771);
   U1014 : AOI22_X1 port map( A1 => n32, A2 => regs(1339), B1 => n30, B2 => 
                           regs(315), ZN => n770);
   U1015 : AOI22_X1 port map( A1 => n13, A2 => regs(2363), B1 => n36, B2 => 
                           regs(1851), ZN => n769);
   U1016 : NAND3_X1 port map( A1 => n771, A2 => n770, A3 => n769, ZN => 
                           curr_proc_regs(315));
   U1017 : NAND2_X1 port map( A1 => regs(828), A2 => n19, ZN => n774);
   U1018 : AOI22_X1 port map( A1 => n32, A2 => regs(1340), B1 => n30, B2 => 
                           regs(316), ZN => n773);
   U1019 : AOI22_X1 port map( A1 => n13, A2 => regs(2364), B1 => n36, B2 => 
                           regs(1852), ZN => n772);
   U1020 : NAND3_X1 port map( A1 => n774, A2 => n773, A3 => n772, ZN => 
                           curr_proc_regs(316));
   U1021 : NAND2_X1 port map( A1 => regs(829), A2 => n6, ZN => n777);
   U1022 : AOI22_X1 port map( A1 => n32, A2 => regs(1341), B1 => n30, B2 => 
                           regs(317), ZN => n776);
   U1023 : AOI22_X1 port map( A1 => n13, A2 => regs(2365), B1 => n36, B2 => 
                           regs(1853), ZN => n775);
   U1024 : NAND3_X1 port map( A1 => n777, A2 => n776, A3 => n775, ZN => 
                           curr_proc_regs(317));
   U1025 : NAND2_X1 port map( A1 => regs(830), A2 => n7, ZN => n780);
   U1026 : AOI22_X1 port map( A1 => n32, A2 => regs(1342), B1 => n30, B2 => 
                           regs(318), ZN => n779);
   U1027 : AOI22_X1 port map( A1 => n13, A2 => regs(2366), B1 => n36, B2 => 
                           regs(1854), ZN => n778);
   U1028 : NAND3_X1 port map( A1 => n780, A2 => n779, A3 => n778, ZN => 
                           curr_proc_regs(318));
   U1029 : NAND2_X1 port map( A1 => regs(831), A2 => n7, ZN => n783);
   U1030 : AOI22_X1 port map( A1 => n32, A2 => regs(1343), B1 => n30, B2 => 
                           regs(319), ZN => n782);
   U1031 : AOI22_X1 port map( A1 => n13, A2 => regs(2367), B1 => n36, B2 => 
                           regs(1855), ZN => n781);
   U1032 : NAND3_X1 port map( A1 => n783, A2 => n782, A3 => n781, ZN => 
                           curr_proc_regs(319));
   U1033 : NAND2_X1 port map( A1 => regs(543), A2 => n7, ZN => n786);
   U1034 : AOI22_X1 port map( A1 => n32, A2 => regs(1055), B1 => n30, B2 => 
                           regs(31), ZN => n785);
   U1035 : AOI22_X1 port map( A1 => n5, A2 => regs(2079), B1 => n36, B2 => 
                           regs(1567), ZN => n784);
   U1036 : NAND3_X1 port map( A1 => n786, A2 => n785, A3 => n784, ZN => 
                           curr_proc_regs(31));
   U1037 : NAND2_X1 port map( A1 => regs(832), A2 => n7, ZN => n789);
   U1038 : AOI22_X1 port map( A1 => n32, A2 => regs(1344), B1 => n30, B2 => 
                           regs(320), ZN => n788);
   U1039 : AOI22_X1 port map( A1 => n5, A2 => regs(2368), B1 => n36, B2 => 
                           regs(1856), ZN => n787);
   U1040 : NAND3_X1 port map( A1 => n789, A2 => n788, A3 => n787, ZN => 
                           curr_proc_regs(320));
   U1041 : NAND2_X1 port map( A1 => regs(833), A2 => n7, ZN => n792);
   U1042 : AOI22_X1 port map( A1 => n32, A2 => regs(1345), B1 => n30, B2 => 
                           regs(321), ZN => n791);
   U1043 : AOI22_X1 port map( A1 => n5, A2 => regs(2369), B1 => n36, B2 => 
                           regs(1857), ZN => n790);
   U1044 : NAND3_X1 port map( A1 => n792, A2 => n791, A3 => n790, ZN => 
                           curr_proc_regs(321));
   U1045 : NAND2_X1 port map( A1 => regs(834), A2 => n7, ZN => n795);
   U1046 : AOI22_X1 port map( A1 => n32, A2 => regs(1346), B1 => n8, B2 => 
                           regs(322), ZN => n794);
   U1047 : AOI22_X1 port map( A1 => n5, A2 => regs(2370), B1 => n4, B2 => 
                           regs(1858), ZN => n793);
   U1048 : NAND3_X1 port map( A1 => n795, A2 => n794, A3 => n793, ZN => 
                           curr_proc_regs(322));
   U1049 : NAND2_X1 port map( A1 => regs(835), A2 => n7, ZN => n798);
   U1050 : AOI22_X1 port map( A1 => n32, A2 => regs(1347), B1 => n30, B2 => 
                           regs(323), ZN => n797);
   U1051 : AOI22_X1 port map( A1 => n13, A2 => regs(2371), B1 => n36, B2 => 
                           regs(1859), ZN => n796);
   U1052 : NAND3_X1 port map( A1 => n798, A2 => n797, A3 => n796, ZN => 
                           curr_proc_regs(323));
   U1053 : NAND2_X1 port map( A1 => regs(836), A2 => n1, ZN => n801);
   U1054 : AOI22_X1 port map( A1 => n32, A2 => regs(1348), B1 => n30, B2 => 
                           regs(324), ZN => n800);
   U1055 : AOI22_X1 port map( A1 => n13, A2 => regs(2372), B1 => n36, B2 => 
                           regs(1860), ZN => n799);
   U1056 : NAND3_X1 port map( A1 => n801, A2 => n800, A3 => n799, ZN => 
                           curr_proc_regs(324));
   U1057 : NAND2_X1 port map( A1 => regs(837), A2 => n1, ZN => n804);
   U1058 : AOI22_X1 port map( A1 => n32, A2 => regs(1349), B1 => n30, B2 => 
                           regs(325), ZN => n803);
   U1059 : AOI22_X1 port map( A1 => n5, A2 => regs(2373), B1 => n36, B2 => 
                           regs(1861), ZN => n802);
   U1060 : NAND3_X1 port map( A1 => n804, A2 => n803, A3 => n802, ZN => 
                           curr_proc_regs(325));
   U1061 : NAND2_X1 port map( A1 => regs(838), A2 => n1, ZN => n807);
   U1062 : AOI22_X1 port map( A1 => n32, A2 => regs(1350), B1 => n30, B2 => 
                           regs(326), ZN => n806);
   U1063 : AOI22_X1 port map( A1 => n5, A2 => regs(2374), B1 => n36, B2 => 
                           regs(1862), ZN => n805);
   U1064 : NAND3_X1 port map( A1 => n807, A2 => n806, A3 => n805, ZN => 
                           curr_proc_regs(326));
   U1065 : NAND2_X1 port map( A1 => regs(839), A2 => n1, ZN => n810);
   U1066 : AOI22_X1 port map( A1 => n32, A2 => regs(1351), B1 => n30, B2 => 
                           regs(327), ZN => n809);
   U1067 : AOI22_X1 port map( A1 => n5, A2 => regs(2375), B1 => n36, B2 => 
                           regs(1863), ZN => n808);
   U1068 : NAND3_X1 port map( A1 => n810, A2 => n809, A3 => n808, ZN => 
                           curr_proc_regs(327));
   U1069 : NAND2_X1 port map( A1 => regs(840), A2 => n19, ZN => n813);
   U1070 : AOI22_X1 port map( A1 => n32, A2 => regs(1352), B1 => n1586, B2 => 
                           regs(328), ZN => n812);
   U1071 : AOI22_X1 port map( A1 => n5, A2 => regs(2376), B1 => n36, B2 => 
                           regs(1864), ZN => n811);
   U1072 : NAND3_X1 port map( A1 => n813, A2 => n812, A3 => n811, ZN => 
                           curr_proc_regs(328));
   U1073 : NAND2_X1 port map( A1 => regs(841), A2 => n1, ZN => n816);
   U1074 : AOI22_X1 port map( A1 => n32, A2 => regs(1353), B1 => n8, B2 => 
                           regs(329), ZN => n815);
   U1075 : AOI22_X1 port map( A1 => n13, A2 => regs(2377), B1 => n35, B2 => 
                           regs(1865), ZN => n814);
   U1076 : NAND3_X1 port map( A1 => n816, A2 => n815, A3 => n814, ZN => 
                           curr_proc_regs(329));
   U1077 : NAND2_X1 port map( A1 => regs(544), A2 => n6, ZN => n819);
   U1078 : AOI22_X1 port map( A1 => n32, A2 => regs(1056), B1 => n31, B2 => 
                           regs(32), ZN => n818);
   U1079 : AOI22_X1 port map( A1 => n40, A2 => regs(2080), B1 => n35, B2 => 
                           regs(1568), ZN => n817);
   U1080 : NAND3_X1 port map( A1 => n819, A2 => n818, A3 => n817, ZN => 
                           curr_proc_regs(32));
   U1081 : NAND2_X1 port map( A1 => regs(842), A2 => n19, ZN => n822);
   U1082 : AOI22_X1 port map( A1 => n32, A2 => regs(1354), B1 => n3, B2 => 
                           regs(330), ZN => n821);
   U1083 : AOI22_X1 port map( A1 => n46, A2 => regs(2378), B1 => n36, B2 => 
                           regs(1866), ZN => n820);
   U1084 : NAND3_X1 port map( A1 => n822, A2 => n821, A3 => n820, ZN => 
                           curr_proc_regs(330));
   U1085 : NAND2_X1 port map( A1 => regs(843), A2 => n7, ZN => n825);
   U1086 : AOI22_X1 port map( A1 => n32, A2 => regs(1355), B1 => n31, B2 => 
                           regs(331), ZN => n824);
   U1087 : AOI22_X1 port map( A1 => n40, A2 => regs(2379), B1 => n35, B2 => 
                           regs(1867), ZN => n823);
   U1088 : NAND3_X1 port map( A1 => n825, A2 => n824, A3 => n823, ZN => 
                           curr_proc_regs(331));
   U1089 : NAND2_X1 port map( A1 => regs(844), A2 => n1, ZN => n828);
   U1090 : AOI22_X1 port map( A1 => n32, A2 => regs(1356), B1 => n31, B2 => 
                           regs(332), ZN => n827);
   U1091 : AOI22_X1 port map( A1 => n46, A2 => regs(2380), B1 => n35, B2 => 
                           regs(1868), ZN => n826);
   U1092 : NAND3_X1 port map( A1 => n828, A2 => n827, A3 => n826, ZN => 
                           curr_proc_regs(332));
   U1093 : NAND2_X1 port map( A1 => regs(845), A2 => n1585, ZN => n831);
   U1094 : AOI22_X1 port map( A1 => n32, A2 => regs(1357), B1 => n31, B2 => 
                           regs(333), ZN => n830);
   U1095 : AOI22_X1 port map( A1 => n40, A2 => regs(2381), B1 => n35, B2 => 
                           regs(1869), ZN => n829);
   U1096 : NAND3_X1 port map( A1 => n831, A2 => n830, A3 => n829, ZN => 
                           curr_proc_regs(333));
   U1097 : NAND2_X1 port map( A1 => regs(846), A2 => n1585, ZN => n834);
   U1098 : AOI22_X1 port map( A1 => n32, A2 => regs(1358), B1 => n31, B2 => 
                           regs(334), ZN => n833);
   U1099 : AOI22_X1 port map( A1 => n46, A2 => regs(2382), B1 => n35, B2 => 
                           regs(1870), ZN => n832);
   U1100 : NAND3_X1 port map( A1 => n834, A2 => n833, A3 => n832, ZN => 
                           curr_proc_regs(334));
   U1101 : NAND2_X1 port map( A1 => regs(847), A2 => n19, ZN => n837);
   U1102 : AOI22_X1 port map( A1 => n32, A2 => regs(1359), B1 => n31, B2 => 
                           regs(335), ZN => n836);
   U1103 : AOI22_X1 port map( A1 => n10, A2 => regs(2383), B1 => n35, B2 => 
                           regs(1871), ZN => n835);
   U1104 : NAND3_X1 port map( A1 => n837, A2 => n836, A3 => n835, ZN => 
                           curr_proc_regs(335));
   U1105 : NAND2_X1 port map( A1 => regs(848), A2 => n1, ZN => n840);
   U1106 : AOI22_X1 port map( A1 => n32, A2 => regs(1360), B1 => n3, B2 => 
                           regs(336), ZN => n839);
   U1107 : AOI22_X1 port map( A1 => n10, A2 => regs(2384), B1 => n34, B2 => 
                           regs(1872), ZN => n838);
   U1108 : NAND3_X1 port map( A1 => n840, A2 => n839, A3 => n838, ZN => 
                           curr_proc_regs(336));
   U1109 : NAND2_X1 port map( A1 => regs(849), A2 => n2, ZN => n843);
   U1110 : AOI22_X1 port map( A1 => n32, A2 => regs(1361), B1 => n31, B2 => 
                           regs(337), ZN => n842);
   U1111 : AOI22_X1 port map( A1 => n46, A2 => regs(2385), B1 => n35, B2 => 
                           regs(1873), ZN => n841);
   U1112 : NAND3_X1 port map( A1 => n843, A2 => n842, A3 => n841, ZN => 
                           curr_proc_regs(337));
   U1113 : NAND2_X1 port map( A1 => regs(850), A2 => n24, ZN => n846);
   U1114 : AOI22_X1 port map( A1 => n32, A2 => regs(1362), B1 => n28, B2 => 
                           regs(338), ZN => n845);
   U1115 : AOI22_X1 port map( A1 => n47, A2 => regs(2386), B1 => n34, B2 => 
                           regs(1874), ZN => n844);
   U1116 : NAND3_X1 port map( A1 => n846, A2 => n845, A3 => n844, ZN => 
                           curr_proc_regs(338));
   U1117 : NAND2_X1 port map( A1 => regs(851), A2 => n18, ZN => n849);
   U1118 : AOI22_X1 port map( A1 => n32, A2 => regs(1363), B1 => n3, B2 => 
                           regs(339), ZN => n848);
   U1119 : AOI22_X1 port map( A1 => n47, A2 => regs(2387), B1 => n37, B2 => 
                           regs(1875), ZN => n847);
   U1120 : NAND3_X1 port map( A1 => n849, A2 => n848, A3 => n847, ZN => 
                           curr_proc_regs(339));
   U1121 : NAND2_X1 port map( A1 => regs(545), A2 => n24, ZN => n852);
   U1122 : AOI22_X1 port map( A1 => n32, A2 => regs(1057), B1 => n31, B2 => 
                           regs(33), ZN => n851);
   U1123 : AOI22_X1 port map( A1 => n47, A2 => regs(2081), B1 => n35, B2 => 
                           regs(1569), ZN => n850);
   U1124 : NAND3_X1 port map( A1 => n852, A2 => n851, A3 => n850, ZN => 
                           curr_proc_regs(33));
   U1125 : NAND2_X1 port map( A1 => regs(852), A2 => n24, ZN => n855);
   U1126 : AOI22_X1 port map( A1 => n32, A2 => regs(1364), B1 => n8, B2 => 
                           regs(340), ZN => n854);
   U1127 : AOI22_X1 port map( A1 => n16, A2 => regs(2388), B1 => n34, B2 => 
                           regs(1876), ZN => n853);
   U1128 : NAND3_X1 port map( A1 => n855, A2 => n854, A3 => n853, ZN => 
                           curr_proc_regs(340));
   U1129 : NAND2_X1 port map( A1 => regs(853), A2 => n18, ZN => n858);
   U1130 : AOI22_X1 port map( A1 => n32, A2 => regs(1365), B1 => n8, B2 => 
                           regs(341), ZN => n857);
   U1131 : AOI22_X1 port map( A1 => n16, A2 => regs(2389), B1 => n35, B2 => 
                           regs(1877), ZN => n856);
   U1132 : NAND3_X1 port map( A1 => n858, A2 => n857, A3 => n856, ZN => 
                           curr_proc_regs(341));
   U1133 : NAND2_X1 port map( A1 => regs(854), A2 => n24, ZN => n861);
   U1134 : AOI22_X1 port map( A1 => n32, A2 => regs(1366), B1 => n8, B2 => 
                           regs(342), ZN => n860);
   U1135 : AOI22_X1 port map( A1 => n47, A2 => regs(2390), B1 => n36, B2 => 
                           regs(1878), ZN => n859);
   U1136 : NAND3_X1 port map( A1 => n861, A2 => n860, A3 => n859, ZN => 
                           curr_proc_regs(342));
   U1137 : NAND2_X1 port map( A1 => regs(855), A2 => n24, ZN => n864);
   U1138 : AOI22_X1 port map( A1 => n32, A2 => regs(1367), B1 => n31, B2 => 
                           regs(343), ZN => n863);
   U1139 : AOI22_X1 port map( A1 => n47, A2 => regs(2391), B1 => n35, B2 => 
                           regs(1879), ZN => n862);
   U1140 : NAND3_X1 port map( A1 => n864, A2 => n863, A3 => n862, ZN => 
                           curr_proc_regs(343));
   U1141 : NAND2_X1 port map( A1 => regs(856), A2 => n18, ZN => n867);
   U1142 : AOI22_X1 port map( A1 => n32, A2 => regs(1368), B1 => n1586, B2 => 
                           regs(344), ZN => n866);
   U1143 : AOI22_X1 port map( A1 => n16, A2 => regs(2392), B1 => n39, B2 => 
                           regs(1880), ZN => n865);
   U1144 : NAND3_X1 port map( A1 => n867, A2 => n866, A3 => n865, ZN => 
                           curr_proc_regs(344));
   U1145 : NAND2_X1 port map( A1 => regs(857), A2 => n24, ZN => n870);
   U1146 : AOI22_X1 port map( A1 => n32, A2 => regs(1369), B1 => n3, B2 => 
                           regs(345), ZN => n869);
   U1147 : AOI22_X1 port map( A1 => n16, A2 => regs(2393), B1 => n9, B2 => 
                           regs(1881), ZN => n868);
   U1148 : NAND3_X1 port map( A1 => n870, A2 => n869, A3 => n868, ZN => 
                           curr_proc_regs(345));
   U1149 : NAND2_X1 port map( A1 => regs(858), A2 => n24, ZN => n873);
   U1150 : AOI22_X1 port map( A1 => n32, A2 => regs(1370), B1 => n28, B2 => 
                           regs(346), ZN => n872);
   U1151 : AOI22_X1 port map( A1 => n16, A2 => regs(2394), B1 => n34, B2 => 
                           regs(1882), ZN => n871);
   U1152 : NAND3_X1 port map( A1 => n873, A2 => n872, A3 => n871, ZN => 
                           curr_proc_regs(346));
   U1153 : NAND2_X1 port map( A1 => regs(859), A2 => n24, ZN => n876);
   U1154 : AOI22_X1 port map( A1 => n32, A2 => regs(1371), B1 => n31, B2 => 
                           regs(347), ZN => n875);
   U1155 : AOI22_X1 port map( A1 => n16, A2 => regs(2395), B1 => n35, B2 => 
                           regs(1883), ZN => n874);
   U1156 : NAND3_X1 port map( A1 => n876, A2 => n875, A3 => n874, ZN => 
                           curr_proc_regs(347));
   U1157 : NAND2_X1 port map( A1 => regs(860), A2 => n2, ZN => n879);
   U1158 : AOI22_X1 port map( A1 => n32, A2 => regs(1372), B1 => n3, B2 => 
                           regs(348), ZN => n878);
   U1159 : AOI22_X1 port map( A1 => n16, A2 => regs(2396), B1 => n35, B2 => 
                           regs(1884), ZN => n877);
   U1160 : NAND3_X1 port map( A1 => n879, A2 => n878, A3 => n877, ZN => 
                           curr_proc_regs(348));
   U1161 : NAND2_X1 port map( A1 => regs(861), A2 => n2, ZN => n882);
   U1162 : AOI22_X1 port map( A1 => n32, A2 => regs(1373), B1 => n28, B2 => 
                           regs(349), ZN => n881);
   U1163 : AOI22_X1 port map( A1 => n47, A2 => regs(2397), B1 => n34, B2 => 
                           regs(1885), ZN => n880);
   U1164 : NAND3_X1 port map( A1 => n882, A2 => n881, A3 => n880, ZN => 
                           curr_proc_regs(349));
   U1165 : NAND2_X1 port map( A1 => regs(546), A2 => n2, ZN => n885);
   U1166 : AOI22_X1 port map( A1 => n32, A2 => regs(1058), B1 => n8, B2 => 
                           regs(34), ZN => n884);
   U1167 : AOI22_X1 port map( A1 => n47, A2 => regs(2082), B1 => n35, B2 => 
                           regs(1570), ZN => n883);
   U1168 : NAND3_X1 port map( A1 => n885, A2 => n884, A3 => n883, ZN => 
                           curr_proc_regs(34));
   U1169 : NAND2_X1 port map( A1 => regs(862), A2 => n2, ZN => n888);
   U1170 : AOI22_X1 port map( A1 => n32, A2 => regs(1374), B1 => n28, B2 => 
                           regs(350), ZN => n887);
   U1171 : AOI22_X1 port map( A1 => n16, A2 => regs(2398), B1 => n35, B2 => 
                           regs(1886), ZN => n886);
   U1172 : NAND3_X1 port map( A1 => n888, A2 => n887, A3 => n886, ZN => 
                           curr_proc_regs(350));
   U1173 : NAND2_X1 port map( A1 => regs(863), A2 => n2, ZN => n891);
   U1174 : AOI22_X1 port map( A1 => n32, A2 => regs(1375), B1 => n26, B2 => 
                           regs(351), ZN => n890);
   U1175 : AOI22_X1 port map( A1 => n16, A2 => regs(2399), B1 => n36, B2 => 
                           regs(1887), ZN => n889);
   U1176 : NAND3_X1 port map( A1 => n891, A2 => n890, A3 => n889, ZN => 
                           curr_proc_regs(351));
   U1177 : NAND2_X1 port map( A1 => regs(864), A2 => n2, ZN => n894);
   U1178 : AOI22_X1 port map( A1 => n32, A2 => regs(1376), B1 => n1586, B2 => 
                           regs(352), ZN => n893);
   U1179 : AOI22_X1 port map( A1 => n16, A2 => regs(2400), B1 => n34, B2 => 
                           regs(1888), ZN => n892);
   U1180 : NAND3_X1 port map( A1 => n894, A2 => n893, A3 => n892, ZN => 
                           curr_proc_regs(352));
   U1181 : NAND2_X1 port map( A1 => regs(865), A2 => n2, ZN => n897);
   U1182 : AOI22_X1 port map( A1 => n32, A2 => regs(1377), B1 => n31, B2 => 
                           regs(353), ZN => n896);
   U1183 : AOI22_X1 port map( A1 => n47, A2 => regs(2401), B1 => n37, B2 => 
                           regs(1889), ZN => n895);
   U1184 : NAND3_X1 port map( A1 => n897, A2 => n896, A3 => n895, ZN => 
                           curr_proc_regs(353));
   U1185 : NAND2_X1 port map( A1 => regs(866), A2 => n2, ZN => n900);
   U1186 : AOI22_X1 port map( A1 => n32, A2 => regs(1378), B1 => n3, B2 => 
                           regs(354), ZN => n899);
   U1187 : AOI22_X1 port map( A1 => n16, A2 => regs(2402), B1 => n34, B2 => 
                           regs(1890), ZN => n898);
   U1188 : NAND3_X1 port map( A1 => n900, A2 => n899, A3 => n898, ZN => 
                           curr_proc_regs(354));
   U1189 : NAND2_X1 port map( A1 => regs(867), A2 => n2, ZN => n903);
   U1190 : AOI22_X1 port map( A1 => n32, A2 => regs(1379), B1 => n8, B2 => 
                           regs(355), ZN => n902);
   U1191 : AOI22_X1 port map( A1 => n16, A2 => regs(2403), B1 => n35, B2 => 
                           regs(1891), ZN => n901);
   U1192 : NAND3_X1 port map( A1 => n903, A2 => n902, A3 => n901, ZN => 
                           curr_proc_regs(355));
   U1193 : NAND2_X1 port map( A1 => regs(868), A2 => n2, ZN => n906);
   U1194 : AOI22_X1 port map( A1 => n32, A2 => regs(1380), B1 => n8, B2 => 
                           regs(356), ZN => n905);
   U1195 : AOI22_X1 port map( A1 => n16, A2 => regs(2404), B1 => n35, B2 => 
                           regs(1892), ZN => n904);
   U1196 : NAND3_X1 port map( A1 => n906, A2 => n905, A3 => n904, ZN => 
                           curr_proc_regs(356));
   U1197 : NAND2_X1 port map( A1 => regs(869), A2 => n2, ZN => n909);
   U1198 : AOI22_X1 port map( A1 => n32, A2 => regs(1381), B1 => n25, B2 => 
                           regs(357), ZN => n908);
   U1199 : AOI22_X1 port map( A1 => n47, A2 => regs(2405), B1 => n39, B2 => 
                           regs(1893), ZN => n907);
   U1200 : NAND3_X1 port map( A1 => n909, A2 => n908, A3 => n907, ZN => 
                           curr_proc_regs(357));
   U1201 : NAND2_X1 port map( A1 => regs(870), A2 => n23, ZN => n912);
   U1202 : AOI22_X1 port map( A1 => n32, A2 => regs(1382), B1 => n8, B2 => 
                           regs(358), ZN => n911);
   U1203 : AOI22_X1 port map( A1 => n47, A2 => regs(2406), B1 => n35, B2 => 
                           regs(1894), ZN => n910);
   U1204 : NAND3_X1 port map( A1 => n912, A2 => n911, A3 => n910, ZN => 
                           curr_proc_regs(358));
   U1205 : NAND2_X1 port map( A1 => regs(871), A2 => n23, ZN => n915);
   U1206 : AOI22_X1 port map( A1 => n32, A2 => regs(1383), B1 => n31, B2 => 
                           regs(359), ZN => n914);
   U1207 : AOI22_X1 port map( A1 => n16, A2 => regs(2407), B1 => n35, B2 => 
                           regs(1895), ZN => n913);
   U1208 : NAND3_X1 port map( A1 => n915, A2 => n914, A3 => n913, ZN => 
                           curr_proc_regs(359));
   U1209 : NAND2_X1 port map( A1 => regs(547), A2 => n17, ZN => n918);
   U1210 : AOI22_X1 port map( A1 => n32, A2 => regs(1059), B1 => n31, B2 => 
                           regs(35), ZN => n917);
   U1211 : AOI22_X1 port map( A1 => n16, A2 => regs(2083), B1 => n35, B2 => 
                           regs(1571), ZN => n916);
   U1212 : NAND3_X1 port map( A1 => n918, A2 => n917, A3 => n916, ZN => 
                           curr_proc_regs(35));
   U1213 : NAND2_X1 port map( A1 => regs(872), A2 => n20, ZN => n921);
   U1214 : AOI22_X1 port map( A1 => n32, A2 => regs(1384), B1 => n28, B2 => 
                           regs(360), ZN => n920);
   U1215 : AOI22_X1 port map( A1 => n47, A2 => regs(2408), B1 => n34, B2 => 
                           regs(1896), ZN => n919);
   U1216 : NAND3_X1 port map( A1 => n921, A2 => n920, A3 => n919, ZN => 
                           curr_proc_regs(360));
   U1217 : NAND2_X1 port map( A1 => regs(873), A2 => n23, ZN => n924);
   U1218 : AOI22_X1 port map( A1 => n32, A2 => regs(1385), B1 => n8, B2 => 
                           regs(361), ZN => n923);
   U1219 : AOI22_X1 port map( A1 => n16, A2 => regs(2409), B1 => n35, B2 => 
                           regs(1897), ZN => n922);
   U1220 : NAND3_X1 port map( A1 => n924, A2 => n923, A3 => n922, ZN => 
                           curr_proc_regs(361));
   U1221 : NAND2_X1 port map( A1 => regs(874), A2 => n17, ZN => n927);
   U1222 : AOI22_X1 port map( A1 => n32, A2 => regs(1386), B1 => n8, B2 => 
                           regs(362), ZN => n926);
   U1223 : AOI22_X1 port map( A1 => n16, A2 => regs(2410), B1 => n4, B2 => 
                           regs(1898), ZN => n925);
   U1224 : NAND3_X1 port map( A1 => n927, A2 => n926, A3 => n925, ZN => 
                           curr_proc_regs(362));
   U1225 : NAND2_X1 port map( A1 => regs(875), A2 => n20, ZN => n930);
   U1226 : AOI22_X1 port map( A1 => n32, A2 => regs(1387), B1 => n31, B2 => 
                           regs(363), ZN => n929);
   U1227 : AOI22_X1 port map( A1 => n47, A2 => regs(2411), B1 => n35, B2 => 
                           regs(1899), ZN => n928);
   U1228 : NAND3_X1 port map( A1 => n930, A2 => n929, A3 => n928, ZN => 
                           curr_proc_regs(363));
   U1229 : NAND2_X1 port map( A1 => regs(876), A2 => n23, ZN => n933);
   U1230 : AOI22_X1 port map( A1 => n32, A2 => regs(1388), B1 => n1586, B2 => 
                           regs(364), ZN => n932);
   U1231 : AOI22_X1 port map( A1 => n16, A2 => regs(2412), B1 => n36, B2 => 
                           regs(1900), ZN => n931);
   U1232 : NAND3_X1 port map( A1 => n933, A2 => n932, A3 => n931, ZN => 
                           curr_proc_regs(364));
   U1233 : NAND2_X1 port map( A1 => regs(877), A2 => n17, ZN => n936);
   U1234 : AOI22_X1 port map( A1 => n32, A2 => regs(1389), B1 => n31, B2 => 
                           regs(365), ZN => n935);
   U1235 : AOI22_X1 port map( A1 => n16, A2 => regs(2413), B1 => n35, B2 => 
                           regs(1901), ZN => n934);
   U1236 : NAND3_X1 port map( A1 => n936, A2 => n935, A3 => n934, ZN => 
                           curr_proc_regs(365));
   U1237 : NAND2_X1 port map( A1 => regs(878), A2 => n20, ZN => n939);
   U1238 : AOI22_X1 port map( A1 => n32, A2 => regs(1390), B1 => n31, B2 => 
                           regs(366), ZN => n938);
   U1239 : AOI22_X1 port map( A1 => n47, A2 => regs(2414), B1 => n35, B2 => 
                           regs(1902), ZN => n937);
   U1240 : NAND3_X1 port map( A1 => n939, A2 => n938, A3 => n937, ZN => 
                           curr_proc_regs(366));
   U1241 : NAND2_X1 port map( A1 => regs(879), A2 => n23, ZN => n942);
   U1242 : AOI22_X1 port map( A1 => n32, A2 => regs(1391), B1 => n31, B2 => 
                           regs(367), ZN => n941);
   U1243 : AOI22_X1 port map( A1 => n40, A2 => regs(2415), B1 => n35, B2 => 
                           regs(1903), ZN => n940);
   U1244 : NAND3_X1 port map( A1 => n942, A2 => n941, A3 => n940, ZN => 
                           curr_proc_regs(367));
   U1245 : NAND2_X1 port map( A1 => regs(880), A2 => n22, ZN => n945);
   U1246 : AOI22_X1 port map( A1 => n32, A2 => regs(1392), B1 => n3, B2 => 
                           regs(368), ZN => n944);
   U1247 : AOI22_X1 port map( A1 => n16, A2 => regs(2416), B1 => n4, B2 => 
                           regs(1904), ZN => n943);
   U1248 : NAND3_X1 port map( A1 => n945, A2 => n944, A3 => n943, ZN => 
                           curr_proc_regs(368));
   U1249 : NAND2_X1 port map( A1 => regs(881), A2 => n1585, ZN => n948);
   U1250 : AOI22_X1 port map( A1 => n32, A2 => regs(1393), B1 => n3, B2 => 
                           regs(369), ZN => n947);
   U1251 : AOI22_X1 port map( A1 => n16, A2 => regs(2417), B1 => n36, B2 => 
                           regs(1905), ZN => n946);
   U1252 : NAND3_X1 port map( A1 => n948, A2 => n947, A3 => n946, ZN => 
                           curr_proc_regs(369));
   U1253 : NAND2_X1 port map( A1 => regs(548), A2 => n22, ZN => n951);
   U1254 : AOI22_X1 port map( A1 => n32, A2 => regs(1060), B1 => n31, B2 => 
                           regs(36), ZN => n950);
   U1255 : AOI22_X1 port map( A1 => n16, A2 => regs(2084), B1 => n4, B2 => 
                           regs(1572), ZN => n949);
   U1256 : NAND3_X1 port map( A1 => n951, A2 => n950, A3 => n949, ZN => 
                           curr_proc_regs(36));
   U1257 : NAND2_X1 port map( A1 => regs(882), A2 => n1585, ZN => n954);
   U1258 : AOI22_X1 port map( A1 => n32, A2 => regs(1394), B1 => n31, B2 => 
                           regs(370), ZN => n953);
   U1259 : AOI22_X1 port map( A1 => n16, A2 => regs(2418), B1 => n35, B2 => 
                           regs(1906), ZN => n952);
   U1260 : NAND3_X1 port map( A1 => n954, A2 => n953, A3 => n952, ZN => 
                           curr_proc_regs(370));
   U1261 : NAND2_X1 port map( A1 => regs(883), A2 => n6, ZN => n957);
   U1262 : AOI22_X1 port map( A1 => n32, A2 => regs(1395), B1 => n31, B2 => 
                           regs(371), ZN => n956);
   U1263 : AOI22_X1 port map( A1 => n16, A2 => regs(2419), B1 => n35, B2 => 
                           regs(1907), ZN => n955);
   U1264 : NAND3_X1 port map( A1 => n957, A2 => n956, A3 => n955, ZN => 
                           curr_proc_regs(371));
   U1265 : NAND2_X1 port map( A1 => regs(884), A2 => n7, ZN => n960);
   U1266 : AOI22_X1 port map( A1 => n32, A2 => regs(1396), B1 => n31, B2 => 
                           regs(372), ZN => n959);
   U1267 : AOI22_X1 port map( A1 => n16, A2 => regs(2420), B1 => n35, B2 => 
                           regs(1908), ZN => n958);
   U1268 : NAND3_X1 port map( A1 => n960, A2 => n959, A3 => n958, ZN => 
                           curr_proc_regs(372));
   U1269 : NAND2_X1 port map( A1 => regs(885), A2 => n6, ZN => n963);
   U1270 : AOI22_X1 port map( A1 => n32, A2 => regs(1397), B1 => n31, B2 => 
                           regs(373), ZN => n962);
   U1271 : AOI22_X1 port map( A1 => n16, A2 => regs(2421), B1 => n35, B2 => 
                           regs(1909), ZN => n961);
   U1272 : NAND3_X1 port map( A1 => n963, A2 => n962, A3 => n961, ZN => 
                           curr_proc_regs(373));
   U1273 : NAND2_X1 port map( A1 => regs(886), A2 => n20, ZN => n966);
   U1274 : AOI22_X1 port map( A1 => n32, A2 => regs(1398), B1 => n31, B2 => 
                           regs(374), ZN => n965);
   U1275 : AOI22_X1 port map( A1 => n16, A2 => regs(2422), B1 => n35, B2 => 
                           regs(1910), ZN => n964);
   U1276 : NAND3_X1 port map( A1 => n966, A2 => n965, A3 => n964, ZN => 
                           curr_proc_regs(374));
   U1277 : NAND2_X1 port map( A1 => regs(887), A2 => n18, ZN => n969);
   U1278 : AOI22_X1 port map( A1 => n32, A2 => regs(1399), B1 => n29, B2 => 
                           regs(375), ZN => n968);
   U1279 : AOI22_X1 port map( A1 => n16, A2 => regs(2423), B1 => n34, B2 => 
                           regs(1911), ZN => n967);
   U1280 : NAND3_X1 port map( A1 => n969, A2 => n968, A3 => n967, ZN => 
                           curr_proc_regs(375));
   U1281 : NAND2_X1 port map( A1 => regs(888), A2 => n2, ZN => n972);
   U1282 : AOI22_X1 port map( A1 => n32, A2 => regs(1400), B1 => n31, B2 => 
                           regs(376), ZN => n971);
   U1283 : AOI22_X1 port map( A1 => n16, A2 => regs(2424), B1 => n35, B2 => 
                           regs(1912), ZN => n970);
   U1284 : NAND3_X1 port map( A1 => n972, A2 => n971, A3 => n970, ZN => 
                           curr_proc_regs(376));
   U1285 : NAND2_X1 port map( A1 => regs(889), A2 => n1585, ZN => n975);
   U1286 : AOI22_X1 port map( A1 => n32, A2 => regs(1401), B1 => n31, B2 => 
                           regs(377), ZN => n974);
   U1287 : AOI22_X1 port map( A1 => n16, A2 => regs(2425), B1 => n35, B2 => 
                           regs(1913), ZN => n973);
   U1288 : NAND3_X1 port map( A1 => n975, A2 => n974, A3 => n973, ZN => 
                           curr_proc_regs(377));
   U1289 : NAND2_X1 port map( A1 => regs(890), A2 => n21, ZN => n978);
   U1290 : AOI22_X1 port map( A1 => n32, A2 => regs(1402), B1 => n8, B2 => 
                           regs(378), ZN => n977);
   U1291 : AOI22_X1 port map( A1 => n16, A2 => regs(2426), B1 => n4, B2 => 
                           regs(1914), ZN => n976);
   U1292 : NAND3_X1 port map( A1 => n978, A2 => n977, A3 => n976, ZN => 
                           curr_proc_regs(378));
   U1293 : NAND2_X1 port map( A1 => regs(891), A2 => n21, ZN => n981);
   U1294 : AOI22_X1 port map( A1 => n32, A2 => regs(1403), B1 => n31, B2 => 
                           regs(379), ZN => n980);
   U1295 : AOI22_X1 port map( A1 => n16, A2 => regs(2427), B1 => n35, B2 => 
                           regs(1915), ZN => n979);
   U1296 : NAND3_X1 port map( A1 => n981, A2 => n980, A3 => n979, ZN => 
                           curr_proc_regs(379));
   U1297 : NAND2_X1 port map( A1 => regs(549), A2 => n21, ZN => n984);
   U1298 : AOI22_X1 port map( A1 => n32, A2 => regs(1061), B1 => n8, B2 => 
                           regs(37), ZN => n983);
   U1299 : AOI22_X1 port map( A1 => n16, A2 => regs(2085), B1 => n4, B2 => 
                           regs(1573), ZN => n982);
   U1300 : NAND3_X1 port map( A1 => n984, A2 => n983, A3 => n982, ZN => 
                           curr_proc_regs(37));
   U1301 : NAND2_X1 port map( A1 => regs(892), A2 => n21, ZN => n987);
   U1302 : AOI22_X1 port map( A1 => n32, A2 => regs(1404), B1 => n31, B2 => 
                           regs(380), ZN => n986);
   U1303 : AOI22_X1 port map( A1 => n16, A2 => regs(2428), B1 => n35, B2 => 
                           regs(1916), ZN => n985);
   U1304 : NAND3_X1 port map( A1 => n987, A2 => n986, A3 => n985, ZN => 
                           curr_proc_regs(380));
   U1305 : NAND2_X1 port map( A1 => regs(893), A2 => n21, ZN => n990);
   U1306 : AOI22_X1 port map( A1 => n32, A2 => regs(1405), B1 => n31, B2 => 
                           regs(381), ZN => n989);
   U1307 : AOI22_X1 port map( A1 => n16, A2 => regs(2429), B1 => n35, B2 => 
                           regs(1917), ZN => n988);
   U1308 : NAND3_X1 port map( A1 => n990, A2 => n989, A3 => n988, ZN => 
                           curr_proc_regs(381));
   U1309 : NAND2_X1 port map( A1 => regs(894), A2 => n21, ZN => n993);
   U1310 : AOI22_X1 port map( A1 => n32, A2 => regs(1406), B1 => n31, B2 => 
                           regs(382), ZN => n992);
   U1311 : AOI22_X1 port map( A1 => n16, A2 => regs(2430), B1 => n35, B2 => 
                           regs(1918), ZN => n991);
   U1312 : NAND3_X1 port map( A1 => n993, A2 => n992, A3 => n991, ZN => 
                           curr_proc_regs(382));
   U1313 : NAND2_X1 port map( A1 => regs(895), A2 => n18, ZN => n996);
   U1314 : AOI22_X1 port map( A1 => n32, A2 => regs(1407), B1 => n3, B2 => 
                           regs(383), ZN => n995);
   U1315 : AOI22_X1 port map( A1 => n16, A2 => regs(2431), B1 => n38, B2 => 
                           regs(1919), ZN => n994);
   U1316 : NAND3_X1 port map( A1 => n996, A2 => n995, A3 => n994, ZN => 
                           curr_proc_regs(383));
   U1317 : NAND2_X1 port map( A1 => regs(896), A2 => n1585, ZN => n999);
   U1318 : AOI22_X1 port map( A1 => n32, A2 => regs(1408), B1 => n3, B2 => 
                           regs(384), ZN => n998);
   U1319 : AOI22_X1 port map( A1 => n16, A2 => regs(2432), B1 => n37, B2 => 
                           regs(1920), ZN => n997);
   U1320 : NAND3_X1 port map( A1 => n999, A2 => n998, A3 => n997, ZN => 
                           curr_proc_regs(384));
   U1321 : NAND2_X1 port map( A1 => regs(897), A2 => n19, ZN => n1002);
   U1322 : AOI22_X1 port map( A1 => n32, A2 => regs(1409), B1 => n29, B2 => 
                           regs(385), ZN => n1001);
   U1323 : AOI22_X1 port map( A1 => n16, A2 => regs(2433), B1 => n34, B2 => 
                           regs(1921), ZN => n1000);
   U1324 : NAND3_X1 port map( A1 => n1002, A2 => n1001, A3 => n1000, ZN => 
                           curr_proc_regs(385));
   U1325 : NAND2_X1 port map( A1 => regs(898), A2 => n6, ZN => n1005);
   U1326 : AOI22_X1 port map( A1 => n32, A2 => regs(1410), B1 => n3, B2 => 
                           regs(386), ZN => n1004);
   U1327 : AOI22_X1 port map( A1 => n16, A2 => regs(2434), B1 => n35, B2 => 
                           regs(1922), ZN => n1003);
   U1328 : NAND3_X1 port map( A1 => n1005, A2 => n1004, A3 => n1003, ZN => 
                           curr_proc_regs(386));
   U1329 : NAND2_X1 port map( A1 => regs(899), A2 => n2, ZN => n1008);
   U1330 : AOI22_X1 port map( A1 => n32, A2 => regs(1411), B1 => n1586, B2 => 
                           regs(387), ZN => n1007);
   U1331 : AOI22_X1 port map( A1 => n16, A2 => regs(2435), B1 => n36, B2 => 
                           regs(1923), ZN => n1006);
   U1332 : NAND3_X1 port map( A1 => n1008, A2 => n1007, A3 => n1006, ZN => 
                           curr_proc_regs(387));
   U1333 : NAND2_X1 port map( A1 => regs(900), A2 => n17, ZN => n1011);
   U1334 : AOI22_X1 port map( A1 => n32, A2 => regs(1412), B1 => n3, B2 => 
                           regs(388), ZN => n1010);
   U1335 : AOI22_X1 port map( A1 => n47, A2 => regs(2436), B1 => n4, B2 => 
                           regs(1924), ZN => n1009);
   U1336 : NAND3_X1 port map( A1 => n1011, A2 => n1010, A3 => n1009, ZN => 
                           curr_proc_regs(388));
   U1337 : NAND2_X1 port map( A1 => regs(901), A2 => n1585, ZN => n1014);
   U1338 : AOI22_X1 port map( A1 => n32, A2 => regs(1413), B1 => n3, B2 => 
                           regs(389), ZN => n1013);
   U1339 : AOI22_X1 port map( A1 => n47, A2 => regs(2437), B1 => n38, B2 => 
                           regs(1925), ZN => n1012);
   U1340 : NAND3_X1 port map( A1 => n1014, A2 => n1013, A3 => n1012, ZN => 
                           curr_proc_regs(389));
   U1341 : NAND2_X1 port map( A1 => regs(550), A2 => n2, ZN => n1017);
   U1342 : AOI22_X1 port map( A1 => n32, A2 => regs(1062), B1 => n29, B2 => 
                           regs(38), ZN => n1016);
   U1343 : AOI22_X1 port map( A1 => n47, A2 => regs(2086), B1 => n38, B2 => 
                           regs(1574), ZN => n1015);
   U1344 : NAND3_X1 port map( A1 => n1017, A2 => n1016, A3 => n1015, ZN => 
                           curr_proc_regs(38));
   U1345 : NAND2_X1 port map( A1 => regs(902), A2 => n7, ZN => n1020);
   U1346 : AOI22_X1 port map( A1 => n32, A2 => regs(1414), B1 => n28, B2 => 
                           regs(390), ZN => n1019);
   U1347 : AOI22_X1 port map( A1 => n16, A2 => regs(2438), B1 => n4, B2 => 
                           regs(1926), ZN => n1018);
   U1348 : NAND3_X1 port map( A1 => n1020, A2 => n1019, A3 => n1018, ZN => 
                           curr_proc_regs(390));
   U1349 : NAND2_X1 port map( A1 => regs(903), A2 => n7, ZN => n1023);
   U1350 : AOI22_X1 port map( A1 => n32, A2 => regs(1415), B1 => n1586, B2 => 
                           regs(391), ZN => n1022);
   U1351 : AOI22_X1 port map( A1 => n16, A2 => regs(2439), B1 => n33, B2 => 
                           regs(1927), ZN => n1021);
   U1352 : NAND3_X1 port map( A1 => n1023, A2 => n1022, A3 => n1021, ZN => 
                           curr_proc_regs(391));
   U1353 : NAND2_X1 port map( A1 => regs(904), A2 => n1, ZN => n1026);
   U1354 : AOI22_X1 port map( A1 => n32, A2 => regs(1416), B1 => n28, B2 => 
                           regs(392), ZN => n1025);
   U1355 : AOI22_X1 port map( A1 => n47, A2 => regs(2440), B1 => n4, B2 => 
                           regs(1928), ZN => n1024);
   U1356 : NAND3_X1 port map( A1 => n1026, A2 => n1025, A3 => n1024, ZN => 
                           curr_proc_regs(392));
   U1357 : NAND2_X1 port map( A1 => regs(905), A2 => n19, ZN => n1029);
   U1358 : AOI22_X1 port map( A1 => n32, A2 => regs(1417), B1 => n8, B2 => 
                           regs(393), ZN => n1028);
   U1359 : AOI22_X1 port map( A1 => n47, A2 => regs(2441), B1 => n4, B2 => 
                           regs(1929), ZN => n1027);
   U1360 : NAND3_X1 port map( A1 => n1029, A2 => n1028, A3 => n1027, ZN => 
                           curr_proc_regs(393));
   U1361 : NAND2_X1 port map( A1 => regs(906), A2 => n22, ZN => n1032);
   U1362 : AOI22_X1 port map( A1 => n32, A2 => regs(1418), B1 => n8, B2 => 
                           regs(394), ZN => n1031);
   U1363 : AOI22_X1 port map( A1 => n47, A2 => regs(2442), B1 => n4, B2 => 
                           regs(1930), ZN => n1030);
   U1364 : NAND3_X1 port map( A1 => n1032, A2 => n1031, A3 => n1030, ZN => 
                           curr_proc_regs(394));
   U1365 : NAND2_X1 port map( A1 => regs(907), A2 => n23, ZN => n1035);
   U1366 : AOI22_X1 port map( A1 => n32, A2 => regs(1419), B1 => n3, B2 => 
                           regs(395), ZN => n1034);
   U1367 : AOI22_X1 port map( A1 => n47, A2 => regs(2443), B1 => n37, B2 => 
                           regs(1931), ZN => n1033);
   U1368 : NAND3_X1 port map( A1 => n1035, A2 => n1034, A3 => n1033, ZN => 
                           curr_proc_regs(395));
   U1369 : NAND2_X1 port map( A1 => regs(908), A2 => n17, ZN => n1038);
   U1370 : AOI22_X1 port map( A1 => n32, A2 => regs(1420), B1 => n29, B2 => 
                           regs(396), ZN => n1037);
   U1371 : AOI22_X1 port map( A1 => n16, A2 => regs(2444), B1 => n37, B2 => 
                           regs(1932), ZN => n1036);
   U1372 : NAND3_X1 port map( A1 => n1038, A2 => n1037, A3 => n1036, ZN => 
                           curr_proc_regs(396));
   U1373 : NAND2_X1 port map( A1 => regs(909), A2 => n1585, ZN => n1041);
   U1374 : AOI22_X1 port map( A1 => n32, A2 => regs(1421), B1 => n28, B2 => 
                           regs(397), ZN => n1040);
   U1375 : AOI22_X1 port map( A1 => n5, A2 => regs(2445), B1 => n4, B2 => 
                           regs(1933), ZN => n1039);
   U1376 : NAND3_X1 port map( A1 => n1041, A2 => n1040, A3 => n1039, ZN => 
                           curr_proc_regs(397));
   U1377 : NAND2_X1 port map( A1 => regs(910), A2 => n19, ZN => n1044);
   U1378 : AOI22_X1 port map( A1 => n32, A2 => regs(1422), B1 => n8, B2 => 
                           regs(398), ZN => n1043);
   U1379 : AOI22_X1 port map( A1 => n5, A2 => regs(2446), B1 => n36, B2 => 
                           regs(1934), ZN => n1042);
   U1380 : NAND3_X1 port map( A1 => n1044, A2 => n1043, A3 => n1042, ZN => 
                           curr_proc_regs(398));
   U1381 : NAND2_X1 port map( A1 => regs(911), A2 => n19, ZN => n1047);
   U1382 : AOI22_X1 port map( A1 => n32, A2 => regs(1423), B1 => n3, B2 => 
                           regs(399), ZN => n1046);
   U1383 : AOI22_X1 port map( A1 => n5, A2 => regs(2447), B1 => n4, B2 => 
                           regs(1935), ZN => n1045);
   U1384 : NAND3_X1 port map( A1 => n1047, A2 => n1046, A3 => n1045, ZN => 
                           curr_proc_regs(399));
   U1385 : NAND2_X1 port map( A1 => regs(551), A2 => n19, ZN => n1050);
   U1386 : AOI22_X1 port map( A1 => n32, A2 => regs(1063), B1 => n3, B2 => 
                           regs(39), ZN => n1049);
   U1387 : AOI22_X1 port map( A1 => n5, A2 => regs(2087), B1 => n38, B2 => 
                           regs(1575), ZN => n1048);
   U1388 : NAND3_X1 port map( A1 => n1050, A2 => n1049, A3 => n1048, ZN => 
                           curr_proc_regs(39));
   U1389 : NAND2_X1 port map( A1 => regs(515), A2 => n19, ZN => n1053);
   U1390 : AOI22_X1 port map( A1 => n32, A2 => regs(1027), B1 => n3, B2 => 
                           regs(3), ZN => n1052);
   U1391 : AOI22_X1 port map( A1 => n5, A2 => regs(2051), B1 => n33, B2 => 
                           regs(1539), ZN => n1051);
   U1392 : NAND3_X1 port map( A1 => n1053, A2 => n1052, A3 => n1051, ZN => 
                           curr_proc_regs(3));
   U1393 : NAND2_X1 port map( A1 => regs(912), A2 => n19, ZN => n1056);
   U1394 : AOI22_X1 port map( A1 => n32, A2 => regs(1424), B1 => n29, B2 => 
                           regs(400), ZN => n1055);
   U1395 : AOI22_X1 port map( A1 => n5, A2 => regs(2448), B1 => n37, B2 => 
                           regs(1936), ZN => n1054);
   U1396 : NAND3_X1 port map( A1 => n1056, A2 => n1055, A3 => n1054, ZN => 
                           curr_proc_regs(400));
   U1397 : NAND2_X1 port map( A1 => regs(913), A2 => n19, ZN => n1059);
   U1398 : AOI22_X1 port map( A1 => n32, A2 => regs(1425), B1 => n3, B2 => 
                           regs(401), ZN => n1058);
   U1399 : AOI22_X1 port map( A1 => n14, A2 => regs(2449), B1 => n38, B2 => 
                           regs(1937), ZN => n1057);
   U1400 : NAND3_X1 port map( A1 => n1059, A2 => n1058, A3 => n1057, ZN => 
                           curr_proc_regs(401));
   U1401 : NAND2_X1 port map( A1 => regs(914), A2 => n19, ZN => n1062);
   U1402 : AOI22_X1 port map( A1 => n32, A2 => regs(1426), B1 => n1586, B2 => 
                           regs(402), ZN => n1061);
   U1403 : AOI22_X1 port map( A1 => n5, A2 => regs(2450), B1 => n4, B2 => 
                           regs(1938), ZN => n1060);
   U1404 : NAND3_X1 port map( A1 => n1062, A2 => n1061, A3 => n1060, ZN => 
                           curr_proc_regs(402));
   U1405 : NAND2_X1 port map( A1 => regs(915), A2 => n19, ZN => n1065);
   U1406 : AOI22_X1 port map( A1 => n32, A2 => regs(1427), B1 => n28, B2 => 
                           regs(403), ZN => n1064);
   U1407 : AOI22_X1 port map( A1 => n5, A2 => regs(2451), B1 => n4, B2 => 
                           regs(1939), ZN => n1063);
   U1408 : NAND3_X1 port map( A1 => n1065, A2 => n1064, A3 => n1063, ZN => 
                           curr_proc_regs(403));
   U1409 : NAND2_X1 port map( A1 => regs(916), A2 => n19, ZN => n1068);
   U1410 : AOI22_X1 port map( A1 => n32, A2 => regs(1428), B1 => n8, B2 => 
                           regs(404), ZN => n1067);
   U1411 : AOI22_X1 port map( A1 => n14, A2 => regs(2452), B1 => n37, B2 => 
                           regs(1940), ZN => n1066);
   U1412 : NAND3_X1 port map( A1 => n1068, A2 => n1067, A3 => n1066, ZN => 
                           curr_proc_regs(404));
   U1413 : NAND2_X1 port map( A1 => regs(917), A2 => n19, ZN => n1071);
   U1414 : AOI22_X1 port map( A1 => n32, A2 => regs(1429), B1 => n8, B2 => 
                           regs(405), ZN => n1070);
   U1415 : AOI22_X1 port map( A1 => n5, A2 => regs(2453), B1 => n36, B2 => 
                           regs(1941), ZN => n1069);
   U1416 : NAND3_X1 port map( A1 => n1071, A2 => n1070, A3 => n1069, ZN => 
                           curr_proc_regs(405));
   U1417 : NAND2_X1 port map( A1 => regs(918), A2 => n19, ZN => n1074);
   U1418 : AOI22_X1 port map( A1 => n32, A2 => regs(1430), B1 => n31, B2 => 
                           regs(406), ZN => n1073);
   U1419 : AOI22_X1 port map( A1 => n5, A2 => regs(2454), B1 => n4, B2 => 
                           regs(1942), ZN => n1072);
   U1420 : NAND3_X1 port map( A1 => n1074, A2 => n1073, A3 => n1072, ZN => 
                           curr_proc_regs(406));
   U1421 : NAND2_X1 port map( A1 => regs(919), A2 => n7, ZN => n1077);
   U1422 : AOI22_X1 port map( A1 => n32, A2 => regs(1431), B1 => n8, B2 => 
                           regs(407), ZN => n1076);
   U1423 : AOI22_X1 port map( A1 => n5, A2 => regs(2455), B1 => n4, B2 => 
                           regs(1943), ZN => n1075);
   U1424 : NAND3_X1 port map( A1 => n1077, A2 => n1076, A3 => n1075, ZN => 
                           curr_proc_regs(407));
   U1425 : NAND2_X1 port map( A1 => regs(920), A2 => n20, ZN => n1080);
   U1426 : AOI22_X1 port map( A1 => n32, A2 => regs(1432), B1 => n8, B2 => 
                           regs(408), ZN => n1079);
   U1427 : AOI22_X1 port map( A1 => n14, A2 => regs(2456), B1 => n4, B2 => 
                           regs(1944), ZN => n1078);
   U1428 : NAND3_X1 port map( A1 => n1080, A2 => n1079, A3 => n1078, ZN => 
                           curr_proc_regs(408));
   U1429 : NAND2_X1 port map( A1 => regs(921), A2 => n1585, ZN => n1083);
   U1430 : AOI22_X1 port map( A1 => n32, A2 => regs(1433), B1 => n8, B2 => 
                           regs(409), ZN => n1082);
   U1431 : AOI22_X1 port map( A1 => n14, A2 => regs(2457), B1 => n4, B2 => 
                           regs(1945), ZN => n1081);
   U1432 : NAND3_X1 port map( A1 => n1083, A2 => n1082, A3 => n1081, ZN => 
                           curr_proc_regs(409));
   U1433 : NAND2_X1 port map( A1 => regs(552), A2 => n19, ZN => n1086);
   U1434 : AOI22_X1 port map( A1 => n32, A2 => regs(1064), B1 => n8, B2 => 
                           regs(40), ZN => n1085);
   U1435 : AOI22_X1 port map( A1 => n14, A2 => regs(2088), B1 => n4, B2 => 
                           regs(1576), ZN => n1084);
   U1436 : NAND3_X1 port map( A1 => n1086, A2 => n1085, A3 => n1084, ZN => 
                           curr_proc_regs(40));
   U1437 : NAND2_X1 port map( A1 => regs(922), A2 => n1, ZN => n1089);
   U1438 : AOI22_X1 port map( A1 => n32, A2 => regs(1434), B1 => n8, B2 => 
                           regs(410), ZN => n1088);
   U1439 : AOI22_X1 port map( A1 => n5, A2 => regs(2458), B1 => n4, B2 => 
                           regs(1946), ZN => n1087);
   U1440 : NAND3_X1 port map( A1 => n1089, A2 => n1088, A3 => n1087, ZN => 
                           curr_proc_regs(410));
   U1441 : NAND2_X1 port map( A1 => regs(923), A2 => n2, ZN => n1092);
   U1442 : AOI22_X1 port map( A1 => n32, A2 => regs(1435), B1 => n8, B2 => 
                           regs(411), ZN => n1091);
   U1443 : AOI22_X1 port map( A1 => n14, A2 => regs(2459), B1 => n4, B2 => 
                           regs(1947), ZN => n1090);
   U1444 : NAND3_X1 port map( A1 => n1092, A2 => n1091, A3 => n1090, ZN => 
                           curr_proc_regs(411));
   U1445 : NAND2_X1 port map( A1 => regs(924), A2 => n21, ZN => n1095);
   U1446 : AOI22_X1 port map( A1 => n32, A2 => regs(1436), B1 => n8, B2 => 
                           regs(412), ZN => n1094);
   U1447 : AOI22_X1 port map( A1 => n5, A2 => regs(2460), B1 => n4, B2 => 
                           regs(1948), ZN => n1093);
   U1448 : NAND3_X1 port map( A1 => n1095, A2 => n1094, A3 => n1093, ZN => 
                           curr_proc_regs(412));
   U1449 : NAND2_X1 port map( A1 => regs(925), A2 => n17, ZN => n1098);
   U1450 : AOI22_X1 port map( A1 => n32, A2 => regs(1437), B1 => n8, B2 => 
                           regs(413), ZN => n1097);
   U1451 : AOI22_X1 port map( A1 => n14, A2 => regs(2461), B1 => n4, B2 => 
                           regs(1949), ZN => n1096);
   U1452 : NAND3_X1 port map( A1 => n1098, A2 => n1097, A3 => n1096, ZN => 
                           curr_proc_regs(413));
   U1453 : NAND2_X1 port map( A1 => regs(926), A2 => n22, ZN => n1101);
   U1454 : AOI22_X1 port map( A1 => n32, A2 => regs(1438), B1 => n8, B2 => 
                           regs(414), ZN => n1100);
   U1455 : AOI22_X1 port map( A1 => n5, A2 => regs(2462), B1 => n4, B2 => 
                           regs(1950), ZN => n1099);
   U1456 : NAND3_X1 port map( A1 => n1101, A2 => n1100, A3 => n1099, ZN => 
                           curr_proc_regs(414));
   U1457 : NAND2_X1 port map( A1 => regs(927), A2 => n23, ZN => n1104);
   U1458 : AOI22_X1 port map( A1 => n32, A2 => regs(1439), B1 => n8, B2 => 
                           regs(415), ZN => n1103);
   U1459 : AOI22_X1 port map( A1 => n14, A2 => regs(2463), B1 => n4, B2 => 
                           regs(1951), ZN => n1102);
   U1460 : NAND3_X1 port map( A1 => n1104, A2 => n1103, A3 => n1102, ZN => 
                           curr_proc_regs(415));
   U1461 : NAND2_X1 port map( A1 => regs(928), A2 => n1, ZN => n1107);
   U1462 : AOI22_X1 port map( A1 => n32, A2 => regs(1440), B1 => n8, B2 => 
                           regs(416), ZN => n1106);
   U1463 : AOI22_X1 port map( A1 => n14, A2 => regs(2464), B1 => n4, B2 => 
                           regs(1952), ZN => n1105);
   U1464 : NAND3_X1 port map( A1 => n1107, A2 => n1106, A3 => n1105, ZN => 
                           curr_proc_regs(416));
   U1465 : NAND2_X1 port map( A1 => regs(929), A2 => n1, ZN => n1110);
   U1466 : AOI22_X1 port map( A1 => n32, A2 => regs(1441), B1 => n28, B2 => 
                           regs(417), ZN => n1109);
   U1467 : AOI22_X1 port map( A1 => n14, A2 => regs(2465), B1 => n34, B2 => 
                           regs(1953), ZN => n1108);
   U1468 : NAND3_X1 port map( A1 => n1110, A2 => n1109, A3 => n1108, ZN => 
                           curr_proc_regs(417));
   U1469 : NAND2_X1 port map( A1 => regs(930), A2 => n1, ZN => n1113);
   U1470 : AOI22_X1 port map( A1 => n32, A2 => regs(1442), B1 => n8, B2 => 
                           regs(418), ZN => n1112);
   U1471 : AOI22_X1 port map( A1 => n5, A2 => regs(2466), B1 => n35, B2 => 
                           regs(1954), ZN => n1111);
   U1472 : NAND3_X1 port map( A1 => n1113, A2 => n1112, A3 => n1111, ZN => 
                           curr_proc_regs(418));
   U1473 : NAND2_X1 port map( A1 => regs(931), A2 => n1, ZN => n1116);
   U1474 : AOI22_X1 port map( A1 => n32, A2 => regs(1443), B1 => n28, B2 => 
                           regs(419), ZN => n1115);
   U1475 : AOI22_X1 port map( A1 => n14, A2 => regs(2467), B1 => n37, B2 => 
                           regs(1955), ZN => n1114);
   U1476 : NAND3_X1 port map( A1 => n1116, A2 => n1115, A3 => n1114, ZN => 
                           curr_proc_regs(419));
   U1477 : NAND2_X1 port map( A1 => regs(553), A2 => n1, ZN => n1119);
   U1478 : AOI22_X1 port map( A1 => n32, A2 => regs(1065), B1 => n8, B2 => 
                           regs(41), ZN => n1118);
   U1479 : AOI22_X1 port map( A1 => n14, A2 => regs(2089), B1 => n34, B2 => 
                           regs(1577), ZN => n1117);
   U1480 : NAND3_X1 port map( A1 => n1119, A2 => n1118, A3 => n1117, ZN => 
                           curr_proc_regs(41));
   U1481 : NAND2_X1 port map( A1 => regs(932), A2 => n1, ZN => n1122);
   U1482 : AOI22_X1 port map( A1 => n32, A2 => regs(1444), B1 => n1586, B2 => 
                           regs(420), ZN => n1121);
   U1483 : AOI22_X1 port map( A1 => n5, A2 => regs(2468), B1 => n35, B2 => 
                           regs(1956), ZN => n1120);
   U1484 : NAND3_X1 port map( A1 => n1122, A2 => n1121, A3 => n1120, ZN => 
                           curr_proc_regs(420));
   U1485 : NAND2_X1 port map( A1 => regs(933), A2 => n1, ZN => n1125);
   U1486 : AOI22_X1 port map( A1 => n32, A2 => regs(1445), B1 => n8, B2 => 
                           regs(421), ZN => n1124);
   U1487 : AOI22_X1 port map( A1 => n14, A2 => regs(2469), B1 => n37, B2 => 
                           regs(1957), ZN => n1123);
   U1488 : NAND3_X1 port map( A1 => n1125, A2 => n1124, A3 => n1123, ZN => 
                           curr_proc_regs(421));
   U1489 : NAND2_X1 port map( A1 => regs(934), A2 => n1, ZN => n1128);
   U1490 : AOI22_X1 port map( A1 => n32, A2 => regs(1446), B1 => n8, B2 => 
                           regs(422), ZN => n1127);
   U1491 : AOI22_X1 port map( A1 => n14, A2 => regs(2470), B1 => n34, B2 => 
                           regs(1958), ZN => n1126);
   U1492 : NAND3_X1 port map( A1 => n1128, A2 => n1127, A3 => n1126, ZN => 
                           curr_proc_regs(422));
   U1493 : NAND2_X1 port map( A1 => regs(935), A2 => n1, ZN => n1131);
   U1494 : AOI22_X1 port map( A1 => n32, A2 => regs(1447), B1 => n28, B2 => 
                           regs(423), ZN => n1130);
   U1495 : AOI22_X1 port map( A1 => n5, A2 => regs(2471), B1 => n35, B2 => 
                           regs(1959), ZN => n1129);
   U1496 : NAND3_X1 port map( A1 => n1131, A2 => n1130, A3 => n1129, ZN => 
                           curr_proc_regs(423));
   U1497 : NAND2_X1 port map( A1 => regs(936), A2 => n1, ZN => n1134);
   U1498 : AOI22_X1 port map( A1 => n32, A2 => regs(1448), B1 => n28, B2 => 
                           regs(424), ZN => n1133);
   U1499 : AOI22_X1 port map( A1 => n14, A2 => regs(2472), B1 => n37, B2 => 
                           regs(1960), ZN => n1132);
   U1500 : NAND3_X1 port map( A1 => n1134, A2 => n1133, A3 => n1132, ZN => 
                           curr_proc_regs(424));
   U1501 : NAND2_X1 port map( A1 => regs(937), A2 => n1, ZN => n1137);
   U1502 : AOI22_X1 port map( A1 => n32, A2 => regs(1449), B1 => n8, B2 => 
                           regs(425), ZN => n1136);
   U1503 : AOI22_X1 port map( A1 => n14, A2 => regs(2473), B1 => n34, B2 => 
                           regs(1961), ZN => n1135);
   U1504 : NAND3_X1 port map( A1 => n1137, A2 => n1136, A3 => n1135, ZN => 
                           curr_proc_regs(425));
   U1505 : NAND2_X1 port map( A1 => regs(938), A2 => n1, ZN => n1140);
   U1506 : AOI22_X1 port map( A1 => n32, A2 => regs(1450), B1 => n8, B2 => 
                           regs(426), ZN => n1139);
   U1507 : AOI22_X1 port map( A1 => n14, A2 => regs(2474), B1 => n35, B2 => 
                           regs(1962), ZN => n1138);
   U1508 : NAND3_X1 port map( A1 => n1140, A2 => n1139, A3 => n1138, ZN => 
                           curr_proc_regs(426));
   U1509 : NAND2_X1 port map( A1 => regs(939), A2 => n6, ZN => n1143);
   U1510 : AOI22_X1 port map( A1 => n32, A2 => regs(1451), B1 => n3, B2 => 
                           regs(427), ZN => n1142);
   U1511 : AOI22_X1 port map( A1 => n14, A2 => regs(2475), B1 => n33, B2 => 
                           regs(1963), ZN => n1141);
   U1512 : NAND3_X1 port map( A1 => n1143, A2 => n1142, A3 => n1141, ZN => 
                           curr_proc_regs(427));
   U1513 : NAND2_X1 port map( A1 => regs(940), A2 => n6, ZN => n1146);
   U1514 : AOI22_X1 port map( A1 => n32, A2 => regs(1452), B1 => n3, B2 => 
                           regs(428), ZN => n1145);
   U1515 : AOI22_X1 port map( A1 => n14, A2 => regs(2476), B1 => n33, B2 => 
                           regs(1964), ZN => n1144);
   U1516 : NAND3_X1 port map( A1 => n1146, A2 => n1145, A3 => n1144, ZN => 
                           curr_proc_regs(428));
   U1517 : NAND2_X1 port map( A1 => regs(941), A2 => n6, ZN => n1149);
   U1518 : AOI22_X1 port map( A1 => n32, A2 => regs(1453), B1 => n29, B2 => 
                           regs(429), ZN => n1148);
   U1519 : AOI22_X1 port map( A1 => n14, A2 => regs(2477), B1 => n38, B2 => 
                           regs(1965), ZN => n1147);
   U1520 : NAND3_X1 port map( A1 => n1149, A2 => n1148, A3 => n1147, ZN => 
                           curr_proc_regs(429));
   U1521 : NAND2_X1 port map( A1 => regs(554), A2 => n6, ZN => n1152);
   U1522 : AOI22_X1 port map( A1 => n32, A2 => regs(1066), B1 => n3, B2 => 
                           regs(42), ZN => n1151);
   U1523 : AOI22_X1 port map( A1 => n14, A2 => regs(2090), B1 => n33, B2 => 
                           regs(1578), ZN => n1150);
   U1524 : NAND3_X1 port map( A1 => n1152, A2 => n1151, A3 => n1150, ZN => 
                           curr_proc_regs(42));
   U1525 : NAND2_X1 port map( A1 => regs(942), A2 => n6, ZN => n1155);
   U1526 : AOI22_X1 port map( A1 => n32, A2 => regs(1454), B1 => n1586, B2 => 
                           regs(430), ZN => n1154);
   U1527 : AOI22_X1 port map( A1 => n14, A2 => regs(2478), B1 => n4, B2 => 
                           regs(1966), ZN => n1153);
   U1528 : NAND3_X1 port map( A1 => n1155, A2 => n1154, A3 => n1153, ZN => 
                           curr_proc_regs(430));
   U1529 : NAND2_X1 port map( A1 => regs(943), A2 => n6, ZN => n1158);
   U1530 : AOI22_X1 port map( A1 => n32, A2 => regs(1455), B1 => n28, B2 => 
                           regs(431), ZN => n1157);
   U1531 : AOI22_X1 port map( A1 => n14, A2 => regs(2479), B1 => n4, B2 => 
                           regs(1967), ZN => n1156);
   U1532 : NAND3_X1 port map( A1 => n1158, A2 => n1157, A3 => n1156, ZN => 
                           curr_proc_regs(431));
   U1533 : NAND2_X1 port map( A1 => regs(944), A2 => n6, ZN => n1161);
   U1534 : AOI22_X1 port map( A1 => n32, A2 => regs(1456), B1 => n8, B2 => 
                           regs(432), ZN => n1160);
   U1535 : AOI22_X1 port map( A1 => n14, A2 => regs(2480), B1 => n4, B2 => 
                           regs(1968), ZN => n1159);
   U1536 : NAND3_X1 port map( A1 => n1161, A2 => n1160, A3 => n1159, ZN => 
                           curr_proc_regs(432));
   U1537 : NAND2_X1 port map( A1 => regs(945), A2 => n6, ZN => n1164);
   U1538 : AOI22_X1 port map( A1 => n32, A2 => regs(1457), B1 => n8, B2 => 
                           regs(433), ZN => n1163);
   U1539 : AOI22_X1 port map( A1 => n14, A2 => regs(2481), B1 => n37, B2 => 
                           regs(1969), ZN => n1162);
   U1540 : NAND3_X1 port map( A1 => n1164, A2 => n1163, A3 => n1162, ZN => 
                           curr_proc_regs(433));
   U1541 : NAND2_X1 port map( A1 => regs(946), A2 => n6, ZN => n1167);
   U1542 : AOI22_X1 port map( A1 => n32, A2 => regs(1458), B1 => n3, B2 => 
                           regs(434), ZN => n1166);
   U1543 : AOI22_X1 port map( A1 => n14, A2 => regs(2482), B1 => n36, B2 => 
                           regs(1970), ZN => n1165);
   U1544 : NAND3_X1 port map( A1 => n1167, A2 => n1166, A3 => n1165, ZN => 
                           curr_proc_regs(434));
   U1545 : NAND2_X1 port map( A1 => regs(947), A2 => n6, ZN => n1170);
   U1546 : AOI22_X1 port map( A1 => n32, A2 => regs(1459), B1 => n3, B2 => 
                           regs(435), ZN => n1169);
   U1547 : AOI22_X1 port map( A1 => n14, A2 => regs(2483), B1 => n33, B2 => 
                           regs(1971), ZN => n1168);
   U1548 : NAND3_X1 port map( A1 => n1170, A2 => n1169, A3 => n1168, ZN => 
                           curr_proc_regs(435));
   U1549 : NAND2_X1 port map( A1 => regs(948), A2 => n6, ZN => n1173);
   U1550 : AOI22_X1 port map( A1 => n32, A2 => regs(1460), B1 => n1586, B2 => 
                           regs(436), ZN => n1172);
   U1551 : AOI22_X1 port map( A1 => n14, A2 => regs(2484), B1 => n36, B2 => 
                           regs(1972), ZN => n1171);
   U1552 : NAND3_X1 port map( A1 => n1173, A2 => n1172, A3 => n1171, ZN => 
                           curr_proc_regs(436));
   U1553 : NAND2_X1 port map( A1 => regs(949), A2 => n17, ZN => n1176);
   U1554 : AOI22_X1 port map( A1 => n32, A2 => regs(1461), B1 => n31, B2 => 
                           regs(437), ZN => n1175);
   U1555 : AOI22_X1 port map( A1 => n14, A2 => regs(2485), B1 => n37, B2 => 
                           regs(1973), ZN => n1174);
   U1556 : NAND3_X1 port map( A1 => n1176, A2 => n1175, A3 => n1174, ZN => 
                           curr_proc_regs(437));
   U1557 : NAND2_X1 port map( A1 => regs(950), A2 => n7, ZN => n1179);
   U1558 : AOI22_X1 port map( A1 => n32, A2 => regs(1462), B1 => n1586, B2 => 
                           regs(438), ZN => n1178);
   U1559 : AOI22_X1 port map( A1 => n14, A2 => regs(2486), B1 => n34, B2 => 
                           regs(1974), ZN => n1177);
   U1560 : NAND3_X1 port map( A1 => n1179, A2 => n1178, A3 => n1177, ZN => 
                           curr_proc_regs(438));
   U1561 : NAND2_X1 port map( A1 => regs(951), A2 => n6, ZN => n1182);
   U1562 : AOI22_X1 port map( A1 => n32, A2 => regs(1463), B1 => n28, B2 => 
                           regs(439), ZN => n1181);
   U1563 : AOI22_X1 port map( A1 => n14, A2 => regs(2487), B1 => n35, B2 => 
                           regs(1975), ZN => n1180);
   U1564 : NAND3_X1 port map( A1 => n1182, A2 => n1181, A3 => n1180, ZN => 
                           curr_proc_regs(439));
   U1565 : NAND2_X1 port map( A1 => regs(555), A2 => n18, ZN => n1185);
   U1566 : AOI22_X1 port map( A1 => n32, A2 => regs(1067), B1 => n8, B2 => 
                           regs(43), ZN => n1184);
   U1567 : AOI22_X1 port map( A1 => n14, A2 => regs(2091), B1 => n37, B2 => 
                           regs(1579), ZN => n1183);
   U1568 : NAND3_X1 port map( A1 => n1185, A2 => n1184, A3 => n1183, ZN => 
                           curr_proc_regs(43));
   U1569 : NAND2_X1 port map( A1 => regs(952), A2 => n2, ZN => n1188);
   U1570 : AOI22_X1 port map( A1 => n32, A2 => regs(1464), B1 => n28, B2 => 
                           regs(440), ZN => n1187);
   U1571 : AOI22_X1 port map( A1 => n14, A2 => regs(2488), B1 => n34, B2 => 
                           regs(1976), ZN => n1186);
   U1572 : NAND3_X1 port map( A1 => n1188, A2 => n1187, A3 => n1186, ZN => 
                           curr_proc_regs(440));
   U1573 : NAND2_X1 port map( A1 => regs(953), A2 => n7, ZN => n1191);
   U1574 : AOI22_X1 port map( A1 => n32, A2 => regs(1465), B1 => n8, B2 => 
                           regs(441), ZN => n1190);
   U1575 : AOI22_X1 port map( A1 => n14, A2 => regs(2489), B1 => n35, B2 => 
                           regs(1977), ZN => n1189);
   U1576 : NAND3_X1 port map( A1 => n1191, A2 => n1190, A3 => n1189, ZN => 
                           curr_proc_regs(441));
   U1577 : NAND2_X1 port map( A1 => regs(954), A2 => n20, ZN => n1194);
   U1578 : AOI22_X1 port map( A1 => n32, A2 => regs(1466), B1 => n3, B2 => 
                           regs(442), ZN => n1193);
   U1579 : AOI22_X1 port map( A1 => n14, A2 => regs(2490), B1 => n37, B2 => 
                           regs(1978), ZN => n1192);
   U1580 : NAND3_X1 port map( A1 => n1194, A2 => n1193, A3 => n1192, ZN => 
                           curr_proc_regs(442));
   U1581 : NAND2_X1 port map( A1 => regs(955), A2 => n22, ZN => n1197);
   U1582 : AOI22_X1 port map( A1 => n32, A2 => regs(1467), B1 => n8, B2 => 
                           regs(443), ZN => n1196);
   U1583 : AOI22_X1 port map( A1 => n14, A2 => regs(2491), B1 => n34, B2 => 
                           regs(1979), ZN => n1195);
   U1584 : NAND3_X1 port map( A1 => n1197, A2 => n1196, A3 => n1195, ZN => 
                           curr_proc_regs(443));
   U1585 : NAND2_X1 port map( A1 => regs(956), A2 => n1585, ZN => n1200);
   U1586 : AOI22_X1 port map( A1 => n32, A2 => regs(1468), B1 => n28, B2 => 
                           regs(444), ZN => n1199);
   U1587 : AOI22_X1 port map( A1 => n47, A2 => regs(2492), B1 => n35, B2 => 
                           regs(1980), ZN => n1198);
   U1588 : NAND3_X1 port map( A1 => n1200, A2 => n1199, A3 => n1198, ZN => 
                           curr_proc_regs(444));
   U1589 : NAND2_X1 port map( A1 => regs(957), A2 => n1585, ZN => n1203);
   U1590 : AOI22_X1 port map( A1 => n32, A2 => regs(1469), B1 => n8, B2 => 
                           regs(445), ZN => n1202);
   U1591 : AOI22_X1 port map( A1 => n44, A2 => regs(2493), B1 => n37, B2 => 
                           regs(1981), ZN => n1201);
   U1592 : NAND3_X1 port map( A1 => n1203, A2 => n1202, A3 => n1201, ZN => 
                           curr_proc_regs(445));
   U1593 : NAND2_X1 port map( A1 => regs(958), A2 => n22, ZN => n1206);
   U1594 : AOI22_X1 port map( A1 => n32, A2 => regs(1470), B1 => n29, B2 => 
                           regs(446), ZN => n1205);
   U1595 : AOI22_X1 port map( A1 => n44, A2 => regs(2494), B1 => n34, B2 => 
                           regs(1982), ZN => n1204);
   U1596 : NAND3_X1 port map( A1 => n1206, A2 => n1205, A3 => n1204, ZN => 
                           curr_proc_regs(446));
   U1597 : NAND2_X1 port map( A1 => regs(959), A2 => n24, ZN => n1209);
   U1598 : AOI22_X1 port map( A1 => n32, A2 => regs(1471), B1 => n31, B2 => 
                           regs(447), ZN => n1208);
   U1599 : AOI22_X1 port map( A1 => n44, A2 => regs(2495), B1 => n38, B2 => 
                           regs(1983), ZN => n1207);
   U1600 : NAND3_X1 port map( A1 => n1209, A2 => n1208, A3 => n1207, ZN => 
                           curr_proc_regs(447));
   U1601 : NAND2_X1 port map( A1 => regs(960), A2 => n18, ZN => n1212);
   U1602 : AOI22_X1 port map( A1 => n32, A2 => regs(1472), B1 => n3, B2 => 
                           regs(448), ZN => n1211);
   U1603 : AOI22_X1 port map( A1 => n11, A2 => regs(2496), B1 => n33, B2 => 
                           regs(1984), ZN => n1210);
   U1604 : NAND3_X1 port map( A1 => n1212, A2 => n1211, A3 => n1210, ZN => 
                           curr_proc_regs(448));
   U1605 : NAND2_X1 port map( A1 => regs(961), A2 => n24, ZN => n1215);
   U1606 : AOI22_X1 port map( A1 => n32, A2 => regs(1473), B1 => n3, B2 => 
                           regs(449), ZN => n1214);
   U1607 : AOI22_X1 port map( A1 => n45, A2 => regs(2497), B1 => n4, B2 => 
                           regs(1985), ZN => n1213);
   U1608 : NAND3_X1 port map( A1 => n1215, A2 => n1214, A3 => n1213, ZN => 
                           curr_proc_regs(449));
   U1609 : NAND2_X1 port map( A1 => regs(556), A2 => n18, ZN => n1218);
   U1610 : AOI22_X1 port map( A1 => n32, A2 => regs(1068), B1 => n3, B2 => 
                           regs(44), ZN => n1217);
   U1611 : AOI22_X1 port map( A1 => n45, A2 => regs(2092), B1 => n33, B2 => 
                           regs(1580), ZN => n1216);
   U1612 : NAND3_X1 port map( A1 => n1218, A2 => n1217, A3 => n1216, ZN => 
                           curr_proc_regs(44));
   U1613 : NAND2_X1 port map( A1 => regs(962), A2 => n18, ZN => n1221);
   U1614 : AOI22_X1 port map( A1 => n32, A2 => regs(1474), B1 => n8, B2 => 
                           regs(450), ZN => n1220);
   U1615 : AOI22_X1 port map( A1 => n45, A2 => regs(2498), B1 => n38, B2 => 
                           regs(1986), ZN => n1219);
   U1616 : NAND3_X1 port map( A1 => n1221, A2 => n1220, A3 => n1219, ZN => 
                           curr_proc_regs(450));
   U1617 : NAND2_X1 port map( A1 => regs(963), A2 => n18, ZN => n1224);
   U1618 : AOI22_X1 port map( A1 => n32, A2 => regs(1475), B1 => n8, B2 => 
                           regs(451), ZN => n1223);
   U1619 : AOI22_X1 port map( A1 => n15, A2 => regs(2499), B1 => n4, B2 => 
                           regs(1987), ZN => n1222);
   U1620 : NAND3_X1 port map( A1 => n1224, A2 => n1223, A3 => n1222, ZN => 
                           curr_proc_regs(451));
   U1621 : NAND2_X1 port map( A1 => regs(964), A2 => n24, ZN => n1227);
   U1622 : AOI22_X1 port map( A1 => n32, A2 => regs(1476), B1 => n1586, B2 => 
                           regs(452), ZN => n1226);
   U1623 : AOI22_X1 port map( A1 => n15, A2 => regs(2500), B1 => n4, B2 => 
                           regs(1988), ZN => n1225);
   U1624 : NAND3_X1 port map( A1 => n1227, A2 => n1226, A3 => n1225, ZN => 
                           curr_proc_regs(452));
   U1625 : NAND2_X1 port map( A1 => regs(965), A2 => n24, ZN => n1230);
   U1626 : AOI22_X1 port map( A1 => n32, A2 => regs(1477), B1 => n3, B2 => 
                           regs(453), ZN => n1229);
   U1627 : AOI22_X1 port map( A1 => n45, A2 => regs(2501), B1 => n37, B2 => 
                           regs(1989), ZN => n1228);
   U1628 : NAND3_X1 port map( A1 => n1230, A2 => n1229, A3 => n1228, ZN => 
                           curr_proc_regs(453));
   U1629 : NAND2_X1 port map( A1 => regs(966), A2 => n18, ZN => n1233);
   U1630 : AOI22_X1 port map( A1 => n32, A2 => regs(1478), B1 => n3, B2 => 
                           regs(454), ZN => n1232);
   U1631 : AOI22_X1 port map( A1 => n45, A2 => regs(2502), B1 => n36, B2 => 
                           regs(1990), ZN => n1231);
   U1632 : NAND3_X1 port map( A1 => n1233, A2 => n1232, A3 => n1231, ZN => 
                           curr_proc_regs(454));
   U1633 : NAND2_X1 port map( A1 => regs(967), A2 => n24, ZN => n1236);
   U1634 : AOI22_X1 port map( A1 => n32, A2 => regs(1479), B1 => n3, B2 => 
                           regs(455), ZN => n1235);
   U1635 : AOI22_X1 port map( A1 => n15, A2 => regs(2503), B1 => n4, B2 => 
                           regs(1991), ZN => n1234);
   U1636 : NAND3_X1 port map( A1 => n1236, A2 => n1235, A3 => n1234, ZN => 
                           curr_proc_regs(455));
   U1637 : NAND2_X1 port map( A1 => regs(968), A2 => n24, ZN => n1239);
   U1638 : AOI22_X1 port map( A1 => n32, A2 => regs(1480), B1 => n29, B2 => 
                           regs(456), ZN => n1238);
   U1639 : AOI22_X1 port map( A1 => n15, A2 => regs(2504), B1 => n4, B2 => 
                           regs(1992), ZN => n1237);
   U1640 : NAND3_X1 port map( A1 => n1239, A2 => n1238, A3 => n1237, ZN => 
                           curr_proc_regs(456));
   U1641 : NAND2_X1 port map( A1 => regs(969), A2 => n18, ZN => n1242);
   U1642 : AOI22_X1 port map( A1 => n32, A2 => regs(1481), B1 => n29, B2 => 
                           regs(457), ZN => n1241);
   U1643 : AOI22_X1 port map( A1 => n15, A2 => regs(2505), B1 => n38, B2 => 
                           regs(1993), ZN => n1240);
   U1644 : NAND3_X1 port map( A1 => n1242, A2 => n1241, A3 => n1240, ZN => 
                           curr_proc_regs(457));
   U1645 : NAND2_X1 port map( A1 => regs(970), A2 => n18, ZN => n1245);
   U1646 : AOI22_X1 port map( A1 => n32, A2 => regs(1482), B1 => n1586, B2 => 
                           regs(458), ZN => n1244);
   U1647 : AOI22_X1 port map( A1 => n15, A2 => regs(2506), B1 => n33, B2 => 
                           regs(1994), ZN => n1243);
   U1648 : NAND3_X1 port map( A1 => n1245, A2 => n1244, A3 => n1243, ZN => 
                           curr_proc_regs(458));
   U1649 : NAND2_X1 port map( A1 => regs(971), A2 => n18, ZN => n1248);
   U1650 : AOI22_X1 port map( A1 => n32, A2 => regs(1483), B1 => n8, B2 => 
                           regs(459), ZN => n1247);
   U1651 : AOI22_X1 port map( A1 => n15, A2 => regs(2507), B1 => n37, B2 => 
                           regs(1995), ZN => n1246);
   U1652 : NAND3_X1 port map( A1 => n1248, A2 => n1247, A3 => n1246, ZN => 
                           curr_proc_regs(459));
   U1653 : NAND2_X1 port map( A1 => regs(557), A2 => n24, ZN => n1251);
   U1654 : AOI22_X1 port map( A1 => n32, A2 => regs(1069), B1 => n8, B2 => 
                           regs(45), ZN => n1250);
   U1655 : AOI22_X1 port map( A1 => n45, A2 => regs(2093), B1 => n33, B2 => 
                           regs(1581), ZN => n1249);
   U1656 : NAND3_X1 port map( A1 => n1251, A2 => n1250, A3 => n1249, ZN => 
                           curr_proc_regs(45));
   U1657 : NAND2_X1 port map( A1 => regs(972), A2 => n18, ZN => n1254);
   U1658 : AOI22_X1 port map( A1 => n32, A2 => regs(1484), B1 => n1586, B2 => 
                           regs(460), ZN => n1253);
   U1659 : AOI22_X1 port map( A1 => n45, A2 => regs(2508), B1 => n33, B2 => 
                           regs(1996), ZN => n1252);
   U1660 : NAND3_X1 port map( A1 => n1254, A2 => n1253, A3 => n1252, ZN => 
                           curr_proc_regs(460));
   U1661 : NAND2_X1 port map( A1 => regs(973), A2 => n24, ZN => n1257);
   U1662 : AOI22_X1 port map( A1 => n32, A2 => regs(1485), B1 => n28, B2 => 
                           regs(461), ZN => n1256);
   U1663 : AOI22_X1 port map( A1 => n15, A2 => regs(2509), B1 => n38, B2 => 
                           regs(1997), ZN => n1255);
   U1664 : NAND3_X1 port map( A1 => n1257, A2 => n1256, A3 => n1255, ZN => 
                           curr_proc_regs(461));
   U1665 : NAND2_X1 port map( A1 => regs(974), A2 => n18, ZN => n1260);
   U1666 : AOI22_X1 port map( A1 => n32, A2 => regs(1486), B1 => n8, B2 => 
                           regs(462), ZN => n1259);
   U1667 : AOI22_X1 port map( A1 => n15, A2 => regs(2510), B1 => n4, B2 => 
                           regs(1998), ZN => n1258);
   U1668 : NAND3_X1 port map( A1 => n1260, A2 => n1259, A3 => n1258, ZN => 
                           curr_proc_regs(462));
   U1669 : NAND2_X1 port map( A1 => regs(975), A2 => n24, ZN => n1263);
   U1670 : AOI22_X1 port map( A1 => n32, A2 => regs(1487), B1 => n8, B2 => 
                           regs(463), ZN => n1262);
   U1671 : AOI22_X1 port map( A1 => n15, A2 => regs(2511), B1 => n4, B2 => 
                           regs(1999), ZN => n1261);
   U1672 : NAND3_X1 port map( A1 => n1263, A2 => n1262, A3 => n1261, ZN => 
                           curr_proc_regs(463));
   U1673 : NAND2_X1 port map( A1 => regs(976), A2 => n18, ZN => n1266);
   U1674 : AOI22_X1 port map( A1 => n32, A2 => regs(1488), B1 => n29, B2 => 
                           regs(464), ZN => n1265);
   U1675 : AOI22_X1 port map( A1 => n45, A2 => regs(2512), B1 => n38, B2 => 
                           regs(2000), ZN => n1264);
   U1676 : NAND3_X1 port map( A1 => n1266, A2 => n1265, A3 => n1264, ZN => 
                           curr_proc_regs(464));
   U1677 : NAND2_X1 port map( A1 => regs(977), A2 => n24, ZN => n1269);
   U1678 : AOI22_X1 port map( A1 => n32, A2 => regs(1489), B1 => n28, B2 => 
                           regs(465), ZN => n1268);
   U1679 : AOI22_X1 port map( A1 => n15, A2 => regs(2513), B1 => n4, B2 => 
                           regs(2001), ZN => n1267);
   U1680 : NAND3_X1 port map( A1 => n1269, A2 => n1268, A3 => n1267, ZN => 
                           curr_proc_regs(465));
   U1681 : NAND2_X1 port map( A1 => regs(978), A2 => n18, ZN => n1272);
   U1682 : AOI22_X1 port map( A1 => n32, A2 => regs(1490), B1 => n8, B2 => 
                           regs(466), ZN => n1271);
   U1683 : AOI22_X1 port map( A1 => n15, A2 => regs(2514), B1 => n4, B2 => 
                           regs(2002), ZN => n1270);
   U1684 : NAND3_X1 port map( A1 => n1272, A2 => n1271, A3 => n1270, ZN => 
                           curr_proc_regs(466));
   U1685 : NAND2_X1 port map( A1 => regs(979), A2 => n7, ZN => n1275);
   U1686 : AOI22_X1 port map( A1 => n32, A2 => regs(1491), B1 => n3, B2 => 
                           regs(467), ZN => n1274);
   U1687 : AOI22_X1 port map( A1 => n15, A2 => regs(2515), B1 => n37, B2 => 
                           regs(2003), ZN => n1273);
   U1688 : NAND3_X1 port map( A1 => n1275, A2 => n1274, A3 => n1273, ZN => 
                           curr_proc_regs(467));
   U1689 : NAND2_X1 port map( A1 => regs(980), A2 => n20, ZN => n1278);
   U1690 : AOI22_X1 port map( A1 => n32, A2 => regs(1492), B1 => n3, B2 => 
                           regs(468), ZN => n1277);
   U1691 : AOI22_X1 port map( A1 => n45, A2 => regs(2516), B1 => n33, B2 => 
                           regs(2004), ZN => n1276);
   U1692 : NAND3_X1 port map( A1 => n1278, A2 => n1277, A3 => n1276, ZN => 
                           curr_proc_regs(468));
   U1693 : NAND2_X1 port map( A1 => regs(981), A2 => n1585, ZN => n1281);
   U1694 : AOI22_X1 port map( A1 => n32, A2 => regs(1493), B1 => n3, B2 => 
                           regs(469), ZN => n1280);
   U1695 : AOI22_X1 port map( A1 => n45, A2 => regs(2517), B1 => n36, B2 => 
                           regs(2005), ZN => n1279);
   U1696 : NAND3_X1 port map( A1 => n1281, A2 => n1280, A3 => n1279, ZN => 
                           curr_proc_regs(469));
   U1697 : NAND2_X1 port map( A1 => regs(558), A2 => n18, ZN => n1284);
   U1698 : AOI22_X1 port map( A1 => n32, A2 => regs(1070), B1 => n3, B2 => 
                           regs(46), ZN => n1283);
   U1699 : AOI22_X1 port map( A1 => n40, A2 => regs(2094), B1 => n4, B2 => 
                           regs(1582), ZN => n1282);
   U1700 : NAND3_X1 port map( A1 => n1284, A2 => n1283, A3 => n1282, ZN => 
                           curr_proc_regs(46));
   U1701 : NAND2_X1 port map( A1 => regs(982), A2 => n1, ZN => n1287);
   U1702 : AOI22_X1 port map( A1 => n32, A2 => regs(1494), B1 => n3, B2 => 
                           regs(470), ZN => n1286);
   U1703 : AOI22_X1 port map( A1 => n15, A2 => regs(2518), B1 => n37, B2 => 
                           regs(2006), ZN => n1285);
   U1704 : NAND3_X1 port map( A1 => n1287, A2 => n1286, A3 => n1285, ZN => 
                           curr_proc_regs(470));
   U1705 : NAND2_X1 port map( A1 => regs(983), A2 => n22, ZN => n1290);
   U1706 : AOI22_X1 port map( A1 => n32, A2 => regs(1495), B1 => n3, B2 => 
                           regs(471), ZN => n1289);
   U1707 : AOI22_X1 port map( A1 => n15, A2 => regs(2519), B1 => n33, B2 => 
                           regs(2007), ZN => n1288);
   U1708 : NAND3_X1 port map( A1 => n1290, A2 => n1289, A3 => n1288, ZN => 
                           curr_proc_regs(471));
   U1709 : NAND2_X1 port map( A1 => regs(984), A2 => n1585, ZN => n1293);
   U1710 : AOI22_X1 port map( A1 => n32, A2 => regs(1496), B1 => n31, B2 => 
                           regs(472), ZN => n1292);
   U1711 : AOI22_X1 port map( A1 => n45, A2 => regs(2520), B1 => n36, B2 => 
                           regs(2008), ZN => n1291);
   U1712 : NAND3_X1 port map( A1 => n1293, A2 => n1292, A3 => n1291, ZN => 
                           curr_proc_regs(472));
   U1713 : NAND2_X1 port map( A1 => regs(985), A2 => n7, ZN => n1296);
   U1714 : AOI22_X1 port map( A1 => n32, A2 => regs(1497), B1 => n1586, B2 => 
                           regs(473), ZN => n1295);
   U1715 : AOI22_X1 port map( A1 => n40, A2 => regs(2521), B1 => n33, B2 => 
                           regs(2009), ZN => n1294);
   U1716 : NAND3_X1 port map( A1 => n1296, A2 => n1295, A3 => n1294, ZN => 
                           curr_proc_regs(473));
   U1717 : NAND2_X1 port map( A1 => regs(986), A2 => n1, ZN => n1299);
   U1718 : AOI22_X1 port map( A1 => n32, A2 => regs(1498), B1 => n1586, B2 => 
                           regs(474), ZN => n1298);
   U1719 : AOI22_X1 port map( A1 => n15, A2 => regs(2522), B1 => n33, B2 => 
                           regs(2010), ZN => n1297);
   U1720 : NAND3_X1 port map( A1 => n1299, A2 => n1298, A3 => n1297, ZN => 
                           curr_proc_regs(474));
   U1721 : NAND2_X1 port map( A1 => regs(987), A2 => n22, ZN => n1302);
   U1722 : AOI22_X1 port map( A1 => n32, A2 => regs(1499), B1 => n1586, B2 => 
                           regs(475), ZN => n1301);
   U1723 : AOI22_X1 port map( A1 => n15, A2 => regs(2523), B1 => n33, B2 => 
                           regs(2011), ZN => n1300);
   U1724 : NAND3_X1 port map( A1 => n1302, A2 => n1301, A3 => n1300, ZN => 
                           curr_proc_regs(475));
   U1725 : NAND2_X1 port map( A1 => regs(988), A2 => n1585, ZN => n1305);
   U1726 : AOI22_X1 port map( A1 => n32, A2 => regs(1500), B1 => n1586, B2 => 
                           regs(476), ZN => n1304);
   U1727 : AOI22_X1 port map( A1 => n45, A2 => regs(2524), B1 => n33, B2 => 
                           regs(2012), ZN => n1303);
   U1728 : NAND3_X1 port map( A1 => n1305, A2 => n1304, A3 => n1303, ZN => 
                           curr_proc_regs(476));
   U1729 : NAND2_X1 port map( A1 => regs(989), A2 => n1, ZN => n1308);
   U1730 : AOI22_X1 port map( A1 => n32, A2 => regs(1501), B1 => n8, B2 => 
                           regs(477), ZN => n1307);
   U1731 : AOI22_X1 port map( A1 => n40, A2 => regs(2525), B1 => n4, B2 => 
                           regs(2013), ZN => n1306);
   U1732 : NAND3_X1 port map( A1 => n1308, A2 => n1307, A3 => n1306, ZN => 
                           curr_proc_regs(477));
   U1733 : NAND2_X1 port map( A1 => regs(990), A2 => n1, ZN => n1311);
   U1734 : AOI22_X1 port map( A1 => n32, A2 => regs(1502), B1 => n8, B2 => 
                           regs(478), ZN => n1310);
   U1735 : AOI22_X1 port map( A1 => n15, A2 => regs(2526), B1 => n4, B2 => 
                           regs(2014), ZN => n1309);
   U1736 : NAND3_X1 port map( A1 => n1311, A2 => n1310, A3 => n1309, ZN => 
                           curr_proc_regs(478));
   U1737 : NAND2_X1 port map( A1 => regs(991), A2 => n1, ZN => n1314);
   U1738 : AOI22_X1 port map( A1 => n32, A2 => regs(1503), B1 => n8, B2 => 
                           regs(479), ZN => n1313);
   U1739 : AOI22_X1 port map( A1 => n15, A2 => regs(2527), B1 => n4, B2 => 
                           regs(2015), ZN => n1312);
   U1740 : NAND3_X1 port map( A1 => n1314, A2 => n1313, A3 => n1312, ZN => 
                           curr_proc_regs(479));
   U1741 : NAND2_X1 port map( A1 => regs(559), A2 => n1, ZN => n1317);
   U1742 : AOI22_X1 port map( A1 => n32, A2 => regs(1071), B1 => n8, B2 => 
                           regs(47), ZN => n1316);
   U1743 : AOI22_X1 port map( A1 => n15, A2 => regs(2095), B1 => n4, B2 => 
                           regs(1583), ZN => n1315);
   U1744 : NAND3_X1 port map( A1 => n1317, A2 => n1316, A3 => n1315, ZN => 
                           curr_proc_regs(47));
   U1745 : NAND2_X1 port map( A1 => regs(992), A2 => n1, ZN => n1320);
   U1746 : AOI22_X1 port map( A1 => n32, A2 => regs(1504), B1 => n8, B2 => 
                           regs(480), ZN => n1319);
   U1747 : AOI22_X1 port map( A1 => n15, A2 => regs(2528), B1 => n4, B2 => 
                           regs(2016), ZN => n1318);
   U1748 : NAND3_X1 port map( A1 => n1320, A2 => n1319, A3 => n1318, ZN => 
                           curr_proc_regs(480));
   U1749 : NAND2_X1 port map( A1 => regs(993), A2 => n1, ZN => n1323);
   U1750 : AOI22_X1 port map( A1 => n32, A2 => regs(1505), B1 => n8, B2 => 
                           regs(481), ZN => n1322);
   U1751 : AOI22_X1 port map( A1 => n15, A2 => regs(2529), B1 => n4, B2 => 
                           regs(2017), ZN => n1321);
   U1752 : NAND3_X1 port map( A1 => n1323, A2 => n1322, A3 => n1321, ZN => 
                           curr_proc_regs(481));
   U1753 : NAND2_X1 port map( A1 => regs(994), A2 => n1, ZN => n1326);
   U1754 : AOI22_X1 port map( A1 => n32, A2 => regs(1506), B1 => n8, B2 => 
                           regs(482), ZN => n1325);
   U1755 : AOI22_X1 port map( A1 => n15, A2 => regs(2530), B1 => n4, B2 => 
                           regs(2018), ZN => n1324);
   U1756 : NAND3_X1 port map( A1 => n1326, A2 => n1325, A3 => n1324, ZN => 
                           curr_proc_regs(482));
   U1757 : NAND2_X1 port map( A1 => regs(995), A2 => n1, ZN => n1329);
   U1758 : AOI22_X1 port map( A1 => n32, A2 => regs(1507), B1 => n8, B2 => 
                           regs(483), ZN => n1328);
   U1759 : AOI22_X1 port map( A1 => n15, A2 => regs(2531), B1 => n4, B2 => 
                           regs(2019), ZN => n1327);
   U1760 : NAND3_X1 port map( A1 => n1329, A2 => n1328, A3 => n1327, ZN => 
                           curr_proc_regs(483));
   U1761 : NAND2_X1 port map( A1 => regs(996), A2 => n1, ZN => n1332);
   U1762 : AOI22_X1 port map( A1 => n32, A2 => regs(1508), B1 => n8, B2 => 
                           regs(484), ZN => n1331);
   U1763 : AOI22_X1 port map( A1 => n15, A2 => regs(2532), B1 => n4, B2 => 
                           regs(2020), ZN => n1330);
   U1764 : NAND3_X1 port map( A1 => n1332, A2 => n1331, A3 => n1330, ZN => 
                           curr_proc_regs(484));
   U1765 : NAND2_X1 port map( A1 => regs(997), A2 => n1, ZN => n1335);
   U1766 : AOI22_X1 port map( A1 => n32, A2 => regs(1509), B1 => n8, B2 => 
                           regs(485), ZN => n1334);
   U1767 : AOI22_X1 port map( A1 => n15, A2 => regs(2533), B1 => n4, B2 => 
                           regs(2021), ZN => n1333);
   U1768 : NAND3_X1 port map( A1 => n1335, A2 => n1334, A3 => n1333, ZN => 
                           curr_proc_regs(485));
   U1769 : NAND2_X1 port map( A1 => regs(998), A2 => n1, ZN => n1338);
   U1770 : AOI22_X1 port map( A1 => n32, A2 => regs(1510), B1 => n8, B2 => 
                           regs(486), ZN => n1337);
   U1771 : AOI22_X1 port map( A1 => n15, A2 => regs(2534), B1 => n4, B2 => 
                           regs(2022), ZN => n1336);
   U1772 : NAND3_X1 port map( A1 => n1338, A2 => n1337, A3 => n1336, ZN => 
                           curr_proc_regs(486));
   U1773 : NAND2_X1 port map( A1 => regs(999), A2 => n18, ZN => n1341);
   U1774 : AOI22_X1 port map( A1 => n32, A2 => regs(1511), B1 => n8, B2 => 
                           regs(487), ZN => n1340);
   U1775 : AOI22_X1 port map( A1 => n15, A2 => regs(2535), B1 => n4, B2 => 
                           regs(2023), ZN => n1339);
   U1776 : NAND3_X1 port map( A1 => n1341, A2 => n1340, A3 => n1339, ZN => 
                           curr_proc_regs(487));
   U1777 : NAND2_X1 port map( A1 => regs(1000), A2 => n18, ZN => n1344);
   U1778 : AOI22_X1 port map( A1 => n32, A2 => regs(1512), B1 => n31, B2 => 
                           regs(488), ZN => n1343);
   U1779 : AOI22_X1 port map( A1 => n15, A2 => regs(2536), B1 => n37, B2 => 
                           regs(2024), ZN => n1342);
   U1780 : NAND3_X1 port map( A1 => n1344, A2 => n1343, A3 => n1342, ZN => 
                           curr_proc_regs(488));
   U1781 : NAND2_X1 port map( A1 => regs(1001), A2 => n18, ZN => n1347);
   U1782 : AOI22_X1 port map( A1 => n32, A2 => regs(1513), B1 => n3, B2 => 
                           regs(489), ZN => n1346);
   U1783 : AOI22_X1 port map( A1 => n15, A2 => regs(2537), B1 => n37, B2 => 
                           regs(2025), ZN => n1345);
   U1784 : NAND3_X1 port map( A1 => n1347, A2 => n1346, A3 => n1345, ZN => 
                           curr_proc_regs(489));
   U1785 : NAND2_X1 port map( A1 => regs(560), A2 => n18, ZN => n1350);
   U1786 : AOI22_X1 port map( A1 => n32, A2 => regs(1072), B1 => n3, B2 => 
                           regs(48), ZN => n1349);
   U1787 : AOI22_X1 port map( A1 => n15, A2 => regs(2096), B1 => n36, B2 => 
                           regs(1584), ZN => n1348);
   U1788 : NAND3_X1 port map( A1 => n1350, A2 => n1349, A3 => n1348, ZN => 
                           curr_proc_regs(48));
   U1789 : NAND2_X1 port map( A1 => regs(1002), A2 => n18, ZN => n1353);
   U1790 : AOI22_X1 port map( A1 => n32, A2 => regs(1514), B1 => n3, B2 => 
                           regs(490), ZN => n1352);
   U1791 : AOI22_X1 port map( A1 => n15, A2 => regs(2538), B1 => n4, B2 => 
                           regs(2026), ZN => n1351);
   U1792 : NAND3_X1 port map( A1 => n1353, A2 => n1352, A3 => n1351, ZN => 
                           curr_proc_regs(490));
   U1793 : NAND2_X1 port map( A1 => regs(1003), A2 => n18, ZN => n1356);
   U1794 : AOI22_X1 port map( A1 => n32, A2 => regs(1515), B1 => n1586, B2 => 
                           regs(491), ZN => n1355);
   U1795 : AOI22_X1 port map( A1 => n15, A2 => regs(2539), B1 => n4, B2 => 
                           regs(2027), ZN => n1354);
   U1796 : NAND3_X1 port map( A1 => n1356, A2 => n1355, A3 => n1354, ZN => 
                           curr_proc_regs(491));
   U1797 : NAND2_X1 port map( A1 => regs(1004), A2 => n18, ZN => n1359);
   U1798 : AOI22_X1 port map( A1 => n32, A2 => regs(1516), B1 => n29, B2 => 
                           regs(492), ZN => n1358);
   U1799 : AOI22_X1 port map( A1 => n15, A2 => regs(2540), B1 => n38, B2 => 
                           regs(2028), ZN => n1357);
   U1800 : NAND3_X1 port map( A1 => n1359, A2 => n1358, A3 => n1357, ZN => 
                           curr_proc_regs(492));
   U1801 : NAND2_X1 port map( A1 => regs(1005), A2 => n18, ZN => n1362);
   U1802 : AOI22_X1 port map( A1 => n32, A2 => regs(1517), B1 => n1586, B2 => 
                           regs(493), ZN => n1361);
   U1803 : AOI22_X1 port map( A1 => n15, A2 => regs(2541), B1 => n33, B2 => 
                           regs(2029), ZN => n1360);
   U1804 : NAND3_X1 port map( A1 => n1362, A2 => n1361, A3 => n1360, ZN => 
                           curr_proc_regs(493));
   U1805 : NAND2_X1 port map( A1 => regs(1006), A2 => n18, ZN => n1365);
   U1806 : AOI22_X1 port map( A1 => n32, A2 => regs(1518), B1 => n29, B2 => 
                           regs(494), ZN => n1364);
   U1807 : AOI22_X1 port map( A1 => n15, A2 => regs(2542), B1 => n38, B2 => 
                           regs(2030), ZN => n1363);
   U1808 : NAND3_X1 port map( A1 => n1365, A2 => n1364, A3 => n1363, ZN => 
                           curr_proc_regs(494));
   U1809 : NAND2_X1 port map( A1 => regs(1007), A2 => n18, ZN => n1368);
   U1810 : AOI22_X1 port map( A1 => n32, A2 => regs(1519), B1 => n1586, B2 => 
                           regs(495), ZN => n1367);
   U1811 : AOI22_X1 port map( A1 => n15, A2 => regs(2543), B1 => n33, B2 => 
                           regs(2031), ZN => n1366);
   U1812 : NAND3_X1 port map( A1 => n1368, A2 => n1367, A3 => n1366, ZN => 
                           curr_proc_regs(495));
   U1813 : NAND2_X1 port map( A1 => regs(1008), A2 => n18, ZN => n1371);
   U1814 : AOI22_X1 port map( A1 => n32, A2 => regs(1520), B1 => n1586, B2 => 
                           regs(496), ZN => n1370);
   U1815 : AOI22_X1 port map( A1 => n15, A2 => regs(2544), B1 => n33, B2 => 
                           regs(2032), ZN => n1369);
   U1816 : NAND3_X1 port map( A1 => n1371, A2 => n1370, A3 => n1369, ZN => 
                           curr_proc_regs(496));
   U1817 : NAND2_X1 port map( A1 => regs(1009), A2 => n6, ZN => n1374);
   U1818 : AOI22_X1 port map( A1 => n32, A2 => regs(1521), B1 => n28, B2 => 
                           regs(497), ZN => n1373);
   U1819 : AOI22_X1 port map( A1 => n15, A2 => regs(2545), B1 => n4, B2 => 
                           regs(2033), ZN => n1372);
   U1820 : NAND3_X1 port map( A1 => n1374, A2 => n1373, A3 => n1372, ZN => 
                           curr_proc_regs(497));
   U1821 : NAND2_X1 port map( A1 => regs(1010), A2 => n7, ZN => n1377);
   U1822 : AOI22_X1 port map( A1 => n32, A2 => regs(1522), B1 => n28, B2 => 
                           regs(498), ZN => n1376);
   U1823 : AOI22_X1 port map( A1 => n15, A2 => regs(2546), B1 => n4, B2 => 
                           regs(2034), ZN => n1375);
   U1824 : NAND3_X1 port map( A1 => n1377, A2 => n1376, A3 => n1375, ZN => 
                           curr_proc_regs(498));
   U1825 : NAND2_X1 port map( A1 => regs(1011), A2 => n2, ZN => n1380);
   U1826 : AOI22_X1 port map( A1 => n32, A2 => regs(1523), B1 => n28, B2 => 
                           regs(499), ZN => n1379);
   U1827 : AOI22_X1 port map( A1 => n45, A2 => regs(2547), B1 => n38, B2 => 
                           regs(2035), ZN => n1378);
   U1828 : NAND3_X1 port map( A1 => n1380, A2 => n1379, A3 => n1378, ZN => 
                           curr_proc_regs(499));
   U1829 : NAND2_X1 port map( A1 => regs(561), A2 => n21, ZN => n1383);
   U1830 : AOI22_X1 port map( A1 => n32, A2 => regs(1073), B1 => n28, B2 => 
                           regs(49), ZN => n1382);
   U1831 : AOI22_X1 port map( A1 => n45, A2 => regs(2097), B1 => n4, B2 => 
                           regs(1585), ZN => n1381);
   U1832 : NAND3_X1 port map( A1 => n1383, A2 => n1382, A3 => n1381, ZN => 
                           curr_proc_regs(49));
   U1833 : NAND2_X1 port map( A1 => regs(516), A2 => n22, ZN => n1386);
   U1834 : AOI22_X1 port map( A1 => n32, A2 => regs(1028), B1 => n28, B2 => 
                           regs(4), ZN => n1385);
   U1835 : AOI22_X1 port map( A1 => n45, A2 => regs(2052), B1 => n4, B2 => 
                           regs(1540), ZN => n1384);
   U1836 : NAND3_X1 port map( A1 => n1386, A2 => n1385, A3 => n1384, ZN => 
                           curr_proc_regs(4));
   U1837 : NAND2_X1 port map( A1 => regs(1012), A2 => n20, ZN => n1389);
   U1838 : AOI22_X1 port map( A1 => n32, A2 => regs(1524), B1 => n28, B2 => 
                           regs(500), ZN => n1388);
   U1839 : AOI22_X1 port map( A1 => n45, A2 => regs(2548), B1 => n38, B2 => 
                           regs(2036), ZN => n1387);
   U1840 : NAND3_X1 port map( A1 => n1389, A2 => n1388, A3 => n1387, ZN => 
                           curr_proc_regs(500));
   U1841 : NAND2_X1 port map( A1 => regs(1013), A2 => n1585, ZN => n1392);
   U1842 : AOI22_X1 port map( A1 => n32, A2 => regs(1525), B1 => n28, B2 => 
                           regs(501), ZN => n1391);
   U1843 : AOI22_X1 port map( A1 => n15, A2 => regs(2549), B1 => n4, B2 => 
                           regs(2037), ZN => n1390);
   U1844 : NAND3_X1 port map( A1 => n1392, A2 => n1391, A3 => n1390, ZN => 
                           curr_proc_regs(501));
   U1845 : NAND2_X1 port map( A1 => regs(1014), A2 => n1585, ZN => n1395);
   U1846 : AOI22_X1 port map( A1 => n32, A2 => regs(1526), B1 => n28, B2 => 
                           regs(502), ZN => n1394);
   U1847 : AOI22_X1 port map( A1 => n45, A2 => regs(2550), B1 => n4, B2 => 
                           regs(2038), ZN => n1393);
   U1848 : NAND3_X1 port map( A1 => n1395, A2 => n1394, A3 => n1393, ZN => 
                           curr_proc_regs(502));
   U1849 : NAND2_X1 port map( A1 => regs(1015), A2 => n19, ZN => n1398);
   U1850 : AOI22_X1 port map( A1 => n32, A2 => regs(1527), B1 => n28, B2 => 
                           regs(503), ZN => n1397);
   U1851 : AOI22_X1 port map( A1 => n45, A2 => regs(2551), B1 => n38, B2 => 
                           regs(2039), ZN => n1396);
   U1852 : NAND3_X1 port map( A1 => n1398, A2 => n1397, A3 => n1396, ZN => 
                           curr_proc_regs(503));
   U1853 : NAND2_X1 port map( A1 => regs(1016), A2 => n23, ZN => n1401);
   U1854 : AOI22_X1 port map( A1 => n32, A2 => regs(1528), B1 => n28, B2 => 
                           regs(504), ZN => n1400);
   U1855 : AOI22_X1 port map( A1 => n45, A2 => regs(2552), B1 => n4, B2 => 
                           regs(2040), ZN => n1399);
   U1856 : NAND3_X1 port map( A1 => n1401, A2 => n1400, A3 => n1399, ZN => 
                           curr_proc_regs(504));
   U1857 : NAND2_X1 port map( A1 => regs(1017), A2 => n6, ZN => n1404);
   U1858 : AOI22_X1 port map( A1 => n32, A2 => regs(1529), B1 => n28, B2 => 
                           regs(505), ZN => n1403);
   U1859 : AOI22_X1 port map( A1 => n45, A2 => regs(2553), B1 => n4, B2 => 
                           regs(2041), ZN => n1402);
   U1860 : NAND3_X1 port map( A1 => n1404, A2 => n1403, A3 => n1402, ZN => 
                           curr_proc_regs(505));
   U1861 : NAND2_X1 port map( A1 => regs(1018), A2 => n1585, ZN => n1407);
   U1862 : AOI22_X1 port map( A1 => n32, A2 => regs(1530), B1 => n28, B2 => 
                           regs(506), ZN => n1406);
   U1863 : AOI22_X1 port map( A1 => n15, A2 => regs(2554), B1 => n36, B2 => 
                           regs(2042), ZN => n1405);
   U1864 : NAND3_X1 port map( A1 => n1407, A2 => n1406, A3 => n1405, ZN => 
                           curr_proc_regs(506));
   U1865 : NAND2_X1 port map( A1 => regs(1019), A2 => n1585, ZN => n1410);
   U1866 : AOI22_X1 port map( A1 => n32, A2 => regs(1531), B1 => n8, B2 => 
                           regs(507), ZN => n1409);
   U1867 : AOI22_X1 port map( A1 => n46, A2 => regs(2555), B1 => n4, B2 => 
                           regs(2043), ZN => n1408);
   U1868 : NAND3_X1 port map( A1 => n1410, A2 => n1409, A3 => n1408, ZN => 
                           curr_proc_regs(507));
   U1869 : NAND2_X1 port map( A1 => regs(1020), A2 => n1585, ZN => n1413);
   U1870 : AOI22_X1 port map( A1 => n32, A2 => regs(1532), B1 => n28, B2 => 
                           regs(508), ZN => n1412);
   U1871 : AOI22_X1 port map( A1 => n46, A2 => regs(2556), B1 => n36, B2 => 
                           regs(2044), ZN => n1411);
   U1872 : NAND3_X1 port map( A1 => n1413, A2 => n1412, A3 => n1411, ZN => 
                           curr_proc_regs(508));
   U1873 : NAND2_X1 port map( A1 => regs(1021), A2 => n1585, ZN => n1416);
   U1874 : AOI22_X1 port map( A1 => n32, A2 => regs(1533), B1 => n8, B2 => 
                           regs(509), ZN => n1415);
   U1875 : AOI22_X1 port map( A1 => n46, A2 => regs(2557), B1 => n4, B2 => 
                           regs(2045), ZN => n1414);
   U1876 : NAND3_X1 port map( A1 => n1416, A2 => n1415, A3 => n1414, ZN => 
                           curr_proc_regs(509));
   U1877 : NAND2_X1 port map( A1 => regs(562), A2 => n1585, ZN => n1419);
   U1878 : AOI22_X1 port map( A1 => n32, A2 => regs(1074), B1 => n28, B2 => 
                           regs(50), ZN => n1418);
   U1879 : AOI22_X1 port map( A1 => n46, A2 => regs(2098), B1 => n36, B2 => 
                           regs(1586), ZN => n1417);
   U1880 : NAND3_X1 port map( A1 => n1419, A2 => n1418, A3 => n1417, ZN => 
                           curr_proc_regs(50));
   U1881 : NAND2_X1 port map( A1 => regs(1022), A2 => n1585, ZN => n1422);
   U1882 : AOI22_X1 port map( A1 => n32, A2 => regs(1534), B1 => n8, B2 => 
                           regs(510), ZN => n1421);
   U1883 : AOI22_X1 port map( A1 => n40, A2 => regs(2558), B1 => n4, B2 => 
                           regs(2046), ZN => n1420);
   U1884 : NAND3_X1 port map( A1 => n1422, A2 => n1421, A3 => n1420, ZN => 
                           curr_proc_regs(510));
   U1885 : NAND2_X1 port map( A1 => regs(1023), A2 => n1585, ZN => n1425);
   U1886 : AOI22_X1 port map( A1 => n32, A2 => regs(1535), B1 => n28, B2 => 
                           regs(511), ZN => n1424);
   U1887 : AOI22_X1 port map( A1 => n46, A2 => regs(2559), B1 => n36, B2 => 
                           regs(2047), ZN => n1423);
   U1888 : NAND3_X1 port map( A1 => n1425, A2 => n1424, A3 => n1423, ZN => 
                           curr_proc_regs(511));
   U1889 : NAND2_X1 port map( A1 => regs(563), A2 => n1585, ZN => n1428);
   U1890 : AOI22_X1 port map( A1 => n32, A2 => regs(1075), B1 => n8, B2 => 
                           regs(51), ZN => n1427);
   U1891 : AOI22_X1 port map( A1 => n46, A2 => regs(2099), B1 => n4, B2 => 
                           regs(1587), ZN => n1426);
   U1892 : NAND3_X1 port map( A1 => n1428, A2 => n1427, A3 => n1426, ZN => 
                           curr_proc_regs(51));
   U1893 : NAND2_X1 port map( A1 => regs(564), A2 => n1585, ZN => n1431);
   U1894 : AOI22_X1 port map( A1 => n32, A2 => regs(1076), B1 => n28, B2 => 
                           regs(52), ZN => n1430);
   U1895 : AOI22_X1 port map( A1 => n40, A2 => regs(2100), B1 => n36, B2 => 
                           regs(1588), ZN => n1429);
   U1896 : NAND3_X1 port map( A1 => n1431, A2 => n1430, A3 => n1429, ZN => 
                           curr_proc_regs(52));
   U1897 : NAND2_X1 port map( A1 => regs(565), A2 => n1585, ZN => n1434);
   U1898 : AOI22_X1 port map( A1 => n32, A2 => regs(1077), B1 => n8, B2 => 
                           regs(53), ZN => n1433);
   U1899 : AOI22_X1 port map( A1 => n10, A2 => regs(2101), B1 => n4, B2 => 
                           regs(1589), ZN => n1432);
   U1900 : NAND3_X1 port map( A1 => n1434, A2 => n1433, A3 => n1432, ZN => 
                           curr_proc_regs(53));
   U1901 : NAND2_X1 port map( A1 => regs(566), A2 => n1585, ZN => n1437);
   U1902 : AOI22_X1 port map( A1 => n32, A2 => regs(1078), B1 => n28, B2 => 
                           regs(54), ZN => n1436);
   U1903 : AOI22_X1 port map( A1 => n10, A2 => regs(2102), B1 => n36, B2 => 
                           regs(1590), ZN => n1435);
   U1904 : NAND3_X1 port map( A1 => n1437, A2 => n1436, A3 => n1435, ZN => 
                           curr_proc_regs(54));
   U1905 : NAND2_X1 port map( A1 => regs(567), A2 => n21, ZN => n1440);
   U1906 : AOI22_X1 port map( A1 => n32, A2 => regs(1079), B1 => n3, B2 => 
                           regs(55), ZN => n1439);
   U1907 : AOI22_X1 port map( A1 => n40, A2 => regs(2103), B1 => n36, B2 => 
                           regs(1591), ZN => n1438);
   U1908 : NAND3_X1 port map( A1 => n1440, A2 => n1439, A3 => n1438, ZN => 
                           curr_proc_regs(55));
   U1909 : NAND2_X1 port map( A1 => regs(568), A2 => n17, ZN => n1443);
   U1910 : AOI22_X1 port map( A1 => n32, A2 => regs(1080), B1 => n3, B2 => 
                           regs(56), ZN => n1442);
   U1911 : AOI22_X1 port map( A1 => n46, A2 => regs(2104), B1 => n36, B2 => 
                           regs(1592), ZN => n1441);
   U1912 : NAND3_X1 port map( A1 => n1443, A2 => n1442, A3 => n1441, ZN => 
                           curr_proc_regs(56));
   U1913 : NAND2_X1 port map( A1 => regs(569), A2 => n6, ZN => n1446);
   U1914 : AOI22_X1 port map( A1 => n32, A2 => regs(1081), B1 => n3, B2 => 
                           regs(57), ZN => n1445);
   U1915 : AOI22_X1 port map( A1 => n40, A2 => regs(2105), B1 => n36, B2 => 
                           regs(1593), ZN => n1444);
   U1916 : NAND3_X1 port map( A1 => n1446, A2 => n1445, A3 => n1444, ZN => 
                           curr_proc_regs(57));
   U1917 : NAND2_X1 port map( A1 => regs(570), A2 => n7, ZN => n1449);
   U1918 : AOI22_X1 port map( A1 => n32, A2 => regs(1082), B1 => n3, B2 => 
                           regs(58), ZN => n1448);
   U1919 : AOI22_X1 port map( A1 => n10, A2 => regs(2106), B1 => n36, B2 => 
                           regs(1594), ZN => n1447);
   U1920 : NAND3_X1 port map( A1 => n1449, A2 => n1448, A3 => n1447, ZN => 
                           curr_proc_regs(58));
   U1921 : NAND2_X1 port map( A1 => regs(571), A2 => n1, ZN => n1452);
   U1922 : AOI22_X1 port map( A1 => n32, A2 => regs(1083), B1 => n3, B2 => 
                           regs(59), ZN => n1451);
   U1923 : AOI22_X1 port map( A1 => n10, A2 => regs(2107), B1 => n36, B2 => 
                           regs(1595), ZN => n1450);
   U1924 : NAND3_X1 port map( A1 => n1452, A2 => n1451, A3 => n1450, ZN => 
                           curr_proc_regs(59));
   U1925 : NAND2_X1 port map( A1 => regs(517), A2 => n20, ZN => n1455);
   U1926 : AOI22_X1 port map( A1 => n32, A2 => regs(1029), B1 => n3, B2 => 
                           regs(5), ZN => n1454);
   U1927 : AOI22_X1 port map( A1 => n10, A2 => regs(2053), B1 => n36, B2 => 
                           regs(1541), ZN => n1453);
   U1928 : NAND3_X1 port map( A1 => n1455, A2 => n1454, A3 => n1453, ZN => 
                           curr_proc_regs(5));
   U1929 : NAND2_X1 port map( A1 => regs(572), A2 => n23, ZN => n1458);
   U1930 : AOI22_X1 port map( A1 => n32, A2 => regs(1084), B1 => n3, B2 => 
                           regs(60), ZN => n1457);
   U1931 : AOI22_X1 port map( A1 => n46, A2 => regs(2108), B1 => n36, B2 => 
                           regs(1596), ZN => n1456);
   U1932 : NAND3_X1 port map( A1 => n1458, A2 => n1457, A3 => n1456, ZN => 
                           curr_proc_regs(60));
   U1933 : NAND2_X1 port map( A1 => regs(573), A2 => n17, ZN => n1461);
   U1934 : AOI22_X1 port map( A1 => n32, A2 => regs(1085), B1 => n3, B2 => 
                           regs(61), ZN => n1460);
   U1935 : AOI22_X1 port map( A1 => n40, A2 => regs(2109), B1 => n36, B2 => 
                           regs(1597), ZN => n1459);
   U1936 : NAND3_X1 port map( A1 => n1461, A2 => n1460, A3 => n1459, ZN => 
                           curr_proc_regs(61));
   U1937 : NAND2_X1 port map( A1 => regs(574), A2 => n22, ZN => n1464);
   U1938 : AOI22_X1 port map( A1 => n32, A2 => regs(1086), B1 => n3, B2 => 
                           regs(62), ZN => n1463);
   U1939 : AOI22_X1 port map( A1 => n10, A2 => regs(2110), B1 => n36, B2 => 
                           regs(1598), ZN => n1462);
   U1940 : NAND3_X1 port map( A1 => n1464, A2 => n1463, A3 => n1462, ZN => 
                           curr_proc_regs(62));
   U1941 : NAND2_X1 port map( A1 => regs(575), A2 => n7, ZN => n1467);
   U1942 : AOI22_X1 port map( A1 => n32, A2 => regs(1087), B1 => n3, B2 => 
                           regs(63), ZN => n1466);
   U1943 : AOI22_X1 port map( A1 => n10, A2 => regs(2111), B1 => n36, B2 => 
                           regs(1599), ZN => n1465);
   U1944 : NAND3_X1 port map( A1 => n1467, A2 => n1466, A3 => n1465, ZN => 
                           curr_proc_regs(63));
   U1945 : NAND2_X1 port map( A1 => regs(576), A2 => n6, ZN => n1470);
   U1946 : AOI22_X1 port map( A1 => n32, A2 => regs(1088), B1 => n3, B2 => 
                           regs(64), ZN => n1469);
   U1947 : AOI22_X1 port map( A1 => n10, A2 => regs(2112), B1 => n36, B2 => 
                           regs(1600), ZN => n1468);
   U1948 : NAND3_X1 port map( A1 => n1470, A2 => n1469, A3 => n1468, ZN => 
                           curr_proc_regs(64));
   U1949 : NAND2_X1 port map( A1 => regs(577), A2 => n18, ZN => n1473);
   U1950 : AOI22_X1 port map( A1 => n32, A2 => regs(1089), B1 => n3, B2 => 
                           regs(65), ZN => n1472);
   U1951 : AOI22_X1 port map( A1 => n46, A2 => regs(2113), B1 => n4, B2 => 
                           regs(1601), ZN => n1471);
   U1952 : NAND3_X1 port map( A1 => n1473, A2 => n1472, A3 => n1471, ZN => 
                           curr_proc_regs(65));
   U1953 : NAND2_X1 port map( A1 => regs(578), A2 => n1585, ZN => n1476);
   U1954 : AOI22_X1 port map( A1 => n32, A2 => regs(1090), B1 => n3, B2 => 
                           regs(66), ZN => n1475);
   U1955 : AOI22_X1 port map( A1 => n46, A2 => regs(2114), B1 => n4, B2 => 
                           regs(1602), ZN => n1474);
   U1956 : NAND3_X1 port map( A1 => n1476, A2 => n1475, A3 => n1474, ZN => 
                           curr_proc_regs(66));
   U1957 : NAND2_X1 port map( A1 => regs(579), A2 => n2, ZN => n1479);
   U1958 : AOI22_X1 port map( A1 => n32, A2 => regs(1091), B1 => n3, B2 => 
                           regs(67), ZN => n1478);
   U1959 : AOI22_X1 port map( A1 => n40, A2 => regs(2115), B1 => n4, B2 => 
                           regs(1603), ZN => n1477);
   U1960 : NAND3_X1 port map( A1 => n1479, A2 => n1478, A3 => n1477, ZN => 
                           curr_proc_regs(67));
   U1961 : NAND2_X1 port map( A1 => regs(580), A2 => n1585, ZN => n1482);
   U1962 : AOI22_X1 port map( A1 => n32, A2 => regs(1092), B1 => n3, B2 => 
                           regs(68), ZN => n1481);
   U1963 : AOI22_X1 port map( A1 => n10, A2 => regs(2116), B1 => n4, B2 => 
                           regs(1604), ZN => n1480);
   U1964 : NAND3_X1 port map( A1 => n1482, A2 => n1481, A3 => n1480, ZN => 
                           curr_proc_regs(68));
   U1965 : NAND2_X1 port map( A1 => regs(581), A2 => n7, ZN => n1485);
   U1966 : AOI22_X1 port map( A1 => n32, A2 => regs(1093), B1 => n3, B2 => 
                           regs(69), ZN => n1484);
   U1967 : AOI22_X1 port map( A1 => n10, A2 => regs(2117), B1 => n4, B2 => 
                           regs(1605), ZN => n1483);
   U1968 : NAND3_X1 port map( A1 => n1485, A2 => n1484, A3 => n1483, ZN => 
                           curr_proc_regs(69));
   U1969 : NAND2_X1 port map( A1 => regs(518), A2 => n1585, ZN => n1488);
   U1970 : AOI22_X1 port map( A1 => n32, A2 => regs(1030), B1 => n3, B2 => 
                           regs(6), ZN => n1487);
   U1971 : AOI22_X1 port map( A1 => n46, A2 => regs(2054), B1 => n4, B2 => 
                           regs(1542), ZN => n1486);
   U1972 : NAND3_X1 port map( A1 => n1488, A2 => n1487, A3 => n1486, ZN => 
                           curr_proc_regs(6));
   U1973 : NAND2_X1 port map( A1 => regs(582), A2 => n21, ZN => n1491);
   U1974 : AOI22_X1 port map( A1 => n32, A2 => regs(1094), B1 => n3, B2 => 
                           regs(70), ZN => n1490);
   U1975 : AOI22_X1 port map( A1 => n40, A2 => regs(2118), B1 => n4, B2 => 
                           regs(1606), ZN => n1489);
   U1976 : NAND3_X1 port map( A1 => n1491, A2 => n1490, A3 => n1489, ZN => 
                           curr_proc_regs(70));
   U1977 : NAND2_X1 port map( A1 => regs(583), A2 => n1585, ZN => n1494);
   U1978 : AOI22_X1 port map( A1 => n32, A2 => regs(1095), B1 => n3, B2 => 
                           regs(71), ZN => n1493);
   U1979 : AOI22_X1 port map( A1 => n10, A2 => regs(2119), B1 => n4, B2 => 
                           regs(1607), ZN => n1492);
   U1980 : NAND3_X1 port map( A1 => n1494, A2 => n1493, A3 => n1492, ZN => 
                           curr_proc_regs(71));
   U1981 : NAND2_X1 port map( A1 => regs(584), A2 => n1585, ZN => n1497);
   U1982 : AOI22_X1 port map( A1 => n32, A2 => regs(1096), B1 => n3, B2 => 
                           regs(72), ZN => n1496);
   U1983 : AOI22_X1 port map( A1 => n10, A2 => regs(2120), B1 => n4, B2 => 
                           regs(1608), ZN => n1495);
   U1984 : NAND3_X1 port map( A1 => n1497, A2 => n1496, A3 => n1495, ZN => 
                           curr_proc_regs(72));
   U1985 : NAND2_X1 port map( A1 => regs(585), A2 => n20, ZN => n1500);
   U1986 : AOI22_X1 port map( A1 => n32, A2 => regs(1097), B1 => n3, B2 => 
                           regs(73), ZN => n1499);
   U1987 : AOI22_X1 port map( A1 => n46, A2 => regs(2121), B1 => n4, B2 => 
                           regs(1609), ZN => n1498);
   U1988 : NAND3_X1 port map( A1 => n1500, A2 => n1499, A3 => n1498, ZN => 
                           curr_proc_regs(73));
   U1989 : NAND2_X1 port map( A1 => regs(586), A2 => n2, ZN => n1503);
   U1990 : AOI22_X1 port map( A1 => n32, A2 => regs(1098), B1 => n3, B2 => 
                           regs(74), ZN => n1502);
   U1991 : AOI22_X1 port map( A1 => n40, A2 => regs(2122), B1 => n4, B2 => 
                           regs(1610), ZN => n1501);
   U1992 : NAND3_X1 port map( A1 => n1503, A2 => n1502, A3 => n1501, ZN => 
                           curr_proc_regs(74));
   U1993 : NAND2_X1 port map( A1 => regs(587), A2 => n7, ZN => n1506);
   U1994 : AOI22_X1 port map( A1 => n32, A2 => regs(1099), B1 => n3, B2 => 
                           regs(75), ZN => n1505);
   U1995 : AOI22_X1 port map( A1 => n10, A2 => regs(2123), B1 => n37, B2 => 
                           regs(1611), ZN => n1504);
   U1996 : NAND3_X1 port map( A1 => n1506, A2 => n1505, A3 => n1504, ZN => 
                           curr_proc_regs(75));
   U1997 : NAND2_X1 port map( A1 => regs(588), A2 => n21, ZN => n1509);
   U1998 : AOI22_X1 port map( A1 => n32, A2 => regs(1100), B1 => n3, B2 => 
                           regs(76), ZN => n1508);
   U1999 : AOI22_X1 port map( A1 => n10, A2 => regs(2124), B1 => n37, B2 => 
                           regs(1612), ZN => n1507);
   U2000 : NAND3_X1 port map( A1 => n1509, A2 => n1508, A3 => n1507, ZN => 
                           curr_proc_regs(76));
   U2001 : NAND2_X1 port map( A1 => regs(589), A2 => n23, ZN => n1512);
   U2002 : AOI22_X1 port map( A1 => n32, A2 => regs(1101), B1 => n3, B2 => 
                           regs(77), ZN => n1511);
   U2003 : AOI22_X1 port map( A1 => n10, A2 => regs(2125), B1 => n37, B2 => 
                           regs(1613), ZN => n1510);
   U2004 : NAND3_X1 port map( A1 => n1512, A2 => n1511, A3 => n1510, ZN => 
                           curr_proc_regs(77));
   U2005 : NAND2_X1 port map( A1 => regs(590), A2 => n22, ZN => n1515);
   U2006 : AOI22_X1 port map( A1 => n32, A2 => regs(1102), B1 => n3, B2 => 
                           regs(78), ZN => n1514);
   U2007 : AOI22_X1 port map( A1 => n10, A2 => regs(2126), B1 => n37, B2 => 
                           regs(1614), ZN => n1513);
   U2008 : NAND3_X1 port map( A1 => n1515, A2 => n1514, A3 => n1513, ZN => 
                           curr_proc_regs(78));
   U2009 : NAND2_X1 port map( A1 => regs(591), A2 => n2, ZN => n1518);
   U2010 : AOI22_X1 port map( A1 => n32, A2 => regs(1103), B1 => n3, B2 => 
                           regs(79), ZN => n1517);
   U2011 : AOI22_X1 port map( A1 => n10, A2 => regs(2127), B1 => n33, B2 => 
                           regs(1615), ZN => n1516);
   U2012 : NAND3_X1 port map( A1 => n1518, A2 => n1517, A3 => n1516, ZN => 
                           curr_proc_regs(79));
   U2013 : NAND2_X1 port map( A1 => regs(519), A2 => n7, ZN => n1521);
   U2014 : AOI22_X1 port map( A1 => n32, A2 => regs(1031), B1 => n3, B2 => 
                           regs(7), ZN => n1520);
   U2015 : AOI22_X1 port map( A1 => n10, A2 => regs(2055), B1 => n37, B2 => 
                           regs(1543), ZN => n1519);
   U2016 : NAND3_X1 port map( A1 => n1521, A2 => n1520, A3 => n1519, ZN => 
                           curr_proc_regs(7));
   U2017 : NAND2_X1 port map( A1 => regs(592), A2 => n7, ZN => n1524);
   U2018 : AOI22_X1 port map( A1 => n32, A2 => regs(1104), B1 => n3, B2 => 
                           regs(80), ZN => n1523);
   U2019 : AOI22_X1 port map( A1 => n10, A2 => regs(2128), B1 => n33, B2 => 
                           regs(1616), ZN => n1522);
   U2020 : NAND3_X1 port map( A1 => n1524, A2 => n1523, A3 => n1522, ZN => 
                           curr_proc_regs(80));
   U2021 : NAND2_X1 port map( A1 => regs(593), A2 => n1, ZN => n1527);
   U2022 : AOI22_X1 port map( A1 => n32, A2 => regs(1105), B1 => n3, B2 => 
                           regs(81), ZN => n1526);
   U2023 : AOI22_X1 port map( A1 => n10, A2 => regs(2129), B1 => n37, B2 => 
                           regs(1617), ZN => n1525);
   U2024 : NAND3_X1 port map( A1 => n1527, A2 => n1526, A3 => n1525, ZN => 
                           curr_proc_regs(81));
   U2025 : NAND2_X1 port map( A1 => regs(594), A2 => n2, ZN => n1530);
   U2026 : AOI22_X1 port map( A1 => n32, A2 => regs(1106), B1 => n3, B2 => 
                           regs(82), ZN => n1529);
   U2027 : AOI22_X1 port map( A1 => n10, A2 => regs(2130), B1 => n33, B2 => 
                           regs(1618), ZN => n1528);
   U2028 : NAND3_X1 port map( A1 => n1530, A2 => n1529, A3 => n1528, ZN => 
                           curr_proc_regs(82));
   U2029 : NAND2_X1 port map( A1 => regs(595), A2 => n23, ZN => n1533);
   U2030 : AOI22_X1 port map( A1 => n32, A2 => regs(1107), B1 => n3, B2 => 
                           regs(83), ZN => n1532);
   U2031 : AOI22_X1 port map( A1 => n10, A2 => regs(2131), B1 => n37, B2 => 
                           regs(1619), ZN => n1531);
   U2032 : NAND3_X1 port map( A1 => n1533, A2 => n1532, A3 => n1531, ZN => 
                           curr_proc_regs(83));
   U2033 : NAND2_X1 port map( A1 => regs(596), A2 => n17, ZN => n1536);
   U2034 : AOI22_X1 port map( A1 => n32, A2 => regs(1108), B1 => n3, B2 => 
                           regs(84), ZN => n1535);
   U2035 : AOI22_X1 port map( A1 => n10, A2 => regs(2132), B1 => n33, B2 => 
                           regs(1620), ZN => n1534);
   U2036 : NAND3_X1 port map( A1 => n1536, A2 => n1535, A3 => n1534, ZN => 
                           curr_proc_regs(84));
   U2037 : NAND2_X1 port map( A1 => regs(597), A2 => n1585, ZN => n1539);
   U2038 : AOI22_X1 port map( A1 => n32, A2 => regs(1109), B1 => n8, B2 => 
                           regs(85), ZN => n1538);
   U2039 : AOI22_X1 port map( A1 => n10, A2 => regs(2133), B1 => n37, B2 => 
                           regs(1621), ZN => n1537);
   U2040 : NAND3_X1 port map( A1 => n1539, A2 => n1538, A3 => n1537, ZN => 
                           curr_proc_regs(85));
   U2041 : NAND2_X1 port map( A1 => regs(598), A2 => n7, ZN => n1542);
   U2042 : AOI22_X1 port map( A1 => n32, A2 => regs(1110), B1 => n3, B2 => 
                           regs(86), ZN => n1541);
   U2043 : AOI22_X1 port map( A1 => n10, A2 => regs(2134), B1 => n37, B2 => 
                           regs(1622), ZN => n1540);
   U2044 : NAND3_X1 port map( A1 => n1542, A2 => n1541, A3 => n1540, ZN => 
                           curr_proc_regs(86));
   U2045 : NAND2_X1 port map( A1 => regs(599), A2 => n1585, ZN => n1545);
   U2046 : AOI22_X1 port map( A1 => n32, A2 => regs(1111), B1 => n31, B2 => 
                           regs(87), ZN => n1544);
   U2047 : AOI22_X1 port map( A1 => n10, A2 => regs(2135), B1 => n37, B2 => 
                           regs(1623), ZN => n1543);
   U2048 : NAND3_X1 port map( A1 => n1545, A2 => n1544, A3 => n1543, ZN => 
                           curr_proc_regs(87));
   U2049 : NAND2_X1 port map( A1 => regs(600), A2 => n22, ZN => n1548);
   U2050 : AOI22_X1 port map( A1 => n32, A2 => regs(1112), B1 => n8, B2 => 
                           regs(88), ZN => n1547);
   U2051 : AOI22_X1 port map( A1 => n10, A2 => regs(2136), B1 => n37, B2 => 
                           regs(1624), ZN => n1546);
   U2052 : NAND3_X1 port map( A1 => n1548, A2 => n1547, A3 => n1546, ZN => 
                           curr_proc_regs(88));
   U2053 : NAND2_X1 port map( A1 => regs(601), A2 => n1585, ZN => n1551);
   U2054 : AOI22_X1 port map( A1 => n32, A2 => regs(1113), B1 => n3, B2 => 
                           regs(89), ZN => n1550);
   U2055 : AOI22_X1 port map( A1 => n10, A2 => regs(2137), B1 => n37, B2 => 
                           regs(1625), ZN => n1549);
   U2056 : NAND3_X1 port map( A1 => n1551, A2 => n1550, A3 => n1549, ZN => 
                           curr_proc_regs(89));
   U2057 : NAND2_X1 port map( A1 => regs(520), A2 => n6, ZN => n1554);
   U2058 : AOI22_X1 port map( A1 => n32, A2 => regs(1032), B1 => n31, B2 => 
                           regs(8), ZN => n1553);
   U2059 : AOI22_X1 port map( A1 => n10, A2 => regs(2056), B1 => n37, B2 => 
                           regs(1544), ZN => n1552);
   U2060 : NAND3_X1 port map( A1 => n1554, A2 => n1553, A3 => n1552, ZN => 
                           curr_proc_regs(8));
   U2061 : NAND2_X1 port map( A1 => regs(602), A2 => n1585, ZN => n1557);
   U2062 : AOI22_X1 port map( A1 => n32, A2 => regs(1114), B1 => n8, B2 => 
                           regs(90), ZN => n1556);
   U2063 : AOI22_X1 port map( A1 => n10, A2 => regs(2138), B1 => n37, B2 => 
                           regs(1626), ZN => n1555);
   U2064 : NAND3_X1 port map( A1 => n1557, A2 => n1556, A3 => n1555, ZN => 
                           curr_proc_regs(90));
   U2065 : NAND2_X1 port map( A1 => regs(603), A2 => n20, ZN => n1560);
   U2066 : AOI22_X1 port map( A1 => n32, A2 => regs(1115), B1 => n3, B2 => 
                           regs(91), ZN => n1559);
   U2067 : AOI22_X1 port map( A1 => n10, A2 => regs(2139), B1 => n37, B2 => 
                           regs(1627), ZN => n1558);
   U2068 : NAND3_X1 port map( A1 => n1560, A2 => n1559, A3 => n1558, ZN => 
                           curr_proc_regs(91));
   U2069 : NAND2_X1 port map( A1 => regs(604), A2 => n18, ZN => n1563);
   U2070 : AOI22_X1 port map( A1 => n32, A2 => regs(1116), B1 => n31, B2 => 
                           regs(92), ZN => n1562);
   U2071 : AOI22_X1 port map( A1 => n10, A2 => regs(2140), B1 => n37, B2 => 
                           regs(1628), ZN => n1561);
   U2072 : NAND3_X1 port map( A1 => n1563, A2 => n1562, A3 => n1561, ZN => 
                           curr_proc_regs(92));
   U2073 : NAND2_X1 port map( A1 => regs(605), A2 => n2, ZN => n1566);
   U2074 : AOI22_X1 port map( A1 => n32, A2 => regs(1117), B1 => n8, B2 => 
                           regs(93), ZN => n1565);
   U2075 : AOI22_X1 port map( A1 => n10, A2 => regs(2141), B1 => n37, B2 => 
                           regs(1629), ZN => n1564);
   U2076 : NAND3_X1 port map( A1 => n1566, A2 => n1565, A3 => n1564, ZN => 
                           curr_proc_regs(93));
   U2077 : NAND2_X1 port map( A1 => regs(606), A2 => n7, ZN => n1569);
   U2078 : AOI22_X1 port map( A1 => n32, A2 => regs(1118), B1 => n3, B2 => 
                           regs(94), ZN => n1568);
   U2079 : AOI22_X1 port map( A1 => n10, A2 => regs(2142), B1 => n37, B2 => 
                           regs(1630), ZN => n1567);
   U2080 : NAND3_X1 port map( A1 => n1569, A2 => n1568, A3 => n1567, ZN => 
                           curr_proc_regs(94));
   U2081 : NAND2_X1 port map( A1 => regs(607), A2 => n24, ZN => n1572);
   U2082 : AOI22_X1 port map( A1 => n32, A2 => regs(1119), B1 => n29, B2 => 
                           regs(95), ZN => n1571);
   U2083 : AOI22_X1 port map( A1 => n10, A2 => regs(2143), B1 => n38, B2 => 
                           regs(1631), ZN => n1570);
   U2084 : NAND3_X1 port map( A1 => n1572, A2 => n1571, A3 => n1570, ZN => 
                           curr_proc_regs(95));
   U2085 : NAND2_X1 port map( A1 => regs(608), A2 => n24, ZN => n1575);
   U2086 : AOI22_X1 port map( A1 => n32, A2 => regs(1120), B1 => n29, B2 => 
                           regs(96), ZN => n1574);
   U2087 : AOI22_X1 port map( A1 => n40, A2 => regs(2144), B1 => n38, B2 => 
                           regs(1632), ZN => n1573);
   U2088 : NAND3_X1 port map( A1 => n1575, A2 => n1574, A3 => n1573, ZN => 
                           curr_proc_regs(96));
   U2089 : NAND2_X1 port map( A1 => regs(609), A2 => n24, ZN => n1578);
   U2090 : AOI22_X1 port map( A1 => n32, A2 => regs(1121), B1 => n29, B2 => 
                           regs(97), ZN => n1577);
   U2091 : AOI22_X1 port map( A1 => n46, A2 => regs(2145), B1 => n38, B2 => 
                           regs(1633), ZN => n1576);
   U2092 : NAND3_X1 port map( A1 => n1578, A2 => n1577, A3 => n1576, ZN => 
                           curr_proc_regs(97));
   U2093 : NAND2_X1 port map( A1 => regs(610), A2 => n24, ZN => n1581);
   U2094 : AOI22_X1 port map( A1 => n32, A2 => regs(1122), B1 => n29, B2 => 
                           regs(98), ZN => n1580);
   U2095 : AOI22_X1 port map( A1 => n15, A2 => regs(2146), B1 => n38, B2 => 
                           regs(1634), ZN => n1579);
   U2096 : NAND3_X1 port map( A1 => n1581, A2 => n1580, A3 => n1579, ZN => 
                           curr_proc_regs(98));
   U2097 : NAND2_X1 port map( A1 => regs(611), A2 => n24, ZN => n1584);
   U2098 : AOI22_X1 port map( A1 => n32, A2 => regs(1123), B1 => n29, B2 => 
                           regs(99), ZN => n1583);
   U2099 : AOI22_X1 port map( A1 => n14, A2 => regs(2147), B1 => n38, B2 => 
                           regs(1635), ZN => n1582);
   U2100 : NAND3_X1 port map( A1 => n1584, A2 => n1583, A3 => n1582, ZN => 
                           curr_proc_regs(99));
   U2101 : NAND2_X1 port map( A1 => regs(521), A2 => n24, ZN => n1591);
   U2102 : AOI22_X1 port map( A1 => n32, A2 => regs(1033), B1 => n29, B2 => 
                           regs(9), ZN => n1590);
   U2103 : AOI22_X1 port map( A1 => n44, A2 => regs(2057), B1 => n38, B2 => 
                           regs(1545), ZN => n1589);
   U2104 : NAND3_X1 port map( A1 => n1591, A2 => n1590, A3 => n1589, ZN => 
                           curr_proc_regs(9));

end SYN_behav;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32.all;

entity hazard_table_N_REGS_LOG5 is

   port( CLK, RST, WR1, WR2 : in std_logic;  ADD_WR1, ADD_WR2, ADD_CHECK1, 
         ADD_CHECK2 : in std_logic_vector (4 downto 0);  BUSY, BUSY_WINDOW : 
         out std_logic);

end hazard_table_N_REGS_LOG5;

architecture SYN_behavioural of hazard_table_N_REGS_LOG5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Table_0_2_port, Table_0_1_port, Table_0_0_port, Table_1_2_port, 
      Table_1_1_port, Table_1_0_port, Table_2_2_port, Table_2_1_port, 
      Table_2_0_port, Table_3_2_port, Table_3_1_port, Table_3_0_port, 
      Table_4_2_port, Table_4_1_port, Table_4_0_port, Table_5_2_port, 
      Table_5_1_port, Table_5_0_port, Table_6_2_port, Table_6_1_port, 
      Table_6_0_port, Table_7_2_port, Table_7_1_port, Table_7_0_port, 
      Table_8_2_port, Table_8_1_port, Table_8_0_port, Table_9_2_port, 
      Table_9_1_port, Table_9_0_port, Table_10_2_port, Table_10_1_port, 
      Table_10_0_port, Table_11_2_port, Table_11_1_port, Table_11_0_port, 
      Table_12_2_port, Table_12_1_port, Table_12_0_port, Table_13_2_port, 
      Table_13_1_port, Table_13_0_port, Table_14_2_port, Table_14_1_port, 
      Table_14_0_port, Table_15_2_port, Table_15_1_port, Table_15_0_port, 
      Table_16_2_port, Table_16_1_port, Table_16_0_port, Table_17_2_port, 
      Table_17_1_port, Table_17_0_port, Table_18_2_port, Table_18_1_port, 
      Table_18_0_port, Table_19_2_port, Table_19_1_port, Table_19_0_port, 
      Table_20_2_port, Table_20_1_port, Table_20_0_port, Table_21_2_port, 
      Table_21_1_port, Table_21_0_port, Table_22_2_port, Table_22_1_port, 
      Table_22_0_port, Table_23_2_port, Table_23_1_port, Table_23_0_port, 
      Table_24_2_port, Table_24_1_port, Table_24_0_port, Table_25_2_port, 
      Table_25_1_port, Table_25_0_port, Table_26_2_port, Table_26_1_port, 
      Table_26_0_port, Table_27_2_port, Table_27_1_port, Table_27_0_port, 
      Table_28_2_port, Table_28_1_port, Table_28_0_port, Table_29_2_port, 
      Table_29_1_port, Table_29_0_port, Table_30_2_port, Table_30_1_port, 
      Table_30_0_port, Table_31_2_port, Table_31_1_port, Table_31_0_port, n702,
      n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, 
      n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, 
      n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n1, n2,
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, 
      n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, 
      n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, 
      n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, 
      n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
      n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, 
      n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, 
      n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, 
      n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, 
      n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, 
      n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, 
      n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, 
      n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, 
      n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, 
      n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, 
      n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, 
      n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, 
      n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, 
      n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, 
      n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, 
      n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, 
      n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, 
      n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, 
      n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, 
      n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, 
      n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, 
      n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, 
      n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, 
      n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, 
      n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, 
      n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, 
      n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, 
      n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, 
      n694, n695, n_1064 : std_logic;

begin
   
   Table_reg_31_2_inst : DFF_X1 port map( D => n795, CK => CLK, Q => 
                           Table_31_2_port, QN => n_1064);
   Table_reg_0_2_inst : DFF_X1 port map( D => n702, CK => CLK, Q => 
                           Table_0_2_port, QN => n12);
   Table_reg_1_2_inst : DFF_X1 port map( D => n705, CK => CLK, Q => 
                           Table_1_2_port, QN => n103);
   Table_reg_2_2_inst : DFF_X1 port map( D => n708, CK => CLK, Q => 
                           Table_2_2_port, QN => n79);
   Table_reg_3_2_inst : DFF_X1 port map( D => n711, CK => CLK, Q => 
                           Table_3_2_port, QN => n15);
   Table_reg_4_2_inst : DFF_X1 port map( D => n714, CK => CLK, Q => 
                           Table_4_2_port, QN => n78);
   Table_reg_5_2_inst : DFF_X1 port map( D => n717, CK => CLK, Q => 
                           Table_5_2_port, QN => n102);
   Table_reg_6_2_inst : DFF_X1 port map( D => n720, CK => CLK, Q => 
                           Table_6_2_port, QN => n77);
   Table_reg_7_2_inst : DFF_X1 port map( D => n723, CK => CLK, Q => 
                           Table_7_2_port, QN => n14);
   Table_reg_8_2_inst : DFF_X1 port map( D => n726, CK => CLK, Q => 
                           Table_8_2_port, QN => n54);
   Table_reg_9_2_inst : DFF_X1 port map( D => n729, CK => CLK, Q => 
                           Table_9_2_port, QN => n42);
   Table_reg_10_2_inst : DFF_X1 port map( D => n732, CK => CLK, Q => 
                           Table_10_2_port, QN => n53);
   Table_reg_11_2_inst : DFF_X1 port map( D => n735, CK => CLK, Q => 
                           Table_11_2_port, QN => n88);
   Table_reg_12_2_inst : DFF_X1 port map( D => n738, CK => CLK, Q => 
                           Table_12_2_port, QN => n52);
   Table_reg_13_2_inst : DFF_X1 port map( D => n741, CK => CLK, Q => 
                           Table_13_2_port, QN => n34);
   Table_reg_14_2_inst : DFF_X1 port map( D => n744, CK => CLK, Q => 
                           Table_14_2_port, QN => n51);
   Table_reg_15_2_inst : DFF_X1 port map( D => n747, CK => CLK, Q => 
                           Table_15_2_port, QN => n87);
   Table_reg_16_2_inst : DFF_X1 port map( D => n750, CK => CLK, Q => 
                           Table_16_2_port, QN => n141);
   Table_reg_17_2_inst : DFF_X1 port map( D => n753, CK => CLK, Q => 
                           Table_17_2_port, QN => n33);
   Table_reg_18_2_inst : DFF_X1 port map( D => n756, CK => CLK, Q => 
                           Table_18_2_port, QN => n50);
   Table_reg_19_2_inst : DFF_X1 port map( D => n759, CK => CLK, Q => 
                           Table_19_2_port, QN => n101);
   Table_reg_20_2_inst : DFF_X1 port map( D => n762, CK => CLK, Q => 
                           Table_20_2_port, QN => n49);
   Table_reg_21_2_inst : DFF_X1 port map( D => n765, CK => CLK, Q => 
                           Table_21_2_port, QN => n10);
   Table_reg_22_2_inst : DFF_X1 port map( D => n768, CK => CLK, Q => 
                           Table_22_2_port, QN => n48);
   Table_reg_23_2_inst : DFF_X1 port map( D => n771, CK => CLK, Q => 
                           Table_23_2_port, QN => n90);
   Table_reg_24_2_inst : DFF_X1 port map( D => n774, CK => CLK, Q => 
                           Table_24_2_port, QN => n11);
   Table_reg_25_2_inst : DFF_X1 port map( D => n777, CK => CLK, Q => 
                           Table_25_2_port, QN => n32);
   Table_reg_26_2_inst : DFF_X1 port map( D => n780, CK => CLK, Q => 
                           Table_26_2_port, QN => n47);
   Table_reg_27_2_inst : DFF_X1 port map( D => n783, CK => CLK, Q => 
                           Table_27_2_port, QN => n85);
   Table_reg_28_2_inst : DFF_X1 port map( D => n786, CK => CLK, Q => 
                           Table_28_2_port, QN => n13);
   Table_reg_29_2_inst : DFF_X1 port map( D => n789, CK => CLK, Q => 
                           Table_29_2_port, QN => n76);
   Table_reg_30_2_inst : DFF_X1 port map( D => n792, CK => CLK, Q => 
                           Table_30_2_port, QN => n75);
   Table_reg_29_0_inst : DFF_X1 port map( D => n791, CK => CLK, Q => 
                           Table_29_0_port, QN => n55);
   Table_reg_21_0_inst : DFF_X1 port map( D => n767, CK => CLK, Q => 
                           Table_21_0_port, QN => n16);
   Table_reg_13_0_inst : DFF_X1 port map( D => n743, CK => CLK, Q => 
                           Table_13_0_port, QN => n38);
   Table_reg_5_0_inst : DFF_X1 port map( D => n719, CK => CLK, Q => 
                           Table_5_0_port, QN => n94);
   Table_reg_23_0_inst : DFF_X1 port map( D => n773, CK => CLK, Q => 
                           Table_23_0_port, QN => n98);
   Table_reg_15_0_inst : DFF_X1 port map( D => n749, CK => CLK, Q => 
                           Table_15_0_port, QN => n99);
   Table_reg_7_0_inst : DFF_X1 port map( D => n725, CK => CLK, Q => 
                           Table_7_0_port, QN => n20);
   Table_reg_27_0_inst : DFF_X1 port map( D => n785, CK => CLK, Q => 
                           Table_27_0_port, QN => n97);
   Table_reg_25_0_inst : DFF_X1 port map( D => n779, CK => CLK, Q => 
                           Table_25_0_port, QN => n36);
   Table_reg_19_0_inst : DFF_X1 port map( D => n761, CK => CLK, Q => 
                           Table_19_0_port, QN => n93);
   Table_reg_17_0_inst : DFF_X1 port map( D => n755, CK => CLK, Q => 
                           Table_17_0_port, QN => n37);
   Table_reg_11_0_inst : DFF_X1 port map( D => n737, CK => CLK, Q => 
                           Table_11_0_port, QN => n100);
   Table_reg_9_0_inst : DFF_X1 port map( D => n731, CK => CLK, Q => 
                           Table_9_0_port, QN => n41);
   Table_reg_3_0_inst : DFF_X1 port map( D => n713, CK => CLK, Q => 
                           Table_3_0_port, QN => n21);
   Table_reg_1_0_inst : DFF_X1 port map( D => n707, CK => CLK, Q => 
                           Table_1_0_port, QN => n95);
   Table_reg_30_0_inst : DFF_X1 port map( D => n794, CK => CLK, Q => 
                           Table_30_0_port, QN => n84);
   Table_reg_22_0_inst : DFF_X1 port map( D => n770, CK => CLK, Q => 
                           Table_22_0_port, QN => n57);
   Table_reg_14_0_inst : DFF_X1 port map( D => n746, CK => CLK, Q => 
                           Table_14_0_port, QN => n60);
   Table_reg_6_0_inst : DFF_X1 port map( D => n722, CK => CLK, Q => 
                           Table_6_0_port, QN => n64);
   Table_reg_28_0_inst : DFF_X1 port map( D => n788, CK => CLK, Q => 
                           Table_28_0_port, QN => n19);
   Table_reg_26_0_inst : DFF_X1 port map( D => n782, CK => CLK, Q => 
                           Table_26_0_port, QN => n67);
   Table_reg_24_0_inst : DFF_X1 port map( D => n776, CK => CLK, Q => 
                           Table_24_0_port, QN => n17);
   Table_reg_20_0_inst : DFF_X1 port map( D => n764, CK => CLK, Q => 
                           Table_20_0_port, QN => n58);
   Table_reg_18_0_inst : DFF_X1 port map( D => n758, CK => CLK, Q => 
                           Table_18_0_port, QN => n59);
   Table_reg_16_0_inst : DFF_X1 port map( D => n752, CK => CLK, Q => 
                           Table_16_0_port, QN => n140);
   Table_reg_12_0_inst : DFF_X1 port map( D => n740, CK => CLK, Q => 
                           Table_12_0_port, QN => n61);
   Table_reg_10_0_inst : DFF_X1 port map( D => n734, CK => CLK, Q => 
                           Table_10_0_port, QN => n62);
   Table_reg_8_0_inst : DFF_X1 port map( D => n728, CK => CLK, Q => 
                           Table_8_0_port, QN => n63);
   Table_reg_4_0_inst : DFF_X1 port map( D => n716, CK => CLK, Q => 
                           Table_4_0_port, QN => n65);
   Table_reg_2_0_inst : DFF_X1 port map( D => n710, CK => CLK, Q => 
                           Table_2_0_port, QN => n66);
   Table_reg_0_0_inst : DFF_X1 port map( D => n704, CK => CLK, Q => 
                           Table_0_0_port, QN => n18);
   Table_reg_31_0_inst : DFF_X1 port map( D => n797, CK => CLK, Q => 
                           Table_31_0_port, QN => n96);
   Table_reg_31_1_inst : DFF_X1 port map( D => n796, CK => CLK, Q => 
                           Table_31_1_port, QN => n80);
   Table_reg_30_1_inst : DFF_X1 port map( D => n793, CK => CLK, Q => 
                           Table_30_1_port, QN => n22);
   Table_reg_29_1_inst : DFF_X1 port map( D => n790, CK => CLK, Q => 
                           Table_29_1_port, QN => n31);
   Table_reg_28_1_inst : DFF_X1 port map( D => n787, CK => CLK, Q => 
                           Table_28_1_port, QN => n27);
   Table_reg_27_1_inst : DFF_X1 port map( D => n784, CK => CLK, Q => 
                           Table_27_1_port, QN => n89);
   Table_reg_26_1_inst : DFF_X1 port map( D => n781, CK => CLK, Q => 
                           Table_26_1_port, QN => n56);
   Table_reg_25_1_inst : DFF_X1 port map( D => n778, CK => CLK, Q => 
                           Table_25_1_port, QN => n39);
   Table_reg_24_1_inst : DFF_X1 port map( D => n775, CK => CLK, Q => 
                           Table_24_1_port, QN => n23);
   Table_reg_23_1_inst : DFF_X1 port map( D => n772, CK => CLK, Q => 
                           Table_23_1_port, QN => n86);
   Table_reg_22_1_inst : DFF_X1 port map( D => n769, CK => CLK, Q => 
                           Table_22_1_port, QN => n68);
   Table_reg_21_1_inst : DFF_X1 port map( D => n766, CK => CLK, Q => 
                           Table_21_1_port, QN => n24);
   Table_reg_20_1_inst : DFF_X1 port map( D => n763, CK => CLK, Q => 
                           Table_20_1_port, QN => n69);
   Table_reg_19_1_inst : DFF_X1 port map( D => n760, CK => CLK, Q => 
                           Table_19_1_port, QN => n81);
   Table_reg_18_1_inst : DFF_X1 port map( D => n757, CK => CLK, Q => 
                           Table_18_1_port, QN => n70);
   Table_reg_17_1_inst : DFF_X1 port map( D => n754, CK => CLK, Q => 
                           Table_17_1_port, QN => n40);
   Table_reg_16_1_inst : DFF_X1 port map( D => n751, CK => CLK, Q => 
                           Table_16_1_port, QN => n139);
   Table_reg_15_1_inst : DFF_X1 port map( D => n748, CK => CLK, Q => 
                           Table_15_1_port, QN => n91);
   Table_reg_14_1_inst : DFF_X1 port map( D => n745, CK => CLK, Q => 
                           Table_14_1_port, QN => n71);
   Table_reg_13_1_inst : DFF_X1 port map( D => n742, CK => CLK, Q => 
                           Table_13_1_port, QN => n35);
   Table_reg_12_1_inst : DFF_X1 port map( D => n739, CK => CLK, Q => 
                           Table_12_1_port, QN => n72);
   Table_reg_11_1_inst : DFF_X1 port map( D => n736, CK => CLK, Q => 
                           Table_11_1_port, QN => n92);
   Table_reg_10_1_inst : DFF_X1 port map( D => n733, CK => CLK, Q => 
                           Table_10_1_port, QN => n73);
   Table_reg_8_1_inst : DFF_X1 port map( D => n727, CK => CLK, Q => 
                           Table_8_1_port, QN => n74);
   Table_reg_7_1_inst : DFF_X1 port map( D => n724, CK => CLK, Q => 
                           Table_7_1_port, QN => n28);
   Table_reg_5_1_inst : DFF_X1 port map( D => n718, CK => CLK, Q => 
                           Table_5_1_port, QN => n82);
   Table_reg_3_1_inst : DFF_X1 port map( D => n712, CK => CLK, Q => 
                           Table_3_1_port, QN => n29);
   Table_reg_1_1_inst : DFF_X1 port map( D => n706, CK => CLK, Q => 
                           Table_1_1_port, QN => n83);
   Table_reg_0_1_inst : DFF_X1 port map( D => n703, CK => CLK, Q => 
                           Table_0_1_port, QN => n26);
   Table_reg_9_1_inst : DFF_X1 port map( D => n730, CK => CLK, Q => 
                           Table_9_1_port, QN => n43);
   Table_reg_6_1_inst : DFF_X1 port map( D => n721, CK => CLK, Q => 
                           Table_6_1_port, QN => n44);
   Table_reg_4_1_inst : DFF_X1 port map( D => n715, CK => CLK, Q => 
                           Table_4_1_port, QN => n45);
   Table_reg_2_1_inst : DFF_X1 port map( D => n709, CK => CLK, Q => 
                           Table_2_1_port, QN => n46);
   U3 : AND2_X2 port map( A1 => n438, A2 => n362, ZN => n684);
   U4 : AOI21_X1 port map( B1 => n271, B2 => WR1, A => n270, ZN => n680);
   U5 : AOI211_X4 port map( C1 => n417, C2 => n416, A => RST, B => n415, ZN => 
                           n692);
   U6 : NOR2_X1 port map( A1 => n6, A2 => Table_12_2_port, ZN => n104);
   U7 : AND2_X1 port map( A1 => n138, A2 => n59, ZN => n164);
   U8 : NOR2_X1 port map( A1 => n4, A2 => Table_8_2_port, ZN => n108);
   U9 : NOR2_X1 port map( A1 => n7, A2 => Table_26_2_port, ZN => n117);
   U10 : BUF_X2 port map( A => n687, Z => n1);
   U11 : BUF_X1 port map( A => n680, Z => n142);
   U12 : BUF_X2 port map( A => n686, Z => n2);
   U13 : BUF_X1 port map( A => n683, Z => n143);
   U14 : INV_X1 port map( A => ADD_WR1(2), ZN => n314);
   U15 : INV_X1 port map( A => ADD_WR1(1), ZN => n313);
   U16 : NOR2_X1 port map( A1 => Table_11_2_port, A2 => n8, ZN => n216);
   U17 : NOR2_X1 port map( A1 => Table_27_2_port, A2 => n9, ZN => n217);
   U18 : NOR3_X1 port map( A1 => Table_19_1_port, A2 => Table_19_0_port, A3 => 
                           Table_19_2_port, ZN => n220);
   U19 : AND3_X1 port map( A1 => n43, A2 => n42, A3 => n41, ZN => n246);
   U20 : AND3_X1 port map( A1 => n24, A2 => n16, A3 => n10, ZN => n195);
   U21 : INV_X1 port map( A => ADD_WR1(0), ZN => n312);
   U22 : BUF_X1 port map( A => n689, Z => n144);
   U23 : NOR2_X2 port map( A1 => ADD_WR1(1), A2 => n311, ZN => n457);
   U24 : AND2_X1 port map( A1 => n75, A2 => n84, ZN => n119);
   U25 : AND2_X1 port map( A1 => n86, A2 => n98, ZN => n120);
   U26 : AND2_X1 port map( A1 => n132, A2 => n80, ZN => n225);
   U27 : NAND2_X1 port map( A1 => n63, A2 => n74, ZN => n4);
   U28 : NOR2_X1 port map( A1 => n5, A2 => n242, ZN => n125);
   U29 : NAND2_X1 port map( A1 => n195, A2 => n220, ZN => n5);
   U30 : AND2_X1 port map( A1 => n33, A2 => n37, ZN => n122);
   U31 : NAND2_X1 port map( A1 => n61, A2 => n72, ZN => n6);
   U32 : AND2_X1 port map( A1 => n135, A2 => n60, ZN => n173);
   U33 : AND4_X1 port map( A1 => n119, A2 => n120, A3 => n90, A4 => n22, ZN => 
                           n118);
   U34 : AND4_X1 port map( A1 => n148, A2 => n118, A3 => n225, A4 => n224, ZN 
                           => n25);
   U35 : AND2_X1 port map( A1 => n137, A2 => n58, ZN => n169);
   U36 : NAND2_X1 port map( A1 => n56, A2 => n67, ZN => n7);
   U37 : AND2_X1 port map( A1 => n134, A2 => n62, ZN => n172);
   U38 : NAND2_X1 port map( A1 => n92, A2 => n100, ZN => n8);
   U39 : AND2_X1 port map( A1 => n55, A2 => n76, ZN => n127);
   U40 : AND2_X1 port map( A1 => n57, A2 => n109, ZN => n165);
   U41 : NAND2_X1 port map( A1 => n89, A2 => n97, ZN => n9);
   U42 : NAND4_X1 port map( A1 => n130, A2 => n124, A3 => n125, A4 => n25, ZN 
                           => BUSY_WINDOW);
   U43 : NOR2_X1 port map( A1 => n115, A2 => n110, ZN => n124);
   U44 : AND2_X1 port map( A1 => n131, A2 => n91, ZN => n224);
   U45 : INV_X1 port map( A => ADD_CHECK2(4), ZN => n218);
   U46 : NOR2_X1 port map( A1 => n136, A2 => n133, ZN => n130);
   U47 : AOI21_X1 port map( B1 => n441, B2 => n440, A => n439, ZN => n689);
   U48 : NOR2_X1 port map( A1 => RST, A2 => n386, ZN => n683);
   U49 : NAND3_X1 port map( A1 => n27, A2 => n19, A3 => n13, ZN => n242);
   U50 : NAND4_X1 port map( A1 => n173, A2 => n172, A3 => n108, A4 => n104, ZN 
                           => n133);
   U51 : NOR2_X1 port map( A1 => Table_15_2_port, A2 => Table_15_0_port, ZN => 
                           n131);
   U52 : NOR2_X1 port map( A1 => Table_31_2_port, A2 => Table_31_0_port, ZN => 
                           n132);
   U53 : INV_X1 port map( A => n489, ZN => n672);
   U54 : INV_X1 port map( A => n457, ZN => n640);
   U55 : INV_X1 port map( A => n481, ZN => n664);
   U56 : INV_X1 port map( A => n465, ZN => n648);
   U57 : INV_X1 port map( A => n447, ZN => n632);
   U58 : INV_X1 port map( A => n473, ZN => n656);
   U59 : INV_X1 port map( A => n405, ZN => n624);
   U60 : INV_X1 port map( A => n497, ZN => n682);
   U61 : INV_X1 port map( A => RST, ZN => n146);
   U62 : INV_X1 port map( A => RST, ZN => n145);
   U63 : INV_X1 port map( A => ADD_WR2(3), ZN => n292);
   U64 : NOR3_X2 port map( A1 => n313, A2 => n314, A3 => n312, ZN => n405);
   U65 : NOR3_X2 port map( A1 => ADD_WR1(0), A2 => n314, A3 => n313, ZN => n447
                           );
   U66 : NOR3_X2 port map( A1 => ADD_WR1(1), A2 => ADD_WR1(0), A3 => n314, ZN 
                           => n465);
   U67 : NOR3_X2 port map( A1 => ADD_WR1(2), A2 => n313, A3 => n312, ZN => n473
                           );
   U68 : NOR3_X2 port map( A1 => ADD_WR1(2), A2 => ADD_WR1(0), A3 => n313, ZN 
                           => n481);
   U69 : NOR3_X2 port map( A1 => ADD_WR1(1), A2 => ADD_WR1(2), A3 => n312, ZN 
                           => n489);
   U70 : INV_X1 port map( A => ADD_WR2(2), ZN => n273);
   U71 : INV_X1 port map( A => ADD_WR2(4), ZN => n293);
   U72 : NOR3_X2 port map( A1 => ADD_WR1(1), A2 => ADD_WR1(2), A3 => ADD_WR1(0)
                           , ZN => n497);
   U73 : OAI21_X1 port map( B1 => n226, B2 => n117, A => n116, ZN => n221);
   U74 : OR2_X1 port map( A1 => n249, A2 => n220, ZN => n116);
   U75 : AND2_X1 port map( A1 => n120, A2 => n90, ZN => n228);
   U76 : AND2_X1 port map( A1 => n129, A2 => n35, ZN => n238);
   U77 : NOR2_X1 port map( A1 => Table_13_0_port, A2 => Table_13_2_port, ZN => 
                           n129);
   U78 : AND2_X1 port map( A1 => n127, A2 => n31, ZN => n239);
   U79 : AND2_X1 port map( A1 => n126, A2 => n39, ZN => n248);
   U80 : NOR2_X1 port map( A1 => Table_25_0_port, A2 => Table_25_2_port, ZN => 
                           n126);
   U81 : AND2_X1 port map( A1 => n128, A2 => n40, ZN => n250);
   U82 : NOR2_X1 port map( A1 => Table_17_0_port, A2 => Table_17_2_port, ZN => 
                           n128);
   U83 : INV_X1 port map( A => n104, ZN => n186);
   U84 : NAND2_X1 port map( A1 => n175, A2 => n106, ZN => n187);
   U85 : INV_X1 port map( A => n107, ZN => n106);
   U86 : OAI21_X1 port map( B1 => n176, B2 => n108, A => ADD_CHECK1(3), ZN => 
                           n107);
   U87 : OAI21_X1 port map( B1 => n177, B2 => n117, A => n30, ZN => n161);
   U88 : AND2_X1 port map( A1 => n119, A2 => n22, ZN => n227);
   U89 : AOI211_X1 port map( C1 => n256, C2 => n108, A => ADD_CHECK2(1), B => 
                           n105, ZN => n159);
   U90 : AND2_X1 port map( A1 => ADD_CHECK2(2), A2 => n104, ZN => n105);
   U91 : AOI211_X1 port map( C1 => n167, C2 => n152, A => n218, B => n149, ZN 
                           => n157);
   U92 : AOI221_X1 port map( B1 => n256, B2 => n164, C1 => ADD_CHECK2(2), C2 =>
                           n165, A => n150, ZN => n149);
   U93 : OR2_X1 port map( A1 => n208, A2 => n227, ZN => n30);
   U94 : NAND4_X1 port map( A1 => n165, A2 => n216, A3 => n217, A4 => n117, ZN 
                           => n115);
   U95 : NOR2_X1 port map( A1 => Table_22_2_port, A2 => Table_22_1_port, ZN => 
                           n109);
   U96 : NAND4_X1 port map( A1 => n112, A2 => n111, A3 => n121, A4 => n123, ZN 
                           => n110);
   U97 : AND2_X1 port map( A1 => n113, A2 => n127, ZN => n111);
   U98 : AND2_X1 port map( A1 => n122, A2 => n114, ZN => n112);
   U99 : NOR2_X1 port map( A1 => Table_29_1_port, A2 => Table_25_1_port, ZN => 
                           n113);
   U100 : NOR2_X1 port map( A1 => Table_13_1_port, A2 => Table_17_1_port, ZN =>
                           n114);
   U101 : NOR2_X1 port map( A1 => Table_25_2_port, A2 => Table_13_0_port, ZN =>
                           n121);
   U102 : NOR2_X1 port map( A1 => Table_13_2_port, A2 => Table_25_0_port, ZN =>
                           n123);
   U103 : NOR2_X1 port map( A1 => Table_10_2_port, A2 => Table_10_1_port, ZN =>
                           n134);
   U104 : NOR2_X1 port map( A1 => Table_14_2_port, A2 => Table_14_1_port, ZN =>
                           n135);
   U105 : NAND4_X1 port map( A1 => n164, A2 => n169, A3 => n246, A4 => n147, ZN
                           => n136);
   U106 : NOR2_X1 port map( A1 => Table_20_2_port, A2 => Table_20_1_port, ZN =>
                           n137);
   U107 : NOR2_X1 port map( A1 => Table_18_2_port, A2 => Table_18_1_port, ZN =>
                           n138);
   U108 : NAND3_X1 port map( A1 => n23, A2 => n17, A3 => n11, ZN => n253);
   U109 : INV_X1 port map( A => n253, ZN => n148);
   U110 : NAND3_X1 port map( A1 => n139, A2 => n140, A3 => n141, ZN => n167);
   U111 : INV_X1 port map( A => n167, ZN => n147);
   U112 : NOR2_X1 port map( A1 => ADD_CHECK2(1), A2 => ADD_CHECK2(2), ZN => 
                           n152);
   U113 : INV_X1 port map( A => ADD_CHECK2(2), ZN => n256);
   U114 : INV_X1 port map( A => ADD_CHECK2(1), ZN => n150);
   U115 : NAND2_X1 port map( A1 => n150, A2 => ADD_CHECK2(2), ZN => n156);
   U116 : NOR3_X1 port map( A1 => Table_4_1_port, A2 => Table_4_0_port, A3 => 
                           Table_4_2_port, ZN => n184);
   U117 : NAND3_X1 port map( A1 => n26, A2 => n18, A3 => n12, ZN => n181);
   U118 : NOR3_X1 port map( A1 => Table_2_1_port, A2 => Table_2_0_port, A3 => 
                           Table_2_2_port, ZN => n178);
   U119 : NAND2_X1 port map( A1 => ADD_CHECK2(1), A2 => n256, ZN => n235);
   U120 : NOR3_X1 port map( A1 => Table_6_1_port, A2 => Table_6_0_port, A3 => 
                           Table_6_2_port, ZN => n179);
   U121 : NAND2_X1 port map( A1 => ADD_CHECK2(1), A2 => ADD_CHECK2(2), ZN => 
                           n233);
   U122 : OAI22_X1 port map( A1 => n178, A2 => n235, B1 => n179, B2 => n233, ZN
                           => n151);
   U123 : AOI211_X1 port map( C1 => n152, C2 => n181, A => ADD_CHECK2(4), B => 
                           n151, ZN => n153);
   U124 : AOI221_X1 port map( B1 => n184, B2 => n153, C1 => n156, C2 => n153, A
                           => ADD_CHECK2(3), ZN => n154);
   U125 : INV_X1 port map( A => n154, ZN => n155);
   U126 : AOI221_X1 port map( B1 => n157, B2 => n156, C1 => n157, C2 => n169, A
                           => n155, ZN => n158);
   U127 : INV_X1 port map( A => n158, ZN => n264);
   U128 : OAI22_X1 port map( A1 => n172, A2 => n235, B1 => n173, B2 => n233, ZN
                           => n160);
   U129 : OAI211_X1 port map( C1 => n160, C2 => n159, A => ADD_CHECK2(3), B => 
                           n218, ZN => n263);
   U130 : NOR2_X1 port map( A1 => ADD_CHECK1(1), A2 => ADD_CHECK1(2), ZN => 
                           n192);
   U131 : INV_X1 port map( A => ADD_CHECK1(3), ZN => n190);
   U132 : NAND2_X1 port map( A1 => ADD_CHECK1(1), A2 => ADD_CHECK1(2), ZN => 
                           n208);
   U133 : INV_X1 port map( A => ADD_CHECK1(1), ZN => n163);
   U134 : NOR2_X1 port map( A1 => ADD_CHECK1(2), A2 => n163, ZN => n200);
   U135 : INV_X1 port map( A => n200, ZN => n177);
   U136 : AOI211_X1 port map( C1 => n253, C2 => n192, A => n190, B => n161, ZN 
                           => n162);
   U137 : INV_X1 port map( A => n162, ZN => n171);
   U138 : NAND2_X1 port map( A1 => n163, A2 => ADD_CHECK1(2), ZN => n183);
   U139 : INV_X1 port map( A => n183, ZN => n196);
   U140 : OAI22_X1 port map( A1 => n165, A2 => n208, B1 => n177, B2 => n164, ZN
                           => n166);
   U141 : AOI211_X1 port map( C1 => n192, C2 => n167, A => ADD_CHECK1(3), B => 
                           n166, ZN => n168);
   U142 : OAI21_X1 port map( B1 => n169, B2 => n183, A => n168, ZN => n170);
   U143 : OAI221_X1 port map( B1 => n171, B2 => n196, C1 => n171, C2 => n242, A
                           => n170, ZN => n189);
   U144 : INV_X1 port map( A => ADD_CHECK1(4), ZN => n191);
   U145 : INV_X1 port map( A => n192, ZN => n176);
   U146 : OAI22_X1 port map( A1 => n208, A2 => n173, B1 => n172, B2 => n177, ZN
                           => n174);
   U147 : INV_X1 port map( A => n174, ZN => n175);
   U148 : OAI22_X1 port map( A1 => n179, A2 => n208, B1 => n178, B2 => n177, ZN
                           => n180);
   U149 : AOI211_X1 port map( C1 => n192, C2 => n181, A => ADD_CHECK1(3), B => 
                           n180, ZN => n182);
   U150 : OAI21_X1 port map( B1 => n184, B2 => n183, A => n182, ZN => n185);
   U151 : OAI221_X1 port map( B1 => n187, B2 => n196, C1 => n187, C2 => n186, A
                           => n185, ZN => n188);
   U152 : AOI221_X1 port map( B1 => ADD_CHECK1(4), B2 => n189, C1 => n191, C2 
                           => n188, A => ADD_CHECK1(0), ZN => n261);
   U153 : NAND3_X1 port map( A1 => ADD_CHECK1(4), A2 => ADD_CHECK1(0), A3 => 
                           n190, ZN => n203);
   U154 : NAND3_X1 port map( A1 => ADD_CHECK1(0), A2 => ADD_CHECK1(4), A3 => 
                           ADD_CHECK1(3), ZN => n204);
   U155 : OAI22_X1 port map( A1 => n250, A2 => n203, B1 => n248, B2 => n204, ZN
                           => n194);
   U156 : NAND3_X1 port map( A1 => ADD_CHECK1(0), A2 => ADD_CHECK1(3), A3 => 
                           n191, ZN => n207);
   U157 : NOR3_X1 port map( A1 => Table_1_1_port, A2 => Table_1_0_port, A3 => 
                           Table_1_2_port, ZN => n244);
   U158 : NAND3_X1 port map( A1 => ADD_CHECK1(0), A2 => n191, A3 => n190, ZN =>
                           n205);
   U159 : OAI22_X1 port map( A1 => n246, A2 => n207, B1 => n244, B2 => n205, ZN
                           => n193);
   U160 : OAI21_X1 port map( B1 => n194, B2 => n193, A => n192, ZN => n215);
   U161 : OAI22_X1 port map( A1 => n239, A2 => n204, B1 => n195, B2 => n203, ZN
                           => n198);
   U162 : NOR3_X1 port map( A1 => Table_5_1_port, A2 => Table_5_0_port, A3 => 
                           Table_5_2_port, ZN => n237);
   U163 : OAI22_X1 port map( A1 => n237, A2 => n205, B1 => n238, B2 => n207, ZN
                           => n197);
   U164 : OAI21_X1 port map( B1 => n198, B2 => n197, A => n196, ZN => n214);
   U165 : OAI22_X1 port map( A1 => n217, A2 => n204, B1 => n203, B2 => n220, ZN
                           => n202);
   U166 : NAND3_X1 port map( A1 => n29, A2 => n21, A3 => n15, ZN => n223);
   U167 : INV_X1 port map( A => n223, ZN => n199);
   U168 : OAI22_X1 port map( A1 => n216, A2 => n207, B1 => n199, B2 => n205, ZN
                           => n201);
   U169 : OAI21_X1 port map( B1 => n202, B2 => n201, A => n200, ZN => n213);
   U170 : OAI22_X1 port map( A1 => n225, A2 => n204, B1 => n228, B2 => n203, ZN
                           => n211);
   U171 : NAND3_X1 port map( A1 => n28, A2 => n20, A3 => n14, ZN => n231);
   U172 : INV_X1 port map( A => n231, ZN => n206);
   U173 : OAI22_X1 port map( A1 => n224, A2 => n207, B1 => n206, B2 => n205, ZN
                           => n210);
   U174 : INV_X1 port map( A => n208, ZN => n209);
   U175 : OAI21_X1 port map( B1 => n211, B2 => n210, A => n209, ZN => n212);
   U176 : NAND4_X1 port map( A1 => n215, A2 => n214, A3 => n213, A4 => n212, ZN
                           => n260);
   U177 : INV_X1 port map( A => ADD_CHECK2(3), ZN => n219);
   U178 : NAND3_X1 port map( A1 => n219, A2 => n218, A3 => ADD_CHECK2(0), ZN =>
                           n243);
   U179 : INV_X1 port map( A => n243, ZN => n232);
   U180 : NAND3_X1 port map( A1 => ADD_CHECK2(0), A2 => ADD_CHECK2(3), A3 => 
                           ADD_CHECK2(4), ZN => n247);
   U181 : NAND3_X1 port map( A1 => ADD_CHECK2(3), A2 => ADD_CHECK2(0), A3 => 
                           n218, ZN => n245);
   U182 : OAI22_X1 port map( A1 => n217, A2 => n247, B1 => n245, B2 => n216, ZN
                           => n222);
   U183 : NAND3_X1 port map( A1 => ADD_CHECK2(0), A2 => ADD_CHECK2(4), A3 => 
                           n219, ZN => n249);
   U184 : NOR3_X1 port map( A1 => n219, A2 => n218, A3 => ADD_CHECK2(0), ZN => 
                           n254);
   U185 : INV_X1 port map( A => n254, ZN => n226);
   U186 : AOI211_X1 port map( C1 => n232, C2 => n223, A => n222, B => n221, ZN 
                           => n236);
   U187 : OAI22_X1 port map( A1 => n225, A2 => n247, B1 => n224, B2 => n245, ZN
                           => n230);
   U188 : OAI22_X1 port map( A1 => n228, A2 => n249, B1 => n227, B2 => n226, ZN
                           => n229);
   U189 : AOI211_X1 port map( C1 => n232, C2 => n231, A => n230, B => n229, ZN 
                           => n234);
   U190 : OAI22_X1 port map( A1 => n236, A2 => n235, B1 => n234, B2 => n233, ZN
                           => n259);
   U191 : OAI22_X1 port map( A1 => n238, A2 => n245, B1 => n237, B2 => n243, ZN
                           => n241);
   U192 : OAI22_X1 port map( A1 => n195, A2 => n249, B1 => n239, B2 => n247, ZN
                           => n240);
   U193 : AOI211_X1 port map( C1 => n254, C2 => n242, A => n241, B => n240, ZN 
                           => n257);
   U194 : OAI22_X1 port map( A1 => n245, A2 => n246, B1 => n244, B2 => n243, ZN
                           => n252);
   U195 : OAI22_X1 port map( A1 => n250, A2 => n249, B1 => n248, B2 => n247, ZN
                           => n251);
   U196 : AOI211_X1 port map( C1 => n254, C2 => n253, A => n252, B => n251, ZN 
                           => n255);
   U197 : AOI221_X1 port map( B1 => ADD_CHECK2(2), B2 => n257, C1 => n256, C2 
                           => n255, A => ADD_CHECK2(1), ZN => n258);
   U198 : NOR4_X1 port map( A1 => n261, A2 => n260, A3 => n259, A4 => n258, ZN 
                           => n262);
   U199 : OAI221_X1 port map( B1 => ADD_CHECK2(0), B2 => n264, C1 => 
                           ADD_CHECK2(0), C2 => n263, A => n262, ZN => BUSY);
   U200 : NAND2_X1 port map( A1 => ADD_WR1(3), A2 => ADD_WR1(4), ZN => n448);
   U201 : NOR2_X1 port map( A1 => n624, A2 => n448, ZN => n399);
   U202 : INV_X1 port map( A => ADD_WR1(4), ZN => n324);
   U203 : INV_X1 port map( A => ADD_WR2(0), ZN => n276);
   U204 : INV_X1 port map( A => ADD_WR1(3), ZN => n329);
   U205 : AOI22_X1 port map( A1 => n313, A2 => ADD_WR2(1), B1 => ADD_WR2(3), B2
                           => n329, ZN => n265);
   U206 : OAI221_X1 port map( B1 => n313, B2 => ADD_WR2(1), C1 => n329, C2 => 
                           ADD_WR2(3), A => n265, ZN => n266);
   U207 : AOI221_X1 port map( B1 => ADD_WR1(0), B2 => n276, C1 => n312, C2 => 
                           ADD_WR2(0), A => n266, ZN => n267);
   U208 : OAI221_X1 port map( B1 => ADD_WR1(2), B2 => n273, C1 => n314, C2 => 
                           ADD_WR2(2), A => n267, ZN => n268);
   U209 : AOI221_X1 port map( B1 => ADD_WR1(4), B2 => n293, C1 => n324, C2 => 
                           ADD_WR2(4), A => n268, ZN => n271);
   U210 : INV_X1 port map( A => WR1, ZN => n269);
   U211 : AOI21_X1 port map( B1 => n271, B2 => WR2, A => n269, ZN => n622);
   U212 : INV_X1 port map( A => WR2, ZN => n270);
   U213 : NAND2_X1 port map( A1 => ADD_WR2(4), A2 => ADD_WR2(3), ZN => n277);
   U214 : NAND3_X1 port map( A1 => ADD_WR2(2), A2 => ADD_WR2(0), A3 => 
                           ADD_WR2(1), ZN => n302);
   U215 : NOR2_X1 port map( A1 => n277, A2 => n302, ZN => n442);
   U216 : NAND2_X1 port map( A1 => n142, A2 => n442, ZN => n443);
   U217 : INV_X1 port map( A => n443, ZN => n272);
   U218 : AOI211_X1 port map( C1 => n399, C2 => n622, A => RST, B => n272, ZN 
                           => n446);
   U219 : NAND2_X1 port map( A1 => n145, A2 => n142, ZN => n360);
   U220 : INV_X1 port map( A => n360, ZN => n438);
   U221 : NOR2_X1 port map( A1 => ADD_WR2(0), A2 => ADD_WR2(1), ZN => n275);
   U222 : NAND2_X1 port map( A1 => n275, A2 => n273, ZN => n294);
   U223 : NOR2_X1 port map( A1 => n277, A2 => n294, ZN => n501);
   U224 : INV_X1 port map( A => ADD_WR2(1), ZN => n274);
   U225 : NAND3_X1 port map( A1 => ADD_WR2(0), A2 => n273, A3 => n274, ZN => 
                           n295);
   U226 : NOR2_X1 port map( A1 => n277, A2 => n295, ZN => n492);
   U227 : AOI22_X1 port map( A1 => Table_24_0_port, A2 => n501, B1 => 
                           Table_25_0_port, B2 => n492, ZN => n281);
   U228 : NAND3_X1 port map( A1 => ADD_WR2(1), A2 => n273, A3 => n276, ZN => 
                           n296);
   U229 : NOR2_X1 port map( A1 => n277, A2 => n296, ZN => n484);
   U230 : NAND3_X1 port map( A1 => ADD_WR2(0), A2 => ADD_WR2(1), A3 => n273, ZN
                           => n297);
   U231 : NOR2_X1 port map( A1 => n277, A2 => n297, ZN => n476);
   U232 : AOI22_X1 port map( A1 => Table_26_0_port, A2 => n484, B1 => 
                           Table_27_0_port, B2 => n476, ZN => n280);
   U233 : NAND3_X1 port map( A1 => ADD_WR2(0), A2 => ADD_WR2(2), A3 => n274, ZN
                           => n299);
   U234 : NOR2_X1 port map( A1 => n277, A2 => n299, ZN => n460);
   U235 : NAND2_X1 port map( A1 => ADD_WR2(2), A2 => n275, ZN => n298);
   U236 : NOR2_X1 port map( A1 => n277, A2 => n298, ZN => n468);
   U237 : AOI22_X1 port map( A1 => Table_29_0_port, A2 => n460, B1 => 
                           Table_28_0_port, B2 => n468, ZN => n279);
   U238 : NAND3_X1 port map( A1 => ADD_WR2(2), A2 => ADD_WR2(1), A3 => n276, ZN
                           => n300);
   U239 : NOR2_X1 port map( A1 => n277, A2 => n300, ZN => n452);
   U240 : AOI22_X1 port map( A1 => Table_30_0_port, A2 => n452, B1 => 
                           Table_31_0_port, B2 => n442, ZN => n278);
   U241 : NAND4_X1 port map( A1 => n281, A2 => n280, A3 => n279, A4 => n278, ZN
                           => n310);
   U242 : NAND2_X1 port map( A1 => ADD_WR2(4), A2 => n292, ZN => n282);
   U243 : NOR2_X1 port map( A1 => n294, A2 => n282, ZN => n559);
   U244 : NOR2_X1 port map( A1 => n295, A2 => n282, ZN => n551);
   U245 : AOI22_X1 port map( A1 => Table_16_0_port, A2 => n559, B1 => 
                           Table_17_0_port, B2 => n551, ZN => n286);
   U246 : NOR2_X1 port map( A1 => n296, A2 => n282, ZN => n544);
   U247 : NOR2_X1 port map( A1 => n297, A2 => n282, ZN => n537);
   U248 : AOI22_X1 port map( A1 => Table_18_0_port, A2 => n544, B1 => 
                           Table_19_0_port, B2 => n537, ZN => n285);
   U249 : NOR2_X1 port map( A1 => n298, A2 => n282, ZN => n530);
   U250 : NOR2_X1 port map( A1 => n299, A2 => n282, ZN => n523);
   U251 : AOI22_X1 port map( A1 => Table_20_0_port, A2 => n530, B1 => 
                           Table_21_0_port, B2 => n523, ZN => n284);
   U252 : NOR2_X1 port map( A1 => n300, A2 => n282, ZN => n516);
   U253 : NOR2_X1 port map( A1 => n302, A2 => n282, ZN => n509);
   U254 : AOI22_X1 port map( A1 => Table_22_0_port, A2 => n516, B1 => 
                           Table_23_0_port, B2 => n509, ZN => n283);
   U255 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => n309);
   U256 : NAND2_X1 port map( A1 => ADD_WR2(3), A2 => n293, ZN => n287);
   U257 : NOR2_X1 port map( A1 => n294, A2 => n287, ZN => n617);
   U258 : NOR2_X1 port map( A1 => n295, A2 => n287, ZN => n609);
   U259 : AOI22_X1 port map( A1 => Table_8_0_port, A2 => n617, B1 => 
                           Table_9_0_port, B2 => n609, ZN => n291);
   U260 : NOR2_X1 port map( A1 => n296, A2 => n287, ZN => n602);
   U261 : NOR2_X1 port map( A1 => n297, A2 => n287, ZN => n595);
   U262 : AOI22_X1 port map( A1 => Table_10_0_port, A2 => n602, B1 => 
                           Table_11_0_port, B2 => n595, ZN => n290);
   U263 : NOR2_X1 port map( A1 => n298, A2 => n287, ZN => n588);
   U264 : NOR2_X1 port map( A1 => n299, A2 => n287, ZN => n581);
   U265 : AOI22_X1 port map( A1 => Table_12_0_port, A2 => n588, B1 => 
                           Table_13_0_port, B2 => n581, ZN => n289);
   U266 : NOR2_X1 port map( A1 => n300, A2 => n287, ZN => n574);
   U267 : NOR2_X1 port map( A1 => n302, A2 => n287, ZN => n567);
   U268 : AOI22_X1 port map( A1 => Table_14_0_port, A2 => n574, B1 => 
                           Table_15_0_port, B2 => n567, ZN => n288);
   U269 : NAND4_X1 port map( A1 => n291, A2 => n290, A3 => n289, A4 => n288, ZN
                           => n308);
   U270 : NAND2_X1 port map( A1 => n293, A2 => n292, ZN => n301);
   U271 : NOR2_X1 port map( A1 => n294, A2 => n301, ZN => n690);
   U272 : NOR2_X1 port map( A1 => n295, A2 => n301, ZN => n675);
   U273 : AOI22_X1 port map( A1 => Table_0_0_port, A2 => n690, B1 => 
                           Table_1_0_port, B2 => n675, ZN => n306);
   U274 : NOR2_X1 port map( A1 => n296, A2 => n301, ZN => n667);
   U275 : NOR2_X1 port map( A1 => n297, A2 => n301, ZN => n659);
   U276 : AOI22_X1 port map( A1 => Table_2_0_port, A2 => n667, B1 => 
                           Table_3_0_port, B2 => n659, ZN => n305);
   U277 : NOR2_X1 port map( A1 => n298, A2 => n301, ZN => n651);
   U278 : NOR2_X1 port map( A1 => n299, A2 => n301, ZN => n643);
   U279 : AOI22_X1 port map( A1 => Table_4_0_port, A2 => n651, B1 => 
                           Table_5_0_port, B2 => n643, ZN => n304);
   U280 : NOR2_X1 port map( A1 => n300, A2 => n301, ZN => n635);
   U281 : NOR2_X1 port map( A1 => n302, A2 => n301, ZN => n627);
   U282 : AOI22_X1 port map( A1 => Table_6_0_port, A2 => n635, B1 => 
                           Table_7_0_port, B2 => n627, ZN => n303);
   U283 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => n307);
   U284 : NOR4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN 
                           => n362);
   U285 : NAND2_X1 port map( A1 => ADD_WR1(2), A2 => ADD_WR1(0), ZN => n311);
   U286 : AOI22_X1 port map( A1 => n497, A2 => Table_24_0_port, B1 => n489, B2 
                           => Table_25_0_port, ZN => n317);
   U287 : AOI22_X1 port map( A1 => n481, A2 => Table_26_0_port, B1 => n473, B2 
                           => Table_27_0_port, ZN => n316);
   U288 : AOI22_X1 port map( A1 => n465, A2 => Table_28_0_port, B1 => n447, B2 
                           => Table_30_0_port, ZN => n315);
   U289 : NAND3_X1 port map( A1 => n317, A2 => n316, A3 => n315, ZN => n318);
   U290 : AOI21_X1 port map( B1 => n457, B2 => Table_29_0_port, A => n318, ZN 
                           => n338);
   U291 : NOR2_X1 port map( A1 => ADD_WR1(3), A2 => ADD_WR1(4), ZN => n623);
   U292 : AOI22_X1 port map( A1 => n497, A2 => Table_0_0_port, B1 => n489, B2 
                           => Table_1_0_port, ZN => n322);
   U293 : AOI22_X1 port map( A1 => n481, A2 => Table_2_0_port, B1 => n473, B2 
                           => Table_3_0_port, ZN => n321);
   U294 : AOI22_X1 port map( A1 => n465, A2 => Table_4_0_port, B1 => n457, B2 
                           => Table_5_0_port, ZN => n320);
   U295 : AOI22_X1 port map( A1 => n447, A2 => Table_6_0_port, B1 => n405, B2 
                           => Table_7_0_port, ZN => n319);
   U296 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => n323);
   U297 : AOI22_X1 port map( A1 => n623, A2 => n323, B1 => n399, B2 => 
                           Table_31_0_port, ZN => n337);
   U298 : NOR2_X1 port map( A1 => ADD_WR1(3), A2 => n324, ZN => n506);
   U299 : AOI22_X1 port map( A1 => n497, A2 => Table_16_0_port, B1 => n489, B2 
                           => Table_17_0_port, ZN => n328);
   U300 : AOI22_X1 port map( A1 => n481, A2 => Table_18_0_port, B1 => n473, B2 
                           => Table_19_0_port, ZN => n327);
   U301 : AOI22_X1 port map( A1 => n465, A2 => Table_20_0_port, B1 => n457, B2 
                           => Table_21_0_port, ZN => n326);
   U302 : AOI22_X1 port map( A1 => n447, A2 => Table_22_0_port, B1 => n405, B2 
                           => Table_23_0_port, ZN => n325);
   U303 : NAND4_X1 port map( A1 => n328, A2 => n327, A3 => n326, A4 => n325, ZN
                           => n335);
   U304 : NOR2_X1 port map( A1 => ADD_WR1(4), A2 => n329, ZN => n564);
   U305 : AOI22_X1 port map( A1 => n497, A2 => Table_8_0_port, B1 => n489, B2 
                           => Table_9_0_port, ZN => n333);
   U306 : AOI22_X1 port map( A1 => n481, A2 => Table_10_0_port, B1 => n473, B2 
                           => Table_11_0_port, ZN => n332);
   U307 : AOI22_X1 port map( A1 => n465, A2 => Table_12_0_port, B1 => n457, B2 
                           => Table_13_0_port, ZN => n331);
   U308 : AOI22_X1 port map( A1 => n447, A2 => Table_14_0_port, B1 => n405, B2 
                           => Table_15_0_port, ZN => n330);
   U309 : NAND4_X1 port map( A1 => n333, A2 => n332, A3 => n331, A4 => n330, ZN
                           => n334);
   U310 : AOI22_X1 port map( A1 => n506, A2 => n335, B1 => n564, B2 => n334, ZN
                           => n336);
   U311 : OAI211_X1 port map( C1 => n338, C2 => n448, A => n337, B => n336, ZN 
                           => n386);
   U312 : AOI22_X1 port map( A1 => n442, A2 => n684, B1 => n143, B2 => n443, ZN
                           => n339);
   U313 : INV_X1 port map( A => n446, ZN => n389);
   U314 : AOI22_X1 port map( A1 => n446, A2 => n96, B1 => n339, B2 => n389, ZN 
                           => n797);
   U315 : AOI22_X1 port map( A1 => Table_24_1_port, A2 => n501, B1 => 
                           Table_25_1_port, B2 => n492, ZN => n343);
   U316 : AOI22_X1 port map( A1 => Table_26_1_port, A2 => n484, B1 => 
                           Table_27_1_port, B2 => n476, ZN => n342);
   U317 : AOI22_X1 port map( A1 => Table_29_1_port, A2 => n460, B1 => 
                           Table_28_1_port, B2 => n468, ZN => n341);
   U318 : AOI22_X1 port map( A1 => Table_30_1_port, A2 => n452, B1 => 
                           Table_31_1_port, B2 => n442, ZN => n340);
   U319 : NAND4_X1 port map( A1 => n343, A2 => n342, A3 => n341, A4 => n340, ZN
                           => n359);
   U320 : AOI22_X1 port map( A1 => Table_16_1_port, A2 => n559, B1 => 
                           Table_17_1_port, B2 => n551, ZN => n347);
   U321 : AOI22_X1 port map( A1 => Table_18_1_port, A2 => n544, B1 => 
                           Table_19_1_port, B2 => n537, ZN => n346);
   U322 : AOI22_X1 port map( A1 => Table_20_1_port, A2 => n530, B1 => 
                           Table_21_1_port, B2 => n523, ZN => n345);
   U323 : AOI22_X1 port map( A1 => Table_22_1_port, A2 => n516, B1 => 
                           Table_23_1_port, B2 => n509, ZN => n344);
   U324 : NAND4_X1 port map( A1 => n347, A2 => n346, A3 => n345, A4 => n344, ZN
                           => n358);
   U325 : AOI22_X1 port map( A1 => Table_8_1_port, A2 => n617, B1 => 
                           Table_9_1_port, B2 => n609, ZN => n351);
   U326 : AOI22_X1 port map( A1 => Table_10_1_port, A2 => n602, B1 => 
                           Table_11_1_port, B2 => n595, ZN => n350);
   U327 : AOI22_X1 port map( A1 => Table_12_1_port, A2 => n588, B1 => 
                           Table_13_1_port, B2 => n581, ZN => n349);
   U328 : AOI22_X1 port map( A1 => Table_14_1_port, A2 => n574, B1 => 
                           Table_15_1_port, B2 => n567, ZN => n348);
   U329 : NAND4_X1 port map( A1 => n351, A2 => n350, A3 => n349, A4 => n348, ZN
                           => n357);
   U330 : AOI22_X1 port map( A1 => Table_0_1_port, A2 => n690, B1 => 
                           Table_1_1_port, B2 => n675, ZN => n355);
   U331 : AOI22_X1 port map( A1 => Table_2_1_port, A2 => n667, B1 => 
                           Table_3_1_port, B2 => n659, ZN => n354);
   U332 : AOI22_X1 port map( A1 => Table_4_1_port, A2 => n651, B1 => 
                           Table_5_1_port, B2 => n643, ZN => n353);
   U333 : AOI22_X1 port map( A1 => Table_6_1_port, A2 => n635, B1 => 
                           Table_7_1_port, B2 => n627, ZN => n352);
   U334 : NAND4_X1 port map( A1 => n355, A2 => n354, A3 => n353, A4 => n352, ZN
                           => n356);
   U335 : NOR4_X1 port map( A1 => n359, A2 => n358, A3 => n357, A4 => n356, ZN 
                           => n361);
   U336 : NAND2_X1 port map( A1 => n361, A2 => n362, ZN => n440);
   U337 : AOI221_X1 port map( B1 => n362, B2 => n440, C1 => n361, C2 => n440, A
                           => n360, ZN => n687);
   U338 : AOI22_X1 port map( A1 => n497, A2 => Table_24_1_port, B1 => n489, B2 
                           => Table_25_1_port, ZN => n365);
   U339 : AOI22_X1 port map( A1 => n481, A2 => Table_26_1_port, B1 => n473, B2 
                           => Table_27_1_port, ZN => n364);
   U340 : AOI22_X1 port map( A1 => n465, A2 => Table_28_1_port, B1 => n447, B2 
                           => Table_30_1_port, ZN => n363);
   U341 : NAND3_X1 port map( A1 => n365, A2 => n364, A3 => n363, ZN => n366);
   U342 : AOI21_X1 port map( B1 => n457, B2 => Table_29_1_port, A => n366, ZN 
                           => n384);
   U343 : AOI22_X1 port map( A1 => n497, A2 => Table_0_1_port, B1 => n489, B2 
                           => Table_1_1_port, ZN => n370);
   U344 : AOI22_X1 port map( A1 => n481, A2 => Table_2_1_port, B1 => n473, B2 
                           => Table_3_1_port, ZN => n369);
   U345 : AOI22_X1 port map( A1 => n465, A2 => Table_4_1_port, B1 => n457, B2 
                           => Table_5_1_port, ZN => n368);
   U346 : AOI22_X1 port map( A1 => n447, A2 => Table_6_1_port, B1 => n405, B2 
                           => Table_7_1_port, ZN => n367);
   U347 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => n371);
   U348 : AOI22_X1 port map( A1 => Table_31_1_port, A2 => n399, B1 => n623, B2 
                           => n371, ZN => n383);
   U349 : AOI22_X1 port map( A1 => n497, A2 => Table_8_1_port, B1 => n489, B2 
                           => Table_9_1_port, ZN => n375);
   U350 : AOI22_X1 port map( A1 => n481, A2 => Table_10_1_port, B1 => n473, B2 
                           => Table_11_1_port, ZN => n374);
   U351 : AOI22_X1 port map( A1 => n465, A2 => Table_12_1_port, B1 => n457, B2 
                           => Table_13_1_port, ZN => n373);
   U352 : AOI22_X1 port map( A1 => n447, A2 => Table_14_1_port, B1 => n405, B2 
                           => Table_15_1_port, ZN => n372);
   U353 : NAND4_X1 port map( A1 => n375, A2 => n374, A3 => n373, A4 => n372, ZN
                           => n381);
   U354 : AOI22_X1 port map( A1 => n497, A2 => Table_16_1_port, B1 => n489, B2 
                           => Table_17_1_port, ZN => n379);
   U355 : AOI22_X1 port map( A1 => n481, A2 => Table_18_1_port, B1 => n473, B2 
                           => Table_19_1_port, ZN => n378);
   U356 : AOI22_X1 port map( A1 => n465, A2 => Table_20_1_port, B1 => n457, B2 
                           => Table_21_1_port, ZN => n377);
   U357 : AOI22_X1 port map( A1 => n447, A2 => Table_22_1_port, B1 => n405, B2 
                           => Table_23_1_port, ZN => n376);
   U358 : NAND4_X1 port map( A1 => n379, A2 => n378, A3 => n377, A4 => n376, ZN
                           => n380);
   U359 : AOI22_X1 port map( A1 => n564, A2 => n381, B1 => n506, B2 => n380, ZN
                           => n382);
   U360 : OAI211_X1 port map( C1 => n384, C2 => n448, A => n383, B => n382, ZN 
                           => n385);
   U361 : INV_X1 port map( A => n385, ZN => n388);
   U362 : INV_X1 port map( A => n386, ZN => n387);
   U363 : NOR2_X1 port map( A1 => n388, A2 => n387, ZN => n417);
   U364 : AOI211_X1 port map( C1 => n388, C2 => n387, A => RST, B => n417, ZN 
                           => n686);
   U365 : AOI22_X1 port map( A1 => n442, A2 => n1, B1 => n2, B2 => n443, ZN => 
                           n390);
   U366 : AOI22_X1 port map( A1 => n446, A2 => n80, B1 => n390, B2 => n389, ZN 
                           => n796);
   U367 : AOI22_X1 port map( A1 => n497, A2 => Table_24_2_port, B1 => n489, B2 
                           => Table_25_2_port, ZN => n393);
   U368 : AOI22_X1 port map( A1 => n481, A2 => Table_26_2_port, B1 => n473, B2 
                           => Table_27_2_port, ZN => n392);
   U369 : AOI22_X1 port map( A1 => n465, A2 => Table_28_2_port, B1 => n447, B2 
                           => Table_30_2_port, ZN => n391);
   U370 : NAND3_X1 port map( A1 => n393, A2 => n392, A3 => n391, ZN => n394);
   U371 : AOI21_X1 port map( B1 => n457, B2 => Table_29_2_port, A => n394, ZN 
                           => n414);
   U372 : AOI22_X1 port map( A1 => n497, A2 => Table_0_2_port, B1 => n489, B2 
                           => Table_1_2_port, ZN => n398);
   U373 : AOI22_X1 port map( A1 => n481, A2 => Table_2_2_port, B1 => n473, B2 
                           => Table_3_2_port, ZN => n397);
   U374 : AOI22_X1 port map( A1 => n465, A2 => Table_4_2_port, B1 => n457, B2 
                           => Table_5_2_port, ZN => n396);
   U375 : AOI22_X1 port map( A1 => n447, A2 => Table_6_2_port, B1 => n405, B2 
                           => Table_7_2_port, ZN => n395);
   U376 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => n400);
   U377 : AOI22_X1 port map( A1 => n623, A2 => n400, B1 => n399, B2 => 
                           Table_31_2_port, ZN => n413);
   U378 : AOI22_X1 port map( A1 => n497, A2 => Table_16_2_port, B1 => n489, B2 
                           => Table_17_2_port, ZN => n404);
   U379 : AOI22_X1 port map( A1 => n481, A2 => Table_18_2_port, B1 => n473, B2 
                           => Table_19_2_port, ZN => n403);
   U380 : AOI22_X1 port map( A1 => n465, A2 => Table_20_2_port, B1 => n457, B2 
                           => Table_21_2_port, ZN => n402);
   U381 : AOI22_X1 port map( A1 => n447, A2 => Table_22_2_port, B1 => n405, B2 
                           => Table_23_2_port, ZN => n401);
   U382 : NAND4_X1 port map( A1 => n404, A2 => n403, A3 => n402, A4 => n401, ZN
                           => n411);
   U383 : AOI22_X1 port map( A1 => n497, A2 => Table_8_2_port, B1 => n489, B2 
                           => Table_9_2_port, ZN => n409);
   U384 : AOI22_X1 port map( A1 => n481, A2 => Table_10_2_port, B1 => n473, B2 
                           => Table_11_2_port, ZN => n408);
   U385 : AOI22_X1 port map( A1 => n465, A2 => Table_12_2_port, B1 => n457, B2 
                           => Table_13_2_port, ZN => n407);
   U386 : AOI22_X1 port map( A1 => n447, A2 => Table_14_2_port, B1 => n405, B2 
                           => Table_15_2_port, ZN => n406);
   U387 : NAND4_X1 port map( A1 => n409, A2 => n408, A3 => n407, A4 => n406, ZN
                           => n410);
   U388 : AOI22_X1 port map( A1 => n506, A2 => n411, B1 => n564, B2 => n410, ZN
                           => n412);
   U389 : OAI211_X1 port map( C1 => n414, C2 => n448, A => n413, B => n412, ZN 
                           => n416);
   U390 : NOR2_X1 port map( A1 => n417, A2 => n416, ZN => n415);
   U391 : AOI22_X1 port map( A1 => Table_24_2_port, A2 => n501, B1 => 
                           Table_25_2_port, B2 => n492, ZN => n421);
   U392 : AOI22_X1 port map( A1 => Table_26_2_port, A2 => n484, B1 => 
                           Table_27_2_port, B2 => n476, ZN => n420);
   U393 : AOI22_X1 port map( A1 => Table_29_2_port, A2 => n460, B1 => 
                           Table_28_2_port, B2 => n468, ZN => n419);
   U394 : AOI22_X1 port map( A1 => Table_30_2_port, A2 => n452, B1 => 
                           Table_31_2_port, B2 => n442, ZN => n418);
   U395 : NAND4_X1 port map( A1 => n421, A2 => n420, A3 => n419, A4 => n418, ZN
                           => n437);
   U396 : AOI22_X1 port map( A1 => Table_16_2_port, A2 => n559, B1 => 
                           Table_17_2_port, B2 => n551, ZN => n425);
   U397 : AOI22_X1 port map( A1 => Table_18_2_port, A2 => n544, B1 => 
                           Table_19_2_port, B2 => n537, ZN => n424);
   U398 : AOI22_X1 port map( A1 => Table_20_2_port, A2 => n530, B1 => 
                           Table_21_2_port, B2 => n523, ZN => n423);
   U399 : AOI22_X1 port map( A1 => Table_22_2_port, A2 => n516, B1 => 
                           Table_23_2_port, B2 => n509, ZN => n422);
   U400 : NAND4_X1 port map( A1 => n425, A2 => n424, A3 => n423, A4 => n422, ZN
                           => n436);
   U401 : AOI22_X1 port map( A1 => Table_8_2_port, A2 => n617, B1 => 
                           Table_9_2_port, B2 => n609, ZN => n429);
   U402 : AOI22_X1 port map( A1 => Table_10_2_port, A2 => n602, B1 => 
                           Table_11_2_port, B2 => n595, ZN => n428);
   U403 : AOI22_X1 port map( A1 => Table_12_2_port, A2 => n588, B1 => 
                           Table_13_2_port, B2 => n581, ZN => n427);
   U404 : AOI22_X1 port map( A1 => Table_14_2_port, A2 => n574, B1 => 
                           Table_15_2_port, B2 => n567, ZN => n426);
   U405 : NAND4_X1 port map( A1 => n429, A2 => n428, A3 => n427, A4 => n426, ZN
                           => n435);
   U406 : AOI22_X1 port map( A1 => Table_0_2_port, A2 => n690, B1 => 
                           Table_1_2_port, B2 => n675, ZN => n433);
   U407 : AOI22_X1 port map( A1 => Table_2_2_port, A2 => n667, B1 => 
                           Table_3_2_port, B2 => n659, ZN => n432);
   U408 : AOI22_X1 port map( A1 => Table_4_2_port, A2 => n651, B1 => 
                           Table_5_2_port, B2 => n643, ZN => n431);
   U409 : AOI22_X1 port map( A1 => Table_6_2_port, A2 => n635, B1 => 
                           Table_7_2_port, B2 => n627, ZN => n430);
   U410 : NAND4_X1 port map( A1 => n433, A2 => n432, A3 => n431, A4 => n430, ZN
                           => n434);
   U411 : NOR4_X1 port map( A1 => n437, A2 => n436, A3 => n435, A4 => n434, ZN 
                           => n441);
   U412 : OAI21_X1 port map( B1 => n441, B2 => n440, A => n438, ZN => n439);
   U413 : AOI22_X1 port map( A1 => n692, A2 => n443, B1 => n442, B2 => n144, ZN
                           => n445);
   U414 : NAND2_X1 port map( A1 => n446, A2 => Table_31_2_port, ZN => n444);
   U415 : OAI21_X1 port map( B1 => n446, B2 => n445, A => n444, ZN => n795);
   U416 : INV_X1 port map( A => n448, ZN => n449);
   U417 : NAND2_X1 port map( A1 => n449, A2 => n622, ZN => n498);
   U418 : NAND2_X1 port map( A1 => n680, A2 => n452, ZN => n453);
   U419 : OAI211_X1 port map( C1 => n632, C2 => n498, A => n146, B => n453, ZN 
                           => n454);
   U420 : INV_X1 port map( A => n454, ZN => n456);
   U421 : AOI22_X1 port map( A1 => n452, A2 => n684, B1 => n143, B2 => n453, ZN
                           => n450);
   U422 : AOI22_X1 port map( A1 => n456, A2 => n84, B1 => n450, B2 => n454, ZN 
                           => n794);
   U423 : AOI22_X1 port map( A1 => n452, A2 => n1, B1 => n2, B2 => n453, ZN => 
                           n451);
   U424 : AOI22_X1 port map( A1 => n456, A2 => n22, B1 => n451, B2 => n454, ZN 
                           => n793);
   U425 : AOI22_X1 port map( A1 => n692, A2 => n453, B1 => n452, B2 => n144, ZN
                           => n455);
   U426 : AOI22_X1 port map( A1 => n456, A2 => n75, B1 => n455, B2 => n454, ZN 
                           => n792);
   U427 : NAND2_X1 port map( A1 => n680, A2 => n460, ZN => n461);
   U428 : OAI211_X1 port map( C1 => n640, C2 => n498, A => n145, B => n461, ZN 
                           => n462);
   U429 : INV_X1 port map( A => n462, ZN => n464);
   U430 : AOI22_X1 port map( A1 => n460, A2 => n684, B1 => n143, B2 => n461, ZN
                           => n458);
   U431 : AOI22_X1 port map( A1 => n464, A2 => n55, B1 => n458, B2 => n462, ZN 
                           => n791);
   U432 : AOI22_X1 port map( A1 => n460, A2 => n1, B1 => n2, B2 => n461, ZN => 
                           n459);
   U433 : AOI22_X1 port map( A1 => n464, A2 => n31, B1 => n459, B2 => n462, ZN 
                           => n790);
   U434 : AOI22_X1 port map( A1 => n692, A2 => n461, B1 => n460, B2 => n144, ZN
                           => n463);
   U435 : AOI22_X1 port map( A1 => n464, A2 => n76, B1 => n463, B2 => n462, ZN 
                           => n789);
   U436 : NAND2_X1 port map( A1 => n680, A2 => n468, ZN => n469);
   U437 : OAI211_X1 port map( C1 => n648, C2 => n498, A => n146, B => n469, ZN 
                           => n470);
   U438 : INV_X1 port map( A => n470, ZN => n472);
   U439 : AOI22_X1 port map( A1 => n468, A2 => n684, B1 => n143, B2 => n469, ZN
                           => n466);
   U440 : AOI22_X1 port map( A1 => n472, A2 => n19, B1 => n466, B2 => n470, ZN 
                           => n788);
   U441 : AOI22_X1 port map( A1 => n468, A2 => n1, B1 => n2, B2 => n469, ZN => 
                           n467);
   U442 : AOI22_X1 port map( A1 => n472, A2 => n27, B1 => n467, B2 => n470, ZN 
                           => n787);
   U443 : AOI22_X1 port map( A1 => n692, A2 => n469, B1 => n468, B2 => n144, ZN
                           => n471);
   U444 : AOI22_X1 port map( A1 => n472, A2 => n13, B1 => n471, B2 => n470, ZN 
                           => n786);
   U445 : NAND2_X1 port map( A1 => n680, A2 => n476, ZN => n477);
   U446 : OAI211_X1 port map( C1 => n656, C2 => n498, A => n145, B => n477, ZN 
                           => n478);
   U447 : INV_X1 port map( A => n478, ZN => n480);
   U448 : AOI22_X1 port map( A1 => n476, A2 => n684, B1 => n143, B2 => n477, ZN
                           => n474);
   U449 : AOI22_X1 port map( A1 => n480, A2 => n97, B1 => n474, B2 => n478, ZN 
                           => n785);
   U450 : AOI22_X1 port map( A1 => n476, A2 => n1, B1 => n2, B2 => n477, ZN => 
                           n475);
   U451 : AOI22_X1 port map( A1 => n480, A2 => n89, B1 => n475, B2 => n478, ZN 
                           => n784);
   U452 : AOI22_X1 port map( A1 => n692, A2 => n477, B1 => n476, B2 => n144, ZN
                           => n479);
   U453 : AOI22_X1 port map( A1 => n480, A2 => n85, B1 => n479, B2 => n478, ZN 
                           => n783);
   U454 : NAND2_X1 port map( A1 => n680, A2 => n484, ZN => n485);
   U455 : OAI211_X1 port map( C1 => n664, C2 => n498, A => n146, B => n485, ZN 
                           => n486);
   U456 : INV_X1 port map( A => n486, ZN => n488);
   U457 : AOI22_X1 port map( A1 => n484, A2 => n684, B1 => n143, B2 => n485, ZN
                           => n482);
   U458 : AOI22_X1 port map( A1 => n488, A2 => n67, B1 => n482, B2 => n486, ZN 
                           => n782);
   U459 : AOI22_X1 port map( A1 => n484, A2 => n1, B1 => n2, B2 => n485, ZN => 
                           n483);
   U460 : AOI22_X1 port map( A1 => n488, A2 => n56, B1 => n483, B2 => n486, ZN 
                           => n781);
   U461 : AOI22_X1 port map( A1 => n692, A2 => n485, B1 => n484, B2 => n144, ZN
                           => n487);
   U462 : AOI22_X1 port map( A1 => n488, A2 => n47, B1 => n487, B2 => n486, ZN 
                           => n780);
   U463 : NAND2_X1 port map( A1 => n680, A2 => n492, ZN => n493);
   U464 : OAI211_X1 port map( C1 => n672, C2 => n498, A => n145, B => n493, ZN 
                           => n494);
   U465 : INV_X1 port map( A => n494, ZN => n496);
   U466 : AOI22_X1 port map( A1 => n492, A2 => n684, B1 => n143, B2 => n493, ZN
                           => n490);
   U467 : AOI22_X1 port map( A1 => n496, A2 => n36, B1 => n490, B2 => n494, ZN 
                           => n779);
   U468 : AOI22_X1 port map( A1 => n492, A2 => n1, B1 => n2, B2 => n493, ZN => 
                           n491);
   U469 : AOI22_X1 port map( A1 => n496, A2 => n39, B1 => n491, B2 => n494, ZN 
                           => n778);
   U470 : AOI22_X1 port map( A1 => n692, A2 => n493, B1 => n492, B2 => n144, ZN
                           => n495);
   U471 : AOI22_X1 port map( A1 => n496, A2 => n32, B1 => n495, B2 => n494, ZN 
                           => n777);
   U472 : NAND2_X1 port map( A1 => n680, A2 => n501, ZN => n502);
   U473 : OAI211_X1 port map( C1 => n682, C2 => n498, A => n146, B => n502, ZN 
                           => n503);
   U474 : INV_X1 port map( A => n503, ZN => n505);
   U475 : AOI22_X1 port map( A1 => n501, A2 => n684, B1 => n143, B2 => n502, ZN
                           => n499);
   U476 : AOI22_X1 port map( A1 => n505, A2 => n17, B1 => n499, B2 => n503, ZN 
                           => n776);
   U477 : AOI22_X1 port map( A1 => n501, A2 => n1, B1 => n2, B2 => n502, ZN => 
                           n500);
   U478 : AOI22_X1 port map( A1 => n505, A2 => n23, B1 => n500, B2 => n503, ZN 
                           => n775);
   U479 : AOI22_X1 port map( A1 => n692, A2 => n502, B1 => n501, B2 => n689, ZN
                           => n504);
   U480 : AOI22_X1 port map( A1 => n505, A2 => n11, B1 => n504, B2 => n503, ZN 
                           => n774);
   U481 : NAND2_X1 port map( A1 => n506, A2 => n622, ZN => n556);
   U482 : NAND2_X1 port map( A1 => n142, A2 => n509, ZN => n510);
   U483 : OAI211_X1 port map( C1 => n624, C2 => n556, A => n145, B => n510, ZN 
                           => n511);
   U484 : INV_X1 port map( A => n511, ZN => n513);
   U485 : AOI22_X1 port map( A1 => n509, A2 => n684, B1 => n143, B2 => n510, ZN
                           => n507);
   U486 : AOI22_X1 port map( A1 => n513, A2 => n98, B1 => n507, B2 => n511, ZN 
                           => n773);
   U487 : AOI22_X1 port map( A1 => n509, A2 => n1, B1 => n2, B2 => n510, ZN => 
                           n508);
   U488 : AOI22_X1 port map( A1 => n513, A2 => n86, B1 => n508, B2 => n511, ZN 
                           => n772);
   U489 : AOI22_X1 port map( A1 => n692, A2 => n510, B1 => n509, B2 => n689, ZN
                           => n512);
   U490 : AOI22_X1 port map( A1 => n513, A2 => n90, B1 => n512, B2 => n511, ZN 
                           => n771);
   U491 : NAND2_X1 port map( A1 => n680, A2 => n516, ZN => n517);
   U492 : OAI211_X1 port map( C1 => n632, C2 => n556, A => n146, B => n517, ZN 
                           => n518);
   U493 : INV_X1 port map( A => n518, ZN => n520);
   U494 : AOI22_X1 port map( A1 => n516, A2 => n684, B1 => n143, B2 => n517, ZN
                           => n514);
   U495 : AOI22_X1 port map( A1 => n520, A2 => n57, B1 => n514, B2 => n518, ZN 
                           => n770);
   U496 : AOI22_X1 port map( A1 => n516, A2 => n1, B1 => n2, B2 => n517, ZN => 
                           n515);
   U497 : AOI22_X1 port map( A1 => n520, A2 => n68, B1 => n515, B2 => n518, ZN 
                           => n769);
   U498 : AOI22_X1 port map( A1 => n692, A2 => n517, B1 => n516, B2 => n144, ZN
                           => n519);
   U499 : AOI22_X1 port map( A1 => n520, A2 => n48, B1 => n519, B2 => n518, ZN 
                           => n768);
   U500 : NAND2_X1 port map( A1 => n142, A2 => n523, ZN => n524);
   U501 : OAI211_X1 port map( C1 => n640, C2 => n556, A => n146, B => n524, ZN 
                           => n525);
   U502 : INV_X1 port map( A => n525, ZN => n527);
   U503 : AOI22_X1 port map( A1 => n523, A2 => n684, B1 => n143, B2 => n524, ZN
                           => n521);
   U504 : AOI22_X1 port map( A1 => n527, A2 => n16, B1 => n521, B2 => n525, ZN 
                           => n767);
   U505 : AOI22_X1 port map( A1 => n523, A2 => n1, B1 => n2, B2 => n524, ZN => 
                           n522);
   U506 : AOI22_X1 port map( A1 => n527, A2 => n24, B1 => n522, B2 => n525, ZN 
                           => n766);
   U507 : AOI22_X1 port map( A1 => n692, A2 => n524, B1 => n523, B2 => n144, ZN
                           => n526);
   U508 : AOI22_X1 port map( A1 => n527, A2 => n10, B1 => n526, B2 => n525, ZN 
                           => n765);
   U509 : NAND2_X1 port map( A1 => n142, A2 => n530, ZN => n531);
   U510 : OAI211_X1 port map( C1 => n648, C2 => n556, A => n146, B => n531, ZN 
                           => n532);
   U511 : INV_X1 port map( A => n532, ZN => n534);
   U512 : AOI22_X1 port map( A1 => n530, A2 => n684, B1 => n143, B2 => n531, ZN
                           => n528);
   U513 : AOI22_X1 port map( A1 => n534, A2 => n58, B1 => n528, B2 => n532, ZN 
                           => n764);
   U514 : AOI22_X1 port map( A1 => n530, A2 => n1, B1 => n2, B2 => n531, ZN => 
                           n529);
   U515 : AOI22_X1 port map( A1 => n534, A2 => n69, B1 => n529, B2 => n532, ZN 
                           => n763);
   U516 : AOI22_X1 port map( A1 => n692, A2 => n531, B1 => n530, B2 => n144, ZN
                           => n533);
   U517 : AOI22_X1 port map( A1 => n534, A2 => n49, B1 => n533, B2 => n532, ZN 
                           => n762);
   U518 : NAND2_X1 port map( A1 => n142, A2 => n537, ZN => n538);
   U519 : OAI211_X1 port map( C1 => n656, C2 => n556, A => n146, B => n538, ZN 
                           => n539);
   U520 : INV_X1 port map( A => n539, ZN => n541);
   U521 : AOI22_X1 port map( A1 => n537, A2 => n684, B1 => n143, B2 => n538, ZN
                           => n535);
   U522 : AOI22_X1 port map( A1 => n541, A2 => n93, B1 => n535, B2 => n539, ZN 
                           => n761);
   U523 : AOI22_X1 port map( A1 => n537, A2 => n1, B1 => n2, B2 => n538, ZN => 
                           n536);
   U524 : AOI22_X1 port map( A1 => n541, A2 => n81, B1 => n536, B2 => n539, ZN 
                           => n760);
   U525 : AOI22_X1 port map( A1 => n692, A2 => n538, B1 => n537, B2 => n144, ZN
                           => n540);
   U526 : AOI22_X1 port map( A1 => n541, A2 => n101, B1 => n540, B2 => n539, ZN
                           => n759);
   U527 : NAND2_X1 port map( A1 => n142, A2 => n544, ZN => n545);
   U528 : OAI211_X1 port map( C1 => n664, C2 => n556, A => n146, B => n545, ZN 
                           => n546);
   U529 : INV_X1 port map( A => n546, ZN => n548);
   U530 : AOI22_X1 port map( A1 => n544, A2 => n684, B1 => n143, B2 => n545, ZN
                           => n542);
   U531 : AOI22_X1 port map( A1 => n548, A2 => n59, B1 => n542, B2 => n546, ZN 
                           => n758);
   U532 : AOI22_X1 port map( A1 => n544, A2 => n1, B1 => n2, B2 => n545, ZN => 
                           n543);
   U533 : AOI22_X1 port map( A1 => n548, A2 => n70, B1 => n543, B2 => n546, ZN 
                           => n757);
   U534 : AOI22_X1 port map( A1 => n692, A2 => n545, B1 => n544, B2 => n144, ZN
                           => n547);
   U535 : AOI22_X1 port map( A1 => n548, A2 => n50, B1 => n547, B2 => n546, ZN 
                           => n756);
   U536 : NAND2_X1 port map( A1 => n142, A2 => n551, ZN => n552);
   U537 : OAI211_X1 port map( C1 => n672, C2 => n556, A => n146, B => n552, ZN 
                           => n553);
   U538 : INV_X1 port map( A => n553, ZN => n555);
   U539 : AOI22_X1 port map( A1 => n551, A2 => n684, B1 => n143, B2 => n552, ZN
                           => n549);
   U540 : AOI22_X1 port map( A1 => n555, A2 => n37, B1 => n549, B2 => n553, ZN 
                           => n755);
   U541 : AOI22_X1 port map( A1 => n551, A2 => n1, B1 => n2, B2 => n552, ZN => 
                           n550);
   U542 : AOI22_X1 port map( A1 => n555, A2 => n40, B1 => n550, B2 => n553, ZN 
                           => n754);
   U543 : AOI22_X1 port map( A1 => n692, A2 => n552, B1 => n551, B2 => n144, ZN
                           => n554);
   U544 : AOI22_X1 port map( A1 => n555, A2 => n33, B1 => n554, B2 => n553, ZN 
                           => n753);
   U545 : NAND2_X1 port map( A1 => n680, A2 => n559, ZN => n560);
   U546 : OAI211_X1 port map( C1 => n682, C2 => n556, A => n146, B => n560, ZN 
                           => n561);
   U547 : INV_X1 port map( A => n561, ZN => n563);
   U548 : AOI22_X1 port map( A1 => n559, A2 => n684, B1 => n683, B2 => n560, ZN
                           => n557);
   U549 : AOI22_X1 port map( A1 => n563, A2 => n140, B1 => n557, B2 => n561, ZN
                           => n752);
   U550 : AOI22_X1 port map( A1 => n559, A2 => n1, B1 => n2, B2 => n560, ZN => 
                           n558);
   U551 : AOI22_X1 port map( A1 => n563, A2 => n139, B1 => n558, B2 => n561, ZN
                           => n751);
   U552 : AOI22_X1 port map( A1 => n692, A2 => n560, B1 => n559, B2 => n144, ZN
                           => n562);
   U553 : AOI22_X1 port map( A1 => n563, A2 => n141, B1 => n562, B2 => n561, ZN
                           => n750);
   U554 : NAND2_X1 port map( A1 => n564, A2 => n622, ZN => n614);
   U555 : NAND2_X1 port map( A1 => n142, A2 => n567, ZN => n568);
   U556 : OAI211_X1 port map( C1 => n624, C2 => n614, A => n146, B => n568, ZN 
                           => n569);
   U557 : INV_X1 port map( A => n569, ZN => n571);
   U558 : AOI22_X1 port map( A1 => n567, A2 => n684, B1 => n683, B2 => n568, ZN
                           => n565);
   U559 : AOI22_X1 port map( A1 => n571, A2 => n99, B1 => n565, B2 => n569, ZN 
                           => n749);
   U560 : AOI22_X1 port map( A1 => n567, A2 => n1, B1 => n2, B2 => n568, ZN => 
                           n566);
   U561 : AOI22_X1 port map( A1 => n571, A2 => n91, B1 => n566, B2 => n569, ZN 
                           => n748);
   U562 : AOI22_X1 port map( A1 => n692, A2 => n568, B1 => n567, B2 => n144, ZN
                           => n570);
   U563 : AOI22_X1 port map( A1 => n571, A2 => n87, B1 => n570, B2 => n569, ZN 
                           => n747);
   U564 : NAND2_X1 port map( A1 => n142, A2 => n574, ZN => n575);
   U565 : OAI211_X1 port map( C1 => n632, C2 => n614, A => n146, B => n575, ZN 
                           => n576);
   U566 : INV_X1 port map( A => n576, ZN => n578);
   U567 : AOI22_X1 port map( A1 => n574, A2 => n684, B1 => n143, B2 => n575, ZN
                           => n572);
   U568 : AOI22_X1 port map( A1 => n578, A2 => n60, B1 => n572, B2 => n576, ZN 
                           => n746);
   U569 : AOI22_X1 port map( A1 => n574, A2 => n1, B1 => n2, B2 => n575, ZN => 
                           n573);
   U570 : AOI22_X1 port map( A1 => n578, A2 => n71, B1 => n573, B2 => n576, ZN 
                           => n745);
   U571 : AOI22_X1 port map( A1 => n692, A2 => n575, B1 => n574, B2 => n144, ZN
                           => n577);
   U572 : AOI22_X1 port map( A1 => n578, A2 => n51, B1 => n577, B2 => n576, ZN 
                           => n744);
   U573 : NAND2_X1 port map( A1 => n142, A2 => n581, ZN => n582);
   U574 : OAI211_X1 port map( C1 => n640, C2 => n614, A => n146, B => n582, ZN 
                           => n583);
   U575 : INV_X1 port map( A => n583, ZN => n585);
   U576 : AOI22_X1 port map( A1 => n581, A2 => n684, B1 => n143, B2 => n582, ZN
                           => n579);
   U577 : AOI22_X1 port map( A1 => n585, A2 => n38, B1 => n579, B2 => n583, ZN 
                           => n743);
   U578 : AOI22_X1 port map( A1 => n581, A2 => n1, B1 => n2, B2 => n582, ZN => 
                           n580);
   U579 : AOI22_X1 port map( A1 => n585, A2 => n35, B1 => n580, B2 => n583, ZN 
                           => n742);
   U580 : AOI22_X1 port map( A1 => n692, A2 => n582, B1 => n581, B2 => n144, ZN
                           => n584);
   U581 : AOI22_X1 port map( A1 => n585, A2 => n34, B1 => n584, B2 => n583, ZN 
                           => n741);
   U582 : NAND2_X1 port map( A1 => n142, A2 => n588, ZN => n589);
   U583 : OAI211_X1 port map( C1 => n648, C2 => n614, A => n146, B => n589, ZN 
                           => n590);
   U584 : INV_X1 port map( A => n590, ZN => n592);
   U585 : AOI22_X1 port map( A1 => n588, A2 => n684, B1 => n143, B2 => n589, ZN
                           => n586);
   U586 : AOI22_X1 port map( A1 => n592, A2 => n61, B1 => n586, B2 => n590, ZN 
                           => n740);
   U587 : AOI22_X1 port map( A1 => n588, A2 => n1, B1 => n2, B2 => n589, ZN => 
                           n587);
   U588 : AOI22_X1 port map( A1 => n592, A2 => n72, B1 => n587, B2 => n590, ZN 
                           => n739);
   U589 : AOI22_X1 port map( A1 => n692, A2 => n589, B1 => n588, B2 => n144, ZN
                           => n591);
   U590 : AOI22_X1 port map( A1 => n592, A2 => n52, B1 => n591, B2 => n590, ZN 
                           => n738);
   U591 : NAND2_X1 port map( A1 => n142, A2 => n595, ZN => n596);
   U592 : OAI211_X1 port map( C1 => n656, C2 => n614, A => n146, B => n596, ZN 
                           => n597);
   U593 : INV_X1 port map( A => n597, ZN => n599);
   U594 : AOI22_X1 port map( A1 => n595, A2 => n684, B1 => n143, B2 => n596, ZN
                           => n593);
   U595 : AOI22_X1 port map( A1 => n599, A2 => n100, B1 => n593, B2 => n597, ZN
                           => n737);
   U596 : AOI22_X1 port map( A1 => n595, A2 => n1, B1 => n2, B2 => n596, ZN => 
                           n594);
   U597 : AOI22_X1 port map( A1 => n599, A2 => n92, B1 => n594, B2 => n597, ZN 
                           => n736);
   U598 : AOI22_X1 port map( A1 => n692, A2 => n596, B1 => n595, B2 => n144, ZN
                           => n598);
   U599 : AOI22_X1 port map( A1 => n599, A2 => n88, B1 => n598, B2 => n597, ZN 
                           => n735);
   U600 : NAND2_X1 port map( A1 => n142, A2 => n602, ZN => n603);
   U601 : OAI211_X1 port map( C1 => n664, C2 => n614, A => n145, B => n603, ZN 
                           => n604);
   U602 : INV_X1 port map( A => n604, ZN => n606);
   U603 : AOI22_X1 port map( A1 => n602, A2 => n684, B1 => n143, B2 => n603, ZN
                           => n600);
   U604 : AOI22_X1 port map( A1 => n606, A2 => n62, B1 => n600, B2 => n604, ZN 
                           => n734);
   U605 : AOI22_X1 port map( A1 => n602, A2 => n1, B1 => n2, B2 => n603, ZN => 
                           n601);
   U606 : AOI22_X1 port map( A1 => n606, A2 => n73, B1 => n601, B2 => n604, ZN 
                           => n733);
   U607 : AOI22_X1 port map( A1 => n692, A2 => n603, B1 => n602, B2 => n144, ZN
                           => n605);
   U608 : AOI22_X1 port map( A1 => n606, A2 => n53, B1 => n605, B2 => n604, ZN 
                           => n732);
   U609 : NAND2_X1 port map( A1 => n142, A2 => n609, ZN => n610);
   U610 : OAI211_X1 port map( C1 => n672, C2 => n614, A => n145, B => n610, ZN 
                           => n611);
   U611 : INV_X1 port map( A => n611, ZN => n613);
   U612 : AOI22_X1 port map( A1 => n609, A2 => n684, B1 => n683, B2 => n610, ZN
                           => n607);
   U613 : AOI22_X1 port map( A1 => n613, A2 => n41, B1 => n607, B2 => n611, ZN 
                           => n731);
   U614 : AOI22_X1 port map( A1 => n609, A2 => n1, B1 => n686, B2 => n610, ZN 
                           => n608);
   U615 : AOI22_X1 port map( A1 => n613, A2 => n43, B1 => n608, B2 => n611, ZN 
                           => n730);
   U616 : AOI22_X1 port map( A1 => n692, A2 => n610, B1 => n609, B2 => n689, ZN
                           => n612);
   U617 : AOI22_X1 port map( A1 => n613, A2 => n42, B1 => n612, B2 => n611, ZN 
                           => n729);
   U618 : NAND2_X1 port map( A1 => n142, A2 => n617, ZN => n618);
   U619 : OAI211_X1 port map( C1 => n682, C2 => n614, A => n145, B => n618, ZN 
                           => n619);
   U620 : INV_X1 port map( A => n619, ZN => n621);
   U621 : AOI22_X1 port map( A1 => n617, A2 => n684, B1 => n683, B2 => n618, ZN
                           => n615);
   U622 : AOI22_X1 port map( A1 => n621, A2 => n63, B1 => n615, B2 => n619, ZN 
                           => n728);
   U623 : AOI22_X1 port map( A1 => n617, A2 => n1, B1 => n2, B2 => n618, ZN => 
                           n616);
   U624 : AOI22_X1 port map( A1 => n621, A2 => n74, B1 => n616, B2 => n619, ZN 
                           => n727);
   U625 : AOI22_X1 port map( A1 => n692, A2 => n618, B1 => n617, B2 => n144, ZN
                           => n620);
   U626 : AOI22_X1 port map( A1 => n621, A2 => n54, B1 => n620, B2 => n619, ZN 
                           => n726);
   U627 : NAND2_X1 port map( A1 => n623, A2 => n622, ZN => n681);
   U628 : NAND2_X1 port map( A1 => n142, A2 => n627, ZN => n628);
   U629 : OAI211_X1 port map( C1 => n624, C2 => n681, A => n145, B => n628, ZN 
                           => n629);
   U630 : INV_X1 port map( A => n629, ZN => n631);
   U631 : AOI22_X1 port map( A1 => n627, A2 => n684, B1 => n143, B2 => n628, ZN
                           => n625);
   U632 : AOI22_X1 port map( A1 => n631, A2 => n20, B1 => n625, B2 => n629, ZN 
                           => n725);
   U633 : AOI22_X1 port map( A1 => n627, A2 => n1, B1 => n2, B2 => n628, ZN => 
                           n626);
   U634 : AOI22_X1 port map( A1 => n631, A2 => n28, B1 => n626, B2 => n629, ZN 
                           => n724);
   U635 : AOI22_X1 port map( A1 => n692, A2 => n628, B1 => n627, B2 => n689, ZN
                           => n630);
   U636 : AOI22_X1 port map( A1 => n631, A2 => n14, B1 => n630, B2 => n629, ZN 
                           => n723);
   U637 : NAND2_X1 port map( A1 => n142, A2 => n635, ZN => n636);
   U638 : OAI211_X1 port map( C1 => n632, C2 => n681, A => n145, B => n636, ZN 
                           => n637);
   U639 : INV_X1 port map( A => n637, ZN => n639);
   U640 : AOI22_X1 port map( A1 => n635, A2 => n684, B1 => n683, B2 => n636, ZN
                           => n633);
   U641 : AOI22_X1 port map( A1 => n639, A2 => n64, B1 => n633, B2 => n637, ZN 
                           => n722);
   U642 : AOI22_X1 port map( A1 => n635, A2 => n1, B1 => n686, B2 => n636, ZN 
                           => n634);
   U643 : AOI22_X1 port map( A1 => n639, A2 => n44, B1 => n634, B2 => n637, ZN 
                           => n721);
   U644 : AOI22_X1 port map( A1 => n692, A2 => n636, B1 => n635, B2 => n689, ZN
                           => n638);
   U645 : AOI22_X1 port map( A1 => n639, A2 => n77, B1 => n638, B2 => n637, ZN 
                           => n720);
   U646 : NAND2_X1 port map( A1 => n142, A2 => n643, ZN => n644);
   U647 : OAI211_X1 port map( C1 => n640, C2 => n681, A => n145, B => n644, ZN 
                           => n645);
   U648 : INV_X1 port map( A => n645, ZN => n647);
   U649 : AOI22_X1 port map( A1 => n643, A2 => n684, B1 => n683, B2 => n644, ZN
                           => n641);
   U650 : AOI22_X1 port map( A1 => n647, A2 => n94, B1 => n641, B2 => n645, ZN 
                           => n719);
   U651 : AOI22_X1 port map( A1 => n643, A2 => n1, B1 => n2, B2 => n644, ZN => 
                           n642);
   U652 : AOI22_X1 port map( A1 => n647, A2 => n82, B1 => n642, B2 => n645, ZN 
                           => n718);
   U653 : AOI22_X1 port map( A1 => n692, A2 => n644, B1 => n643, B2 => n689, ZN
                           => n646);
   U654 : AOI22_X1 port map( A1 => n647, A2 => n102, B1 => n646, B2 => n645, ZN
                           => n717);
   U655 : NAND2_X1 port map( A1 => n142, A2 => n651, ZN => n652);
   U656 : OAI211_X1 port map( C1 => n648, C2 => n681, A => n145, B => n652, ZN 
                           => n653);
   U657 : INV_X1 port map( A => n653, ZN => n655);
   U658 : AOI22_X1 port map( A1 => n651, A2 => n684, B1 => n683, B2 => n652, ZN
                           => n649);
   U659 : AOI22_X1 port map( A1 => n655, A2 => n65, B1 => n649, B2 => n653, ZN 
                           => n716);
   U660 : AOI22_X1 port map( A1 => n651, A2 => n1, B1 => n686, B2 => n652, ZN 
                           => n650);
   U661 : AOI22_X1 port map( A1 => n655, A2 => n45, B1 => n650, B2 => n653, ZN 
                           => n715);
   U662 : AOI22_X1 port map( A1 => n692, A2 => n652, B1 => n651, B2 => n689, ZN
                           => n654);
   U663 : AOI22_X1 port map( A1 => n655, A2 => n78, B1 => n654, B2 => n653, ZN 
                           => n714);
   U664 : NAND2_X1 port map( A1 => n142, A2 => n659, ZN => n660);
   U665 : OAI211_X1 port map( C1 => n656, C2 => n681, A => n145, B => n660, ZN 
                           => n661);
   U666 : INV_X1 port map( A => n661, ZN => n663);
   U667 : AOI22_X1 port map( A1 => n659, A2 => n684, B1 => n683, B2 => n660, ZN
                           => n657);
   U668 : AOI22_X1 port map( A1 => n663, A2 => n21, B1 => n657, B2 => n661, ZN 
                           => n713);
   U669 : AOI22_X1 port map( A1 => n659, A2 => n1, B1 => n2, B2 => n660, ZN => 
                           n658);
   U670 : AOI22_X1 port map( A1 => n663, A2 => n29, B1 => n658, B2 => n661, ZN 
                           => n712);
   U671 : AOI22_X1 port map( A1 => n692, A2 => n660, B1 => n659, B2 => n689, ZN
                           => n662);
   U672 : AOI22_X1 port map( A1 => n663, A2 => n15, B1 => n662, B2 => n661, ZN 
                           => n711);
   U673 : NAND2_X1 port map( A1 => n142, A2 => n667, ZN => n668);
   U674 : OAI211_X1 port map( C1 => n664, C2 => n681, A => n145, B => n668, ZN 
                           => n669);
   U675 : INV_X1 port map( A => n669, ZN => n671);
   U676 : AOI22_X1 port map( A1 => n667, A2 => n684, B1 => n683, B2 => n668, ZN
                           => n665);
   U677 : AOI22_X1 port map( A1 => n671, A2 => n66, B1 => n665, B2 => n669, ZN 
                           => n710);
   U678 : AOI22_X1 port map( A1 => n667, A2 => n1, B1 => n686, B2 => n668, ZN 
                           => n666);
   U679 : AOI22_X1 port map( A1 => n671, A2 => n46, B1 => n666, B2 => n669, ZN 
                           => n709);
   U680 : AOI22_X1 port map( A1 => n692, A2 => n668, B1 => n667, B2 => n689, ZN
                           => n670);
   U681 : AOI22_X1 port map( A1 => n671, A2 => n79, B1 => n670, B2 => n669, ZN 
                           => n708);
   U682 : NAND2_X1 port map( A1 => n142, A2 => n675, ZN => n676);
   U683 : OAI211_X1 port map( C1 => n672, C2 => n681, A => n145, B => n676, ZN 
                           => n677);
   U684 : INV_X1 port map( A => n677, ZN => n679);
   U685 : AOI22_X1 port map( A1 => n675, A2 => n684, B1 => n683, B2 => n676, ZN
                           => n673);
   U686 : AOI22_X1 port map( A1 => n679, A2 => n95, B1 => n673, B2 => n677, ZN 
                           => n707);
   U687 : AOI22_X1 port map( A1 => n675, A2 => n1, B1 => n2, B2 => n676, ZN => 
                           n674);
   U688 : AOI22_X1 port map( A1 => n679, A2 => n83, B1 => n674, B2 => n677, ZN 
                           => n706);
   U689 : AOI22_X1 port map( A1 => n692, A2 => n676, B1 => n675, B2 => n689, ZN
                           => n678);
   U690 : AOI22_X1 port map( A1 => n679, A2 => n103, B1 => n678, B2 => n677, ZN
                           => n705);
   U691 : NAND2_X1 port map( A1 => n680, A2 => n690, ZN => n691);
   U692 : OAI211_X1 port map( C1 => n682, C2 => n681, A => n145, B => n691, ZN 
                           => n693);
   U693 : INV_X1 port map( A => n693, ZN => n695);
   U694 : AOI22_X1 port map( A1 => n690, A2 => n684, B1 => n143, B2 => n691, ZN
                           => n685);
   U695 : AOI22_X1 port map( A1 => n695, A2 => n18, B1 => n685, B2 => n693, ZN 
                           => n704);
   U696 : AOI22_X1 port map( A1 => n690, A2 => n1, B1 => n2, B2 => n691, ZN => 
                           n688);
   U697 : AOI22_X1 port map( A1 => n695, A2 => n26, B1 => n688, B2 => n693, ZN 
                           => n703);
   U698 : AOI22_X1 port map( A1 => n692, A2 => n691, B1 => n690, B2 => n144, ZN
                           => n694);
   U699 : AOI22_X1 port map( A1 => n695, A2 => n12, B1 => n694, B2 => n693, ZN 
                           => n702);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32.all;

entity DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32 is

   port( CLK, RST : in std_logic;  IRAM_ADDRESS : out std_logic_vector (31 
         downto 0);  IRAM_ISSUE : out std_logic;  IRAM_READY : in std_logic;  
         IRAM_DATA : in std_logic_vector (31 downto 0);  DRAM_ADDRESS : out 
         std_logic_vector (31 downto 0);  DRAM_ISSUE, DRAM_READNOTWRITE : out 
         std_logic;  DRAM_READY : in std_logic;  DRAM_DATA_IN : in 
         std_logic_vector (31 downto 0);  DRAM_DATA_OUT : out std_logic_vector 
         (31 downto 0);  DATA_SIZE : out std_logic_vector (1 downto 0);  
         DRAMRF_ADDRESS : out std_logic_vector (31 downto 0);  DRAMRF_ISSUE, 
         DRAMRF_READNOTWRITE : out std_logic;  DRAMRF_READY : in std_logic;  
         DRAMRF_DATA_IN : in std_logic_vector (31 downto 0);  DRAMRF_DATA_OUT :
         out std_logic_vector (31 downto 0);  DATA_SIZE_RF : out 
         std_logic_vector (1 downto 0));

end DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32_RAM_DEPTH32 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X4
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X2
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X4
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X2
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component select_block_NBIT_DATA32_N8_F5
      port( regs : in std_logic_vector (2559 downto 0);  win : in 
            std_logic_vector (4 downto 0);  curr_proc_regs : out 
            std_logic_vector (767 downto 0));
   end component;
   
   component mux_N32_M5_0
      port( S : in std_logic_vector (4 downto 0);  Q : in std_logic_vector 
            (1023 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component mux_N32_M5_1
      port( S : in std_logic_vector (4 downto 0);  Q : in std_logic_vector 
            (1023 downto 0);  Y : out std_logic_vector (31 downto 0));
   end component;
   
   component in_loc_selblock_NBIT_DATA32_N8_F5
      port( regs : in std_logic_vector (2559 downto 0);  win : in 
            std_logic_vector (4 downto 0);  curr_proc_regs : out 
            std_logic_vector (511 downto 0));
   end component;
   
   component hazard_table_N_REGS_LOG5
      port( CLK, RST, WR1, WR2 : in std_logic;  ADD_WR1, ADD_WR2, ADD_CHECK1, 
            ADD_CHECK2 : in std_logic_vector (4 downto 0);  BUSY, BUSY_WINDOW :
            out std_logic);
   end component;
   
   signal IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, IRAM_ADDRESS_29_port, 
      IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, IRAM_ADDRESS_26_port, 
      IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, IRAM_ADDRESS_23_port, 
      IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, IRAM_ADDRESS_20_port, 
      IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, IRAM_ADDRESS_17_port, 
      IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, IRAM_ADDRESS_14_port, 
      IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, IRAM_ADDRESS_11_port, 
      IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, IRAM_ADDRESS_8_port, 
      IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, IRAM_ADDRESS_5_port, 
      IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, IRAM_ADDRESS_2_port, 
      IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port, DRAM_ADDRESS_31_port, 
      DRAM_ADDRESS_30_port, DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, 
      DRAM_ADDRESS_27_port, DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, 
      DRAM_ADDRESS_24_port, DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, 
      DRAM_ADDRESS_21_port, DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, 
      DRAM_ADDRESS_18_port, DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, 
      DRAM_ADDRESS_15_port, DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, 
      DRAM_ADDRESS_12_port, DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, 
      DRAM_ADDRESS_9_port, DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, 
      DRAM_ADDRESS_6_port, DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, 
      DRAM_ADDRESS_3_port, DRAM_ADDRESS_2_port, DRAM_ADDRESS_1_port, 
      DRAM_ADDRESS_0_port, DRAM_DATA_OUT_31_port, DRAM_DATA_OUT_30_port, 
      DRAM_DATA_OUT_29_port, DRAM_DATA_OUT_28_port, DRAM_DATA_OUT_27_port, 
      DRAM_DATA_OUT_26_port, DRAM_DATA_OUT_25_port, DRAM_DATA_OUT_24_port, 
      DRAM_DATA_OUT_23_port, DRAM_DATA_OUT_22_port, DRAM_DATA_OUT_21_port, 
      DRAM_DATA_OUT_20_port, DRAM_DATA_OUT_19_port, DRAM_DATA_OUT_18_port, 
      DRAM_DATA_OUT_17_port, DRAM_DATA_OUT_16_port, DRAM_DATA_OUT_15_port, 
      DRAM_DATA_OUT_14_port, DRAM_DATA_OUT_13_port, DRAM_DATA_OUT_12_port, 
      DRAM_DATA_OUT_11_port, DRAM_DATA_OUT_10_port, DRAM_DATA_OUT_9_port, 
      DRAM_DATA_OUT_8_port, DRAM_DATA_OUT_7_port, DRAM_DATA_OUT_6_port, 
      DRAM_DATA_OUT_5_port, DRAM_DATA_OUT_4_port, DRAM_DATA_OUT_3_port, 
      DRAM_DATA_OUT_2_port, DRAM_DATA_OUT_1_port, DRAM_DATA_OUT_0_port, 
      DATA_SIZE_1_port, DATA_SIZE_0_port, DRAMRF_ADDRESS_31_port, 
      DRAMRF_ADDRESS_30_port, DRAMRF_ADDRESS_29_port, DRAMRF_ADDRESS_28_port, 
      DRAMRF_ADDRESS_27_port, DRAMRF_ADDRESS_26_port, DRAMRF_ADDRESS_25_port, 
      DRAMRF_ADDRESS_24_port, DRAMRF_ADDRESS_23_port, DRAMRF_ADDRESS_22_port, 
      DRAMRF_ADDRESS_21_port, DRAMRF_ADDRESS_20_port, DRAMRF_ADDRESS_19_port, 
      DRAMRF_ADDRESS_18_port, DRAMRF_ADDRESS_17_port, DRAMRF_ADDRESS_16_port, 
      DRAMRF_ADDRESS_15_port, DRAMRF_ADDRESS_14_port, DRAMRF_ADDRESS_13_port, 
      DRAMRF_ADDRESS_12_port, DRAMRF_ADDRESS_11_port, DRAMRF_ADDRESS_10_port, 
      DRAMRF_ADDRESS_9_port, DRAMRF_ADDRESS_8_port, DRAMRF_ADDRESS_7_port, 
      DRAMRF_ADDRESS_6_port, DRAMRF_ADDRESS_5_port, DRAMRF_ADDRESS_4_port, 
      DRAMRF_ADDRESS_3_port, DRAMRF_ADDRESS_2_port, DRAMRF_ADDRESS_1_port, 
      i_DATAMEM_WM, IR_29_port, IR_26_port, IR_24_port, IR_21_port, IR_13_port,
      IR_10_port, IR_9_port, IR_8_port, IR_7_port, IR_6_port, IR_5_port, 
      IR_4_port, IR_3_port, IR_2_port, IR_1_port, i_HAZARD_SIG_CU, 
      i_BUSY_WINDOW, i_SEL_CMPB, i_NPC_SEL, i_ALU_OP_4_port, i_ALU_OP_3_port, 
      i_ALU_OP_2_port, i_ALU_OP_1_port, i_ALU_OP_0_port, i_SEL_LGET_1_port, 
      i_SEL_LGET_0_port, i_DATAMEM_RM, i_S3, i_WF, i_RF1, i_RF2, 
      i_ADD_WB_4_port, i_ADD_WB_3_port, i_ADD_WB_2_port, i_ADD_WB_1_port, 
      i_ADD_WB_0_port, i_RD1_31_port, i_RD1_30_port, i_RD1_29_port, 
      i_RD1_28_port, i_RD1_27_port, i_RD1_26_port, i_RD1_25_port, i_RD1_24_port
      , i_RD1_23_port, i_RD1_22_port, i_RD1_21_port, i_RD1_20_port, 
      i_RD1_19_port, i_RD1_18_port, i_RD1_17_port, i_RD1_16_port, i_RD1_15_port
      , i_RD1_14_port, i_RD1_13_port, i_RD1_12_port, i_RD1_11_port, 
      i_RD1_10_port, i_RD1_9_port, i_RD1_8_port, i_RD1_7_port, i_RD1_6_port, 
      i_RD1_5_port, i_RD1_4_port, i_RD1_3_port, i_RD1_2_port, i_RD1_1_port, 
      i_RD1_0_port, i_RD2_31_port, i_RD2_30_port, i_RD2_29_port, i_RD2_28_port,
      i_RD2_27_port, i_RD2_26_port, i_RD2_25_port, i_RD2_24_port, i_RD2_23_port
      , i_RD2_22_port, i_RD2_21_port, i_RD2_20_port, i_RD2_19_port, 
      i_RD2_18_port, i_RD2_17_port, i_RD2_16_port, i_RD2_15_port, i_RD2_14_port
      , i_RD2_13_port, i_RD2_12_port, i_RD2_11_port, i_RD2_10_port, 
      i_RD2_9_port, i_RD2_8_port, i_RD2_7_port, i_RD2_6_port, i_RD2_5_port, 
      i_RD2_4_port, i_RD2_3_port, i_RD2_2_port, i_RD2_1_port, i_RD2_0_port, 
      i_ADD_RS1_4_port, i_ADD_RS1_3_port, i_ADD_RS1_2_port, i_ADD_RS1_1_port, 
      i_ADD_RS1_0_port, i_ADD_RS2_4_port, i_ADD_RS2_3_port, i_ADD_RS2_2_port, 
      i_ADD_RS2_1_port, i_ADD_RS2_0_port, i_ADD_WS1_4_port, i_ADD_WS1_3_port, 
      i_ADD_WS1_2_port, i_ADD_WS1_1_port, i_ADD_WS1_0_port, CU_I_N318, 
      CU_I_N317, CU_I_N305, CU_I_N304, CU_I_i_FILL_delay, 
      CU_I_CW_MEM_WB_EN_port, CU_I_CW_MEM_WB_MUX_SEL_port, 
      CU_I_CW_MEM_MEM_EN_port, CU_I_CW_EX_WB_EN_port, 
      CU_I_CW_EX_WB_MUX_SEL_port, CU_I_CW_EX_MEM_EN_port, 
      CU_I_CW_EX_DATA_SIZE_0_port, CU_I_CW_EX_DATA_SIZE_1_port, 
      CU_I_CW_EX_DRAM_RE_port, CU_I_CW_EX_DRAM_WE_port, CU_I_CW_EX_EX_EN_port, 
      CU_I_CW_ID_WB_EN_port, CU_I_CW_ID_WB_MUX_SEL_port, CU_I_CW_ID_MEM_EN_port
      , CU_I_CW_ID_DATA_SIZE_0_port, CU_I_CW_ID_DATA_SIZE_1_port, 
      CU_I_CW_ID_DRAM_RE_port, CU_I_CW_ID_DRAM_WE_port, 
      CU_I_CW_ID_MUXB_SEL_port, CU_I_CW_ID_MUXA_SEL_port, CU_I_CW_ID_EX_EN_port
      , CU_I_CW_ID_ID_EN_port, CU_I_CW_ID_UNSIGNED_ID_port, 
      CU_I_CW_IF_WB_EN_port, CU_I_CW_IF_MEM_EN_port, CU_I_CW_WB_MUX_SEL_port, 
      CU_I_CW_DATA_SIZE_0_port, CU_I_CW_DATA_SIZE_1_port, CU_I_CW_MUXB_SEL_port
      , CU_I_CW_MUXA_SEL_port, CU_I_CW_NPC_SEL_port, CU_I_CW_UNSIGNED_ID_port, 
      CU_I_CW_SEL_CMPB_port, CU_I_CW_RF_RD2_EN_port, CU_I_CW_RF_RD1_EN_port, 
      DECODEhw_i_tickcounter_2_port, DECODEhw_i_tickcounter_4_port, 
      DECODEhw_i_tickcounter_6_port, DECODEhw_i_tickcounter_8_port, 
      DECODEhw_i_tickcounter_10_port, DECODEhw_i_tickcounter_12_port, 
      DECODEhw_i_tickcounter_14_port, DECODEhw_i_tickcounter_16_port, 
      DECODEhw_i_tickcounter_18_port, DECODEhw_i_tickcounter_20_port, 
      DECODEhw_i_tickcounter_22_port, DECODEhw_i_tickcounter_24_port, 
      DECODEhw_i_tickcounter_26_port, DECODEhw_i_tickcounter_29_port, 
      DECODEhw_i_tickcounter_31_port, DECODEhw_i_WR1, 
      DataPath_i_PIPLIN_WRB2_0_port, DataPath_i_PIPLIN_WRB2_1_port, 
      DataPath_i_PIPLIN_WRB2_2_port, DataPath_i_PIPLIN_WRB2_3_port, 
      DataPath_i_PIPLIN_WRB2_4_port, DataPath_i_PIPLIN_WRB1_0_port, 
      DataPath_i_PIPLIN_WRB1_1_port, DataPath_i_PIPLIN_WRB1_2_port, 
      DataPath_i_PIPLIN_WRB1_3_port, DataPath_i_PIPLIN_WRB1_4_port, 
      DataPath_i_REG_MEM_ALUOUT_0_port, DataPath_i_REG_MEM_ALUOUT_1_port, 
      DataPath_i_REG_MEM_ALUOUT_2_port, DataPath_i_REG_MEM_ALUOUT_3_port, 
      DataPath_i_REG_MEM_ALUOUT_4_port, DataPath_i_REG_MEM_ALUOUT_5_port, 
      DataPath_i_REG_MEM_ALUOUT_6_port, DataPath_i_REG_MEM_ALUOUT_7_port, 
      DataPath_i_REG_MEM_ALUOUT_8_port, DataPath_i_REG_MEM_ALUOUT_9_port, 
      DataPath_i_REG_MEM_ALUOUT_10_port, DataPath_i_REG_MEM_ALUOUT_11_port, 
      DataPath_i_REG_MEM_ALUOUT_12_port, DataPath_i_REG_MEM_ALUOUT_13_port, 
      DataPath_i_REG_MEM_ALUOUT_14_port, DataPath_i_REG_MEM_ALUOUT_15_port, 
      DataPath_i_REG_MEM_ALUOUT_16_port, DataPath_i_REG_MEM_ALUOUT_17_port, 
      DataPath_i_REG_MEM_ALUOUT_18_port, DataPath_i_REG_MEM_ALUOUT_19_port, 
      DataPath_i_REG_MEM_ALUOUT_20_port, DataPath_i_REG_MEM_ALUOUT_21_port, 
      DataPath_i_REG_MEM_ALUOUT_22_port, DataPath_i_REG_MEM_ALUOUT_23_port, 
      DataPath_i_REG_MEM_ALUOUT_24_port, DataPath_i_REG_MEM_ALUOUT_25_port, 
      DataPath_i_REG_MEM_ALUOUT_26_port, DataPath_i_REG_MEM_ALUOUT_27_port, 
      DataPath_i_REG_MEM_ALUOUT_28_port, DataPath_i_REG_MEM_ALUOUT_29_port, 
      DataPath_i_REG_MEM_ALUOUT_30_port, DataPath_i_REG_MEM_ALUOUT_31_port, 
      DataPath_i_REG_LDSTR_OUT_0_port, DataPath_i_REG_LDSTR_OUT_1_port, 
      DataPath_i_REG_LDSTR_OUT_2_port, DataPath_i_REG_LDSTR_OUT_3_port, 
      DataPath_i_REG_LDSTR_OUT_4_port, DataPath_i_REG_LDSTR_OUT_5_port, 
      DataPath_i_REG_LDSTR_OUT_6_port, DataPath_i_REG_LDSTR_OUT_7_port, 
      DataPath_i_REG_LDSTR_OUT_8_port, DataPath_i_REG_LDSTR_OUT_9_port, 
      DataPath_i_REG_LDSTR_OUT_10_port, DataPath_i_REG_LDSTR_OUT_11_port, 
      DataPath_i_REG_LDSTR_OUT_12_port, DataPath_i_REG_LDSTR_OUT_13_port, 
      DataPath_i_REG_LDSTR_OUT_14_port, DataPath_i_REG_LDSTR_OUT_15_port, 
      DataPath_i_REG_LDSTR_OUT_16_port, DataPath_i_REG_LDSTR_OUT_17_port, 
      DataPath_i_REG_LDSTR_OUT_18_port, DataPath_i_REG_LDSTR_OUT_19_port, 
      DataPath_i_REG_LDSTR_OUT_20_port, DataPath_i_REG_LDSTR_OUT_21_port, 
      DataPath_i_REG_LDSTR_OUT_22_port, DataPath_i_REG_LDSTR_OUT_23_port, 
      DataPath_i_REG_LDSTR_OUT_24_port, DataPath_i_REG_LDSTR_OUT_25_port, 
      DataPath_i_REG_LDSTR_OUT_26_port, DataPath_i_REG_LDSTR_OUT_27_port, 
      DataPath_i_REG_LDSTR_OUT_28_port, DataPath_i_REG_LDSTR_OUT_29_port, 
      DataPath_i_REG_LDSTR_OUT_30_port, DataPath_i_REG_LDSTR_OUT_31_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_0_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_1_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_2_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_3_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_4_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_5_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_6_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_7_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_8_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_9_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_10_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_11_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_12_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_13_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_14_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_15_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_16_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_17_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_18_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_19_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_20_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_21_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_22_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_23_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_24_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_25_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_26_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_27_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_28_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_29_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_30_port, 
      DataPath_i_REG_ME_DATA_DATAMEM_31_port, DataPath_i_PIPLIN_IN2_0_port, 
      DataPath_i_PIPLIN_IN2_1_port, DataPath_i_PIPLIN_IN2_2_port, 
      DataPath_i_PIPLIN_IN2_3_port, DataPath_i_PIPLIN_IN2_4_port, 
      DataPath_i_PIPLIN_IN2_5_port, DataPath_i_PIPLIN_IN2_7_port, 
      DataPath_i_PIPLIN_IN2_8_port, DataPath_i_PIPLIN_IN2_9_port, 
      DataPath_i_PIPLIN_IN2_10_port, DataPath_i_PIPLIN_IN2_11_port, 
      DataPath_i_PIPLIN_IN2_12_port, DataPath_i_PIPLIN_IN2_13_port, 
      DataPath_i_PIPLIN_IN2_14_port, DataPath_i_PIPLIN_IN2_15_port, 
      DataPath_i_PIPLIN_IN2_16_port, DataPath_i_PIPLIN_IN2_17_port, 
      DataPath_i_PIPLIN_IN2_18_port, DataPath_i_PIPLIN_IN2_19_port, 
      DataPath_i_PIPLIN_IN2_20_port, DataPath_i_PIPLIN_IN2_21_port, 
      DataPath_i_PIPLIN_IN2_22_port, DataPath_i_PIPLIN_IN2_23_port, 
      DataPath_i_PIPLIN_IN2_24_port, DataPath_i_PIPLIN_IN2_25_port, 
      DataPath_i_PIPLIN_IN2_26_port, DataPath_i_PIPLIN_IN2_27_port, 
      DataPath_i_PIPLIN_IN2_28_port, DataPath_i_PIPLIN_IN2_29_port, 
      DataPath_i_PIPLIN_IN2_30_port, DataPath_i_PIPLIN_IN2_31_port, 
      DataPath_i_PIPLIN_IN1_0_port, DataPath_i_PIPLIN_IN1_1_port, 
      DataPath_i_PIPLIN_IN1_2_port, DataPath_i_PIPLIN_IN1_3_port, 
      DataPath_i_PIPLIN_IN1_4_port, DataPath_i_PIPLIN_IN1_5_port, 
      DataPath_i_PIPLIN_IN1_6_port, DataPath_i_PIPLIN_IN1_7_port, 
      DataPath_i_PIPLIN_IN1_8_port, DataPath_i_PIPLIN_IN1_9_port, 
      DataPath_i_PIPLIN_IN1_10_port, DataPath_i_PIPLIN_IN1_11_port, 
      DataPath_i_PIPLIN_IN1_12_port, DataPath_i_PIPLIN_IN1_13_port, 
      DataPath_i_PIPLIN_IN1_14_port, DataPath_i_PIPLIN_IN1_15_port, 
      DataPath_i_PIPLIN_B_0_port, DataPath_i_PIPLIN_B_1_port, 
      DataPath_i_PIPLIN_B_2_port, DataPath_i_PIPLIN_B_3_port, 
      DataPath_i_PIPLIN_B_4_port, DataPath_i_PIPLIN_B_5_port, 
      DataPath_i_PIPLIN_B_7_port, DataPath_i_PIPLIN_B_8_port, 
      DataPath_i_PIPLIN_B_9_port, DataPath_i_PIPLIN_B_10_port, 
      DataPath_i_PIPLIN_B_11_port, DataPath_i_PIPLIN_B_12_port, 
      DataPath_i_PIPLIN_B_13_port, DataPath_i_PIPLIN_B_14_port, 
      DataPath_i_PIPLIN_B_15_port, DataPath_i_PIPLIN_B_16_port, 
      DataPath_i_PIPLIN_B_17_port, DataPath_i_PIPLIN_B_18_port, 
      DataPath_i_PIPLIN_B_19_port, DataPath_i_PIPLIN_B_20_port, 
      DataPath_i_PIPLIN_B_21_port, DataPath_i_PIPLIN_B_22_port, 
      DataPath_i_PIPLIN_B_23_port, DataPath_i_PIPLIN_B_24_port, 
      DataPath_i_PIPLIN_B_25_port, DataPath_i_PIPLIN_B_26_port, 
      DataPath_i_PIPLIN_B_27_port, DataPath_i_PIPLIN_B_28_port, 
      DataPath_i_PIPLIN_B_29_port, DataPath_i_PIPLIN_B_30_port, 
      DataPath_i_PIPLIN_B_31_port, DataPath_i_PIPLIN_A_0_port, 
      DataPath_i_PIPLIN_A_1_port, DataPath_i_PIPLIN_A_2_port, 
      DataPath_i_PIPLIN_A_3_port, DataPath_i_PIPLIN_A_4_port, 
      DataPath_i_PIPLIN_A_5_port, DataPath_i_PIPLIN_A_6_port, 
      DataPath_i_PIPLIN_A_7_port, DataPath_i_PIPLIN_A_8_port, 
      DataPath_i_PIPLIN_A_9_port, DataPath_i_PIPLIN_A_10_port, 
      DataPath_i_PIPLIN_A_11_port, DataPath_i_PIPLIN_A_12_port, 
      DataPath_i_PIPLIN_A_13_port, DataPath_i_PIPLIN_A_14_port, 
      DataPath_i_PIPLIN_A_15_port, DataPath_i_PIPLIN_A_16_port, 
      DataPath_i_PIPLIN_A_17_port, DataPath_i_PIPLIN_A_18_port, 
      DataPath_i_PIPLIN_A_19_port, DataPath_i_PIPLIN_A_20_port, 
      DataPath_i_PIPLIN_A_21_port, DataPath_i_PIPLIN_A_22_port, 
      DataPath_i_PIPLIN_A_23_port, DataPath_i_PIPLIN_A_24_port, 
      DataPath_i_PIPLIN_A_25_port, DataPath_i_PIPLIN_A_26_port, 
      DataPath_i_PIPLIN_A_27_port, DataPath_i_PIPLIN_A_28_port, 
      DataPath_i_PIPLIN_A_29_port, DataPath_i_PIPLIN_A_30_port, 
      DataPath_i_PIPLIN_A_31_port, DataPath_RF_bus_sel_savedwin_data_0_port, 
      DataPath_RF_bus_sel_savedwin_data_1_port, 
      DataPath_RF_bus_sel_savedwin_data_2_port, 
      DataPath_RF_bus_sel_savedwin_data_3_port, 
      DataPath_RF_bus_sel_savedwin_data_4_port, 
      DataPath_RF_bus_sel_savedwin_data_5_port, 
      DataPath_RF_bus_sel_savedwin_data_6_port, 
      DataPath_RF_bus_sel_savedwin_data_7_port, 
      DataPath_RF_bus_sel_savedwin_data_8_port, 
      DataPath_RF_bus_sel_savedwin_data_9_port, 
      DataPath_RF_bus_sel_savedwin_data_10_port, 
      DataPath_RF_bus_sel_savedwin_data_11_port, 
      DataPath_RF_bus_sel_savedwin_data_12_port, 
      DataPath_RF_bus_sel_savedwin_data_13_port, 
      DataPath_RF_bus_sel_savedwin_data_14_port, 
      DataPath_RF_bus_sel_savedwin_data_15_port, 
      DataPath_RF_bus_sel_savedwin_data_16_port, 
      DataPath_RF_bus_sel_savedwin_data_17_port, 
      DataPath_RF_bus_sel_savedwin_data_18_port, 
      DataPath_RF_bus_sel_savedwin_data_19_port, 
      DataPath_RF_bus_sel_savedwin_data_20_port, 
      DataPath_RF_bus_sel_savedwin_data_21_port, 
      DataPath_RF_bus_sel_savedwin_data_22_port, 
      DataPath_RF_bus_sel_savedwin_data_23_port, 
      DataPath_RF_bus_sel_savedwin_data_24_port, 
      DataPath_RF_bus_sel_savedwin_data_25_port, 
      DataPath_RF_bus_sel_savedwin_data_26_port, 
      DataPath_RF_bus_sel_savedwin_data_27_port, 
      DataPath_RF_bus_sel_savedwin_data_28_port, 
      DataPath_RF_bus_sel_savedwin_data_29_port, 
      DataPath_RF_bus_sel_savedwin_data_30_port, 
      DataPath_RF_bus_sel_savedwin_data_31_port, 
      DataPath_RF_bus_sel_savedwin_data_32_port, 
      DataPath_RF_bus_sel_savedwin_data_33_port, 
      DataPath_RF_bus_sel_savedwin_data_34_port, 
      DataPath_RF_bus_sel_savedwin_data_35_port, 
      DataPath_RF_bus_sel_savedwin_data_36_port, 
      DataPath_RF_bus_sel_savedwin_data_37_port, 
      DataPath_RF_bus_sel_savedwin_data_38_port, 
      DataPath_RF_bus_sel_savedwin_data_39_port, 
      DataPath_RF_bus_sel_savedwin_data_40_port, 
      DataPath_RF_bus_sel_savedwin_data_41_port, 
      DataPath_RF_bus_sel_savedwin_data_42_port, 
      DataPath_RF_bus_sel_savedwin_data_43_port, 
      DataPath_RF_bus_sel_savedwin_data_44_port, 
      DataPath_RF_bus_sel_savedwin_data_45_port, 
      DataPath_RF_bus_sel_savedwin_data_46_port, 
      DataPath_RF_bus_sel_savedwin_data_47_port, 
      DataPath_RF_bus_sel_savedwin_data_48_port, 
      DataPath_RF_bus_sel_savedwin_data_49_port, 
      DataPath_RF_bus_sel_savedwin_data_50_port, 
      DataPath_RF_bus_sel_savedwin_data_51_port, 
      DataPath_RF_bus_sel_savedwin_data_52_port, 
      DataPath_RF_bus_sel_savedwin_data_53_port, 
      DataPath_RF_bus_sel_savedwin_data_54_port, 
      DataPath_RF_bus_sel_savedwin_data_55_port, 
      DataPath_RF_bus_sel_savedwin_data_56_port, 
      DataPath_RF_bus_sel_savedwin_data_57_port, 
      DataPath_RF_bus_sel_savedwin_data_58_port, 
      DataPath_RF_bus_sel_savedwin_data_59_port, 
      DataPath_RF_bus_sel_savedwin_data_60_port, 
      DataPath_RF_bus_sel_savedwin_data_61_port, 
      DataPath_RF_bus_sel_savedwin_data_62_port, 
      DataPath_RF_bus_sel_savedwin_data_63_port, 
      DataPath_RF_bus_sel_savedwin_data_64_port, 
      DataPath_RF_bus_sel_savedwin_data_65_port, 
      DataPath_RF_bus_sel_savedwin_data_66_port, 
      DataPath_RF_bus_sel_savedwin_data_67_port, 
      DataPath_RF_bus_sel_savedwin_data_68_port, 
      DataPath_RF_bus_sel_savedwin_data_69_port, 
      DataPath_RF_bus_sel_savedwin_data_70_port, 
      DataPath_RF_bus_sel_savedwin_data_71_port, 
      DataPath_RF_bus_sel_savedwin_data_72_port, 
      DataPath_RF_bus_sel_savedwin_data_73_port, 
      DataPath_RF_bus_sel_savedwin_data_74_port, 
      DataPath_RF_bus_sel_savedwin_data_75_port, 
      DataPath_RF_bus_sel_savedwin_data_76_port, 
      DataPath_RF_bus_sel_savedwin_data_77_port, 
      DataPath_RF_bus_sel_savedwin_data_78_port, 
      DataPath_RF_bus_sel_savedwin_data_79_port, 
      DataPath_RF_bus_sel_savedwin_data_80_port, 
      DataPath_RF_bus_sel_savedwin_data_81_port, 
      DataPath_RF_bus_sel_savedwin_data_82_port, 
      DataPath_RF_bus_sel_savedwin_data_83_port, 
      DataPath_RF_bus_sel_savedwin_data_84_port, 
      DataPath_RF_bus_sel_savedwin_data_85_port, 
      DataPath_RF_bus_sel_savedwin_data_86_port, 
      DataPath_RF_bus_sel_savedwin_data_87_port, 
      DataPath_RF_bus_sel_savedwin_data_88_port, 
      DataPath_RF_bus_sel_savedwin_data_89_port, 
      DataPath_RF_bus_sel_savedwin_data_90_port, 
      DataPath_RF_bus_sel_savedwin_data_91_port, 
      DataPath_RF_bus_sel_savedwin_data_92_port, 
      DataPath_RF_bus_sel_savedwin_data_93_port, 
      DataPath_RF_bus_sel_savedwin_data_94_port, 
      DataPath_RF_bus_sel_savedwin_data_95_port, 
      DataPath_RF_bus_sel_savedwin_data_96_port, 
      DataPath_RF_bus_sel_savedwin_data_97_port, 
      DataPath_RF_bus_sel_savedwin_data_98_port, 
      DataPath_RF_bus_sel_savedwin_data_99_port, 
      DataPath_RF_bus_sel_savedwin_data_100_port, 
      DataPath_RF_bus_sel_savedwin_data_101_port, 
      DataPath_RF_bus_sel_savedwin_data_102_port, 
      DataPath_RF_bus_sel_savedwin_data_103_port, 
      DataPath_RF_bus_sel_savedwin_data_104_port, 
      DataPath_RF_bus_sel_savedwin_data_105_port, 
      DataPath_RF_bus_sel_savedwin_data_106_port, 
      DataPath_RF_bus_sel_savedwin_data_107_port, 
      DataPath_RF_bus_sel_savedwin_data_108_port, 
      DataPath_RF_bus_sel_savedwin_data_109_port, 
      DataPath_RF_bus_sel_savedwin_data_110_port, 
      DataPath_RF_bus_sel_savedwin_data_111_port, 
      DataPath_RF_bus_sel_savedwin_data_112_port, 
      DataPath_RF_bus_sel_savedwin_data_113_port, 
      DataPath_RF_bus_sel_savedwin_data_114_port, 
      DataPath_RF_bus_sel_savedwin_data_115_port, 
      DataPath_RF_bus_sel_savedwin_data_116_port, 
      DataPath_RF_bus_sel_savedwin_data_117_port, 
      DataPath_RF_bus_sel_savedwin_data_118_port, 
      DataPath_RF_bus_sel_savedwin_data_119_port, 
      DataPath_RF_bus_sel_savedwin_data_120_port, 
      DataPath_RF_bus_sel_savedwin_data_121_port, 
      DataPath_RF_bus_sel_savedwin_data_122_port, 
      DataPath_RF_bus_sel_savedwin_data_123_port, 
      DataPath_RF_bus_sel_savedwin_data_124_port, 
      DataPath_RF_bus_sel_savedwin_data_125_port, 
      DataPath_RF_bus_sel_savedwin_data_126_port, 
      DataPath_RF_bus_sel_savedwin_data_127_port, 
      DataPath_RF_bus_sel_savedwin_data_128_port, 
      DataPath_RF_bus_sel_savedwin_data_129_port, 
      DataPath_RF_bus_sel_savedwin_data_130_port, 
      DataPath_RF_bus_sel_savedwin_data_131_port, 
      DataPath_RF_bus_sel_savedwin_data_132_port, 
      DataPath_RF_bus_sel_savedwin_data_133_port, 
      DataPath_RF_bus_sel_savedwin_data_134_port, 
      DataPath_RF_bus_sel_savedwin_data_135_port, 
      DataPath_RF_bus_sel_savedwin_data_136_port, 
      DataPath_RF_bus_sel_savedwin_data_137_port, 
      DataPath_RF_bus_sel_savedwin_data_138_port, 
      DataPath_RF_bus_sel_savedwin_data_139_port, 
      DataPath_RF_bus_sel_savedwin_data_140_port, 
      DataPath_RF_bus_sel_savedwin_data_141_port, 
      DataPath_RF_bus_sel_savedwin_data_142_port, 
      DataPath_RF_bus_sel_savedwin_data_143_port, 
      DataPath_RF_bus_sel_savedwin_data_144_port, 
      DataPath_RF_bus_sel_savedwin_data_145_port, 
      DataPath_RF_bus_sel_savedwin_data_146_port, 
      DataPath_RF_bus_sel_savedwin_data_147_port, 
      DataPath_RF_bus_sel_savedwin_data_148_port, 
      DataPath_RF_bus_sel_savedwin_data_149_port, 
      DataPath_RF_bus_sel_savedwin_data_150_port, 
      DataPath_RF_bus_sel_savedwin_data_151_port, 
      DataPath_RF_bus_sel_savedwin_data_152_port, 
      DataPath_RF_bus_sel_savedwin_data_153_port, 
      DataPath_RF_bus_sel_savedwin_data_154_port, 
      DataPath_RF_bus_sel_savedwin_data_155_port, 
      DataPath_RF_bus_sel_savedwin_data_156_port, 
      DataPath_RF_bus_sel_savedwin_data_157_port, 
      DataPath_RF_bus_sel_savedwin_data_158_port, 
      DataPath_RF_bus_sel_savedwin_data_159_port, 
      DataPath_RF_bus_sel_savedwin_data_160_port, 
      DataPath_RF_bus_sel_savedwin_data_161_port, 
      DataPath_RF_bus_sel_savedwin_data_162_port, 
      DataPath_RF_bus_sel_savedwin_data_163_port, 
      DataPath_RF_bus_sel_savedwin_data_164_port, 
      DataPath_RF_bus_sel_savedwin_data_165_port, 
      DataPath_RF_bus_sel_savedwin_data_166_port, 
      DataPath_RF_bus_sel_savedwin_data_167_port, 
      DataPath_RF_bus_sel_savedwin_data_168_port, 
      DataPath_RF_bus_sel_savedwin_data_169_port, 
      DataPath_RF_bus_sel_savedwin_data_170_port, 
      DataPath_RF_bus_sel_savedwin_data_171_port, 
      DataPath_RF_bus_sel_savedwin_data_172_port, 
      DataPath_RF_bus_sel_savedwin_data_173_port, 
      DataPath_RF_bus_sel_savedwin_data_174_port, 
      DataPath_RF_bus_sel_savedwin_data_175_port, 
      DataPath_RF_bus_sel_savedwin_data_176_port, 
      DataPath_RF_bus_sel_savedwin_data_177_port, 
      DataPath_RF_bus_sel_savedwin_data_178_port, 
      DataPath_RF_bus_sel_savedwin_data_179_port, 
      DataPath_RF_bus_sel_savedwin_data_180_port, 
      DataPath_RF_bus_sel_savedwin_data_181_port, 
      DataPath_RF_bus_sel_savedwin_data_182_port, 
      DataPath_RF_bus_sel_savedwin_data_183_port, 
      DataPath_RF_bus_sel_savedwin_data_184_port, 
      DataPath_RF_bus_sel_savedwin_data_185_port, 
      DataPath_RF_bus_sel_savedwin_data_186_port, 
      DataPath_RF_bus_sel_savedwin_data_187_port, 
      DataPath_RF_bus_sel_savedwin_data_188_port, 
      DataPath_RF_bus_sel_savedwin_data_189_port, 
      DataPath_RF_bus_sel_savedwin_data_190_port, 
      DataPath_RF_bus_sel_savedwin_data_191_port, 
      DataPath_RF_bus_sel_savedwin_data_192_port, 
      DataPath_RF_bus_sel_savedwin_data_193_port, 
      DataPath_RF_bus_sel_savedwin_data_194_port, 
      DataPath_RF_bus_sel_savedwin_data_195_port, 
      DataPath_RF_bus_sel_savedwin_data_196_port, 
      DataPath_RF_bus_sel_savedwin_data_197_port, 
      DataPath_RF_bus_sel_savedwin_data_198_port, 
      DataPath_RF_bus_sel_savedwin_data_199_port, 
      DataPath_RF_bus_sel_savedwin_data_200_port, 
      DataPath_RF_bus_sel_savedwin_data_201_port, 
      DataPath_RF_bus_sel_savedwin_data_202_port, 
      DataPath_RF_bus_sel_savedwin_data_203_port, 
      DataPath_RF_bus_sel_savedwin_data_204_port, 
      DataPath_RF_bus_sel_savedwin_data_205_port, 
      DataPath_RF_bus_sel_savedwin_data_206_port, 
      DataPath_RF_bus_sel_savedwin_data_207_port, 
      DataPath_RF_bus_sel_savedwin_data_208_port, 
      DataPath_RF_bus_sel_savedwin_data_209_port, 
      DataPath_RF_bus_sel_savedwin_data_210_port, 
      DataPath_RF_bus_sel_savedwin_data_211_port, 
      DataPath_RF_bus_sel_savedwin_data_212_port, 
      DataPath_RF_bus_sel_savedwin_data_213_port, 
      DataPath_RF_bus_sel_savedwin_data_214_port, 
      DataPath_RF_bus_sel_savedwin_data_215_port, 
      DataPath_RF_bus_sel_savedwin_data_216_port, 
      DataPath_RF_bus_sel_savedwin_data_217_port, 
      DataPath_RF_bus_sel_savedwin_data_218_port, 
      DataPath_RF_bus_sel_savedwin_data_219_port, 
      DataPath_RF_bus_sel_savedwin_data_220_port, 
      DataPath_RF_bus_sel_savedwin_data_221_port, 
      DataPath_RF_bus_sel_savedwin_data_222_port, 
      DataPath_RF_bus_sel_savedwin_data_223_port, 
      DataPath_RF_bus_sel_savedwin_data_224_port, 
      DataPath_RF_bus_sel_savedwin_data_225_port, 
      DataPath_RF_bus_sel_savedwin_data_226_port, 
      DataPath_RF_bus_sel_savedwin_data_227_port, 
      DataPath_RF_bus_sel_savedwin_data_228_port, 
      DataPath_RF_bus_sel_savedwin_data_229_port, 
      DataPath_RF_bus_sel_savedwin_data_230_port, 
      DataPath_RF_bus_sel_savedwin_data_231_port, 
      DataPath_RF_bus_sel_savedwin_data_232_port, 
      DataPath_RF_bus_sel_savedwin_data_233_port, 
      DataPath_RF_bus_sel_savedwin_data_234_port, 
      DataPath_RF_bus_sel_savedwin_data_235_port, 
      DataPath_RF_bus_sel_savedwin_data_236_port, 
      DataPath_RF_bus_sel_savedwin_data_237_port, 
      DataPath_RF_bus_sel_savedwin_data_238_port, 
      DataPath_RF_bus_sel_savedwin_data_239_port, 
      DataPath_RF_bus_sel_savedwin_data_240_port, 
      DataPath_RF_bus_sel_savedwin_data_241_port, 
      DataPath_RF_bus_sel_savedwin_data_242_port, 
      DataPath_RF_bus_sel_savedwin_data_243_port, 
      DataPath_RF_bus_sel_savedwin_data_244_port, 
      DataPath_RF_bus_sel_savedwin_data_245_port, 
      DataPath_RF_bus_sel_savedwin_data_246_port, 
      DataPath_RF_bus_sel_savedwin_data_247_port, 
      DataPath_RF_bus_sel_savedwin_data_248_port, 
      DataPath_RF_bus_sel_savedwin_data_249_port, 
      DataPath_RF_bus_sel_savedwin_data_250_port, 
      DataPath_RF_bus_sel_savedwin_data_251_port, 
      DataPath_RF_bus_sel_savedwin_data_252_port, 
      DataPath_RF_bus_sel_savedwin_data_253_port, 
      DataPath_RF_bus_sel_savedwin_data_254_port, 
      DataPath_RF_bus_sel_savedwin_data_255_port, 
      DataPath_RF_bus_sel_savedwin_data_256_port, 
      DataPath_RF_bus_sel_savedwin_data_257_port, 
      DataPath_RF_bus_sel_savedwin_data_258_port, 
      DataPath_RF_bus_sel_savedwin_data_259_port, 
      DataPath_RF_bus_sel_savedwin_data_260_port, 
      DataPath_RF_bus_sel_savedwin_data_261_port, 
      DataPath_RF_bus_sel_savedwin_data_262_port, 
      DataPath_RF_bus_sel_savedwin_data_263_port, 
      DataPath_RF_bus_sel_savedwin_data_264_port, 
      DataPath_RF_bus_sel_savedwin_data_265_port, 
      DataPath_RF_bus_sel_savedwin_data_266_port, 
      DataPath_RF_bus_sel_savedwin_data_267_port, 
      DataPath_RF_bus_sel_savedwin_data_268_port, 
      DataPath_RF_bus_sel_savedwin_data_269_port, 
      DataPath_RF_bus_sel_savedwin_data_270_port, 
      DataPath_RF_bus_sel_savedwin_data_271_port, 
      DataPath_RF_bus_sel_savedwin_data_272_port, 
      DataPath_RF_bus_sel_savedwin_data_273_port, 
      DataPath_RF_bus_sel_savedwin_data_274_port, 
      DataPath_RF_bus_sel_savedwin_data_275_port, 
      DataPath_RF_bus_sel_savedwin_data_276_port, 
      DataPath_RF_bus_sel_savedwin_data_277_port, 
      DataPath_RF_bus_sel_savedwin_data_278_port, 
      DataPath_RF_bus_sel_savedwin_data_279_port, 
      DataPath_RF_bus_sel_savedwin_data_280_port, 
      DataPath_RF_bus_sel_savedwin_data_281_port, 
      DataPath_RF_bus_sel_savedwin_data_282_port, 
      DataPath_RF_bus_sel_savedwin_data_283_port, 
      DataPath_RF_bus_sel_savedwin_data_284_port, 
      DataPath_RF_bus_sel_savedwin_data_285_port, 
      DataPath_RF_bus_sel_savedwin_data_286_port, 
      DataPath_RF_bus_sel_savedwin_data_287_port, 
      DataPath_RF_bus_sel_savedwin_data_288_port, 
      DataPath_RF_bus_sel_savedwin_data_289_port, 
      DataPath_RF_bus_sel_savedwin_data_290_port, 
      DataPath_RF_bus_sel_savedwin_data_291_port, 
      DataPath_RF_bus_sel_savedwin_data_292_port, 
      DataPath_RF_bus_sel_savedwin_data_293_port, 
      DataPath_RF_bus_sel_savedwin_data_294_port, 
      DataPath_RF_bus_sel_savedwin_data_295_port, 
      DataPath_RF_bus_sel_savedwin_data_296_port, 
      DataPath_RF_bus_sel_savedwin_data_297_port, 
      DataPath_RF_bus_sel_savedwin_data_298_port, 
      DataPath_RF_bus_sel_savedwin_data_299_port, 
      DataPath_RF_bus_sel_savedwin_data_300_port, 
      DataPath_RF_bus_sel_savedwin_data_301_port, 
      DataPath_RF_bus_sel_savedwin_data_302_port, 
      DataPath_RF_bus_sel_savedwin_data_303_port, 
      DataPath_RF_bus_sel_savedwin_data_304_port, 
      DataPath_RF_bus_sel_savedwin_data_305_port, 
      DataPath_RF_bus_sel_savedwin_data_306_port, 
      DataPath_RF_bus_sel_savedwin_data_307_port, 
      DataPath_RF_bus_sel_savedwin_data_308_port, 
      DataPath_RF_bus_sel_savedwin_data_309_port, 
      DataPath_RF_bus_sel_savedwin_data_310_port, 
      DataPath_RF_bus_sel_savedwin_data_311_port, 
      DataPath_RF_bus_sel_savedwin_data_312_port, 
      DataPath_RF_bus_sel_savedwin_data_313_port, 
      DataPath_RF_bus_sel_savedwin_data_314_port, 
      DataPath_RF_bus_sel_savedwin_data_315_port, 
      DataPath_RF_bus_sel_savedwin_data_316_port, 
      DataPath_RF_bus_sel_savedwin_data_317_port, 
      DataPath_RF_bus_sel_savedwin_data_318_port, 
      DataPath_RF_bus_sel_savedwin_data_319_port, 
      DataPath_RF_bus_sel_savedwin_data_320_port, 
      DataPath_RF_bus_sel_savedwin_data_321_port, 
      DataPath_RF_bus_sel_savedwin_data_322_port, 
      DataPath_RF_bus_sel_savedwin_data_323_port, 
      DataPath_RF_bus_sel_savedwin_data_324_port, 
      DataPath_RF_bus_sel_savedwin_data_325_port, 
      DataPath_RF_bus_sel_savedwin_data_326_port, 
      DataPath_RF_bus_sel_savedwin_data_327_port, 
      DataPath_RF_bus_sel_savedwin_data_328_port, 
      DataPath_RF_bus_sel_savedwin_data_329_port, 
      DataPath_RF_bus_sel_savedwin_data_330_port, 
      DataPath_RF_bus_sel_savedwin_data_331_port, 
      DataPath_RF_bus_sel_savedwin_data_332_port, 
      DataPath_RF_bus_sel_savedwin_data_333_port, 
      DataPath_RF_bus_sel_savedwin_data_334_port, 
      DataPath_RF_bus_sel_savedwin_data_335_port, 
      DataPath_RF_bus_sel_savedwin_data_336_port, 
      DataPath_RF_bus_sel_savedwin_data_337_port, 
      DataPath_RF_bus_sel_savedwin_data_338_port, 
      DataPath_RF_bus_sel_savedwin_data_339_port, 
      DataPath_RF_bus_sel_savedwin_data_340_port, 
      DataPath_RF_bus_sel_savedwin_data_341_port, 
      DataPath_RF_bus_sel_savedwin_data_342_port, 
      DataPath_RF_bus_sel_savedwin_data_343_port, 
      DataPath_RF_bus_sel_savedwin_data_344_port, 
      DataPath_RF_bus_sel_savedwin_data_345_port, 
      DataPath_RF_bus_sel_savedwin_data_346_port, 
      DataPath_RF_bus_sel_savedwin_data_347_port, 
      DataPath_RF_bus_sel_savedwin_data_348_port, 
      DataPath_RF_bus_sel_savedwin_data_349_port, 
      DataPath_RF_bus_sel_savedwin_data_350_port, 
      DataPath_RF_bus_sel_savedwin_data_351_port, 
      DataPath_RF_bus_sel_savedwin_data_352_port, 
      DataPath_RF_bus_sel_savedwin_data_353_port, 
      DataPath_RF_bus_sel_savedwin_data_354_port, 
      DataPath_RF_bus_sel_savedwin_data_355_port, 
      DataPath_RF_bus_sel_savedwin_data_356_port, 
      DataPath_RF_bus_sel_savedwin_data_357_port, 
      DataPath_RF_bus_sel_savedwin_data_358_port, 
      DataPath_RF_bus_sel_savedwin_data_359_port, 
      DataPath_RF_bus_sel_savedwin_data_360_port, 
      DataPath_RF_bus_sel_savedwin_data_361_port, 
      DataPath_RF_bus_sel_savedwin_data_362_port, 
      DataPath_RF_bus_sel_savedwin_data_363_port, 
      DataPath_RF_bus_sel_savedwin_data_364_port, 
      DataPath_RF_bus_sel_savedwin_data_365_port, 
      DataPath_RF_bus_sel_savedwin_data_366_port, 
      DataPath_RF_bus_sel_savedwin_data_367_port, 
      DataPath_RF_bus_sel_savedwin_data_368_port, 
      DataPath_RF_bus_sel_savedwin_data_369_port, 
      DataPath_RF_bus_sel_savedwin_data_370_port, 
      DataPath_RF_bus_sel_savedwin_data_371_port, 
      DataPath_RF_bus_sel_savedwin_data_372_port, 
      DataPath_RF_bus_sel_savedwin_data_373_port, 
      DataPath_RF_bus_sel_savedwin_data_374_port, 
      DataPath_RF_bus_sel_savedwin_data_375_port, 
      DataPath_RF_bus_sel_savedwin_data_376_port, 
      DataPath_RF_bus_sel_savedwin_data_377_port, 
      DataPath_RF_bus_sel_savedwin_data_378_port, 
      DataPath_RF_bus_sel_savedwin_data_379_port, 
      DataPath_RF_bus_sel_savedwin_data_380_port, 
      DataPath_RF_bus_sel_savedwin_data_381_port, 
      DataPath_RF_bus_sel_savedwin_data_382_port, 
      DataPath_RF_bus_sel_savedwin_data_383_port, 
      DataPath_RF_bus_sel_savedwin_data_384_port, 
      DataPath_RF_bus_sel_savedwin_data_385_port, 
      DataPath_RF_bus_sel_savedwin_data_386_port, 
      DataPath_RF_bus_sel_savedwin_data_387_port, 
      DataPath_RF_bus_sel_savedwin_data_388_port, 
      DataPath_RF_bus_sel_savedwin_data_389_port, 
      DataPath_RF_bus_sel_savedwin_data_390_port, 
      DataPath_RF_bus_sel_savedwin_data_391_port, 
      DataPath_RF_bus_sel_savedwin_data_392_port, 
      DataPath_RF_bus_sel_savedwin_data_393_port, 
      DataPath_RF_bus_sel_savedwin_data_394_port, 
      DataPath_RF_bus_sel_savedwin_data_395_port, 
      DataPath_RF_bus_sel_savedwin_data_396_port, 
      DataPath_RF_bus_sel_savedwin_data_397_port, 
      DataPath_RF_bus_sel_savedwin_data_398_port, 
      DataPath_RF_bus_sel_savedwin_data_399_port, 
      DataPath_RF_bus_sel_savedwin_data_400_port, 
      DataPath_RF_bus_sel_savedwin_data_401_port, 
      DataPath_RF_bus_sel_savedwin_data_402_port, 
      DataPath_RF_bus_sel_savedwin_data_403_port, 
      DataPath_RF_bus_sel_savedwin_data_404_port, 
      DataPath_RF_bus_sel_savedwin_data_405_port, 
      DataPath_RF_bus_sel_savedwin_data_406_port, 
      DataPath_RF_bus_sel_savedwin_data_407_port, 
      DataPath_RF_bus_sel_savedwin_data_408_port, 
      DataPath_RF_bus_sel_savedwin_data_409_port, 
      DataPath_RF_bus_sel_savedwin_data_410_port, 
      DataPath_RF_bus_sel_savedwin_data_411_port, 
      DataPath_RF_bus_sel_savedwin_data_412_port, 
      DataPath_RF_bus_sel_savedwin_data_413_port, 
      DataPath_RF_bus_sel_savedwin_data_414_port, 
      DataPath_RF_bus_sel_savedwin_data_415_port, 
      DataPath_RF_bus_sel_savedwin_data_416_port, 
      DataPath_RF_bus_sel_savedwin_data_417_port, 
      DataPath_RF_bus_sel_savedwin_data_418_port, 
      DataPath_RF_bus_sel_savedwin_data_419_port, 
      DataPath_RF_bus_sel_savedwin_data_420_port, 
      DataPath_RF_bus_sel_savedwin_data_421_port, 
      DataPath_RF_bus_sel_savedwin_data_422_port, 
      DataPath_RF_bus_sel_savedwin_data_423_port, 
      DataPath_RF_bus_sel_savedwin_data_424_port, 
      DataPath_RF_bus_sel_savedwin_data_425_port, 
      DataPath_RF_bus_sel_savedwin_data_426_port, 
      DataPath_RF_bus_sel_savedwin_data_427_port, 
      DataPath_RF_bus_sel_savedwin_data_428_port, 
      DataPath_RF_bus_sel_savedwin_data_429_port, 
      DataPath_RF_bus_sel_savedwin_data_430_port, 
      DataPath_RF_bus_sel_savedwin_data_431_port, 
      DataPath_RF_bus_sel_savedwin_data_432_port, 
      DataPath_RF_bus_sel_savedwin_data_433_port, 
      DataPath_RF_bus_sel_savedwin_data_434_port, 
      DataPath_RF_bus_sel_savedwin_data_435_port, 
      DataPath_RF_bus_sel_savedwin_data_436_port, 
      DataPath_RF_bus_sel_savedwin_data_437_port, 
      DataPath_RF_bus_sel_savedwin_data_438_port, 
      DataPath_RF_bus_sel_savedwin_data_439_port, 
      DataPath_RF_bus_sel_savedwin_data_440_port, 
      DataPath_RF_bus_sel_savedwin_data_441_port, 
      DataPath_RF_bus_sel_savedwin_data_442_port, 
      DataPath_RF_bus_sel_savedwin_data_443_port, 
      DataPath_RF_bus_sel_savedwin_data_444_port, 
      DataPath_RF_bus_sel_savedwin_data_445_port, 
      DataPath_RF_bus_sel_savedwin_data_446_port, 
      DataPath_RF_bus_sel_savedwin_data_447_port, 
      DataPath_RF_bus_sel_savedwin_data_448_port, 
      DataPath_RF_bus_sel_savedwin_data_449_port, 
      DataPath_RF_bus_sel_savedwin_data_450_port, 
      DataPath_RF_bus_sel_savedwin_data_451_port, 
      DataPath_RF_bus_sel_savedwin_data_452_port, 
      DataPath_RF_bus_sel_savedwin_data_453_port, 
      DataPath_RF_bus_sel_savedwin_data_454_port, 
      DataPath_RF_bus_sel_savedwin_data_455_port, 
      DataPath_RF_bus_sel_savedwin_data_456_port, 
      DataPath_RF_bus_sel_savedwin_data_457_port, 
      DataPath_RF_bus_sel_savedwin_data_458_port, 
      DataPath_RF_bus_sel_savedwin_data_459_port, 
      DataPath_RF_bus_sel_savedwin_data_460_port, 
      DataPath_RF_bus_sel_savedwin_data_461_port, 
      DataPath_RF_bus_sel_savedwin_data_462_port, 
      DataPath_RF_bus_sel_savedwin_data_463_port, 
      DataPath_RF_bus_sel_savedwin_data_464_port, 
      DataPath_RF_bus_sel_savedwin_data_465_port, 
      DataPath_RF_bus_sel_savedwin_data_466_port, 
      DataPath_RF_bus_sel_savedwin_data_467_port, 
      DataPath_RF_bus_sel_savedwin_data_468_port, 
      DataPath_RF_bus_sel_savedwin_data_469_port, 
      DataPath_RF_bus_sel_savedwin_data_470_port, 
      DataPath_RF_bus_sel_savedwin_data_471_port, 
      DataPath_RF_bus_sel_savedwin_data_472_port, 
      DataPath_RF_bus_sel_savedwin_data_473_port, 
      DataPath_RF_bus_sel_savedwin_data_474_port, 
      DataPath_RF_bus_sel_savedwin_data_475_port, 
      DataPath_RF_bus_sel_savedwin_data_476_port, 
      DataPath_RF_bus_sel_savedwin_data_477_port, 
      DataPath_RF_bus_sel_savedwin_data_478_port, 
      DataPath_RF_bus_sel_savedwin_data_479_port, 
      DataPath_RF_bus_sel_savedwin_data_480_port, 
      DataPath_RF_bus_sel_savedwin_data_481_port, 
      DataPath_RF_bus_sel_savedwin_data_482_port, 
      DataPath_RF_bus_sel_savedwin_data_483_port, 
      DataPath_RF_bus_sel_savedwin_data_484_port, 
      DataPath_RF_bus_sel_savedwin_data_485_port, 
      DataPath_RF_bus_sel_savedwin_data_486_port, 
      DataPath_RF_bus_sel_savedwin_data_487_port, 
      DataPath_RF_bus_sel_savedwin_data_488_port, 
      DataPath_RF_bus_sel_savedwin_data_489_port, 
      DataPath_RF_bus_sel_savedwin_data_490_port, 
      DataPath_RF_bus_sel_savedwin_data_491_port, 
      DataPath_RF_bus_sel_savedwin_data_492_port, 
      DataPath_RF_bus_sel_savedwin_data_493_port, 
      DataPath_RF_bus_sel_savedwin_data_494_port, 
      DataPath_RF_bus_sel_savedwin_data_495_port, 
      DataPath_RF_bus_sel_savedwin_data_496_port, 
      DataPath_RF_bus_sel_savedwin_data_497_port, 
      DataPath_RF_bus_sel_savedwin_data_498_port, 
      DataPath_RF_bus_sel_savedwin_data_499_port, 
      DataPath_RF_bus_sel_savedwin_data_500_port, 
      DataPath_RF_bus_sel_savedwin_data_501_port, 
      DataPath_RF_bus_sel_savedwin_data_502_port, 
      DataPath_RF_bus_sel_savedwin_data_503_port, 
      DataPath_RF_bus_sel_savedwin_data_504_port, 
      DataPath_RF_bus_sel_savedwin_data_505_port, 
      DataPath_RF_bus_sel_savedwin_data_506_port, 
      DataPath_RF_bus_sel_savedwin_data_507_port, 
      DataPath_RF_bus_sel_savedwin_data_508_port, 
      DataPath_RF_bus_sel_savedwin_data_509_port, 
      DataPath_RF_bus_sel_savedwin_data_510_port, 
      DataPath_RF_bus_sel_savedwin_data_511_port, DataPath_RF_c_swin_0_port, 
      DataPath_RF_c_swin_1_port, DataPath_RF_c_swin_2_port, 
      DataPath_RF_c_swin_3_port, DataPath_RF_c_swin_4_port, 
      DataPath_RF_internal_out2_0_port, DataPath_RF_internal_out2_1_port, 
      DataPath_RF_internal_out2_2_port, DataPath_RF_internal_out2_3_port, 
      DataPath_RF_internal_out2_4_port, DataPath_RF_internal_out2_5_port, 
      DataPath_RF_internal_out2_6_port, DataPath_RF_internal_out2_7_port, 
      DataPath_RF_internal_out2_8_port, DataPath_RF_internal_out2_9_port, 
      DataPath_RF_internal_out2_10_port, DataPath_RF_internal_out2_11_port, 
      DataPath_RF_internal_out2_12_port, DataPath_RF_internal_out2_13_port, 
      DataPath_RF_internal_out2_14_port, DataPath_RF_internal_out2_15_port, 
      DataPath_RF_internal_out2_16_port, DataPath_RF_internal_out2_17_port, 
      DataPath_RF_internal_out2_18_port, DataPath_RF_internal_out2_19_port, 
      DataPath_RF_internal_out2_20_port, DataPath_RF_internal_out2_21_port, 
      DataPath_RF_internal_out2_22_port, DataPath_RF_internal_out2_23_port, 
      DataPath_RF_internal_out2_24_port, DataPath_RF_internal_out2_25_port, 
      DataPath_RF_internal_out2_26_port, DataPath_RF_internal_out2_27_port, 
      DataPath_RF_internal_out2_28_port, DataPath_RF_internal_out2_29_port, 
      DataPath_RF_internal_out2_30_port, DataPath_RF_internal_out2_31_port, 
      DataPath_RF_internal_out1_0_port, DataPath_RF_internal_out1_1_port, 
      DataPath_RF_internal_out1_2_port, DataPath_RF_internal_out1_3_port, 
      DataPath_RF_internal_out1_4_port, DataPath_RF_internal_out1_5_port, 
      DataPath_RF_internal_out1_6_port, DataPath_RF_internal_out1_7_port, 
      DataPath_RF_internal_out1_8_port, DataPath_RF_internal_out1_9_port, 
      DataPath_RF_internal_out1_10_port, DataPath_RF_internal_out1_11_port, 
      DataPath_RF_internal_out1_12_port, DataPath_RF_internal_out1_13_port, 
      DataPath_RF_internal_out1_14_port, DataPath_RF_internal_out1_15_port, 
      DataPath_RF_internal_out1_16_port, DataPath_RF_internal_out1_17_port, 
      DataPath_RF_internal_out1_18_port, DataPath_RF_internal_out1_19_port, 
      DataPath_RF_internal_out1_20_port, DataPath_RF_internal_out1_21_port, 
      DataPath_RF_internal_out1_22_port, DataPath_RF_internal_out1_23_port, 
      DataPath_RF_internal_out1_24_port, DataPath_RF_internal_out1_25_port, 
      DataPath_RF_internal_out1_26_port, DataPath_RF_internal_out1_27_port, 
      DataPath_RF_internal_out1_28_port, DataPath_RF_internal_out1_29_port, 
      DataPath_RF_internal_out1_30_port, DataPath_RF_internal_out1_31_port, 
      DataPath_RF_bus_complete_win_data_0_port, 
      DataPath_RF_bus_complete_win_data_32_port, 
      DataPath_RF_bus_complete_win_data_33_port, 
      DataPath_RF_bus_complete_win_data_34_port, 
      DataPath_RF_bus_complete_win_data_35_port, 
      DataPath_RF_bus_complete_win_data_36_port, 
      DataPath_RF_bus_complete_win_data_37_port, 
      DataPath_RF_bus_complete_win_data_38_port, 
      DataPath_RF_bus_complete_win_data_39_port, 
      DataPath_RF_bus_complete_win_data_40_port, 
      DataPath_RF_bus_complete_win_data_41_port, 
      DataPath_RF_bus_complete_win_data_42_port, 
      DataPath_RF_bus_complete_win_data_43_port, 
      DataPath_RF_bus_complete_win_data_44_port, 
      DataPath_RF_bus_complete_win_data_45_port, 
      DataPath_RF_bus_complete_win_data_46_port, 
      DataPath_RF_bus_complete_win_data_47_port, 
      DataPath_RF_bus_complete_win_data_48_port, 
      DataPath_RF_bus_complete_win_data_49_port, 
      DataPath_RF_bus_complete_win_data_50_port, 
      DataPath_RF_bus_complete_win_data_51_port, 
      DataPath_RF_bus_complete_win_data_52_port, 
      DataPath_RF_bus_complete_win_data_53_port, 
      DataPath_RF_bus_complete_win_data_54_port, 
      DataPath_RF_bus_complete_win_data_55_port, 
      DataPath_RF_bus_complete_win_data_56_port, 
      DataPath_RF_bus_complete_win_data_57_port, 
      DataPath_RF_bus_complete_win_data_58_port, 
      DataPath_RF_bus_complete_win_data_59_port, 
      DataPath_RF_bus_complete_win_data_60_port, 
      DataPath_RF_bus_complete_win_data_61_port, 
      DataPath_RF_bus_complete_win_data_62_port, 
      DataPath_RF_bus_complete_win_data_63_port, 
      DataPath_RF_bus_complete_win_data_64_port, 
      DataPath_RF_bus_complete_win_data_65_port, 
      DataPath_RF_bus_complete_win_data_66_port, 
      DataPath_RF_bus_complete_win_data_67_port, 
      DataPath_RF_bus_complete_win_data_68_port, 
      DataPath_RF_bus_complete_win_data_69_port, 
      DataPath_RF_bus_complete_win_data_70_port, 
      DataPath_RF_bus_complete_win_data_71_port, 
      DataPath_RF_bus_complete_win_data_72_port, 
      DataPath_RF_bus_complete_win_data_73_port, 
      DataPath_RF_bus_complete_win_data_74_port, 
      DataPath_RF_bus_complete_win_data_75_port, 
      DataPath_RF_bus_complete_win_data_76_port, 
      DataPath_RF_bus_complete_win_data_77_port, 
      DataPath_RF_bus_complete_win_data_78_port, 
      DataPath_RF_bus_complete_win_data_79_port, 
      DataPath_RF_bus_complete_win_data_80_port, 
      DataPath_RF_bus_complete_win_data_81_port, 
      DataPath_RF_bus_complete_win_data_82_port, 
      DataPath_RF_bus_complete_win_data_83_port, 
      DataPath_RF_bus_complete_win_data_84_port, 
      DataPath_RF_bus_complete_win_data_85_port, 
      DataPath_RF_bus_complete_win_data_86_port, 
      DataPath_RF_bus_complete_win_data_87_port, 
      DataPath_RF_bus_complete_win_data_88_port, 
      DataPath_RF_bus_complete_win_data_89_port, 
      DataPath_RF_bus_complete_win_data_90_port, 
      DataPath_RF_bus_complete_win_data_91_port, 
      DataPath_RF_bus_complete_win_data_92_port, 
      DataPath_RF_bus_complete_win_data_93_port, 
      DataPath_RF_bus_complete_win_data_94_port, 
      DataPath_RF_bus_complete_win_data_95_port, 
      DataPath_RF_bus_complete_win_data_96_port, 
      DataPath_RF_bus_complete_win_data_97_port, 
      DataPath_RF_bus_complete_win_data_98_port, 
      DataPath_RF_bus_complete_win_data_99_port, 
      DataPath_RF_bus_complete_win_data_100_port, 
      DataPath_RF_bus_complete_win_data_101_port, 
      DataPath_RF_bus_complete_win_data_102_port, 
      DataPath_RF_bus_complete_win_data_103_port, 
      DataPath_RF_bus_complete_win_data_104_port, 
      DataPath_RF_bus_complete_win_data_105_port, 
      DataPath_RF_bus_complete_win_data_106_port, 
      DataPath_RF_bus_complete_win_data_107_port, 
      DataPath_RF_bus_complete_win_data_108_port, 
      DataPath_RF_bus_complete_win_data_109_port, 
      DataPath_RF_bus_complete_win_data_110_port, 
      DataPath_RF_bus_complete_win_data_111_port, 
      DataPath_RF_bus_complete_win_data_112_port, 
      DataPath_RF_bus_complete_win_data_113_port, 
      DataPath_RF_bus_complete_win_data_114_port, 
      DataPath_RF_bus_complete_win_data_115_port, 
      DataPath_RF_bus_complete_win_data_116_port, 
      DataPath_RF_bus_complete_win_data_117_port, 
      DataPath_RF_bus_complete_win_data_118_port, 
      DataPath_RF_bus_complete_win_data_119_port, 
      DataPath_RF_bus_complete_win_data_120_port, 
      DataPath_RF_bus_complete_win_data_121_port, 
      DataPath_RF_bus_complete_win_data_122_port, 
      DataPath_RF_bus_complete_win_data_123_port, 
      DataPath_RF_bus_complete_win_data_124_port, 
      DataPath_RF_bus_complete_win_data_125_port, 
      DataPath_RF_bus_complete_win_data_126_port, 
      DataPath_RF_bus_complete_win_data_127_port, 
      DataPath_RF_bus_complete_win_data_128_port, 
      DataPath_RF_bus_complete_win_data_129_port, 
      DataPath_RF_bus_complete_win_data_130_port, 
      DataPath_RF_bus_complete_win_data_131_port, 
      DataPath_RF_bus_complete_win_data_132_port, 
      DataPath_RF_bus_complete_win_data_133_port, 
      DataPath_RF_bus_complete_win_data_134_port, 
      DataPath_RF_bus_complete_win_data_135_port, 
      DataPath_RF_bus_complete_win_data_136_port, 
      DataPath_RF_bus_complete_win_data_137_port, 
      DataPath_RF_bus_complete_win_data_138_port, 
      DataPath_RF_bus_complete_win_data_139_port, 
      DataPath_RF_bus_complete_win_data_140_port, 
      DataPath_RF_bus_complete_win_data_141_port, 
      DataPath_RF_bus_complete_win_data_142_port, 
      DataPath_RF_bus_complete_win_data_143_port, 
      DataPath_RF_bus_complete_win_data_144_port, 
      DataPath_RF_bus_complete_win_data_145_port, 
      DataPath_RF_bus_complete_win_data_146_port, 
      DataPath_RF_bus_complete_win_data_147_port, 
      DataPath_RF_bus_complete_win_data_148_port, 
      DataPath_RF_bus_complete_win_data_149_port, 
      DataPath_RF_bus_complete_win_data_150_port, 
      DataPath_RF_bus_complete_win_data_151_port, 
      DataPath_RF_bus_complete_win_data_152_port, 
      DataPath_RF_bus_complete_win_data_153_port, 
      DataPath_RF_bus_complete_win_data_154_port, 
      DataPath_RF_bus_complete_win_data_155_port, 
      DataPath_RF_bus_complete_win_data_156_port, 
      DataPath_RF_bus_complete_win_data_157_port, 
      DataPath_RF_bus_complete_win_data_158_port, 
      DataPath_RF_bus_complete_win_data_159_port, 
      DataPath_RF_bus_complete_win_data_160_port, 
      DataPath_RF_bus_complete_win_data_161_port, 
      DataPath_RF_bus_complete_win_data_162_port, 
      DataPath_RF_bus_complete_win_data_163_port, 
      DataPath_RF_bus_complete_win_data_164_port, 
      DataPath_RF_bus_complete_win_data_165_port, 
      DataPath_RF_bus_complete_win_data_166_port, 
      DataPath_RF_bus_complete_win_data_167_port, 
      DataPath_RF_bus_complete_win_data_168_port, 
      DataPath_RF_bus_complete_win_data_169_port, 
      DataPath_RF_bus_complete_win_data_170_port, 
      DataPath_RF_bus_complete_win_data_171_port, 
      DataPath_RF_bus_complete_win_data_172_port, 
      DataPath_RF_bus_complete_win_data_173_port, 
      DataPath_RF_bus_complete_win_data_174_port, 
      DataPath_RF_bus_complete_win_data_175_port, 
      DataPath_RF_bus_complete_win_data_176_port, 
      DataPath_RF_bus_complete_win_data_177_port, 
      DataPath_RF_bus_complete_win_data_178_port, 
      DataPath_RF_bus_complete_win_data_179_port, 
      DataPath_RF_bus_complete_win_data_180_port, 
      DataPath_RF_bus_complete_win_data_181_port, 
      DataPath_RF_bus_complete_win_data_182_port, 
      DataPath_RF_bus_complete_win_data_183_port, 
      DataPath_RF_bus_complete_win_data_184_port, 
      DataPath_RF_bus_complete_win_data_185_port, 
      DataPath_RF_bus_complete_win_data_186_port, 
      DataPath_RF_bus_complete_win_data_187_port, 
      DataPath_RF_bus_complete_win_data_188_port, 
      DataPath_RF_bus_complete_win_data_189_port, 
      DataPath_RF_bus_complete_win_data_190_port, 
      DataPath_RF_bus_complete_win_data_191_port, 
      DataPath_RF_bus_complete_win_data_192_port, 
      DataPath_RF_bus_complete_win_data_193_port, 
      DataPath_RF_bus_complete_win_data_194_port, 
      DataPath_RF_bus_complete_win_data_195_port, 
      DataPath_RF_bus_complete_win_data_196_port, 
      DataPath_RF_bus_complete_win_data_197_port, 
      DataPath_RF_bus_complete_win_data_198_port, 
      DataPath_RF_bus_complete_win_data_199_port, 
      DataPath_RF_bus_complete_win_data_200_port, 
      DataPath_RF_bus_complete_win_data_201_port, 
      DataPath_RF_bus_complete_win_data_202_port, 
      DataPath_RF_bus_complete_win_data_203_port, 
      DataPath_RF_bus_complete_win_data_204_port, 
      DataPath_RF_bus_complete_win_data_205_port, 
      DataPath_RF_bus_complete_win_data_206_port, 
      DataPath_RF_bus_complete_win_data_207_port, 
      DataPath_RF_bus_complete_win_data_208_port, 
      DataPath_RF_bus_complete_win_data_209_port, 
      DataPath_RF_bus_complete_win_data_210_port, 
      DataPath_RF_bus_complete_win_data_211_port, 
      DataPath_RF_bus_complete_win_data_212_port, 
      DataPath_RF_bus_complete_win_data_213_port, 
      DataPath_RF_bus_complete_win_data_214_port, 
      DataPath_RF_bus_complete_win_data_215_port, 
      DataPath_RF_bus_complete_win_data_216_port, 
      DataPath_RF_bus_complete_win_data_217_port, 
      DataPath_RF_bus_complete_win_data_218_port, 
      DataPath_RF_bus_complete_win_data_219_port, 
      DataPath_RF_bus_complete_win_data_220_port, 
      DataPath_RF_bus_complete_win_data_221_port, 
      DataPath_RF_bus_complete_win_data_222_port, 
      DataPath_RF_bus_complete_win_data_223_port, 
      DataPath_RF_bus_complete_win_data_224_port, 
      DataPath_RF_bus_complete_win_data_225_port, 
      DataPath_RF_bus_complete_win_data_226_port, 
      DataPath_RF_bus_complete_win_data_227_port, 
      DataPath_RF_bus_complete_win_data_228_port, 
      DataPath_RF_bus_complete_win_data_229_port, 
      DataPath_RF_bus_complete_win_data_230_port, 
      DataPath_RF_bus_complete_win_data_231_port, 
      DataPath_RF_bus_complete_win_data_232_port, 
      DataPath_RF_bus_complete_win_data_233_port, 
      DataPath_RF_bus_complete_win_data_234_port, 
      DataPath_RF_bus_complete_win_data_235_port, 
      DataPath_RF_bus_complete_win_data_236_port, 
      DataPath_RF_bus_complete_win_data_237_port, 
      DataPath_RF_bus_complete_win_data_238_port, 
      DataPath_RF_bus_complete_win_data_239_port, 
      DataPath_RF_bus_complete_win_data_240_port, 
      DataPath_RF_bus_complete_win_data_241_port, 
      DataPath_RF_bus_complete_win_data_242_port, 
      DataPath_RF_bus_complete_win_data_243_port, 
      DataPath_RF_bus_complete_win_data_244_port, 
      DataPath_RF_bus_complete_win_data_245_port, 
      DataPath_RF_bus_complete_win_data_246_port, 
      DataPath_RF_bus_complete_win_data_247_port, 
      DataPath_RF_bus_complete_win_data_248_port, 
      DataPath_RF_bus_complete_win_data_249_port, 
      DataPath_RF_bus_complete_win_data_250_port, 
      DataPath_RF_bus_complete_win_data_251_port, 
      DataPath_RF_bus_complete_win_data_252_port, 
      DataPath_RF_bus_complete_win_data_253_port, 
      DataPath_RF_bus_complete_win_data_254_port, 
      DataPath_RF_bus_complete_win_data_255_port, 
      DataPath_RF_bus_selected_win_data_0_port, 
      DataPath_RF_bus_selected_win_data_1_port, 
      DataPath_RF_bus_selected_win_data_2_port, 
      DataPath_RF_bus_selected_win_data_3_port, 
      DataPath_RF_bus_selected_win_data_4_port, 
      DataPath_RF_bus_selected_win_data_5_port, 
      DataPath_RF_bus_selected_win_data_6_port, 
      DataPath_RF_bus_selected_win_data_7_port, 
      DataPath_RF_bus_selected_win_data_8_port, 
      DataPath_RF_bus_selected_win_data_9_port, 
      DataPath_RF_bus_selected_win_data_10_port, 
      DataPath_RF_bus_selected_win_data_11_port, 
      DataPath_RF_bus_selected_win_data_12_port, 
      DataPath_RF_bus_selected_win_data_13_port, 
      DataPath_RF_bus_selected_win_data_14_port, 
      DataPath_RF_bus_selected_win_data_15_port, 
      DataPath_RF_bus_selected_win_data_16_port, 
      DataPath_RF_bus_selected_win_data_17_port, 
      DataPath_RF_bus_selected_win_data_18_port, 
      DataPath_RF_bus_selected_win_data_19_port, 
      DataPath_RF_bus_selected_win_data_20_port, 
      DataPath_RF_bus_selected_win_data_21_port, 
      DataPath_RF_bus_selected_win_data_22_port, 
      DataPath_RF_bus_selected_win_data_23_port, 
      DataPath_RF_bus_selected_win_data_24_port, 
      DataPath_RF_bus_selected_win_data_25_port, 
      DataPath_RF_bus_selected_win_data_26_port, 
      DataPath_RF_bus_selected_win_data_27_port, 
      DataPath_RF_bus_selected_win_data_28_port, 
      DataPath_RF_bus_selected_win_data_29_port, 
      DataPath_RF_bus_selected_win_data_30_port, 
      DataPath_RF_bus_selected_win_data_31_port, 
      DataPath_RF_bus_selected_win_data_32_port, 
      DataPath_RF_bus_selected_win_data_33_port, 
      DataPath_RF_bus_selected_win_data_34_port, 
      DataPath_RF_bus_selected_win_data_35_port, 
      DataPath_RF_bus_selected_win_data_36_port, 
      DataPath_RF_bus_selected_win_data_37_port, 
      DataPath_RF_bus_selected_win_data_38_port, 
      DataPath_RF_bus_selected_win_data_39_port, 
      DataPath_RF_bus_selected_win_data_40_port, 
      DataPath_RF_bus_selected_win_data_41_port, 
      DataPath_RF_bus_selected_win_data_42_port, 
      DataPath_RF_bus_selected_win_data_43_port, 
      DataPath_RF_bus_selected_win_data_44_port, 
      DataPath_RF_bus_selected_win_data_45_port, 
      DataPath_RF_bus_selected_win_data_46_port, 
      DataPath_RF_bus_selected_win_data_47_port, 
      DataPath_RF_bus_selected_win_data_48_port, 
      DataPath_RF_bus_selected_win_data_49_port, 
      DataPath_RF_bus_selected_win_data_50_port, 
      DataPath_RF_bus_selected_win_data_51_port, 
      DataPath_RF_bus_selected_win_data_52_port, 
      DataPath_RF_bus_selected_win_data_53_port, 
      DataPath_RF_bus_selected_win_data_54_port, 
      DataPath_RF_bus_selected_win_data_55_port, 
      DataPath_RF_bus_selected_win_data_56_port, 
      DataPath_RF_bus_selected_win_data_57_port, 
      DataPath_RF_bus_selected_win_data_58_port, 
      DataPath_RF_bus_selected_win_data_59_port, 
      DataPath_RF_bus_selected_win_data_60_port, 
      DataPath_RF_bus_selected_win_data_61_port, 
      DataPath_RF_bus_selected_win_data_62_port, 
      DataPath_RF_bus_selected_win_data_63_port, 
      DataPath_RF_bus_selected_win_data_64_port, 
      DataPath_RF_bus_selected_win_data_65_port, 
      DataPath_RF_bus_selected_win_data_66_port, 
      DataPath_RF_bus_selected_win_data_67_port, 
      DataPath_RF_bus_selected_win_data_68_port, 
      DataPath_RF_bus_selected_win_data_69_port, 
      DataPath_RF_bus_selected_win_data_70_port, 
      DataPath_RF_bus_selected_win_data_71_port, 
      DataPath_RF_bus_selected_win_data_72_port, 
      DataPath_RF_bus_selected_win_data_73_port, 
      DataPath_RF_bus_selected_win_data_74_port, 
      DataPath_RF_bus_selected_win_data_75_port, 
      DataPath_RF_bus_selected_win_data_76_port, 
      DataPath_RF_bus_selected_win_data_77_port, 
      DataPath_RF_bus_selected_win_data_78_port, 
      DataPath_RF_bus_selected_win_data_79_port, 
      DataPath_RF_bus_selected_win_data_80_port, 
      DataPath_RF_bus_selected_win_data_81_port, 
      DataPath_RF_bus_selected_win_data_82_port, 
      DataPath_RF_bus_selected_win_data_83_port, 
      DataPath_RF_bus_selected_win_data_84_port, 
      DataPath_RF_bus_selected_win_data_85_port, 
      DataPath_RF_bus_selected_win_data_86_port, 
      DataPath_RF_bus_selected_win_data_87_port, 
      DataPath_RF_bus_selected_win_data_88_port, 
      DataPath_RF_bus_selected_win_data_89_port, 
      DataPath_RF_bus_selected_win_data_90_port, 
      DataPath_RF_bus_selected_win_data_91_port, 
      DataPath_RF_bus_selected_win_data_92_port, 
      DataPath_RF_bus_selected_win_data_93_port, 
      DataPath_RF_bus_selected_win_data_94_port, 
      DataPath_RF_bus_selected_win_data_95_port, 
      DataPath_RF_bus_selected_win_data_96_port, 
      DataPath_RF_bus_selected_win_data_97_port, 
      DataPath_RF_bus_selected_win_data_98_port, 
      DataPath_RF_bus_selected_win_data_99_port, 
      DataPath_RF_bus_selected_win_data_100_port, 
      DataPath_RF_bus_selected_win_data_101_port, 
      DataPath_RF_bus_selected_win_data_102_port, 
      DataPath_RF_bus_selected_win_data_103_port, 
      DataPath_RF_bus_selected_win_data_104_port, 
      DataPath_RF_bus_selected_win_data_105_port, 
      DataPath_RF_bus_selected_win_data_106_port, 
      DataPath_RF_bus_selected_win_data_107_port, 
      DataPath_RF_bus_selected_win_data_108_port, 
      DataPath_RF_bus_selected_win_data_109_port, 
      DataPath_RF_bus_selected_win_data_110_port, 
      DataPath_RF_bus_selected_win_data_111_port, 
      DataPath_RF_bus_selected_win_data_112_port, 
      DataPath_RF_bus_selected_win_data_113_port, 
      DataPath_RF_bus_selected_win_data_114_port, 
      DataPath_RF_bus_selected_win_data_115_port, 
      DataPath_RF_bus_selected_win_data_116_port, 
      DataPath_RF_bus_selected_win_data_117_port, 
      DataPath_RF_bus_selected_win_data_118_port, 
      DataPath_RF_bus_selected_win_data_119_port, 
      DataPath_RF_bus_selected_win_data_120_port, 
      DataPath_RF_bus_selected_win_data_121_port, 
      DataPath_RF_bus_selected_win_data_122_port, 
      DataPath_RF_bus_selected_win_data_123_port, 
      DataPath_RF_bus_selected_win_data_124_port, 
      DataPath_RF_bus_selected_win_data_125_port, 
      DataPath_RF_bus_selected_win_data_126_port, 
      DataPath_RF_bus_selected_win_data_127_port, 
      DataPath_RF_bus_selected_win_data_128_port, 
      DataPath_RF_bus_selected_win_data_129_port, 
      DataPath_RF_bus_selected_win_data_130_port, 
      DataPath_RF_bus_selected_win_data_131_port, 
      DataPath_RF_bus_selected_win_data_132_port, 
      DataPath_RF_bus_selected_win_data_133_port, 
      DataPath_RF_bus_selected_win_data_134_port, 
      DataPath_RF_bus_selected_win_data_135_port, 
      DataPath_RF_bus_selected_win_data_136_port, 
      DataPath_RF_bus_selected_win_data_137_port, 
      DataPath_RF_bus_selected_win_data_138_port, 
      DataPath_RF_bus_selected_win_data_139_port, 
      DataPath_RF_bus_selected_win_data_140_port, 
      DataPath_RF_bus_selected_win_data_141_port, 
      DataPath_RF_bus_selected_win_data_142_port, 
      DataPath_RF_bus_selected_win_data_143_port, 
      DataPath_RF_bus_selected_win_data_144_port, 
      DataPath_RF_bus_selected_win_data_145_port, 
      DataPath_RF_bus_selected_win_data_146_port, 
      DataPath_RF_bus_selected_win_data_147_port, 
      DataPath_RF_bus_selected_win_data_148_port, 
      DataPath_RF_bus_selected_win_data_149_port, 
      DataPath_RF_bus_selected_win_data_150_port, 
      DataPath_RF_bus_selected_win_data_151_port, 
      DataPath_RF_bus_selected_win_data_152_port, 
      DataPath_RF_bus_selected_win_data_153_port, 
      DataPath_RF_bus_selected_win_data_154_port, 
      DataPath_RF_bus_selected_win_data_155_port, 
      DataPath_RF_bus_selected_win_data_156_port, 
      DataPath_RF_bus_selected_win_data_157_port, 
      DataPath_RF_bus_selected_win_data_158_port, 
      DataPath_RF_bus_selected_win_data_159_port, 
      DataPath_RF_bus_selected_win_data_160_port, 
      DataPath_RF_bus_selected_win_data_161_port, 
      DataPath_RF_bus_selected_win_data_162_port, 
      DataPath_RF_bus_selected_win_data_163_port, 
      DataPath_RF_bus_selected_win_data_164_port, 
      DataPath_RF_bus_selected_win_data_165_port, 
      DataPath_RF_bus_selected_win_data_166_port, 
      DataPath_RF_bus_selected_win_data_167_port, 
      DataPath_RF_bus_selected_win_data_168_port, 
      DataPath_RF_bus_selected_win_data_169_port, 
      DataPath_RF_bus_selected_win_data_170_port, 
      DataPath_RF_bus_selected_win_data_171_port, 
      DataPath_RF_bus_selected_win_data_172_port, 
      DataPath_RF_bus_selected_win_data_173_port, 
      DataPath_RF_bus_selected_win_data_174_port, 
      DataPath_RF_bus_selected_win_data_175_port, 
      DataPath_RF_bus_selected_win_data_176_port, 
      DataPath_RF_bus_selected_win_data_177_port, 
      DataPath_RF_bus_selected_win_data_178_port, 
      DataPath_RF_bus_selected_win_data_179_port, 
      DataPath_RF_bus_selected_win_data_180_port, 
      DataPath_RF_bus_selected_win_data_181_port, 
      DataPath_RF_bus_selected_win_data_182_port, 
      DataPath_RF_bus_selected_win_data_183_port, 
      DataPath_RF_bus_selected_win_data_184_port, 
      DataPath_RF_bus_selected_win_data_185_port, 
      DataPath_RF_bus_selected_win_data_186_port, 
      DataPath_RF_bus_selected_win_data_187_port, 
      DataPath_RF_bus_selected_win_data_188_port, 
      DataPath_RF_bus_selected_win_data_189_port, 
      DataPath_RF_bus_selected_win_data_190_port, 
      DataPath_RF_bus_selected_win_data_191_port, 
      DataPath_RF_bus_selected_win_data_192_port, 
      DataPath_RF_bus_selected_win_data_193_port, 
      DataPath_RF_bus_selected_win_data_194_port, 
      DataPath_RF_bus_selected_win_data_195_port, 
      DataPath_RF_bus_selected_win_data_196_port, 
      DataPath_RF_bus_selected_win_data_197_port, 
      DataPath_RF_bus_selected_win_data_198_port, 
      DataPath_RF_bus_selected_win_data_199_port, 
      DataPath_RF_bus_selected_win_data_200_port, 
      DataPath_RF_bus_selected_win_data_201_port, 
      DataPath_RF_bus_selected_win_data_202_port, 
      DataPath_RF_bus_selected_win_data_203_port, 
      DataPath_RF_bus_selected_win_data_204_port, 
      DataPath_RF_bus_selected_win_data_205_port, 
      DataPath_RF_bus_selected_win_data_206_port, 
      DataPath_RF_bus_selected_win_data_207_port, 
      DataPath_RF_bus_selected_win_data_208_port, 
      DataPath_RF_bus_selected_win_data_209_port, 
      DataPath_RF_bus_selected_win_data_210_port, 
      DataPath_RF_bus_selected_win_data_211_port, 
      DataPath_RF_bus_selected_win_data_212_port, 
      DataPath_RF_bus_selected_win_data_213_port, 
      DataPath_RF_bus_selected_win_data_214_port, 
      DataPath_RF_bus_selected_win_data_215_port, 
      DataPath_RF_bus_selected_win_data_216_port, 
      DataPath_RF_bus_selected_win_data_217_port, 
      DataPath_RF_bus_selected_win_data_218_port, 
      DataPath_RF_bus_selected_win_data_219_port, 
      DataPath_RF_bus_selected_win_data_220_port, 
      DataPath_RF_bus_selected_win_data_221_port, 
      DataPath_RF_bus_selected_win_data_222_port, 
      DataPath_RF_bus_selected_win_data_223_port, 
      DataPath_RF_bus_selected_win_data_224_port, 
      DataPath_RF_bus_selected_win_data_225_port, 
      DataPath_RF_bus_selected_win_data_226_port, 
      DataPath_RF_bus_selected_win_data_227_port, 
      DataPath_RF_bus_selected_win_data_228_port, 
      DataPath_RF_bus_selected_win_data_229_port, 
      DataPath_RF_bus_selected_win_data_230_port, 
      DataPath_RF_bus_selected_win_data_231_port, 
      DataPath_RF_bus_selected_win_data_232_port, 
      DataPath_RF_bus_selected_win_data_233_port, 
      DataPath_RF_bus_selected_win_data_234_port, 
      DataPath_RF_bus_selected_win_data_235_port, 
      DataPath_RF_bus_selected_win_data_236_port, 
      DataPath_RF_bus_selected_win_data_237_port, 
      DataPath_RF_bus_selected_win_data_238_port, 
      DataPath_RF_bus_selected_win_data_239_port, 
      DataPath_RF_bus_selected_win_data_240_port, 
      DataPath_RF_bus_selected_win_data_241_port, 
      DataPath_RF_bus_selected_win_data_242_port, 
      DataPath_RF_bus_selected_win_data_243_port, 
      DataPath_RF_bus_selected_win_data_244_port, 
      DataPath_RF_bus_selected_win_data_245_port, 
      DataPath_RF_bus_selected_win_data_246_port, 
      DataPath_RF_bus_selected_win_data_247_port, 
      DataPath_RF_bus_selected_win_data_248_port, 
      DataPath_RF_bus_selected_win_data_249_port, 
      DataPath_RF_bus_selected_win_data_250_port, 
      DataPath_RF_bus_selected_win_data_251_port, 
      DataPath_RF_bus_selected_win_data_252_port, 
      DataPath_RF_bus_selected_win_data_253_port, 
      DataPath_RF_bus_selected_win_data_254_port, 
      DataPath_RF_bus_selected_win_data_255_port, 
      DataPath_RF_bus_selected_win_data_256_port, 
      DataPath_RF_bus_selected_win_data_257_port, 
      DataPath_RF_bus_selected_win_data_258_port, 
      DataPath_RF_bus_selected_win_data_259_port, 
      DataPath_RF_bus_selected_win_data_260_port, 
      DataPath_RF_bus_selected_win_data_261_port, 
      DataPath_RF_bus_selected_win_data_262_port, 
      DataPath_RF_bus_selected_win_data_263_port, 
      DataPath_RF_bus_selected_win_data_264_port, 
      DataPath_RF_bus_selected_win_data_265_port, 
      DataPath_RF_bus_selected_win_data_266_port, 
      DataPath_RF_bus_selected_win_data_267_port, 
      DataPath_RF_bus_selected_win_data_268_port, 
      DataPath_RF_bus_selected_win_data_269_port, 
      DataPath_RF_bus_selected_win_data_270_port, 
      DataPath_RF_bus_selected_win_data_271_port, 
      DataPath_RF_bus_selected_win_data_272_port, 
      DataPath_RF_bus_selected_win_data_273_port, 
      DataPath_RF_bus_selected_win_data_274_port, 
      DataPath_RF_bus_selected_win_data_275_port, 
      DataPath_RF_bus_selected_win_data_276_port, 
      DataPath_RF_bus_selected_win_data_277_port, 
      DataPath_RF_bus_selected_win_data_278_port, 
      DataPath_RF_bus_selected_win_data_279_port, 
      DataPath_RF_bus_selected_win_data_280_port, 
      DataPath_RF_bus_selected_win_data_281_port, 
      DataPath_RF_bus_selected_win_data_282_port, 
      DataPath_RF_bus_selected_win_data_283_port, 
      DataPath_RF_bus_selected_win_data_284_port, 
      DataPath_RF_bus_selected_win_data_285_port, 
      DataPath_RF_bus_selected_win_data_286_port, 
      DataPath_RF_bus_selected_win_data_287_port, 
      DataPath_RF_bus_selected_win_data_288_port, 
      DataPath_RF_bus_selected_win_data_289_port, 
      DataPath_RF_bus_selected_win_data_290_port, 
      DataPath_RF_bus_selected_win_data_291_port, 
      DataPath_RF_bus_selected_win_data_292_port, 
      DataPath_RF_bus_selected_win_data_293_port, 
      DataPath_RF_bus_selected_win_data_294_port, 
      DataPath_RF_bus_selected_win_data_295_port, 
      DataPath_RF_bus_selected_win_data_296_port, 
      DataPath_RF_bus_selected_win_data_297_port, 
      DataPath_RF_bus_selected_win_data_298_port, 
      DataPath_RF_bus_selected_win_data_299_port, 
      DataPath_RF_bus_selected_win_data_300_port, 
      DataPath_RF_bus_selected_win_data_301_port, 
      DataPath_RF_bus_selected_win_data_302_port, 
      DataPath_RF_bus_selected_win_data_303_port, 
      DataPath_RF_bus_selected_win_data_304_port, 
      DataPath_RF_bus_selected_win_data_305_port, 
      DataPath_RF_bus_selected_win_data_306_port, 
      DataPath_RF_bus_selected_win_data_307_port, 
      DataPath_RF_bus_selected_win_data_308_port, 
      DataPath_RF_bus_selected_win_data_309_port, 
      DataPath_RF_bus_selected_win_data_310_port, 
      DataPath_RF_bus_selected_win_data_311_port, 
      DataPath_RF_bus_selected_win_data_312_port, 
      DataPath_RF_bus_selected_win_data_313_port, 
      DataPath_RF_bus_selected_win_data_314_port, 
      DataPath_RF_bus_selected_win_data_315_port, 
      DataPath_RF_bus_selected_win_data_316_port, 
      DataPath_RF_bus_selected_win_data_317_port, 
      DataPath_RF_bus_selected_win_data_318_port, 
      DataPath_RF_bus_selected_win_data_319_port, 
      DataPath_RF_bus_selected_win_data_320_port, 
      DataPath_RF_bus_selected_win_data_321_port, 
      DataPath_RF_bus_selected_win_data_322_port, 
      DataPath_RF_bus_selected_win_data_323_port, 
      DataPath_RF_bus_selected_win_data_324_port, 
      DataPath_RF_bus_selected_win_data_325_port, 
      DataPath_RF_bus_selected_win_data_326_port, 
      DataPath_RF_bus_selected_win_data_327_port, 
      DataPath_RF_bus_selected_win_data_328_port, 
      DataPath_RF_bus_selected_win_data_329_port, 
      DataPath_RF_bus_selected_win_data_330_port, 
      DataPath_RF_bus_selected_win_data_331_port, 
      DataPath_RF_bus_selected_win_data_332_port, 
      DataPath_RF_bus_selected_win_data_333_port, 
      DataPath_RF_bus_selected_win_data_334_port, 
      DataPath_RF_bus_selected_win_data_335_port, 
      DataPath_RF_bus_selected_win_data_336_port, 
      DataPath_RF_bus_selected_win_data_337_port, 
      DataPath_RF_bus_selected_win_data_338_port, 
      DataPath_RF_bus_selected_win_data_339_port, 
      DataPath_RF_bus_selected_win_data_340_port, 
      DataPath_RF_bus_selected_win_data_341_port, 
      DataPath_RF_bus_selected_win_data_342_port, 
      DataPath_RF_bus_selected_win_data_343_port, 
      DataPath_RF_bus_selected_win_data_344_port, 
      DataPath_RF_bus_selected_win_data_345_port, 
      DataPath_RF_bus_selected_win_data_346_port, 
      DataPath_RF_bus_selected_win_data_347_port, 
      DataPath_RF_bus_selected_win_data_348_port, 
      DataPath_RF_bus_selected_win_data_349_port, 
      DataPath_RF_bus_selected_win_data_350_port, 
      DataPath_RF_bus_selected_win_data_351_port, 
      DataPath_RF_bus_selected_win_data_352_port, 
      DataPath_RF_bus_selected_win_data_353_port, 
      DataPath_RF_bus_selected_win_data_354_port, 
      DataPath_RF_bus_selected_win_data_355_port, 
      DataPath_RF_bus_selected_win_data_356_port, 
      DataPath_RF_bus_selected_win_data_357_port, 
      DataPath_RF_bus_selected_win_data_358_port, 
      DataPath_RF_bus_selected_win_data_359_port, 
      DataPath_RF_bus_selected_win_data_360_port, 
      DataPath_RF_bus_selected_win_data_361_port, 
      DataPath_RF_bus_selected_win_data_362_port, 
      DataPath_RF_bus_selected_win_data_363_port, 
      DataPath_RF_bus_selected_win_data_364_port, 
      DataPath_RF_bus_selected_win_data_365_port, 
      DataPath_RF_bus_selected_win_data_366_port, 
      DataPath_RF_bus_selected_win_data_367_port, 
      DataPath_RF_bus_selected_win_data_368_port, 
      DataPath_RF_bus_selected_win_data_369_port, 
      DataPath_RF_bus_selected_win_data_370_port, 
      DataPath_RF_bus_selected_win_data_371_port, 
      DataPath_RF_bus_selected_win_data_372_port, 
      DataPath_RF_bus_selected_win_data_373_port, 
      DataPath_RF_bus_selected_win_data_374_port, 
      DataPath_RF_bus_selected_win_data_375_port, 
      DataPath_RF_bus_selected_win_data_376_port, 
      DataPath_RF_bus_selected_win_data_377_port, 
      DataPath_RF_bus_selected_win_data_378_port, 
      DataPath_RF_bus_selected_win_data_379_port, 
      DataPath_RF_bus_selected_win_data_380_port, 
      DataPath_RF_bus_selected_win_data_381_port, 
      DataPath_RF_bus_selected_win_data_382_port, 
      DataPath_RF_bus_selected_win_data_383_port, 
      DataPath_RF_bus_selected_win_data_384_port, 
      DataPath_RF_bus_selected_win_data_385_port, 
      DataPath_RF_bus_selected_win_data_386_port, 
      DataPath_RF_bus_selected_win_data_387_port, 
      DataPath_RF_bus_selected_win_data_388_port, 
      DataPath_RF_bus_selected_win_data_389_port, 
      DataPath_RF_bus_selected_win_data_390_port, 
      DataPath_RF_bus_selected_win_data_391_port, 
      DataPath_RF_bus_selected_win_data_392_port, 
      DataPath_RF_bus_selected_win_data_393_port, 
      DataPath_RF_bus_selected_win_data_394_port, 
      DataPath_RF_bus_selected_win_data_395_port, 
      DataPath_RF_bus_selected_win_data_396_port, 
      DataPath_RF_bus_selected_win_data_397_port, 
      DataPath_RF_bus_selected_win_data_398_port, 
      DataPath_RF_bus_selected_win_data_399_port, 
      DataPath_RF_bus_selected_win_data_400_port, 
      DataPath_RF_bus_selected_win_data_401_port, 
      DataPath_RF_bus_selected_win_data_402_port, 
      DataPath_RF_bus_selected_win_data_403_port, 
      DataPath_RF_bus_selected_win_data_404_port, 
      DataPath_RF_bus_selected_win_data_405_port, 
      DataPath_RF_bus_selected_win_data_406_port, 
      DataPath_RF_bus_selected_win_data_407_port, 
      DataPath_RF_bus_selected_win_data_408_port, 
      DataPath_RF_bus_selected_win_data_409_port, 
      DataPath_RF_bus_selected_win_data_410_port, 
      DataPath_RF_bus_selected_win_data_411_port, 
      DataPath_RF_bus_selected_win_data_412_port, 
      DataPath_RF_bus_selected_win_data_413_port, 
      DataPath_RF_bus_selected_win_data_414_port, 
      DataPath_RF_bus_selected_win_data_415_port, 
      DataPath_RF_bus_selected_win_data_416_port, 
      DataPath_RF_bus_selected_win_data_417_port, 
      DataPath_RF_bus_selected_win_data_418_port, 
      DataPath_RF_bus_selected_win_data_419_port, 
      DataPath_RF_bus_selected_win_data_420_port, 
      DataPath_RF_bus_selected_win_data_421_port, 
      DataPath_RF_bus_selected_win_data_422_port, 
      DataPath_RF_bus_selected_win_data_423_port, 
      DataPath_RF_bus_selected_win_data_424_port, 
      DataPath_RF_bus_selected_win_data_425_port, 
      DataPath_RF_bus_selected_win_data_426_port, 
      DataPath_RF_bus_selected_win_data_427_port, 
      DataPath_RF_bus_selected_win_data_428_port, 
      DataPath_RF_bus_selected_win_data_429_port, 
      DataPath_RF_bus_selected_win_data_430_port, 
      DataPath_RF_bus_selected_win_data_431_port, 
      DataPath_RF_bus_selected_win_data_432_port, 
      DataPath_RF_bus_selected_win_data_433_port, 
      DataPath_RF_bus_selected_win_data_434_port, 
      DataPath_RF_bus_selected_win_data_435_port, 
      DataPath_RF_bus_selected_win_data_436_port, 
      DataPath_RF_bus_selected_win_data_437_port, 
      DataPath_RF_bus_selected_win_data_438_port, 
      DataPath_RF_bus_selected_win_data_439_port, 
      DataPath_RF_bus_selected_win_data_440_port, 
      DataPath_RF_bus_selected_win_data_441_port, 
      DataPath_RF_bus_selected_win_data_442_port, 
      DataPath_RF_bus_selected_win_data_443_port, 
      DataPath_RF_bus_selected_win_data_444_port, 
      DataPath_RF_bus_selected_win_data_445_port, 
      DataPath_RF_bus_selected_win_data_446_port, 
      DataPath_RF_bus_selected_win_data_447_port, 
      DataPath_RF_bus_selected_win_data_448_port, 
      DataPath_RF_bus_selected_win_data_449_port, 
      DataPath_RF_bus_selected_win_data_450_port, 
      DataPath_RF_bus_selected_win_data_451_port, 
      DataPath_RF_bus_selected_win_data_452_port, 
      DataPath_RF_bus_selected_win_data_453_port, 
      DataPath_RF_bus_selected_win_data_454_port, 
      DataPath_RF_bus_selected_win_data_455_port, 
      DataPath_RF_bus_selected_win_data_456_port, 
      DataPath_RF_bus_selected_win_data_457_port, 
      DataPath_RF_bus_selected_win_data_458_port, 
      DataPath_RF_bus_selected_win_data_459_port, 
      DataPath_RF_bus_selected_win_data_460_port, 
      DataPath_RF_bus_selected_win_data_461_port, 
      DataPath_RF_bus_selected_win_data_462_port, 
      DataPath_RF_bus_selected_win_data_463_port, 
      DataPath_RF_bus_selected_win_data_464_port, 
      DataPath_RF_bus_selected_win_data_465_port, 
      DataPath_RF_bus_selected_win_data_466_port, 
      DataPath_RF_bus_selected_win_data_467_port, 
      DataPath_RF_bus_selected_win_data_468_port, 
      DataPath_RF_bus_selected_win_data_469_port, 
      DataPath_RF_bus_selected_win_data_470_port, 
      DataPath_RF_bus_selected_win_data_471_port, 
      DataPath_RF_bus_selected_win_data_472_port, 
      DataPath_RF_bus_selected_win_data_473_port, 
      DataPath_RF_bus_selected_win_data_474_port, 
      DataPath_RF_bus_selected_win_data_475_port, 
      DataPath_RF_bus_selected_win_data_476_port, 
      DataPath_RF_bus_selected_win_data_477_port, 
      DataPath_RF_bus_selected_win_data_478_port, 
      DataPath_RF_bus_selected_win_data_479_port, 
      DataPath_RF_bus_selected_win_data_480_port, 
      DataPath_RF_bus_selected_win_data_481_port, 
      DataPath_RF_bus_selected_win_data_482_port, 
      DataPath_RF_bus_selected_win_data_483_port, 
      DataPath_RF_bus_selected_win_data_484_port, 
      DataPath_RF_bus_selected_win_data_485_port, 
      DataPath_RF_bus_selected_win_data_486_port, 
      DataPath_RF_bus_selected_win_data_487_port, 
      DataPath_RF_bus_selected_win_data_488_port, 
      DataPath_RF_bus_selected_win_data_489_port, 
      DataPath_RF_bus_selected_win_data_490_port, 
      DataPath_RF_bus_selected_win_data_491_port, 
      DataPath_RF_bus_selected_win_data_492_port, 
      DataPath_RF_bus_selected_win_data_493_port, 
      DataPath_RF_bus_selected_win_data_494_port, 
      DataPath_RF_bus_selected_win_data_495_port, 
      DataPath_RF_bus_selected_win_data_496_port, 
      DataPath_RF_bus_selected_win_data_497_port, 
      DataPath_RF_bus_selected_win_data_498_port, 
      DataPath_RF_bus_selected_win_data_499_port, 
      DataPath_RF_bus_selected_win_data_500_port, 
      DataPath_RF_bus_selected_win_data_501_port, 
      DataPath_RF_bus_selected_win_data_502_port, 
      DataPath_RF_bus_selected_win_data_503_port, 
      DataPath_RF_bus_selected_win_data_504_port, 
      DataPath_RF_bus_selected_win_data_505_port, 
      DataPath_RF_bus_selected_win_data_506_port, 
      DataPath_RF_bus_selected_win_data_507_port, 
      DataPath_RF_bus_selected_win_data_508_port, 
      DataPath_RF_bus_selected_win_data_509_port, 
      DataPath_RF_bus_selected_win_data_510_port, 
      DataPath_RF_bus_selected_win_data_511_port, 
      DataPath_RF_bus_selected_win_data_512_port, 
      DataPath_RF_bus_selected_win_data_513_port, 
      DataPath_RF_bus_selected_win_data_514_port, 
      DataPath_RF_bus_selected_win_data_515_port, 
      DataPath_RF_bus_selected_win_data_516_port, 
      DataPath_RF_bus_selected_win_data_517_port, 
      DataPath_RF_bus_selected_win_data_518_port, 
      DataPath_RF_bus_selected_win_data_519_port, 
      DataPath_RF_bus_selected_win_data_520_port, 
      DataPath_RF_bus_selected_win_data_521_port, 
      DataPath_RF_bus_selected_win_data_522_port, 
      DataPath_RF_bus_selected_win_data_523_port, 
      DataPath_RF_bus_selected_win_data_524_port, 
      DataPath_RF_bus_selected_win_data_525_port, 
      DataPath_RF_bus_selected_win_data_526_port, 
      DataPath_RF_bus_selected_win_data_527_port, 
      DataPath_RF_bus_selected_win_data_528_port, 
      DataPath_RF_bus_selected_win_data_529_port, 
      DataPath_RF_bus_selected_win_data_530_port, 
      DataPath_RF_bus_selected_win_data_531_port, 
      DataPath_RF_bus_selected_win_data_532_port, 
      DataPath_RF_bus_selected_win_data_533_port, 
      DataPath_RF_bus_selected_win_data_534_port, 
      DataPath_RF_bus_selected_win_data_535_port, 
      DataPath_RF_bus_selected_win_data_536_port, 
      DataPath_RF_bus_selected_win_data_537_port, 
      DataPath_RF_bus_selected_win_data_538_port, 
      DataPath_RF_bus_selected_win_data_539_port, 
      DataPath_RF_bus_selected_win_data_540_port, 
      DataPath_RF_bus_selected_win_data_541_port, 
      DataPath_RF_bus_selected_win_data_542_port, 
      DataPath_RF_bus_selected_win_data_543_port, 
      DataPath_RF_bus_selected_win_data_544_port, 
      DataPath_RF_bus_selected_win_data_545_port, 
      DataPath_RF_bus_selected_win_data_546_port, 
      DataPath_RF_bus_selected_win_data_547_port, 
      DataPath_RF_bus_selected_win_data_548_port, 
      DataPath_RF_bus_selected_win_data_549_port, 
      DataPath_RF_bus_selected_win_data_550_port, 
      DataPath_RF_bus_selected_win_data_551_port, 
      DataPath_RF_bus_selected_win_data_552_port, 
      DataPath_RF_bus_selected_win_data_553_port, 
      DataPath_RF_bus_selected_win_data_554_port, 
      DataPath_RF_bus_selected_win_data_555_port, 
      DataPath_RF_bus_selected_win_data_556_port, 
      DataPath_RF_bus_selected_win_data_557_port, 
      DataPath_RF_bus_selected_win_data_558_port, 
      DataPath_RF_bus_selected_win_data_559_port, 
      DataPath_RF_bus_selected_win_data_560_port, 
      DataPath_RF_bus_selected_win_data_561_port, 
      DataPath_RF_bus_selected_win_data_562_port, 
      DataPath_RF_bus_selected_win_data_563_port, 
      DataPath_RF_bus_selected_win_data_564_port, 
      DataPath_RF_bus_selected_win_data_565_port, 
      DataPath_RF_bus_selected_win_data_566_port, 
      DataPath_RF_bus_selected_win_data_567_port, 
      DataPath_RF_bus_selected_win_data_568_port, 
      DataPath_RF_bus_selected_win_data_569_port, 
      DataPath_RF_bus_selected_win_data_570_port, 
      DataPath_RF_bus_selected_win_data_571_port, 
      DataPath_RF_bus_selected_win_data_572_port, 
      DataPath_RF_bus_selected_win_data_573_port, 
      DataPath_RF_bus_selected_win_data_574_port, 
      DataPath_RF_bus_selected_win_data_575_port, 
      DataPath_RF_bus_selected_win_data_576_port, 
      DataPath_RF_bus_selected_win_data_577_port, 
      DataPath_RF_bus_selected_win_data_578_port, 
      DataPath_RF_bus_selected_win_data_579_port, 
      DataPath_RF_bus_selected_win_data_580_port, 
      DataPath_RF_bus_selected_win_data_581_port, 
      DataPath_RF_bus_selected_win_data_582_port, 
      DataPath_RF_bus_selected_win_data_583_port, 
      DataPath_RF_bus_selected_win_data_584_port, 
      DataPath_RF_bus_selected_win_data_585_port, 
      DataPath_RF_bus_selected_win_data_586_port, 
      DataPath_RF_bus_selected_win_data_587_port, 
      DataPath_RF_bus_selected_win_data_588_port, 
      DataPath_RF_bus_selected_win_data_589_port, 
      DataPath_RF_bus_selected_win_data_590_port, 
      DataPath_RF_bus_selected_win_data_591_port, 
      DataPath_RF_bus_selected_win_data_592_port, 
      DataPath_RF_bus_selected_win_data_593_port, 
      DataPath_RF_bus_selected_win_data_594_port, 
      DataPath_RF_bus_selected_win_data_595_port, 
      DataPath_RF_bus_selected_win_data_596_port, 
      DataPath_RF_bus_selected_win_data_597_port, 
      DataPath_RF_bus_selected_win_data_598_port, 
      DataPath_RF_bus_selected_win_data_599_port, 
      DataPath_RF_bus_selected_win_data_600_port, 
      DataPath_RF_bus_selected_win_data_601_port, 
      DataPath_RF_bus_selected_win_data_602_port, 
      DataPath_RF_bus_selected_win_data_603_port, 
      DataPath_RF_bus_selected_win_data_604_port, 
      DataPath_RF_bus_selected_win_data_605_port, 
      DataPath_RF_bus_selected_win_data_606_port, 
      DataPath_RF_bus_selected_win_data_607_port, 
      DataPath_RF_bus_selected_win_data_608_port, 
      DataPath_RF_bus_selected_win_data_609_port, 
      DataPath_RF_bus_selected_win_data_610_port, 
      DataPath_RF_bus_selected_win_data_611_port, 
      DataPath_RF_bus_selected_win_data_612_port, 
      DataPath_RF_bus_selected_win_data_613_port, 
      DataPath_RF_bus_selected_win_data_614_port, 
      DataPath_RF_bus_selected_win_data_615_port, 
      DataPath_RF_bus_selected_win_data_616_port, 
      DataPath_RF_bus_selected_win_data_617_port, 
      DataPath_RF_bus_selected_win_data_618_port, 
      DataPath_RF_bus_selected_win_data_619_port, 
      DataPath_RF_bus_selected_win_data_620_port, 
      DataPath_RF_bus_selected_win_data_621_port, 
      DataPath_RF_bus_selected_win_data_622_port, 
      DataPath_RF_bus_selected_win_data_623_port, 
      DataPath_RF_bus_selected_win_data_624_port, 
      DataPath_RF_bus_selected_win_data_625_port, 
      DataPath_RF_bus_selected_win_data_626_port, 
      DataPath_RF_bus_selected_win_data_627_port, 
      DataPath_RF_bus_selected_win_data_628_port, 
      DataPath_RF_bus_selected_win_data_629_port, 
      DataPath_RF_bus_selected_win_data_630_port, 
      DataPath_RF_bus_selected_win_data_631_port, 
      DataPath_RF_bus_selected_win_data_632_port, 
      DataPath_RF_bus_selected_win_data_633_port, 
      DataPath_RF_bus_selected_win_data_634_port, 
      DataPath_RF_bus_selected_win_data_635_port, 
      DataPath_RF_bus_selected_win_data_636_port, 
      DataPath_RF_bus_selected_win_data_637_port, 
      DataPath_RF_bus_selected_win_data_638_port, 
      DataPath_RF_bus_selected_win_data_639_port, 
      DataPath_RF_bus_selected_win_data_640_port, 
      DataPath_RF_bus_selected_win_data_641_port, 
      DataPath_RF_bus_selected_win_data_642_port, 
      DataPath_RF_bus_selected_win_data_643_port, 
      DataPath_RF_bus_selected_win_data_644_port, 
      DataPath_RF_bus_selected_win_data_645_port, 
      DataPath_RF_bus_selected_win_data_646_port, 
      DataPath_RF_bus_selected_win_data_647_port, 
      DataPath_RF_bus_selected_win_data_648_port, 
      DataPath_RF_bus_selected_win_data_649_port, 
      DataPath_RF_bus_selected_win_data_650_port, 
      DataPath_RF_bus_selected_win_data_651_port, 
      DataPath_RF_bus_selected_win_data_652_port, 
      DataPath_RF_bus_selected_win_data_653_port, 
      DataPath_RF_bus_selected_win_data_654_port, 
      DataPath_RF_bus_selected_win_data_655_port, 
      DataPath_RF_bus_selected_win_data_656_port, 
      DataPath_RF_bus_selected_win_data_657_port, 
      DataPath_RF_bus_selected_win_data_658_port, 
      DataPath_RF_bus_selected_win_data_659_port, 
      DataPath_RF_bus_selected_win_data_660_port, 
      DataPath_RF_bus_selected_win_data_661_port, 
      DataPath_RF_bus_selected_win_data_662_port, 
      DataPath_RF_bus_selected_win_data_663_port, 
      DataPath_RF_bus_selected_win_data_664_port, 
      DataPath_RF_bus_selected_win_data_665_port, 
      DataPath_RF_bus_selected_win_data_666_port, 
      DataPath_RF_bus_selected_win_data_667_port, 
      DataPath_RF_bus_selected_win_data_668_port, 
      DataPath_RF_bus_selected_win_data_669_port, 
      DataPath_RF_bus_selected_win_data_670_port, 
      DataPath_RF_bus_selected_win_data_671_port, 
      DataPath_RF_bus_selected_win_data_672_port, 
      DataPath_RF_bus_selected_win_data_673_port, 
      DataPath_RF_bus_selected_win_data_674_port, 
      DataPath_RF_bus_selected_win_data_675_port, 
      DataPath_RF_bus_selected_win_data_676_port, 
      DataPath_RF_bus_selected_win_data_677_port, 
      DataPath_RF_bus_selected_win_data_678_port, 
      DataPath_RF_bus_selected_win_data_679_port, 
      DataPath_RF_bus_selected_win_data_680_port, 
      DataPath_RF_bus_selected_win_data_681_port, 
      DataPath_RF_bus_selected_win_data_682_port, 
      DataPath_RF_bus_selected_win_data_683_port, 
      DataPath_RF_bus_selected_win_data_684_port, 
      DataPath_RF_bus_selected_win_data_685_port, 
      DataPath_RF_bus_selected_win_data_686_port, 
      DataPath_RF_bus_selected_win_data_687_port, 
      DataPath_RF_bus_selected_win_data_688_port, 
      DataPath_RF_bus_selected_win_data_689_port, 
      DataPath_RF_bus_selected_win_data_690_port, 
      DataPath_RF_bus_selected_win_data_691_port, 
      DataPath_RF_bus_selected_win_data_692_port, 
      DataPath_RF_bus_selected_win_data_693_port, 
      DataPath_RF_bus_selected_win_data_694_port, 
      DataPath_RF_bus_selected_win_data_695_port, 
      DataPath_RF_bus_selected_win_data_696_port, 
      DataPath_RF_bus_selected_win_data_697_port, 
      DataPath_RF_bus_selected_win_data_698_port, 
      DataPath_RF_bus_selected_win_data_699_port, 
      DataPath_RF_bus_selected_win_data_700_port, 
      DataPath_RF_bus_selected_win_data_701_port, 
      DataPath_RF_bus_selected_win_data_702_port, 
      DataPath_RF_bus_selected_win_data_703_port, 
      DataPath_RF_bus_selected_win_data_704_port, 
      DataPath_RF_bus_selected_win_data_705_port, 
      DataPath_RF_bus_selected_win_data_706_port, 
      DataPath_RF_bus_selected_win_data_707_port, 
      DataPath_RF_bus_selected_win_data_708_port, 
      DataPath_RF_bus_selected_win_data_709_port, 
      DataPath_RF_bus_selected_win_data_710_port, 
      DataPath_RF_bus_selected_win_data_711_port, 
      DataPath_RF_bus_selected_win_data_712_port, 
      DataPath_RF_bus_selected_win_data_713_port, 
      DataPath_RF_bus_selected_win_data_714_port, 
      DataPath_RF_bus_selected_win_data_715_port, 
      DataPath_RF_bus_selected_win_data_716_port, 
      DataPath_RF_bus_selected_win_data_717_port, 
      DataPath_RF_bus_selected_win_data_718_port, 
      DataPath_RF_bus_selected_win_data_719_port, 
      DataPath_RF_bus_selected_win_data_720_port, 
      DataPath_RF_bus_selected_win_data_721_port, 
      DataPath_RF_bus_selected_win_data_722_port, 
      DataPath_RF_bus_selected_win_data_723_port, 
      DataPath_RF_bus_selected_win_data_724_port, 
      DataPath_RF_bus_selected_win_data_725_port, 
      DataPath_RF_bus_selected_win_data_726_port, 
      DataPath_RF_bus_selected_win_data_727_port, 
      DataPath_RF_bus_selected_win_data_728_port, 
      DataPath_RF_bus_selected_win_data_729_port, 
      DataPath_RF_bus_selected_win_data_730_port, 
      DataPath_RF_bus_selected_win_data_731_port, 
      DataPath_RF_bus_selected_win_data_732_port, 
      DataPath_RF_bus_selected_win_data_733_port, 
      DataPath_RF_bus_selected_win_data_734_port, 
      DataPath_RF_bus_selected_win_data_735_port, 
      DataPath_RF_bus_selected_win_data_736_port, 
      DataPath_RF_bus_selected_win_data_737_port, 
      DataPath_RF_bus_selected_win_data_738_port, 
      DataPath_RF_bus_selected_win_data_739_port, 
      DataPath_RF_bus_selected_win_data_740_port, 
      DataPath_RF_bus_selected_win_data_741_port, 
      DataPath_RF_bus_selected_win_data_742_port, 
      DataPath_RF_bus_selected_win_data_743_port, 
      DataPath_RF_bus_selected_win_data_744_port, 
      DataPath_RF_bus_selected_win_data_745_port, 
      DataPath_RF_bus_selected_win_data_746_port, 
      DataPath_RF_bus_selected_win_data_747_port, 
      DataPath_RF_bus_selected_win_data_748_port, 
      DataPath_RF_bus_selected_win_data_749_port, 
      DataPath_RF_bus_selected_win_data_750_port, 
      DataPath_RF_bus_selected_win_data_751_port, 
      DataPath_RF_bus_selected_win_data_752_port, 
      DataPath_RF_bus_selected_win_data_753_port, 
      DataPath_RF_bus_selected_win_data_754_port, 
      DataPath_RF_bus_selected_win_data_755_port, 
      DataPath_RF_bus_selected_win_data_756_port, 
      DataPath_RF_bus_selected_win_data_757_port, 
      DataPath_RF_bus_selected_win_data_758_port, 
      DataPath_RF_bus_selected_win_data_759_port, 
      DataPath_RF_bus_selected_win_data_760_port, 
      DataPath_RF_bus_selected_win_data_761_port, 
      DataPath_RF_bus_selected_win_data_762_port, 
      DataPath_RF_bus_selected_win_data_763_port, 
      DataPath_RF_bus_selected_win_data_764_port, 
      DataPath_RF_bus_selected_win_data_765_port, 
      DataPath_RF_bus_selected_win_data_766_port, 
      DataPath_RF_bus_selected_win_data_767_port, 
      DataPath_RF_bus_reg_dataout_0_port, DataPath_RF_bus_reg_dataout_1_port, 
      DataPath_RF_bus_reg_dataout_2_port, DataPath_RF_bus_reg_dataout_3_port, 
      DataPath_RF_bus_reg_dataout_4_port, DataPath_RF_bus_reg_dataout_5_port, 
      DataPath_RF_bus_reg_dataout_6_port, DataPath_RF_bus_reg_dataout_7_port, 
      DataPath_RF_bus_reg_dataout_8_port, DataPath_RF_bus_reg_dataout_9_port, 
      DataPath_RF_bus_reg_dataout_10_port, DataPath_RF_bus_reg_dataout_11_port,
      DataPath_RF_bus_reg_dataout_12_port, DataPath_RF_bus_reg_dataout_13_port,
      DataPath_RF_bus_reg_dataout_14_port, DataPath_RF_bus_reg_dataout_15_port,
      DataPath_RF_bus_reg_dataout_16_port, DataPath_RF_bus_reg_dataout_17_port,
      DataPath_RF_bus_reg_dataout_18_port, DataPath_RF_bus_reg_dataout_19_port,
      DataPath_RF_bus_reg_dataout_20_port, DataPath_RF_bus_reg_dataout_21_port,
      DataPath_RF_bus_reg_dataout_22_port, DataPath_RF_bus_reg_dataout_23_port,
      DataPath_RF_bus_reg_dataout_24_port, DataPath_RF_bus_reg_dataout_25_port,
      DataPath_RF_bus_reg_dataout_26_port, DataPath_RF_bus_reg_dataout_27_port,
      DataPath_RF_bus_reg_dataout_28_port, DataPath_RF_bus_reg_dataout_29_port,
      DataPath_RF_bus_reg_dataout_30_port, DataPath_RF_bus_reg_dataout_31_port,
      DataPath_RF_bus_reg_dataout_32_port, DataPath_RF_bus_reg_dataout_33_port,
      DataPath_RF_bus_reg_dataout_34_port, DataPath_RF_bus_reg_dataout_35_port,
      DataPath_RF_bus_reg_dataout_36_port, DataPath_RF_bus_reg_dataout_37_port,
      DataPath_RF_bus_reg_dataout_38_port, DataPath_RF_bus_reg_dataout_39_port,
      DataPath_RF_bus_reg_dataout_40_port, DataPath_RF_bus_reg_dataout_41_port,
      DataPath_RF_bus_reg_dataout_42_port, DataPath_RF_bus_reg_dataout_43_port,
      DataPath_RF_bus_reg_dataout_44_port, DataPath_RF_bus_reg_dataout_45_port,
      DataPath_RF_bus_reg_dataout_46_port, DataPath_RF_bus_reg_dataout_47_port,
      DataPath_RF_bus_reg_dataout_48_port, DataPath_RF_bus_reg_dataout_49_port,
      DataPath_RF_bus_reg_dataout_50_port, DataPath_RF_bus_reg_dataout_51_port,
      DataPath_RF_bus_reg_dataout_52_port, DataPath_RF_bus_reg_dataout_53_port,
      DataPath_RF_bus_reg_dataout_54_port, DataPath_RF_bus_reg_dataout_55_port,
      DataPath_RF_bus_reg_dataout_56_port, DataPath_RF_bus_reg_dataout_57_port,
      DataPath_RF_bus_reg_dataout_58_port, DataPath_RF_bus_reg_dataout_59_port,
      DataPath_RF_bus_reg_dataout_60_port, DataPath_RF_bus_reg_dataout_61_port,
      DataPath_RF_bus_reg_dataout_62_port, DataPath_RF_bus_reg_dataout_63_port,
      DataPath_RF_bus_reg_dataout_64_port, DataPath_RF_bus_reg_dataout_65_port,
      DataPath_RF_bus_reg_dataout_66_port, DataPath_RF_bus_reg_dataout_67_port,
      DataPath_RF_bus_reg_dataout_68_port, DataPath_RF_bus_reg_dataout_69_port,
      DataPath_RF_bus_reg_dataout_70_port, DataPath_RF_bus_reg_dataout_71_port,
      DataPath_RF_bus_reg_dataout_72_port, DataPath_RF_bus_reg_dataout_73_port,
      DataPath_RF_bus_reg_dataout_74_port, DataPath_RF_bus_reg_dataout_75_port,
      DataPath_RF_bus_reg_dataout_76_port, DataPath_RF_bus_reg_dataout_77_port,
      DataPath_RF_bus_reg_dataout_78_port, DataPath_RF_bus_reg_dataout_79_port,
      DataPath_RF_bus_reg_dataout_80_port, DataPath_RF_bus_reg_dataout_81_port,
      DataPath_RF_bus_reg_dataout_82_port, DataPath_RF_bus_reg_dataout_83_port,
      DataPath_RF_bus_reg_dataout_84_port, DataPath_RF_bus_reg_dataout_85_port,
      DataPath_RF_bus_reg_dataout_86_port, DataPath_RF_bus_reg_dataout_87_port,
      DataPath_RF_bus_reg_dataout_88_port, DataPath_RF_bus_reg_dataout_89_port,
      DataPath_RF_bus_reg_dataout_90_port, DataPath_RF_bus_reg_dataout_91_port,
      DataPath_RF_bus_reg_dataout_92_port, DataPath_RF_bus_reg_dataout_93_port,
      DataPath_RF_bus_reg_dataout_94_port, DataPath_RF_bus_reg_dataout_95_port,
      DataPath_RF_bus_reg_dataout_96_port, DataPath_RF_bus_reg_dataout_97_port,
      DataPath_RF_bus_reg_dataout_98_port, DataPath_RF_bus_reg_dataout_99_port,
      DataPath_RF_bus_reg_dataout_100_port, 
      DataPath_RF_bus_reg_dataout_101_port, 
      DataPath_RF_bus_reg_dataout_102_port, 
      DataPath_RF_bus_reg_dataout_103_port, 
      DataPath_RF_bus_reg_dataout_104_port, 
      DataPath_RF_bus_reg_dataout_105_port, 
      DataPath_RF_bus_reg_dataout_106_port, 
      DataPath_RF_bus_reg_dataout_107_port, 
      DataPath_RF_bus_reg_dataout_108_port, 
      DataPath_RF_bus_reg_dataout_109_port, 
      DataPath_RF_bus_reg_dataout_110_port, 
      DataPath_RF_bus_reg_dataout_111_port, 
      DataPath_RF_bus_reg_dataout_112_port, 
      DataPath_RF_bus_reg_dataout_113_port, 
      DataPath_RF_bus_reg_dataout_114_port, 
      DataPath_RF_bus_reg_dataout_115_port, 
      DataPath_RF_bus_reg_dataout_116_port, 
      DataPath_RF_bus_reg_dataout_117_port, 
      DataPath_RF_bus_reg_dataout_118_port, 
      DataPath_RF_bus_reg_dataout_119_port, 
      DataPath_RF_bus_reg_dataout_120_port, 
      DataPath_RF_bus_reg_dataout_121_port, 
      DataPath_RF_bus_reg_dataout_122_port, 
      DataPath_RF_bus_reg_dataout_123_port, 
      DataPath_RF_bus_reg_dataout_124_port, 
      DataPath_RF_bus_reg_dataout_125_port, 
      DataPath_RF_bus_reg_dataout_126_port, 
      DataPath_RF_bus_reg_dataout_127_port, 
      DataPath_RF_bus_reg_dataout_128_port, 
      DataPath_RF_bus_reg_dataout_129_port, 
      DataPath_RF_bus_reg_dataout_130_port, 
      DataPath_RF_bus_reg_dataout_131_port, 
      DataPath_RF_bus_reg_dataout_132_port, 
      DataPath_RF_bus_reg_dataout_133_port, 
      DataPath_RF_bus_reg_dataout_134_port, 
      DataPath_RF_bus_reg_dataout_135_port, 
      DataPath_RF_bus_reg_dataout_136_port, 
      DataPath_RF_bus_reg_dataout_137_port, 
      DataPath_RF_bus_reg_dataout_138_port, 
      DataPath_RF_bus_reg_dataout_139_port, 
      DataPath_RF_bus_reg_dataout_140_port, 
      DataPath_RF_bus_reg_dataout_141_port, 
      DataPath_RF_bus_reg_dataout_142_port, 
      DataPath_RF_bus_reg_dataout_143_port, 
      DataPath_RF_bus_reg_dataout_144_port, 
      DataPath_RF_bus_reg_dataout_145_port, 
      DataPath_RF_bus_reg_dataout_146_port, 
      DataPath_RF_bus_reg_dataout_147_port, 
      DataPath_RF_bus_reg_dataout_148_port, 
      DataPath_RF_bus_reg_dataout_149_port, 
      DataPath_RF_bus_reg_dataout_150_port, 
      DataPath_RF_bus_reg_dataout_151_port, 
      DataPath_RF_bus_reg_dataout_152_port, 
      DataPath_RF_bus_reg_dataout_153_port, 
      DataPath_RF_bus_reg_dataout_154_port, 
      DataPath_RF_bus_reg_dataout_155_port, 
      DataPath_RF_bus_reg_dataout_156_port, 
      DataPath_RF_bus_reg_dataout_157_port, 
      DataPath_RF_bus_reg_dataout_158_port, 
      DataPath_RF_bus_reg_dataout_159_port, 
      DataPath_RF_bus_reg_dataout_160_port, 
      DataPath_RF_bus_reg_dataout_161_port, 
      DataPath_RF_bus_reg_dataout_162_port, 
      DataPath_RF_bus_reg_dataout_163_port, 
      DataPath_RF_bus_reg_dataout_164_port, 
      DataPath_RF_bus_reg_dataout_165_port, 
      DataPath_RF_bus_reg_dataout_166_port, 
      DataPath_RF_bus_reg_dataout_167_port, 
      DataPath_RF_bus_reg_dataout_168_port, 
      DataPath_RF_bus_reg_dataout_169_port, 
      DataPath_RF_bus_reg_dataout_170_port, 
      DataPath_RF_bus_reg_dataout_171_port, 
      DataPath_RF_bus_reg_dataout_172_port, 
      DataPath_RF_bus_reg_dataout_173_port, 
      DataPath_RF_bus_reg_dataout_174_port, 
      DataPath_RF_bus_reg_dataout_175_port, 
      DataPath_RF_bus_reg_dataout_176_port, 
      DataPath_RF_bus_reg_dataout_177_port, 
      DataPath_RF_bus_reg_dataout_178_port, 
      DataPath_RF_bus_reg_dataout_179_port, 
      DataPath_RF_bus_reg_dataout_180_port, 
      DataPath_RF_bus_reg_dataout_181_port, 
      DataPath_RF_bus_reg_dataout_182_port, 
      DataPath_RF_bus_reg_dataout_183_port, 
      DataPath_RF_bus_reg_dataout_184_port, 
      DataPath_RF_bus_reg_dataout_185_port, 
      DataPath_RF_bus_reg_dataout_186_port, 
      DataPath_RF_bus_reg_dataout_187_port, 
      DataPath_RF_bus_reg_dataout_188_port, 
      DataPath_RF_bus_reg_dataout_189_port, 
      DataPath_RF_bus_reg_dataout_190_port, 
      DataPath_RF_bus_reg_dataout_191_port, 
      DataPath_RF_bus_reg_dataout_192_port, 
      DataPath_RF_bus_reg_dataout_193_port, 
      DataPath_RF_bus_reg_dataout_194_port, 
      DataPath_RF_bus_reg_dataout_195_port, 
      DataPath_RF_bus_reg_dataout_196_port, 
      DataPath_RF_bus_reg_dataout_197_port, 
      DataPath_RF_bus_reg_dataout_198_port, 
      DataPath_RF_bus_reg_dataout_199_port, 
      DataPath_RF_bus_reg_dataout_200_port, 
      DataPath_RF_bus_reg_dataout_201_port, 
      DataPath_RF_bus_reg_dataout_202_port, 
      DataPath_RF_bus_reg_dataout_203_port, 
      DataPath_RF_bus_reg_dataout_204_port, 
      DataPath_RF_bus_reg_dataout_205_port, 
      DataPath_RF_bus_reg_dataout_206_port, 
      DataPath_RF_bus_reg_dataout_207_port, 
      DataPath_RF_bus_reg_dataout_208_port, 
      DataPath_RF_bus_reg_dataout_209_port, 
      DataPath_RF_bus_reg_dataout_210_port, 
      DataPath_RF_bus_reg_dataout_211_port, 
      DataPath_RF_bus_reg_dataout_212_port, 
      DataPath_RF_bus_reg_dataout_213_port, 
      DataPath_RF_bus_reg_dataout_214_port, 
      DataPath_RF_bus_reg_dataout_215_port, 
      DataPath_RF_bus_reg_dataout_216_port, 
      DataPath_RF_bus_reg_dataout_217_port, 
      DataPath_RF_bus_reg_dataout_218_port, 
      DataPath_RF_bus_reg_dataout_219_port, 
      DataPath_RF_bus_reg_dataout_220_port, 
      DataPath_RF_bus_reg_dataout_221_port, 
      DataPath_RF_bus_reg_dataout_222_port, 
      DataPath_RF_bus_reg_dataout_223_port, 
      DataPath_RF_bus_reg_dataout_224_port, 
      DataPath_RF_bus_reg_dataout_225_port, 
      DataPath_RF_bus_reg_dataout_226_port, 
      DataPath_RF_bus_reg_dataout_227_port, 
      DataPath_RF_bus_reg_dataout_228_port, 
      DataPath_RF_bus_reg_dataout_229_port, 
      DataPath_RF_bus_reg_dataout_230_port, 
      DataPath_RF_bus_reg_dataout_231_port, 
      DataPath_RF_bus_reg_dataout_232_port, 
      DataPath_RF_bus_reg_dataout_233_port, 
      DataPath_RF_bus_reg_dataout_234_port, 
      DataPath_RF_bus_reg_dataout_235_port, 
      DataPath_RF_bus_reg_dataout_236_port, 
      DataPath_RF_bus_reg_dataout_237_port, 
      DataPath_RF_bus_reg_dataout_238_port, 
      DataPath_RF_bus_reg_dataout_239_port, 
      DataPath_RF_bus_reg_dataout_240_port, 
      DataPath_RF_bus_reg_dataout_241_port, 
      DataPath_RF_bus_reg_dataout_242_port, 
      DataPath_RF_bus_reg_dataout_243_port, 
      DataPath_RF_bus_reg_dataout_244_port, 
      DataPath_RF_bus_reg_dataout_245_port, 
      DataPath_RF_bus_reg_dataout_246_port, 
      DataPath_RF_bus_reg_dataout_247_port, 
      DataPath_RF_bus_reg_dataout_248_port, 
      DataPath_RF_bus_reg_dataout_249_port, 
      DataPath_RF_bus_reg_dataout_250_port, 
      DataPath_RF_bus_reg_dataout_251_port, 
      DataPath_RF_bus_reg_dataout_252_port, 
      DataPath_RF_bus_reg_dataout_253_port, 
      DataPath_RF_bus_reg_dataout_254_port, 
      DataPath_RF_bus_reg_dataout_255_port, 
      DataPath_RF_bus_reg_dataout_256_port, 
      DataPath_RF_bus_reg_dataout_257_port, 
      DataPath_RF_bus_reg_dataout_258_port, 
      DataPath_RF_bus_reg_dataout_259_port, 
      DataPath_RF_bus_reg_dataout_260_port, 
      DataPath_RF_bus_reg_dataout_261_port, 
      DataPath_RF_bus_reg_dataout_262_port, 
      DataPath_RF_bus_reg_dataout_263_port, 
      DataPath_RF_bus_reg_dataout_264_port, 
      DataPath_RF_bus_reg_dataout_265_port, 
      DataPath_RF_bus_reg_dataout_266_port, 
      DataPath_RF_bus_reg_dataout_267_port, 
      DataPath_RF_bus_reg_dataout_268_port, 
      DataPath_RF_bus_reg_dataout_269_port, 
      DataPath_RF_bus_reg_dataout_270_port, 
      DataPath_RF_bus_reg_dataout_271_port, 
      DataPath_RF_bus_reg_dataout_272_port, 
      DataPath_RF_bus_reg_dataout_273_port, 
      DataPath_RF_bus_reg_dataout_274_port, 
      DataPath_RF_bus_reg_dataout_275_port, 
      DataPath_RF_bus_reg_dataout_276_port, 
      DataPath_RF_bus_reg_dataout_277_port, 
      DataPath_RF_bus_reg_dataout_278_port, 
      DataPath_RF_bus_reg_dataout_279_port, 
      DataPath_RF_bus_reg_dataout_280_port, 
      DataPath_RF_bus_reg_dataout_281_port, 
      DataPath_RF_bus_reg_dataout_282_port, 
      DataPath_RF_bus_reg_dataout_283_port, 
      DataPath_RF_bus_reg_dataout_284_port, 
      DataPath_RF_bus_reg_dataout_285_port, 
      DataPath_RF_bus_reg_dataout_286_port, 
      DataPath_RF_bus_reg_dataout_287_port, 
      DataPath_RF_bus_reg_dataout_288_port, 
      DataPath_RF_bus_reg_dataout_289_port, 
      DataPath_RF_bus_reg_dataout_290_port, 
      DataPath_RF_bus_reg_dataout_291_port, 
      DataPath_RF_bus_reg_dataout_292_port, 
      DataPath_RF_bus_reg_dataout_293_port, 
      DataPath_RF_bus_reg_dataout_294_port, 
      DataPath_RF_bus_reg_dataout_295_port, 
      DataPath_RF_bus_reg_dataout_296_port, 
      DataPath_RF_bus_reg_dataout_297_port, 
      DataPath_RF_bus_reg_dataout_298_port, 
      DataPath_RF_bus_reg_dataout_299_port, 
      DataPath_RF_bus_reg_dataout_300_port, 
      DataPath_RF_bus_reg_dataout_301_port, 
      DataPath_RF_bus_reg_dataout_302_port, 
      DataPath_RF_bus_reg_dataout_303_port, 
      DataPath_RF_bus_reg_dataout_304_port, 
      DataPath_RF_bus_reg_dataout_305_port, 
      DataPath_RF_bus_reg_dataout_306_port, 
      DataPath_RF_bus_reg_dataout_307_port, 
      DataPath_RF_bus_reg_dataout_308_port, 
      DataPath_RF_bus_reg_dataout_309_port, 
      DataPath_RF_bus_reg_dataout_310_port, 
      DataPath_RF_bus_reg_dataout_311_port, 
      DataPath_RF_bus_reg_dataout_312_port, 
      DataPath_RF_bus_reg_dataout_313_port, 
      DataPath_RF_bus_reg_dataout_314_port, 
      DataPath_RF_bus_reg_dataout_315_port, 
      DataPath_RF_bus_reg_dataout_316_port, 
      DataPath_RF_bus_reg_dataout_317_port, 
      DataPath_RF_bus_reg_dataout_318_port, 
      DataPath_RF_bus_reg_dataout_319_port, 
      DataPath_RF_bus_reg_dataout_320_port, 
      DataPath_RF_bus_reg_dataout_321_port, 
      DataPath_RF_bus_reg_dataout_322_port, 
      DataPath_RF_bus_reg_dataout_323_port, 
      DataPath_RF_bus_reg_dataout_324_port, 
      DataPath_RF_bus_reg_dataout_325_port, 
      DataPath_RF_bus_reg_dataout_326_port, 
      DataPath_RF_bus_reg_dataout_327_port, 
      DataPath_RF_bus_reg_dataout_328_port, 
      DataPath_RF_bus_reg_dataout_329_port, 
      DataPath_RF_bus_reg_dataout_330_port, 
      DataPath_RF_bus_reg_dataout_331_port, 
      DataPath_RF_bus_reg_dataout_332_port, 
      DataPath_RF_bus_reg_dataout_333_port, 
      DataPath_RF_bus_reg_dataout_334_port, 
      DataPath_RF_bus_reg_dataout_335_port, 
      DataPath_RF_bus_reg_dataout_336_port, 
      DataPath_RF_bus_reg_dataout_337_port, 
      DataPath_RF_bus_reg_dataout_338_port, 
      DataPath_RF_bus_reg_dataout_339_port, 
      DataPath_RF_bus_reg_dataout_340_port, 
      DataPath_RF_bus_reg_dataout_341_port, 
      DataPath_RF_bus_reg_dataout_342_port, 
      DataPath_RF_bus_reg_dataout_343_port, 
      DataPath_RF_bus_reg_dataout_344_port, 
      DataPath_RF_bus_reg_dataout_345_port, 
      DataPath_RF_bus_reg_dataout_346_port, 
      DataPath_RF_bus_reg_dataout_347_port, 
      DataPath_RF_bus_reg_dataout_348_port, 
      DataPath_RF_bus_reg_dataout_349_port, 
      DataPath_RF_bus_reg_dataout_350_port, 
      DataPath_RF_bus_reg_dataout_351_port, 
      DataPath_RF_bus_reg_dataout_352_port, 
      DataPath_RF_bus_reg_dataout_353_port, 
      DataPath_RF_bus_reg_dataout_354_port, 
      DataPath_RF_bus_reg_dataout_355_port, 
      DataPath_RF_bus_reg_dataout_356_port, 
      DataPath_RF_bus_reg_dataout_357_port, 
      DataPath_RF_bus_reg_dataout_358_port, 
      DataPath_RF_bus_reg_dataout_359_port, 
      DataPath_RF_bus_reg_dataout_360_port, 
      DataPath_RF_bus_reg_dataout_361_port, 
      DataPath_RF_bus_reg_dataout_362_port, 
      DataPath_RF_bus_reg_dataout_363_port, 
      DataPath_RF_bus_reg_dataout_364_port, 
      DataPath_RF_bus_reg_dataout_365_port, 
      DataPath_RF_bus_reg_dataout_366_port, 
      DataPath_RF_bus_reg_dataout_367_port, 
      DataPath_RF_bus_reg_dataout_368_port, 
      DataPath_RF_bus_reg_dataout_369_port, 
      DataPath_RF_bus_reg_dataout_370_port, 
      DataPath_RF_bus_reg_dataout_371_port, 
      DataPath_RF_bus_reg_dataout_372_port, 
      DataPath_RF_bus_reg_dataout_373_port, 
      DataPath_RF_bus_reg_dataout_374_port, 
      DataPath_RF_bus_reg_dataout_375_port, 
      DataPath_RF_bus_reg_dataout_376_port, 
      DataPath_RF_bus_reg_dataout_377_port, 
      DataPath_RF_bus_reg_dataout_378_port, 
      DataPath_RF_bus_reg_dataout_379_port, 
      DataPath_RF_bus_reg_dataout_380_port, 
      DataPath_RF_bus_reg_dataout_381_port, 
      DataPath_RF_bus_reg_dataout_382_port, 
      DataPath_RF_bus_reg_dataout_383_port, 
      DataPath_RF_bus_reg_dataout_384_port, 
      DataPath_RF_bus_reg_dataout_385_port, 
      DataPath_RF_bus_reg_dataout_386_port, 
      DataPath_RF_bus_reg_dataout_387_port, 
      DataPath_RF_bus_reg_dataout_388_port, 
      DataPath_RF_bus_reg_dataout_389_port, 
      DataPath_RF_bus_reg_dataout_390_port, 
      DataPath_RF_bus_reg_dataout_391_port, 
      DataPath_RF_bus_reg_dataout_392_port, 
      DataPath_RF_bus_reg_dataout_393_port, 
      DataPath_RF_bus_reg_dataout_394_port, 
      DataPath_RF_bus_reg_dataout_395_port, 
      DataPath_RF_bus_reg_dataout_396_port, 
      DataPath_RF_bus_reg_dataout_397_port, 
      DataPath_RF_bus_reg_dataout_398_port, 
      DataPath_RF_bus_reg_dataout_399_port, 
      DataPath_RF_bus_reg_dataout_400_port, 
      DataPath_RF_bus_reg_dataout_401_port, 
      DataPath_RF_bus_reg_dataout_402_port, 
      DataPath_RF_bus_reg_dataout_403_port, 
      DataPath_RF_bus_reg_dataout_404_port, 
      DataPath_RF_bus_reg_dataout_405_port, 
      DataPath_RF_bus_reg_dataout_406_port, 
      DataPath_RF_bus_reg_dataout_407_port, 
      DataPath_RF_bus_reg_dataout_408_port, 
      DataPath_RF_bus_reg_dataout_409_port, 
      DataPath_RF_bus_reg_dataout_410_port, 
      DataPath_RF_bus_reg_dataout_411_port, 
      DataPath_RF_bus_reg_dataout_412_port, 
      DataPath_RF_bus_reg_dataout_413_port, 
      DataPath_RF_bus_reg_dataout_414_port, 
      DataPath_RF_bus_reg_dataout_415_port, 
      DataPath_RF_bus_reg_dataout_416_port, 
      DataPath_RF_bus_reg_dataout_417_port, 
      DataPath_RF_bus_reg_dataout_418_port, 
      DataPath_RF_bus_reg_dataout_419_port, 
      DataPath_RF_bus_reg_dataout_420_port, 
      DataPath_RF_bus_reg_dataout_421_port, 
      DataPath_RF_bus_reg_dataout_422_port, 
      DataPath_RF_bus_reg_dataout_423_port, 
      DataPath_RF_bus_reg_dataout_424_port, 
      DataPath_RF_bus_reg_dataout_425_port, 
      DataPath_RF_bus_reg_dataout_426_port, 
      DataPath_RF_bus_reg_dataout_427_port, 
      DataPath_RF_bus_reg_dataout_428_port, 
      DataPath_RF_bus_reg_dataout_429_port, 
      DataPath_RF_bus_reg_dataout_430_port, 
      DataPath_RF_bus_reg_dataout_431_port, 
      DataPath_RF_bus_reg_dataout_432_port, 
      DataPath_RF_bus_reg_dataout_433_port, 
      DataPath_RF_bus_reg_dataout_434_port, 
      DataPath_RF_bus_reg_dataout_435_port, 
      DataPath_RF_bus_reg_dataout_436_port, 
      DataPath_RF_bus_reg_dataout_437_port, 
      DataPath_RF_bus_reg_dataout_438_port, 
      DataPath_RF_bus_reg_dataout_439_port, 
      DataPath_RF_bus_reg_dataout_440_port, 
      DataPath_RF_bus_reg_dataout_441_port, 
      DataPath_RF_bus_reg_dataout_442_port, 
      DataPath_RF_bus_reg_dataout_443_port, 
      DataPath_RF_bus_reg_dataout_444_port, 
      DataPath_RF_bus_reg_dataout_445_port, 
      DataPath_RF_bus_reg_dataout_446_port, 
      DataPath_RF_bus_reg_dataout_447_port, 
      DataPath_RF_bus_reg_dataout_448_port, 
      DataPath_RF_bus_reg_dataout_449_port, 
      DataPath_RF_bus_reg_dataout_450_port, 
      DataPath_RF_bus_reg_dataout_451_port, 
      DataPath_RF_bus_reg_dataout_452_port, 
      DataPath_RF_bus_reg_dataout_453_port, 
      DataPath_RF_bus_reg_dataout_454_port, 
      DataPath_RF_bus_reg_dataout_455_port, 
      DataPath_RF_bus_reg_dataout_456_port, 
      DataPath_RF_bus_reg_dataout_457_port, 
      DataPath_RF_bus_reg_dataout_458_port, 
      DataPath_RF_bus_reg_dataout_459_port, 
      DataPath_RF_bus_reg_dataout_460_port, 
      DataPath_RF_bus_reg_dataout_461_port, 
      DataPath_RF_bus_reg_dataout_462_port, 
      DataPath_RF_bus_reg_dataout_463_port, 
      DataPath_RF_bus_reg_dataout_464_port, 
      DataPath_RF_bus_reg_dataout_465_port, 
      DataPath_RF_bus_reg_dataout_466_port, 
      DataPath_RF_bus_reg_dataout_467_port, 
      DataPath_RF_bus_reg_dataout_468_port, 
      DataPath_RF_bus_reg_dataout_469_port, 
      DataPath_RF_bus_reg_dataout_470_port, 
      DataPath_RF_bus_reg_dataout_471_port, 
      DataPath_RF_bus_reg_dataout_472_port, 
      DataPath_RF_bus_reg_dataout_473_port, 
      DataPath_RF_bus_reg_dataout_474_port, 
      DataPath_RF_bus_reg_dataout_475_port, 
      DataPath_RF_bus_reg_dataout_476_port, 
      DataPath_RF_bus_reg_dataout_477_port, 
      DataPath_RF_bus_reg_dataout_478_port, 
      DataPath_RF_bus_reg_dataout_479_port, 
      DataPath_RF_bus_reg_dataout_480_port, 
      DataPath_RF_bus_reg_dataout_481_port, 
      DataPath_RF_bus_reg_dataout_482_port, 
      DataPath_RF_bus_reg_dataout_483_port, 
      DataPath_RF_bus_reg_dataout_484_port, 
      DataPath_RF_bus_reg_dataout_485_port, 
      DataPath_RF_bus_reg_dataout_486_port, 
      DataPath_RF_bus_reg_dataout_487_port, 
      DataPath_RF_bus_reg_dataout_488_port, 
      DataPath_RF_bus_reg_dataout_489_port, 
      DataPath_RF_bus_reg_dataout_490_port, 
      DataPath_RF_bus_reg_dataout_491_port, 
      DataPath_RF_bus_reg_dataout_492_port, 
      DataPath_RF_bus_reg_dataout_493_port, 
      DataPath_RF_bus_reg_dataout_494_port, 
      DataPath_RF_bus_reg_dataout_495_port, 
      DataPath_RF_bus_reg_dataout_496_port, 
      DataPath_RF_bus_reg_dataout_497_port, 
      DataPath_RF_bus_reg_dataout_498_port, 
      DataPath_RF_bus_reg_dataout_499_port, 
      DataPath_RF_bus_reg_dataout_500_port, 
      DataPath_RF_bus_reg_dataout_501_port, 
      DataPath_RF_bus_reg_dataout_502_port, 
      DataPath_RF_bus_reg_dataout_503_port, 
      DataPath_RF_bus_reg_dataout_504_port, 
      DataPath_RF_bus_reg_dataout_505_port, 
      DataPath_RF_bus_reg_dataout_506_port, 
      DataPath_RF_bus_reg_dataout_507_port, 
      DataPath_RF_bus_reg_dataout_508_port, 
      DataPath_RF_bus_reg_dataout_509_port, 
      DataPath_RF_bus_reg_dataout_510_port, 
      DataPath_RF_bus_reg_dataout_511_port, 
      DataPath_RF_bus_reg_dataout_512_port, 
      DataPath_RF_bus_reg_dataout_513_port, 
      DataPath_RF_bus_reg_dataout_514_port, 
      DataPath_RF_bus_reg_dataout_515_port, 
      DataPath_RF_bus_reg_dataout_516_port, 
      DataPath_RF_bus_reg_dataout_517_port, 
      DataPath_RF_bus_reg_dataout_518_port, 
      DataPath_RF_bus_reg_dataout_519_port, 
      DataPath_RF_bus_reg_dataout_520_port, 
      DataPath_RF_bus_reg_dataout_521_port, 
      DataPath_RF_bus_reg_dataout_522_port, 
      DataPath_RF_bus_reg_dataout_523_port, 
      DataPath_RF_bus_reg_dataout_524_port, 
      DataPath_RF_bus_reg_dataout_525_port, 
      DataPath_RF_bus_reg_dataout_526_port, 
      DataPath_RF_bus_reg_dataout_527_port, 
      DataPath_RF_bus_reg_dataout_528_port, 
      DataPath_RF_bus_reg_dataout_529_port, 
      DataPath_RF_bus_reg_dataout_530_port, 
      DataPath_RF_bus_reg_dataout_531_port, 
      DataPath_RF_bus_reg_dataout_532_port, 
      DataPath_RF_bus_reg_dataout_533_port, 
      DataPath_RF_bus_reg_dataout_534_port, 
      DataPath_RF_bus_reg_dataout_535_port, 
      DataPath_RF_bus_reg_dataout_536_port, 
      DataPath_RF_bus_reg_dataout_537_port, 
      DataPath_RF_bus_reg_dataout_538_port, 
      DataPath_RF_bus_reg_dataout_539_port, 
      DataPath_RF_bus_reg_dataout_540_port, 
      DataPath_RF_bus_reg_dataout_541_port, 
      DataPath_RF_bus_reg_dataout_542_port, 
      DataPath_RF_bus_reg_dataout_543_port, 
      DataPath_RF_bus_reg_dataout_544_port, 
      DataPath_RF_bus_reg_dataout_545_port, 
      DataPath_RF_bus_reg_dataout_546_port, 
      DataPath_RF_bus_reg_dataout_547_port, 
      DataPath_RF_bus_reg_dataout_548_port, 
      DataPath_RF_bus_reg_dataout_549_port, 
      DataPath_RF_bus_reg_dataout_550_port, 
      DataPath_RF_bus_reg_dataout_551_port, 
      DataPath_RF_bus_reg_dataout_552_port, 
      DataPath_RF_bus_reg_dataout_553_port, 
      DataPath_RF_bus_reg_dataout_554_port, 
      DataPath_RF_bus_reg_dataout_555_port, 
      DataPath_RF_bus_reg_dataout_556_port, 
      DataPath_RF_bus_reg_dataout_557_port, 
      DataPath_RF_bus_reg_dataout_558_port, 
      DataPath_RF_bus_reg_dataout_559_port, 
      DataPath_RF_bus_reg_dataout_560_port, 
      DataPath_RF_bus_reg_dataout_561_port, 
      DataPath_RF_bus_reg_dataout_562_port, 
      DataPath_RF_bus_reg_dataout_563_port, 
      DataPath_RF_bus_reg_dataout_564_port, 
      DataPath_RF_bus_reg_dataout_565_port, 
      DataPath_RF_bus_reg_dataout_566_port, 
      DataPath_RF_bus_reg_dataout_567_port, 
      DataPath_RF_bus_reg_dataout_568_port, 
      DataPath_RF_bus_reg_dataout_569_port, 
      DataPath_RF_bus_reg_dataout_570_port, 
      DataPath_RF_bus_reg_dataout_571_port, 
      DataPath_RF_bus_reg_dataout_572_port, 
      DataPath_RF_bus_reg_dataout_573_port, 
      DataPath_RF_bus_reg_dataout_574_port, 
      DataPath_RF_bus_reg_dataout_575_port, 
      DataPath_RF_bus_reg_dataout_576_port, 
      DataPath_RF_bus_reg_dataout_577_port, 
      DataPath_RF_bus_reg_dataout_578_port, 
      DataPath_RF_bus_reg_dataout_579_port, 
      DataPath_RF_bus_reg_dataout_580_port, 
      DataPath_RF_bus_reg_dataout_581_port, 
      DataPath_RF_bus_reg_dataout_582_port, 
      DataPath_RF_bus_reg_dataout_583_port, 
      DataPath_RF_bus_reg_dataout_584_port, 
      DataPath_RF_bus_reg_dataout_585_port, 
      DataPath_RF_bus_reg_dataout_586_port, 
      DataPath_RF_bus_reg_dataout_587_port, 
      DataPath_RF_bus_reg_dataout_588_port, 
      DataPath_RF_bus_reg_dataout_589_port, 
      DataPath_RF_bus_reg_dataout_590_port, 
      DataPath_RF_bus_reg_dataout_591_port, 
      DataPath_RF_bus_reg_dataout_592_port, 
      DataPath_RF_bus_reg_dataout_593_port, 
      DataPath_RF_bus_reg_dataout_594_port, 
      DataPath_RF_bus_reg_dataout_595_port, 
      DataPath_RF_bus_reg_dataout_596_port, 
      DataPath_RF_bus_reg_dataout_597_port, 
      DataPath_RF_bus_reg_dataout_598_port, 
      DataPath_RF_bus_reg_dataout_599_port, 
      DataPath_RF_bus_reg_dataout_600_port, 
      DataPath_RF_bus_reg_dataout_601_port, 
      DataPath_RF_bus_reg_dataout_602_port, 
      DataPath_RF_bus_reg_dataout_603_port, 
      DataPath_RF_bus_reg_dataout_604_port, 
      DataPath_RF_bus_reg_dataout_605_port, 
      DataPath_RF_bus_reg_dataout_606_port, 
      DataPath_RF_bus_reg_dataout_607_port, 
      DataPath_RF_bus_reg_dataout_608_port, 
      DataPath_RF_bus_reg_dataout_609_port, 
      DataPath_RF_bus_reg_dataout_610_port, 
      DataPath_RF_bus_reg_dataout_611_port, 
      DataPath_RF_bus_reg_dataout_612_port, 
      DataPath_RF_bus_reg_dataout_613_port, 
      DataPath_RF_bus_reg_dataout_614_port, 
      DataPath_RF_bus_reg_dataout_615_port, 
      DataPath_RF_bus_reg_dataout_616_port, 
      DataPath_RF_bus_reg_dataout_617_port, 
      DataPath_RF_bus_reg_dataout_618_port, 
      DataPath_RF_bus_reg_dataout_619_port, 
      DataPath_RF_bus_reg_dataout_620_port, 
      DataPath_RF_bus_reg_dataout_621_port, 
      DataPath_RF_bus_reg_dataout_622_port, 
      DataPath_RF_bus_reg_dataout_623_port, 
      DataPath_RF_bus_reg_dataout_624_port, 
      DataPath_RF_bus_reg_dataout_625_port, 
      DataPath_RF_bus_reg_dataout_626_port, 
      DataPath_RF_bus_reg_dataout_627_port, 
      DataPath_RF_bus_reg_dataout_628_port, 
      DataPath_RF_bus_reg_dataout_629_port, 
      DataPath_RF_bus_reg_dataout_630_port, 
      DataPath_RF_bus_reg_dataout_631_port, 
      DataPath_RF_bus_reg_dataout_632_port, 
      DataPath_RF_bus_reg_dataout_633_port, 
      DataPath_RF_bus_reg_dataout_634_port, 
      DataPath_RF_bus_reg_dataout_635_port, 
      DataPath_RF_bus_reg_dataout_636_port, 
      DataPath_RF_bus_reg_dataout_637_port, 
      DataPath_RF_bus_reg_dataout_638_port, 
      DataPath_RF_bus_reg_dataout_639_port, 
      DataPath_RF_bus_reg_dataout_640_port, 
      DataPath_RF_bus_reg_dataout_641_port, 
      DataPath_RF_bus_reg_dataout_642_port, 
      DataPath_RF_bus_reg_dataout_643_port, 
      DataPath_RF_bus_reg_dataout_644_port, 
      DataPath_RF_bus_reg_dataout_645_port, 
      DataPath_RF_bus_reg_dataout_646_port, 
      DataPath_RF_bus_reg_dataout_647_port, 
      DataPath_RF_bus_reg_dataout_648_port, 
      DataPath_RF_bus_reg_dataout_649_port, 
      DataPath_RF_bus_reg_dataout_650_port, 
      DataPath_RF_bus_reg_dataout_651_port, 
      DataPath_RF_bus_reg_dataout_652_port, 
      DataPath_RF_bus_reg_dataout_653_port, 
      DataPath_RF_bus_reg_dataout_654_port, 
      DataPath_RF_bus_reg_dataout_655_port, 
      DataPath_RF_bus_reg_dataout_656_port, 
      DataPath_RF_bus_reg_dataout_657_port, 
      DataPath_RF_bus_reg_dataout_658_port, 
      DataPath_RF_bus_reg_dataout_659_port, 
      DataPath_RF_bus_reg_dataout_660_port, 
      DataPath_RF_bus_reg_dataout_661_port, 
      DataPath_RF_bus_reg_dataout_662_port, 
      DataPath_RF_bus_reg_dataout_663_port, 
      DataPath_RF_bus_reg_dataout_664_port, 
      DataPath_RF_bus_reg_dataout_665_port, 
      DataPath_RF_bus_reg_dataout_666_port, 
      DataPath_RF_bus_reg_dataout_667_port, 
      DataPath_RF_bus_reg_dataout_668_port, 
      DataPath_RF_bus_reg_dataout_669_port, 
      DataPath_RF_bus_reg_dataout_670_port, 
      DataPath_RF_bus_reg_dataout_671_port, 
      DataPath_RF_bus_reg_dataout_672_port, 
      DataPath_RF_bus_reg_dataout_673_port, 
      DataPath_RF_bus_reg_dataout_674_port, 
      DataPath_RF_bus_reg_dataout_675_port, 
      DataPath_RF_bus_reg_dataout_676_port, 
      DataPath_RF_bus_reg_dataout_677_port, 
      DataPath_RF_bus_reg_dataout_678_port, 
      DataPath_RF_bus_reg_dataout_679_port, 
      DataPath_RF_bus_reg_dataout_680_port, 
      DataPath_RF_bus_reg_dataout_681_port, 
      DataPath_RF_bus_reg_dataout_682_port, 
      DataPath_RF_bus_reg_dataout_683_port, 
      DataPath_RF_bus_reg_dataout_684_port, 
      DataPath_RF_bus_reg_dataout_685_port, 
      DataPath_RF_bus_reg_dataout_686_port, 
      DataPath_RF_bus_reg_dataout_687_port, 
      DataPath_RF_bus_reg_dataout_688_port, 
      DataPath_RF_bus_reg_dataout_689_port, 
      DataPath_RF_bus_reg_dataout_690_port, 
      DataPath_RF_bus_reg_dataout_691_port, 
      DataPath_RF_bus_reg_dataout_692_port, 
      DataPath_RF_bus_reg_dataout_693_port, 
      DataPath_RF_bus_reg_dataout_694_port, 
      DataPath_RF_bus_reg_dataout_695_port, 
      DataPath_RF_bus_reg_dataout_696_port, 
      DataPath_RF_bus_reg_dataout_697_port, 
      DataPath_RF_bus_reg_dataout_698_port, 
      DataPath_RF_bus_reg_dataout_699_port, 
      DataPath_RF_bus_reg_dataout_700_port, 
      DataPath_RF_bus_reg_dataout_701_port, 
      DataPath_RF_bus_reg_dataout_702_port, 
      DataPath_RF_bus_reg_dataout_703_port, 
      DataPath_RF_bus_reg_dataout_704_port, 
      DataPath_RF_bus_reg_dataout_705_port, 
      DataPath_RF_bus_reg_dataout_706_port, 
      DataPath_RF_bus_reg_dataout_707_port, 
      DataPath_RF_bus_reg_dataout_708_port, 
      DataPath_RF_bus_reg_dataout_709_port, 
      DataPath_RF_bus_reg_dataout_710_port, 
      DataPath_RF_bus_reg_dataout_711_port, 
      DataPath_RF_bus_reg_dataout_712_port, 
      DataPath_RF_bus_reg_dataout_713_port, 
      DataPath_RF_bus_reg_dataout_714_port, 
      DataPath_RF_bus_reg_dataout_715_port, 
      DataPath_RF_bus_reg_dataout_716_port, 
      DataPath_RF_bus_reg_dataout_717_port, 
      DataPath_RF_bus_reg_dataout_718_port, 
      DataPath_RF_bus_reg_dataout_719_port, 
      DataPath_RF_bus_reg_dataout_720_port, 
      DataPath_RF_bus_reg_dataout_721_port, 
      DataPath_RF_bus_reg_dataout_722_port, 
      DataPath_RF_bus_reg_dataout_723_port, 
      DataPath_RF_bus_reg_dataout_724_port, 
      DataPath_RF_bus_reg_dataout_725_port, 
      DataPath_RF_bus_reg_dataout_726_port, 
      DataPath_RF_bus_reg_dataout_727_port, 
      DataPath_RF_bus_reg_dataout_728_port, 
      DataPath_RF_bus_reg_dataout_729_port, 
      DataPath_RF_bus_reg_dataout_730_port, 
      DataPath_RF_bus_reg_dataout_731_port, 
      DataPath_RF_bus_reg_dataout_732_port, 
      DataPath_RF_bus_reg_dataout_733_port, 
      DataPath_RF_bus_reg_dataout_734_port, 
      DataPath_RF_bus_reg_dataout_735_port, 
      DataPath_RF_bus_reg_dataout_736_port, 
      DataPath_RF_bus_reg_dataout_737_port, 
      DataPath_RF_bus_reg_dataout_738_port, 
      DataPath_RF_bus_reg_dataout_739_port, 
      DataPath_RF_bus_reg_dataout_740_port, 
      DataPath_RF_bus_reg_dataout_741_port, 
      DataPath_RF_bus_reg_dataout_742_port, 
      DataPath_RF_bus_reg_dataout_743_port, 
      DataPath_RF_bus_reg_dataout_744_port, 
      DataPath_RF_bus_reg_dataout_745_port, 
      DataPath_RF_bus_reg_dataout_746_port, 
      DataPath_RF_bus_reg_dataout_747_port, 
      DataPath_RF_bus_reg_dataout_748_port, 
      DataPath_RF_bus_reg_dataout_749_port, 
      DataPath_RF_bus_reg_dataout_750_port, 
      DataPath_RF_bus_reg_dataout_751_port, 
      DataPath_RF_bus_reg_dataout_752_port, 
      DataPath_RF_bus_reg_dataout_753_port, 
      DataPath_RF_bus_reg_dataout_754_port, 
      DataPath_RF_bus_reg_dataout_755_port, 
      DataPath_RF_bus_reg_dataout_756_port, 
      DataPath_RF_bus_reg_dataout_757_port, 
      DataPath_RF_bus_reg_dataout_758_port, 
      DataPath_RF_bus_reg_dataout_759_port, 
      DataPath_RF_bus_reg_dataout_760_port, 
      DataPath_RF_bus_reg_dataout_761_port, 
      DataPath_RF_bus_reg_dataout_762_port, 
      DataPath_RF_bus_reg_dataout_763_port, 
      DataPath_RF_bus_reg_dataout_764_port, 
      DataPath_RF_bus_reg_dataout_765_port, 
      DataPath_RF_bus_reg_dataout_766_port, 
      DataPath_RF_bus_reg_dataout_767_port, 
      DataPath_RF_bus_reg_dataout_768_port, 
      DataPath_RF_bus_reg_dataout_769_port, 
      DataPath_RF_bus_reg_dataout_770_port, 
      DataPath_RF_bus_reg_dataout_771_port, 
      DataPath_RF_bus_reg_dataout_772_port, 
      DataPath_RF_bus_reg_dataout_773_port, 
      DataPath_RF_bus_reg_dataout_774_port, 
      DataPath_RF_bus_reg_dataout_775_port, 
      DataPath_RF_bus_reg_dataout_776_port, 
      DataPath_RF_bus_reg_dataout_777_port, 
      DataPath_RF_bus_reg_dataout_778_port, 
      DataPath_RF_bus_reg_dataout_779_port, 
      DataPath_RF_bus_reg_dataout_780_port, 
      DataPath_RF_bus_reg_dataout_781_port, 
      DataPath_RF_bus_reg_dataout_782_port, 
      DataPath_RF_bus_reg_dataout_783_port, 
      DataPath_RF_bus_reg_dataout_784_port, 
      DataPath_RF_bus_reg_dataout_785_port, 
      DataPath_RF_bus_reg_dataout_786_port, 
      DataPath_RF_bus_reg_dataout_787_port, 
      DataPath_RF_bus_reg_dataout_788_port, 
      DataPath_RF_bus_reg_dataout_789_port, 
      DataPath_RF_bus_reg_dataout_790_port, 
      DataPath_RF_bus_reg_dataout_791_port, 
      DataPath_RF_bus_reg_dataout_792_port, 
      DataPath_RF_bus_reg_dataout_793_port, 
      DataPath_RF_bus_reg_dataout_794_port, 
      DataPath_RF_bus_reg_dataout_795_port, 
      DataPath_RF_bus_reg_dataout_796_port, 
      DataPath_RF_bus_reg_dataout_797_port, 
      DataPath_RF_bus_reg_dataout_798_port, 
      DataPath_RF_bus_reg_dataout_799_port, 
      DataPath_RF_bus_reg_dataout_800_port, 
      DataPath_RF_bus_reg_dataout_801_port, 
      DataPath_RF_bus_reg_dataout_802_port, 
      DataPath_RF_bus_reg_dataout_803_port, 
      DataPath_RF_bus_reg_dataout_804_port, 
      DataPath_RF_bus_reg_dataout_805_port, 
      DataPath_RF_bus_reg_dataout_806_port, 
      DataPath_RF_bus_reg_dataout_807_port, 
      DataPath_RF_bus_reg_dataout_808_port, 
      DataPath_RF_bus_reg_dataout_809_port, 
      DataPath_RF_bus_reg_dataout_810_port, 
      DataPath_RF_bus_reg_dataout_811_port, 
      DataPath_RF_bus_reg_dataout_812_port, 
      DataPath_RF_bus_reg_dataout_813_port, 
      DataPath_RF_bus_reg_dataout_814_port, 
      DataPath_RF_bus_reg_dataout_815_port, 
      DataPath_RF_bus_reg_dataout_816_port, 
      DataPath_RF_bus_reg_dataout_817_port, 
      DataPath_RF_bus_reg_dataout_818_port, 
      DataPath_RF_bus_reg_dataout_819_port, 
      DataPath_RF_bus_reg_dataout_820_port, 
      DataPath_RF_bus_reg_dataout_821_port, 
      DataPath_RF_bus_reg_dataout_822_port, 
      DataPath_RF_bus_reg_dataout_823_port, 
      DataPath_RF_bus_reg_dataout_824_port, 
      DataPath_RF_bus_reg_dataout_825_port, 
      DataPath_RF_bus_reg_dataout_826_port, 
      DataPath_RF_bus_reg_dataout_827_port, 
      DataPath_RF_bus_reg_dataout_828_port, 
      DataPath_RF_bus_reg_dataout_829_port, 
      DataPath_RF_bus_reg_dataout_830_port, 
      DataPath_RF_bus_reg_dataout_831_port, 
      DataPath_RF_bus_reg_dataout_832_port, 
      DataPath_RF_bus_reg_dataout_833_port, 
      DataPath_RF_bus_reg_dataout_834_port, 
      DataPath_RF_bus_reg_dataout_835_port, 
      DataPath_RF_bus_reg_dataout_836_port, 
      DataPath_RF_bus_reg_dataout_837_port, 
      DataPath_RF_bus_reg_dataout_838_port, 
      DataPath_RF_bus_reg_dataout_839_port, 
      DataPath_RF_bus_reg_dataout_840_port, 
      DataPath_RF_bus_reg_dataout_841_port, 
      DataPath_RF_bus_reg_dataout_842_port, 
      DataPath_RF_bus_reg_dataout_843_port, 
      DataPath_RF_bus_reg_dataout_844_port, 
      DataPath_RF_bus_reg_dataout_845_port, 
      DataPath_RF_bus_reg_dataout_846_port, 
      DataPath_RF_bus_reg_dataout_847_port, 
      DataPath_RF_bus_reg_dataout_848_port, 
      DataPath_RF_bus_reg_dataout_849_port, 
      DataPath_RF_bus_reg_dataout_850_port, 
      DataPath_RF_bus_reg_dataout_851_port, 
      DataPath_RF_bus_reg_dataout_852_port, 
      DataPath_RF_bus_reg_dataout_853_port, 
      DataPath_RF_bus_reg_dataout_854_port, 
      DataPath_RF_bus_reg_dataout_855_port, 
      DataPath_RF_bus_reg_dataout_856_port, 
      DataPath_RF_bus_reg_dataout_857_port, 
      DataPath_RF_bus_reg_dataout_858_port, 
      DataPath_RF_bus_reg_dataout_859_port, 
      DataPath_RF_bus_reg_dataout_860_port, 
      DataPath_RF_bus_reg_dataout_861_port, 
      DataPath_RF_bus_reg_dataout_862_port, 
      DataPath_RF_bus_reg_dataout_863_port, 
      DataPath_RF_bus_reg_dataout_864_port, 
      DataPath_RF_bus_reg_dataout_865_port, 
      DataPath_RF_bus_reg_dataout_866_port, 
      DataPath_RF_bus_reg_dataout_867_port, 
      DataPath_RF_bus_reg_dataout_868_port, 
      DataPath_RF_bus_reg_dataout_869_port, 
      DataPath_RF_bus_reg_dataout_870_port, 
      DataPath_RF_bus_reg_dataout_871_port, 
      DataPath_RF_bus_reg_dataout_872_port, 
      DataPath_RF_bus_reg_dataout_873_port, 
      DataPath_RF_bus_reg_dataout_874_port, 
      DataPath_RF_bus_reg_dataout_875_port, 
      DataPath_RF_bus_reg_dataout_876_port, 
      DataPath_RF_bus_reg_dataout_877_port, 
      DataPath_RF_bus_reg_dataout_878_port, 
      DataPath_RF_bus_reg_dataout_879_port, 
      DataPath_RF_bus_reg_dataout_880_port, 
      DataPath_RF_bus_reg_dataout_881_port, 
      DataPath_RF_bus_reg_dataout_882_port, 
      DataPath_RF_bus_reg_dataout_883_port, 
      DataPath_RF_bus_reg_dataout_884_port, 
      DataPath_RF_bus_reg_dataout_885_port, 
      DataPath_RF_bus_reg_dataout_886_port, 
      DataPath_RF_bus_reg_dataout_887_port, 
      DataPath_RF_bus_reg_dataout_888_port, 
      DataPath_RF_bus_reg_dataout_889_port, 
      DataPath_RF_bus_reg_dataout_890_port, 
      DataPath_RF_bus_reg_dataout_891_port, 
      DataPath_RF_bus_reg_dataout_892_port, 
      DataPath_RF_bus_reg_dataout_893_port, 
      DataPath_RF_bus_reg_dataout_894_port, 
      DataPath_RF_bus_reg_dataout_895_port, 
      DataPath_RF_bus_reg_dataout_896_port, 
      DataPath_RF_bus_reg_dataout_897_port, 
      DataPath_RF_bus_reg_dataout_898_port, 
      DataPath_RF_bus_reg_dataout_899_port, 
      DataPath_RF_bus_reg_dataout_900_port, 
      DataPath_RF_bus_reg_dataout_901_port, 
      DataPath_RF_bus_reg_dataout_902_port, 
      DataPath_RF_bus_reg_dataout_903_port, 
      DataPath_RF_bus_reg_dataout_904_port, 
      DataPath_RF_bus_reg_dataout_905_port, 
      DataPath_RF_bus_reg_dataout_906_port, 
      DataPath_RF_bus_reg_dataout_907_port, 
      DataPath_RF_bus_reg_dataout_908_port, 
      DataPath_RF_bus_reg_dataout_909_port, 
      DataPath_RF_bus_reg_dataout_910_port, 
      DataPath_RF_bus_reg_dataout_911_port, 
      DataPath_RF_bus_reg_dataout_912_port, 
      DataPath_RF_bus_reg_dataout_913_port, 
      DataPath_RF_bus_reg_dataout_914_port, 
      DataPath_RF_bus_reg_dataout_915_port, 
      DataPath_RF_bus_reg_dataout_916_port, 
      DataPath_RF_bus_reg_dataout_917_port, 
      DataPath_RF_bus_reg_dataout_918_port, 
      DataPath_RF_bus_reg_dataout_919_port, 
      DataPath_RF_bus_reg_dataout_920_port, 
      DataPath_RF_bus_reg_dataout_921_port, 
      DataPath_RF_bus_reg_dataout_922_port, 
      DataPath_RF_bus_reg_dataout_923_port, 
      DataPath_RF_bus_reg_dataout_924_port, 
      DataPath_RF_bus_reg_dataout_925_port, 
      DataPath_RF_bus_reg_dataout_926_port, 
      DataPath_RF_bus_reg_dataout_927_port, 
      DataPath_RF_bus_reg_dataout_928_port, 
      DataPath_RF_bus_reg_dataout_929_port, 
      DataPath_RF_bus_reg_dataout_930_port, 
      DataPath_RF_bus_reg_dataout_931_port, 
      DataPath_RF_bus_reg_dataout_932_port, 
      DataPath_RF_bus_reg_dataout_933_port, 
      DataPath_RF_bus_reg_dataout_934_port, 
      DataPath_RF_bus_reg_dataout_935_port, 
      DataPath_RF_bus_reg_dataout_936_port, 
      DataPath_RF_bus_reg_dataout_937_port, 
      DataPath_RF_bus_reg_dataout_938_port, 
      DataPath_RF_bus_reg_dataout_939_port, 
      DataPath_RF_bus_reg_dataout_940_port, 
      DataPath_RF_bus_reg_dataout_941_port, 
      DataPath_RF_bus_reg_dataout_942_port, 
      DataPath_RF_bus_reg_dataout_943_port, 
      DataPath_RF_bus_reg_dataout_944_port, 
      DataPath_RF_bus_reg_dataout_945_port, 
      DataPath_RF_bus_reg_dataout_946_port, 
      DataPath_RF_bus_reg_dataout_947_port, 
      DataPath_RF_bus_reg_dataout_948_port, 
      DataPath_RF_bus_reg_dataout_949_port, 
      DataPath_RF_bus_reg_dataout_950_port, 
      DataPath_RF_bus_reg_dataout_951_port, 
      DataPath_RF_bus_reg_dataout_952_port, 
      DataPath_RF_bus_reg_dataout_953_port, 
      DataPath_RF_bus_reg_dataout_954_port, 
      DataPath_RF_bus_reg_dataout_955_port, 
      DataPath_RF_bus_reg_dataout_956_port, 
      DataPath_RF_bus_reg_dataout_957_port, 
      DataPath_RF_bus_reg_dataout_958_port, 
      DataPath_RF_bus_reg_dataout_959_port, 
      DataPath_RF_bus_reg_dataout_960_port, 
      DataPath_RF_bus_reg_dataout_961_port, 
      DataPath_RF_bus_reg_dataout_962_port, 
      DataPath_RF_bus_reg_dataout_963_port, 
      DataPath_RF_bus_reg_dataout_964_port, 
      DataPath_RF_bus_reg_dataout_965_port, 
      DataPath_RF_bus_reg_dataout_966_port, 
      DataPath_RF_bus_reg_dataout_967_port, 
      DataPath_RF_bus_reg_dataout_968_port, 
      DataPath_RF_bus_reg_dataout_969_port, 
      DataPath_RF_bus_reg_dataout_970_port, 
      DataPath_RF_bus_reg_dataout_971_port, 
      DataPath_RF_bus_reg_dataout_972_port, 
      DataPath_RF_bus_reg_dataout_973_port, 
      DataPath_RF_bus_reg_dataout_974_port, 
      DataPath_RF_bus_reg_dataout_975_port, 
      DataPath_RF_bus_reg_dataout_976_port, 
      DataPath_RF_bus_reg_dataout_977_port, 
      DataPath_RF_bus_reg_dataout_978_port, 
      DataPath_RF_bus_reg_dataout_979_port, 
      DataPath_RF_bus_reg_dataout_980_port, 
      DataPath_RF_bus_reg_dataout_981_port, 
      DataPath_RF_bus_reg_dataout_982_port, 
      DataPath_RF_bus_reg_dataout_983_port, 
      DataPath_RF_bus_reg_dataout_984_port, 
      DataPath_RF_bus_reg_dataout_985_port, 
      DataPath_RF_bus_reg_dataout_986_port, 
      DataPath_RF_bus_reg_dataout_987_port, 
      DataPath_RF_bus_reg_dataout_988_port, 
      DataPath_RF_bus_reg_dataout_989_port, 
      DataPath_RF_bus_reg_dataout_990_port, 
      DataPath_RF_bus_reg_dataout_991_port, 
      DataPath_RF_bus_reg_dataout_992_port, 
      DataPath_RF_bus_reg_dataout_993_port, 
      DataPath_RF_bus_reg_dataout_994_port, 
      DataPath_RF_bus_reg_dataout_995_port, 
      DataPath_RF_bus_reg_dataout_996_port, 
      DataPath_RF_bus_reg_dataout_997_port, 
      DataPath_RF_bus_reg_dataout_998_port, 
      DataPath_RF_bus_reg_dataout_999_port, 
      DataPath_RF_bus_reg_dataout_1000_port, 
      DataPath_RF_bus_reg_dataout_1001_port, 
      DataPath_RF_bus_reg_dataout_1002_port, 
      DataPath_RF_bus_reg_dataout_1003_port, 
      DataPath_RF_bus_reg_dataout_1004_port, 
      DataPath_RF_bus_reg_dataout_1005_port, 
      DataPath_RF_bus_reg_dataout_1006_port, 
      DataPath_RF_bus_reg_dataout_1007_port, 
      DataPath_RF_bus_reg_dataout_1008_port, 
      DataPath_RF_bus_reg_dataout_1009_port, 
      DataPath_RF_bus_reg_dataout_1010_port, 
      DataPath_RF_bus_reg_dataout_1011_port, 
      DataPath_RF_bus_reg_dataout_1012_port, 
      DataPath_RF_bus_reg_dataout_1013_port, 
      DataPath_RF_bus_reg_dataout_1014_port, 
      DataPath_RF_bus_reg_dataout_1015_port, 
      DataPath_RF_bus_reg_dataout_1016_port, 
      DataPath_RF_bus_reg_dataout_1017_port, 
      DataPath_RF_bus_reg_dataout_1018_port, 
      DataPath_RF_bus_reg_dataout_1019_port, 
      DataPath_RF_bus_reg_dataout_1020_port, 
      DataPath_RF_bus_reg_dataout_1021_port, 
      DataPath_RF_bus_reg_dataout_1022_port, 
      DataPath_RF_bus_reg_dataout_1023_port, 
      DataPath_RF_bus_reg_dataout_1024_port, 
      DataPath_RF_bus_reg_dataout_1025_port, 
      DataPath_RF_bus_reg_dataout_1026_port, 
      DataPath_RF_bus_reg_dataout_1027_port, 
      DataPath_RF_bus_reg_dataout_1028_port, 
      DataPath_RF_bus_reg_dataout_1029_port, 
      DataPath_RF_bus_reg_dataout_1030_port, 
      DataPath_RF_bus_reg_dataout_1031_port, 
      DataPath_RF_bus_reg_dataout_1032_port, 
      DataPath_RF_bus_reg_dataout_1033_port, 
      DataPath_RF_bus_reg_dataout_1034_port, 
      DataPath_RF_bus_reg_dataout_1035_port, 
      DataPath_RF_bus_reg_dataout_1036_port, 
      DataPath_RF_bus_reg_dataout_1037_port, 
      DataPath_RF_bus_reg_dataout_1038_port, 
      DataPath_RF_bus_reg_dataout_1039_port, 
      DataPath_RF_bus_reg_dataout_1040_port, 
      DataPath_RF_bus_reg_dataout_1041_port, 
      DataPath_RF_bus_reg_dataout_1042_port, 
      DataPath_RF_bus_reg_dataout_1043_port, 
      DataPath_RF_bus_reg_dataout_1044_port, 
      DataPath_RF_bus_reg_dataout_1045_port, 
      DataPath_RF_bus_reg_dataout_1046_port, 
      DataPath_RF_bus_reg_dataout_1047_port, 
      DataPath_RF_bus_reg_dataout_1048_port, 
      DataPath_RF_bus_reg_dataout_1049_port, 
      DataPath_RF_bus_reg_dataout_1050_port, 
      DataPath_RF_bus_reg_dataout_1051_port, 
      DataPath_RF_bus_reg_dataout_1052_port, 
      DataPath_RF_bus_reg_dataout_1053_port, 
      DataPath_RF_bus_reg_dataout_1054_port, 
      DataPath_RF_bus_reg_dataout_1055_port, 
      DataPath_RF_bus_reg_dataout_1056_port, 
      DataPath_RF_bus_reg_dataout_1057_port, 
      DataPath_RF_bus_reg_dataout_1058_port, 
      DataPath_RF_bus_reg_dataout_1059_port, 
      DataPath_RF_bus_reg_dataout_1060_port, 
      DataPath_RF_bus_reg_dataout_1061_port, 
      DataPath_RF_bus_reg_dataout_1062_port, 
      DataPath_RF_bus_reg_dataout_1063_port, 
      DataPath_RF_bus_reg_dataout_1064_port, 
      DataPath_RF_bus_reg_dataout_1065_port, 
      DataPath_RF_bus_reg_dataout_1066_port, 
      DataPath_RF_bus_reg_dataout_1067_port, 
      DataPath_RF_bus_reg_dataout_1068_port, 
      DataPath_RF_bus_reg_dataout_1069_port, 
      DataPath_RF_bus_reg_dataout_1070_port, 
      DataPath_RF_bus_reg_dataout_1071_port, 
      DataPath_RF_bus_reg_dataout_1072_port, 
      DataPath_RF_bus_reg_dataout_1073_port, 
      DataPath_RF_bus_reg_dataout_1074_port, 
      DataPath_RF_bus_reg_dataout_1075_port, 
      DataPath_RF_bus_reg_dataout_1076_port, 
      DataPath_RF_bus_reg_dataout_1077_port, 
      DataPath_RF_bus_reg_dataout_1078_port, 
      DataPath_RF_bus_reg_dataout_1079_port, 
      DataPath_RF_bus_reg_dataout_1080_port, 
      DataPath_RF_bus_reg_dataout_1081_port, 
      DataPath_RF_bus_reg_dataout_1082_port, 
      DataPath_RF_bus_reg_dataout_1083_port, 
      DataPath_RF_bus_reg_dataout_1084_port, 
      DataPath_RF_bus_reg_dataout_1085_port, 
      DataPath_RF_bus_reg_dataout_1086_port, 
      DataPath_RF_bus_reg_dataout_1087_port, 
      DataPath_RF_bus_reg_dataout_1088_port, 
      DataPath_RF_bus_reg_dataout_1089_port, 
      DataPath_RF_bus_reg_dataout_1090_port, 
      DataPath_RF_bus_reg_dataout_1091_port, 
      DataPath_RF_bus_reg_dataout_1092_port, 
      DataPath_RF_bus_reg_dataout_1093_port, 
      DataPath_RF_bus_reg_dataout_1094_port, 
      DataPath_RF_bus_reg_dataout_1095_port, 
      DataPath_RF_bus_reg_dataout_1096_port, 
      DataPath_RF_bus_reg_dataout_1097_port, 
      DataPath_RF_bus_reg_dataout_1098_port, 
      DataPath_RF_bus_reg_dataout_1099_port, 
      DataPath_RF_bus_reg_dataout_1100_port, 
      DataPath_RF_bus_reg_dataout_1101_port, 
      DataPath_RF_bus_reg_dataout_1102_port, 
      DataPath_RF_bus_reg_dataout_1103_port, 
      DataPath_RF_bus_reg_dataout_1104_port, 
      DataPath_RF_bus_reg_dataout_1105_port, 
      DataPath_RF_bus_reg_dataout_1106_port, 
      DataPath_RF_bus_reg_dataout_1107_port, 
      DataPath_RF_bus_reg_dataout_1108_port, 
      DataPath_RF_bus_reg_dataout_1109_port, 
      DataPath_RF_bus_reg_dataout_1110_port, 
      DataPath_RF_bus_reg_dataout_1111_port, 
      DataPath_RF_bus_reg_dataout_1112_port, 
      DataPath_RF_bus_reg_dataout_1113_port, 
      DataPath_RF_bus_reg_dataout_1114_port, 
      DataPath_RF_bus_reg_dataout_1115_port, 
      DataPath_RF_bus_reg_dataout_1116_port, 
      DataPath_RF_bus_reg_dataout_1117_port, 
      DataPath_RF_bus_reg_dataout_1118_port, 
      DataPath_RF_bus_reg_dataout_1119_port, 
      DataPath_RF_bus_reg_dataout_1120_port, 
      DataPath_RF_bus_reg_dataout_1121_port, 
      DataPath_RF_bus_reg_dataout_1122_port, 
      DataPath_RF_bus_reg_dataout_1123_port, 
      DataPath_RF_bus_reg_dataout_1124_port, 
      DataPath_RF_bus_reg_dataout_1125_port, 
      DataPath_RF_bus_reg_dataout_1126_port, 
      DataPath_RF_bus_reg_dataout_1127_port, 
      DataPath_RF_bus_reg_dataout_1128_port, 
      DataPath_RF_bus_reg_dataout_1129_port, 
      DataPath_RF_bus_reg_dataout_1130_port, 
      DataPath_RF_bus_reg_dataout_1131_port, 
      DataPath_RF_bus_reg_dataout_1132_port, 
      DataPath_RF_bus_reg_dataout_1133_port, 
      DataPath_RF_bus_reg_dataout_1134_port, 
      DataPath_RF_bus_reg_dataout_1135_port, 
      DataPath_RF_bus_reg_dataout_1136_port, 
      DataPath_RF_bus_reg_dataout_1137_port, 
      DataPath_RF_bus_reg_dataout_1138_port, 
      DataPath_RF_bus_reg_dataout_1139_port, 
      DataPath_RF_bus_reg_dataout_1140_port, 
      DataPath_RF_bus_reg_dataout_1141_port, 
      DataPath_RF_bus_reg_dataout_1142_port, 
      DataPath_RF_bus_reg_dataout_1143_port, 
      DataPath_RF_bus_reg_dataout_1144_port, 
      DataPath_RF_bus_reg_dataout_1145_port, 
      DataPath_RF_bus_reg_dataout_1146_port, 
      DataPath_RF_bus_reg_dataout_1147_port, 
      DataPath_RF_bus_reg_dataout_1148_port, 
      DataPath_RF_bus_reg_dataout_1149_port, 
      DataPath_RF_bus_reg_dataout_1150_port, 
      DataPath_RF_bus_reg_dataout_1151_port, 
      DataPath_RF_bus_reg_dataout_1152_port, 
      DataPath_RF_bus_reg_dataout_1153_port, 
      DataPath_RF_bus_reg_dataout_1154_port, 
      DataPath_RF_bus_reg_dataout_1155_port, 
      DataPath_RF_bus_reg_dataout_1156_port, 
      DataPath_RF_bus_reg_dataout_1157_port, 
      DataPath_RF_bus_reg_dataout_1158_port, 
      DataPath_RF_bus_reg_dataout_1159_port, 
      DataPath_RF_bus_reg_dataout_1160_port, 
      DataPath_RF_bus_reg_dataout_1161_port, 
      DataPath_RF_bus_reg_dataout_1162_port, 
      DataPath_RF_bus_reg_dataout_1163_port, 
      DataPath_RF_bus_reg_dataout_1164_port, 
      DataPath_RF_bus_reg_dataout_1165_port, 
      DataPath_RF_bus_reg_dataout_1166_port, 
      DataPath_RF_bus_reg_dataout_1167_port, 
      DataPath_RF_bus_reg_dataout_1168_port, 
      DataPath_RF_bus_reg_dataout_1169_port, 
      DataPath_RF_bus_reg_dataout_1170_port, 
      DataPath_RF_bus_reg_dataout_1171_port, 
      DataPath_RF_bus_reg_dataout_1172_port, 
      DataPath_RF_bus_reg_dataout_1173_port, 
      DataPath_RF_bus_reg_dataout_1174_port, 
      DataPath_RF_bus_reg_dataout_1175_port, 
      DataPath_RF_bus_reg_dataout_1176_port, 
      DataPath_RF_bus_reg_dataout_1177_port, 
      DataPath_RF_bus_reg_dataout_1178_port, 
      DataPath_RF_bus_reg_dataout_1179_port, 
      DataPath_RF_bus_reg_dataout_1180_port, 
      DataPath_RF_bus_reg_dataout_1181_port, 
      DataPath_RF_bus_reg_dataout_1182_port, 
      DataPath_RF_bus_reg_dataout_1183_port, 
      DataPath_RF_bus_reg_dataout_1184_port, 
      DataPath_RF_bus_reg_dataout_1185_port, 
      DataPath_RF_bus_reg_dataout_1186_port, 
      DataPath_RF_bus_reg_dataout_1187_port, 
      DataPath_RF_bus_reg_dataout_1188_port, 
      DataPath_RF_bus_reg_dataout_1189_port, 
      DataPath_RF_bus_reg_dataout_1190_port, 
      DataPath_RF_bus_reg_dataout_1191_port, 
      DataPath_RF_bus_reg_dataout_1192_port, 
      DataPath_RF_bus_reg_dataout_1193_port, 
      DataPath_RF_bus_reg_dataout_1194_port, 
      DataPath_RF_bus_reg_dataout_1195_port, 
      DataPath_RF_bus_reg_dataout_1196_port, 
      DataPath_RF_bus_reg_dataout_1197_port, 
      DataPath_RF_bus_reg_dataout_1198_port, 
      DataPath_RF_bus_reg_dataout_1199_port, 
      DataPath_RF_bus_reg_dataout_1200_port, 
      DataPath_RF_bus_reg_dataout_1201_port, 
      DataPath_RF_bus_reg_dataout_1202_port, 
      DataPath_RF_bus_reg_dataout_1203_port, 
      DataPath_RF_bus_reg_dataout_1204_port, 
      DataPath_RF_bus_reg_dataout_1205_port, 
      DataPath_RF_bus_reg_dataout_1206_port, 
      DataPath_RF_bus_reg_dataout_1207_port, 
      DataPath_RF_bus_reg_dataout_1208_port, 
      DataPath_RF_bus_reg_dataout_1209_port, 
      DataPath_RF_bus_reg_dataout_1210_port, 
      DataPath_RF_bus_reg_dataout_1211_port, 
      DataPath_RF_bus_reg_dataout_1212_port, 
      DataPath_RF_bus_reg_dataout_1213_port, 
      DataPath_RF_bus_reg_dataout_1214_port, 
      DataPath_RF_bus_reg_dataout_1215_port, 
      DataPath_RF_bus_reg_dataout_1216_port, 
      DataPath_RF_bus_reg_dataout_1217_port, 
      DataPath_RF_bus_reg_dataout_1218_port, 
      DataPath_RF_bus_reg_dataout_1219_port, 
      DataPath_RF_bus_reg_dataout_1220_port, 
      DataPath_RF_bus_reg_dataout_1221_port, 
      DataPath_RF_bus_reg_dataout_1222_port, 
      DataPath_RF_bus_reg_dataout_1223_port, 
      DataPath_RF_bus_reg_dataout_1224_port, 
      DataPath_RF_bus_reg_dataout_1225_port, 
      DataPath_RF_bus_reg_dataout_1226_port, 
      DataPath_RF_bus_reg_dataout_1227_port, 
      DataPath_RF_bus_reg_dataout_1228_port, 
      DataPath_RF_bus_reg_dataout_1229_port, 
      DataPath_RF_bus_reg_dataout_1230_port, 
      DataPath_RF_bus_reg_dataout_1231_port, 
      DataPath_RF_bus_reg_dataout_1232_port, 
      DataPath_RF_bus_reg_dataout_1233_port, 
      DataPath_RF_bus_reg_dataout_1234_port, 
      DataPath_RF_bus_reg_dataout_1235_port, 
      DataPath_RF_bus_reg_dataout_1236_port, 
      DataPath_RF_bus_reg_dataout_1237_port, 
      DataPath_RF_bus_reg_dataout_1238_port, 
      DataPath_RF_bus_reg_dataout_1239_port, 
      DataPath_RF_bus_reg_dataout_1240_port, 
      DataPath_RF_bus_reg_dataout_1241_port, 
      DataPath_RF_bus_reg_dataout_1242_port, 
      DataPath_RF_bus_reg_dataout_1243_port, 
      DataPath_RF_bus_reg_dataout_1244_port, 
      DataPath_RF_bus_reg_dataout_1245_port, 
      DataPath_RF_bus_reg_dataout_1246_port, 
      DataPath_RF_bus_reg_dataout_1247_port, 
      DataPath_RF_bus_reg_dataout_1248_port, 
      DataPath_RF_bus_reg_dataout_1249_port, 
      DataPath_RF_bus_reg_dataout_1250_port, 
      DataPath_RF_bus_reg_dataout_1251_port, 
      DataPath_RF_bus_reg_dataout_1252_port, 
      DataPath_RF_bus_reg_dataout_1253_port, 
      DataPath_RF_bus_reg_dataout_1254_port, 
      DataPath_RF_bus_reg_dataout_1255_port, 
      DataPath_RF_bus_reg_dataout_1256_port, 
      DataPath_RF_bus_reg_dataout_1257_port, 
      DataPath_RF_bus_reg_dataout_1258_port, 
      DataPath_RF_bus_reg_dataout_1259_port, 
      DataPath_RF_bus_reg_dataout_1260_port, 
      DataPath_RF_bus_reg_dataout_1261_port, 
      DataPath_RF_bus_reg_dataout_1262_port, 
      DataPath_RF_bus_reg_dataout_1263_port, 
      DataPath_RF_bus_reg_dataout_1264_port, 
      DataPath_RF_bus_reg_dataout_1265_port, 
      DataPath_RF_bus_reg_dataout_1266_port, 
      DataPath_RF_bus_reg_dataout_1267_port, 
      DataPath_RF_bus_reg_dataout_1268_port, 
      DataPath_RF_bus_reg_dataout_1269_port, 
      DataPath_RF_bus_reg_dataout_1270_port, 
      DataPath_RF_bus_reg_dataout_1271_port, 
      DataPath_RF_bus_reg_dataout_1272_port, 
      DataPath_RF_bus_reg_dataout_1273_port, 
      DataPath_RF_bus_reg_dataout_1274_port, 
      DataPath_RF_bus_reg_dataout_1275_port, 
      DataPath_RF_bus_reg_dataout_1276_port, 
      DataPath_RF_bus_reg_dataout_1277_port, 
      DataPath_RF_bus_reg_dataout_1278_port, 
      DataPath_RF_bus_reg_dataout_1279_port, 
      DataPath_RF_bus_reg_dataout_1280_port, 
      DataPath_RF_bus_reg_dataout_1281_port, 
      DataPath_RF_bus_reg_dataout_1282_port, 
      DataPath_RF_bus_reg_dataout_1283_port, 
      DataPath_RF_bus_reg_dataout_1284_port, 
      DataPath_RF_bus_reg_dataout_1285_port, 
      DataPath_RF_bus_reg_dataout_1286_port, 
      DataPath_RF_bus_reg_dataout_1287_port, 
      DataPath_RF_bus_reg_dataout_1288_port, 
      DataPath_RF_bus_reg_dataout_1289_port, 
      DataPath_RF_bus_reg_dataout_1290_port, 
      DataPath_RF_bus_reg_dataout_1291_port, 
      DataPath_RF_bus_reg_dataout_1292_port, 
      DataPath_RF_bus_reg_dataout_1293_port, 
      DataPath_RF_bus_reg_dataout_1294_port, 
      DataPath_RF_bus_reg_dataout_1295_port, 
      DataPath_RF_bus_reg_dataout_1296_port, 
      DataPath_RF_bus_reg_dataout_1297_port, 
      DataPath_RF_bus_reg_dataout_1298_port, 
      DataPath_RF_bus_reg_dataout_1299_port, 
      DataPath_RF_bus_reg_dataout_1300_port, 
      DataPath_RF_bus_reg_dataout_1301_port, 
      DataPath_RF_bus_reg_dataout_1302_port, 
      DataPath_RF_bus_reg_dataout_1303_port, 
      DataPath_RF_bus_reg_dataout_1304_port, 
      DataPath_RF_bus_reg_dataout_1305_port, 
      DataPath_RF_bus_reg_dataout_1306_port, 
      DataPath_RF_bus_reg_dataout_1307_port, 
      DataPath_RF_bus_reg_dataout_1308_port, 
      DataPath_RF_bus_reg_dataout_1309_port, 
      DataPath_RF_bus_reg_dataout_1310_port, 
      DataPath_RF_bus_reg_dataout_1311_port, 
      DataPath_RF_bus_reg_dataout_1312_port, 
      DataPath_RF_bus_reg_dataout_1313_port, 
      DataPath_RF_bus_reg_dataout_1314_port, 
      DataPath_RF_bus_reg_dataout_1315_port, 
      DataPath_RF_bus_reg_dataout_1316_port, 
      DataPath_RF_bus_reg_dataout_1317_port, 
      DataPath_RF_bus_reg_dataout_1318_port, 
      DataPath_RF_bus_reg_dataout_1319_port, 
      DataPath_RF_bus_reg_dataout_1320_port, 
      DataPath_RF_bus_reg_dataout_1321_port, 
      DataPath_RF_bus_reg_dataout_1322_port, 
      DataPath_RF_bus_reg_dataout_1323_port, 
      DataPath_RF_bus_reg_dataout_1324_port, 
      DataPath_RF_bus_reg_dataout_1325_port, 
      DataPath_RF_bus_reg_dataout_1326_port, 
      DataPath_RF_bus_reg_dataout_1327_port, 
      DataPath_RF_bus_reg_dataout_1328_port, 
      DataPath_RF_bus_reg_dataout_1329_port, 
      DataPath_RF_bus_reg_dataout_1330_port, 
      DataPath_RF_bus_reg_dataout_1331_port, 
      DataPath_RF_bus_reg_dataout_1332_port, 
      DataPath_RF_bus_reg_dataout_1333_port, 
      DataPath_RF_bus_reg_dataout_1334_port, 
      DataPath_RF_bus_reg_dataout_1335_port, 
      DataPath_RF_bus_reg_dataout_1336_port, 
      DataPath_RF_bus_reg_dataout_1337_port, 
      DataPath_RF_bus_reg_dataout_1338_port, 
      DataPath_RF_bus_reg_dataout_1339_port, 
      DataPath_RF_bus_reg_dataout_1340_port, 
      DataPath_RF_bus_reg_dataout_1341_port, 
      DataPath_RF_bus_reg_dataout_1342_port, 
      DataPath_RF_bus_reg_dataout_1343_port, 
      DataPath_RF_bus_reg_dataout_1344_port, 
      DataPath_RF_bus_reg_dataout_1345_port, 
      DataPath_RF_bus_reg_dataout_1346_port, 
      DataPath_RF_bus_reg_dataout_1347_port, 
      DataPath_RF_bus_reg_dataout_1348_port, 
      DataPath_RF_bus_reg_dataout_1349_port, 
      DataPath_RF_bus_reg_dataout_1350_port, 
      DataPath_RF_bus_reg_dataout_1351_port, 
      DataPath_RF_bus_reg_dataout_1352_port, 
      DataPath_RF_bus_reg_dataout_1353_port, 
      DataPath_RF_bus_reg_dataout_1354_port, 
      DataPath_RF_bus_reg_dataout_1355_port, 
      DataPath_RF_bus_reg_dataout_1356_port, 
      DataPath_RF_bus_reg_dataout_1357_port, 
      DataPath_RF_bus_reg_dataout_1358_port, 
      DataPath_RF_bus_reg_dataout_1359_port, 
      DataPath_RF_bus_reg_dataout_1360_port, 
      DataPath_RF_bus_reg_dataout_1361_port, 
      DataPath_RF_bus_reg_dataout_1362_port, 
      DataPath_RF_bus_reg_dataout_1363_port, 
      DataPath_RF_bus_reg_dataout_1364_port, 
      DataPath_RF_bus_reg_dataout_1365_port, 
      DataPath_RF_bus_reg_dataout_1366_port, 
      DataPath_RF_bus_reg_dataout_1367_port, 
      DataPath_RF_bus_reg_dataout_1368_port, 
      DataPath_RF_bus_reg_dataout_1369_port, 
      DataPath_RF_bus_reg_dataout_1370_port, 
      DataPath_RF_bus_reg_dataout_1371_port, 
      DataPath_RF_bus_reg_dataout_1372_port, 
      DataPath_RF_bus_reg_dataout_1373_port, 
      DataPath_RF_bus_reg_dataout_1374_port, 
      DataPath_RF_bus_reg_dataout_1375_port, 
      DataPath_RF_bus_reg_dataout_1376_port, 
      DataPath_RF_bus_reg_dataout_1377_port, 
      DataPath_RF_bus_reg_dataout_1378_port, 
      DataPath_RF_bus_reg_dataout_1379_port, 
      DataPath_RF_bus_reg_dataout_1380_port, 
      DataPath_RF_bus_reg_dataout_1381_port, 
      DataPath_RF_bus_reg_dataout_1382_port, 
      DataPath_RF_bus_reg_dataout_1383_port, 
      DataPath_RF_bus_reg_dataout_1384_port, 
      DataPath_RF_bus_reg_dataout_1385_port, 
      DataPath_RF_bus_reg_dataout_1386_port, 
      DataPath_RF_bus_reg_dataout_1387_port, 
      DataPath_RF_bus_reg_dataout_1388_port, 
      DataPath_RF_bus_reg_dataout_1389_port, 
      DataPath_RF_bus_reg_dataout_1390_port, 
      DataPath_RF_bus_reg_dataout_1391_port, 
      DataPath_RF_bus_reg_dataout_1392_port, 
      DataPath_RF_bus_reg_dataout_1393_port, 
      DataPath_RF_bus_reg_dataout_1394_port, 
      DataPath_RF_bus_reg_dataout_1395_port, 
      DataPath_RF_bus_reg_dataout_1396_port, 
      DataPath_RF_bus_reg_dataout_1397_port, 
      DataPath_RF_bus_reg_dataout_1398_port, 
      DataPath_RF_bus_reg_dataout_1399_port, 
      DataPath_RF_bus_reg_dataout_1400_port, 
      DataPath_RF_bus_reg_dataout_1401_port, 
      DataPath_RF_bus_reg_dataout_1402_port, 
      DataPath_RF_bus_reg_dataout_1403_port, 
      DataPath_RF_bus_reg_dataout_1404_port, 
      DataPath_RF_bus_reg_dataout_1405_port, 
      DataPath_RF_bus_reg_dataout_1406_port, 
      DataPath_RF_bus_reg_dataout_1407_port, 
      DataPath_RF_bus_reg_dataout_1408_port, 
      DataPath_RF_bus_reg_dataout_1409_port, 
      DataPath_RF_bus_reg_dataout_1410_port, 
      DataPath_RF_bus_reg_dataout_1411_port, 
      DataPath_RF_bus_reg_dataout_1412_port, 
      DataPath_RF_bus_reg_dataout_1413_port, 
      DataPath_RF_bus_reg_dataout_1414_port, 
      DataPath_RF_bus_reg_dataout_1415_port, 
      DataPath_RF_bus_reg_dataout_1416_port, 
      DataPath_RF_bus_reg_dataout_1417_port, 
      DataPath_RF_bus_reg_dataout_1418_port, 
      DataPath_RF_bus_reg_dataout_1419_port, 
      DataPath_RF_bus_reg_dataout_1420_port, 
      DataPath_RF_bus_reg_dataout_1421_port, 
      DataPath_RF_bus_reg_dataout_1422_port, 
      DataPath_RF_bus_reg_dataout_1423_port, 
      DataPath_RF_bus_reg_dataout_1424_port, 
      DataPath_RF_bus_reg_dataout_1425_port, 
      DataPath_RF_bus_reg_dataout_1426_port, 
      DataPath_RF_bus_reg_dataout_1427_port, 
      DataPath_RF_bus_reg_dataout_1428_port, 
      DataPath_RF_bus_reg_dataout_1429_port, 
      DataPath_RF_bus_reg_dataout_1430_port, 
      DataPath_RF_bus_reg_dataout_1431_port, 
      DataPath_RF_bus_reg_dataout_1432_port, 
      DataPath_RF_bus_reg_dataout_1433_port, 
      DataPath_RF_bus_reg_dataout_1434_port, 
      DataPath_RF_bus_reg_dataout_1435_port, 
      DataPath_RF_bus_reg_dataout_1436_port, 
      DataPath_RF_bus_reg_dataout_1437_port, 
      DataPath_RF_bus_reg_dataout_1438_port, 
      DataPath_RF_bus_reg_dataout_1439_port, 
      DataPath_RF_bus_reg_dataout_1440_port, 
      DataPath_RF_bus_reg_dataout_1441_port, 
      DataPath_RF_bus_reg_dataout_1442_port, 
      DataPath_RF_bus_reg_dataout_1443_port, 
      DataPath_RF_bus_reg_dataout_1444_port, 
      DataPath_RF_bus_reg_dataout_1445_port, 
      DataPath_RF_bus_reg_dataout_1446_port, 
      DataPath_RF_bus_reg_dataout_1447_port, 
      DataPath_RF_bus_reg_dataout_1448_port, 
      DataPath_RF_bus_reg_dataout_1449_port, 
      DataPath_RF_bus_reg_dataout_1450_port, 
      DataPath_RF_bus_reg_dataout_1451_port, 
      DataPath_RF_bus_reg_dataout_1452_port, 
      DataPath_RF_bus_reg_dataout_1453_port, 
      DataPath_RF_bus_reg_dataout_1454_port, 
      DataPath_RF_bus_reg_dataout_1455_port, 
      DataPath_RF_bus_reg_dataout_1456_port, 
      DataPath_RF_bus_reg_dataout_1457_port, 
      DataPath_RF_bus_reg_dataout_1458_port, 
      DataPath_RF_bus_reg_dataout_1459_port, 
      DataPath_RF_bus_reg_dataout_1460_port, 
      DataPath_RF_bus_reg_dataout_1461_port, 
      DataPath_RF_bus_reg_dataout_1462_port, 
      DataPath_RF_bus_reg_dataout_1463_port, 
      DataPath_RF_bus_reg_dataout_1464_port, 
      DataPath_RF_bus_reg_dataout_1465_port, 
      DataPath_RF_bus_reg_dataout_1466_port, 
      DataPath_RF_bus_reg_dataout_1467_port, 
      DataPath_RF_bus_reg_dataout_1468_port, 
      DataPath_RF_bus_reg_dataout_1469_port, 
      DataPath_RF_bus_reg_dataout_1470_port, 
      DataPath_RF_bus_reg_dataout_1471_port, 
      DataPath_RF_bus_reg_dataout_1472_port, 
      DataPath_RF_bus_reg_dataout_1473_port, 
      DataPath_RF_bus_reg_dataout_1474_port, 
      DataPath_RF_bus_reg_dataout_1475_port, 
      DataPath_RF_bus_reg_dataout_1476_port, 
      DataPath_RF_bus_reg_dataout_1477_port, 
      DataPath_RF_bus_reg_dataout_1478_port, 
      DataPath_RF_bus_reg_dataout_1479_port, 
      DataPath_RF_bus_reg_dataout_1480_port, 
      DataPath_RF_bus_reg_dataout_1481_port, 
      DataPath_RF_bus_reg_dataout_1482_port, 
      DataPath_RF_bus_reg_dataout_1483_port, 
      DataPath_RF_bus_reg_dataout_1484_port, 
      DataPath_RF_bus_reg_dataout_1485_port, 
      DataPath_RF_bus_reg_dataout_1486_port, 
      DataPath_RF_bus_reg_dataout_1487_port, 
      DataPath_RF_bus_reg_dataout_1488_port, 
      DataPath_RF_bus_reg_dataout_1489_port, 
      DataPath_RF_bus_reg_dataout_1490_port, 
      DataPath_RF_bus_reg_dataout_1491_port, 
      DataPath_RF_bus_reg_dataout_1492_port, 
      DataPath_RF_bus_reg_dataout_1493_port, 
      DataPath_RF_bus_reg_dataout_1494_port, 
      DataPath_RF_bus_reg_dataout_1495_port, 
      DataPath_RF_bus_reg_dataout_1496_port, 
      DataPath_RF_bus_reg_dataout_1497_port, 
      DataPath_RF_bus_reg_dataout_1498_port, 
      DataPath_RF_bus_reg_dataout_1499_port, 
      DataPath_RF_bus_reg_dataout_1500_port, 
      DataPath_RF_bus_reg_dataout_1501_port, 
      DataPath_RF_bus_reg_dataout_1502_port, 
      DataPath_RF_bus_reg_dataout_1503_port, 
      DataPath_RF_bus_reg_dataout_1504_port, 
      DataPath_RF_bus_reg_dataout_1505_port, 
      DataPath_RF_bus_reg_dataout_1506_port, 
      DataPath_RF_bus_reg_dataout_1507_port, 
      DataPath_RF_bus_reg_dataout_1508_port, 
      DataPath_RF_bus_reg_dataout_1509_port, 
      DataPath_RF_bus_reg_dataout_1510_port, 
      DataPath_RF_bus_reg_dataout_1511_port, 
      DataPath_RF_bus_reg_dataout_1512_port, 
      DataPath_RF_bus_reg_dataout_1513_port, 
      DataPath_RF_bus_reg_dataout_1514_port, 
      DataPath_RF_bus_reg_dataout_1515_port, 
      DataPath_RF_bus_reg_dataout_1516_port, 
      DataPath_RF_bus_reg_dataout_1517_port, 
      DataPath_RF_bus_reg_dataout_1518_port, 
      DataPath_RF_bus_reg_dataout_1519_port, 
      DataPath_RF_bus_reg_dataout_1520_port, 
      DataPath_RF_bus_reg_dataout_1521_port, 
      DataPath_RF_bus_reg_dataout_1522_port, 
      DataPath_RF_bus_reg_dataout_1523_port, 
      DataPath_RF_bus_reg_dataout_1524_port, 
      DataPath_RF_bus_reg_dataout_1525_port, 
      DataPath_RF_bus_reg_dataout_1526_port, 
      DataPath_RF_bus_reg_dataout_1527_port, 
      DataPath_RF_bus_reg_dataout_1528_port, 
      DataPath_RF_bus_reg_dataout_1529_port, 
      DataPath_RF_bus_reg_dataout_1530_port, 
      DataPath_RF_bus_reg_dataout_1531_port, 
      DataPath_RF_bus_reg_dataout_1532_port, 
      DataPath_RF_bus_reg_dataout_1533_port, 
      DataPath_RF_bus_reg_dataout_1534_port, 
      DataPath_RF_bus_reg_dataout_1535_port, 
      DataPath_RF_bus_reg_dataout_1536_port, 
      DataPath_RF_bus_reg_dataout_1537_port, 
      DataPath_RF_bus_reg_dataout_1538_port, 
      DataPath_RF_bus_reg_dataout_1539_port, 
      DataPath_RF_bus_reg_dataout_1540_port, 
      DataPath_RF_bus_reg_dataout_1541_port, 
      DataPath_RF_bus_reg_dataout_1542_port, 
      DataPath_RF_bus_reg_dataout_1543_port, 
      DataPath_RF_bus_reg_dataout_1544_port, 
      DataPath_RF_bus_reg_dataout_1545_port, 
      DataPath_RF_bus_reg_dataout_1546_port, 
      DataPath_RF_bus_reg_dataout_1547_port, 
      DataPath_RF_bus_reg_dataout_1548_port, 
      DataPath_RF_bus_reg_dataout_1549_port, 
      DataPath_RF_bus_reg_dataout_1550_port, 
      DataPath_RF_bus_reg_dataout_1551_port, 
      DataPath_RF_bus_reg_dataout_1552_port, 
      DataPath_RF_bus_reg_dataout_1553_port, 
      DataPath_RF_bus_reg_dataout_1554_port, 
      DataPath_RF_bus_reg_dataout_1555_port, 
      DataPath_RF_bus_reg_dataout_1556_port, 
      DataPath_RF_bus_reg_dataout_1557_port, 
      DataPath_RF_bus_reg_dataout_1558_port, 
      DataPath_RF_bus_reg_dataout_1559_port, 
      DataPath_RF_bus_reg_dataout_1560_port, 
      DataPath_RF_bus_reg_dataout_1561_port, 
      DataPath_RF_bus_reg_dataout_1562_port, 
      DataPath_RF_bus_reg_dataout_1563_port, 
      DataPath_RF_bus_reg_dataout_1564_port, 
      DataPath_RF_bus_reg_dataout_1565_port, 
      DataPath_RF_bus_reg_dataout_1566_port, 
      DataPath_RF_bus_reg_dataout_1567_port, 
      DataPath_RF_bus_reg_dataout_1568_port, 
      DataPath_RF_bus_reg_dataout_1569_port, 
      DataPath_RF_bus_reg_dataout_1570_port, 
      DataPath_RF_bus_reg_dataout_1571_port, 
      DataPath_RF_bus_reg_dataout_1572_port, 
      DataPath_RF_bus_reg_dataout_1573_port, 
      DataPath_RF_bus_reg_dataout_1574_port, 
      DataPath_RF_bus_reg_dataout_1575_port, 
      DataPath_RF_bus_reg_dataout_1576_port, 
      DataPath_RF_bus_reg_dataout_1577_port, 
      DataPath_RF_bus_reg_dataout_1578_port, 
      DataPath_RF_bus_reg_dataout_1579_port, 
      DataPath_RF_bus_reg_dataout_1580_port, 
      DataPath_RF_bus_reg_dataout_1581_port, 
      DataPath_RF_bus_reg_dataout_1582_port, 
      DataPath_RF_bus_reg_dataout_1583_port, 
      DataPath_RF_bus_reg_dataout_1584_port, 
      DataPath_RF_bus_reg_dataout_1585_port, 
      DataPath_RF_bus_reg_dataout_1586_port, 
      DataPath_RF_bus_reg_dataout_1587_port, 
      DataPath_RF_bus_reg_dataout_1588_port, 
      DataPath_RF_bus_reg_dataout_1589_port, 
      DataPath_RF_bus_reg_dataout_1590_port, 
      DataPath_RF_bus_reg_dataout_1591_port, 
      DataPath_RF_bus_reg_dataout_1592_port, 
      DataPath_RF_bus_reg_dataout_1593_port, 
      DataPath_RF_bus_reg_dataout_1594_port, 
      DataPath_RF_bus_reg_dataout_1595_port, 
      DataPath_RF_bus_reg_dataout_1596_port, 
      DataPath_RF_bus_reg_dataout_1597_port, 
      DataPath_RF_bus_reg_dataout_1598_port, 
      DataPath_RF_bus_reg_dataout_1599_port, 
      DataPath_RF_bus_reg_dataout_1600_port, 
      DataPath_RF_bus_reg_dataout_1601_port, 
      DataPath_RF_bus_reg_dataout_1602_port, 
      DataPath_RF_bus_reg_dataout_1603_port, 
      DataPath_RF_bus_reg_dataout_1604_port, 
      DataPath_RF_bus_reg_dataout_1605_port, 
      DataPath_RF_bus_reg_dataout_1606_port, 
      DataPath_RF_bus_reg_dataout_1607_port, 
      DataPath_RF_bus_reg_dataout_1608_port, 
      DataPath_RF_bus_reg_dataout_1609_port, 
      DataPath_RF_bus_reg_dataout_1610_port, 
      DataPath_RF_bus_reg_dataout_1611_port, 
      DataPath_RF_bus_reg_dataout_1612_port, 
      DataPath_RF_bus_reg_dataout_1613_port, 
      DataPath_RF_bus_reg_dataout_1614_port, 
      DataPath_RF_bus_reg_dataout_1615_port, 
      DataPath_RF_bus_reg_dataout_1616_port, 
      DataPath_RF_bus_reg_dataout_1617_port, 
      DataPath_RF_bus_reg_dataout_1618_port, 
      DataPath_RF_bus_reg_dataout_1619_port, 
      DataPath_RF_bus_reg_dataout_1620_port, 
      DataPath_RF_bus_reg_dataout_1621_port, 
      DataPath_RF_bus_reg_dataout_1622_port, 
      DataPath_RF_bus_reg_dataout_1623_port, 
      DataPath_RF_bus_reg_dataout_1624_port, 
      DataPath_RF_bus_reg_dataout_1625_port, 
      DataPath_RF_bus_reg_dataout_1626_port, 
      DataPath_RF_bus_reg_dataout_1627_port, 
      DataPath_RF_bus_reg_dataout_1628_port, 
      DataPath_RF_bus_reg_dataout_1629_port, 
      DataPath_RF_bus_reg_dataout_1630_port, 
      DataPath_RF_bus_reg_dataout_1631_port, 
      DataPath_RF_bus_reg_dataout_1632_port, 
      DataPath_RF_bus_reg_dataout_1633_port, 
      DataPath_RF_bus_reg_dataout_1634_port, 
      DataPath_RF_bus_reg_dataout_1635_port, 
      DataPath_RF_bus_reg_dataout_1636_port, 
      DataPath_RF_bus_reg_dataout_1637_port, 
      DataPath_RF_bus_reg_dataout_1638_port, 
      DataPath_RF_bus_reg_dataout_1639_port, 
      DataPath_RF_bus_reg_dataout_1640_port, 
      DataPath_RF_bus_reg_dataout_1641_port, 
      DataPath_RF_bus_reg_dataout_1642_port, 
      DataPath_RF_bus_reg_dataout_1643_port, 
      DataPath_RF_bus_reg_dataout_1644_port, 
      DataPath_RF_bus_reg_dataout_1645_port, 
      DataPath_RF_bus_reg_dataout_1646_port, 
      DataPath_RF_bus_reg_dataout_1647_port, 
      DataPath_RF_bus_reg_dataout_1648_port, 
      DataPath_RF_bus_reg_dataout_1649_port, 
      DataPath_RF_bus_reg_dataout_1650_port, 
      DataPath_RF_bus_reg_dataout_1651_port, 
      DataPath_RF_bus_reg_dataout_1652_port, 
      DataPath_RF_bus_reg_dataout_1653_port, 
      DataPath_RF_bus_reg_dataout_1654_port, 
      DataPath_RF_bus_reg_dataout_1655_port, 
      DataPath_RF_bus_reg_dataout_1656_port, 
      DataPath_RF_bus_reg_dataout_1657_port, 
      DataPath_RF_bus_reg_dataout_1658_port, 
      DataPath_RF_bus_reg_dataout_1659_port, 
      DataPath_RF_bus_reg_dataout_1660_port, 
      DataPath_RF_bus_reg_dataout_1661_port, 
      DataPath_RF_bus_reg_dataout_1662_port, 
      DataPath_RF_bus_reg_dataout_1663_port, 
      DataPath_RF_bus_reg_dataout_1664_port, 
      DataPath_RF_bus_reg_dataout_1665_port, 
      DataPath_RF_bus_reg_dataout_1666_port, 
      DataPath_RF_bus_reg_dataout_1667_port, 
      DataPath_RF_bus_reg_dataout_1668_port, 
      DataPath_RF_bus_reg_dataout_1669_port, 
      DataPath_RF_bus_reg_dataout_1670_port, 
      DataPath_RF_bus_reg_dataout_1671_port, 
      DataPath_RF_bus_reg_dataout_1672_port, 
      DataPath_RF_bus_reg_dataout_1673_port, 
      DataPath_RF_bus_reg_dataout_1674_port, 
      DataPath_RF_bus_reg_dataout_1675_port, 
      DataPath_RF_bus_reg_dataout_1676_port, 
      DataPath_RF_bus_reg_dataout_1677_port, 
      DataPath_RF_bus_reg_dataout_1678_port, 
      DataPath_RF_bus_reg_dataout_1679_port, 
      DataPath_RF_bus_reg_dataout_1680_port, 
      DataPath_RF_bus_reg_dataout_1681_port, 
      DataPath_RF_bus_reg_dataout_1682_port, 
      DataPath_RF_bus_reg_dataout_1683_port, 
      DataPath_RF_bus_reg_dataout_1684_port, 
      DataPath_RF_bus_reg_dataout_1685_port, 
      DataPath_RF_bus_reg_dataout_1686_port, 
      DataPath_RF_bus_reg_dataout_1687_port, 
      DataPath_RF_bus_reg_dataout_1688_port, 
      DataPath_RF_bus_reg_dataout_1689_port, 
      DataPath_RF_bus_reg_dataout_1690_port, 
      DataPath_RF_bus_reg_dataout_1691_port, 
      DataPath_RF_bus_reg_dataout_1692_port, 
      DataPath_RF_bus_reg_dataout_1693_port, 
      DataPath_RF_bus_reg_dataout_1694_port, 
      DataPath_RF_bus_reg_dataout_1695_port, 
      DataPath_RF_bus_reg_dataout_1696_port, 
      DataPath_RF_bus_reg_dataout_1697_port, 
      DataPath_RF_bus_reg_dataout_1698_port, 
      DataPath_RF_bus_reg_dataout_1699_port, 
      DataPath_RF_bus_reg_dataout_1700_port, 
      DataPath_RF_bus_reg_dataout_1701_port, 
      DataPath_RF_bus_reg_dataout_1702_port, 
      DataPath_RF_bus_reg_dataout_1703_port, 
      DataPath_RF_bus_reg_dataout_1704_port, 
      DataPath_RF_bus_reg_dataout_1705_port, 
      DataPath_RF_bus_reg_dataout_1706_port, 
      DataPath_RF_bus_reg_dataout_1707_port, 
      DataPath_RF_bus_reg_dataout_1708_port, 
      DataPath_RF_bus_reg_dataout_1709_port, 
      DataPath_RF_bus_reg_dataout_1710_port, 
      DataPath_RF_bus_reg_dataout_1711_port, 
      DataPath_RF_bus_reg_dataout_1712_port, 
      DataPath_RF_bus_reg_dataout_1713_port, 
      DataPath_RF_bus_reg_dataout_1714_port, 
      DataPath_RF_bus_reg_dataout_1715_port, 
      DataPath_RF_bus_reg_dataout_1716_port, 
      DataPath_RF_bus_reg_dataout_1717_port, 
      DataPath_RF_bus_reg_dataout_1718_port, 
      DataPath_RF_bus_reg_dataout_1719_port, 
      DataPath_RF_bus_reg_dataout_1720_port, 
      DataPath_RF_bus_reg_dataout_1721_port, 
      DataPath_RF_bus_reg_dataout_1722_port, 
      DataPath_RF_bus_reg_dataout_1723_port, 
      DataPath_RF_bus_reg_dataout_1724_port, 
      DataPath_RF_bus_reg_dataout_1725_port, 
      DataPath_RF_bus_reg_dataout_1726_port, 
      DataPath_RF_bus_reg_dataout_1727_port, 
      DataPath_RF_bus_reg_dataout_1728_port, 
      DataPath_RF_bus_reg_dataout_1729_port, 
      DataPath_RF_bus_reg_dataout_1730_port, 
      DataPath_RF_bus_reg_dataout_1731_port, 
      DataPath_RF_bus_reg_dataout_1732_port, 
      DataPath_RF_bus_reg_dataout_1733_port, 
      DataPath_RF_bus_reg_dataout_1734_port, 
      DataPath_RF_bus_reg_dataout_1735_port, 
      DataPath_RF_bus_reg_dataout_1736_port, 
      DataPath_RF_bus_reg_dataout_1737_port, 
      DataPath_RF_bus_reg_dataout_1738_port, 
      DataPath_RF_bus_reg_dataout_1739_port, 
      DataPath_RF_bus_reg_dataout_1740_port, 
      DataPath_RF_bus_reg_dataout_1741_port, 
      DataPath_RF_bus_reg_dataout_1742_port, 
      DataPath_RF_bus_reg_dataout_1743_port, 
      DataPath_RF_bus_reg_dataout_1744_port, 
      DataPath_RF_bus_reg_dataout_1745_port, 
      DataPath_RF_bus_reg_dataout_1746_port, 
      DataPath_RF_bus_reg_dataout_1747_port, 
      DataPath_RF_bus_reg_dataout_1748_port, 
      DataPath_RF_bus_reg_dataout_1749_port, 
      DataPath_RF_bus_reg_dataout_1750_port, 
      DataPath_RF_bus_reg_dataout_1751_port, 
      DataPath_RF_bus_reg_dataout_1752_port, 
      DataPath_RF_bus_reg_dataout_1753_port, 
      DataPath_RF_bus_reg_dataout_1754_port, 
      DataPath_RF_bus_reg_dataout_1755_port, 
      DataPath_RF_bus_reg_dataout_1756_port, 
      DataPath_RF_bus_reg_dataout_1757_port, 
      DataPath_RF_bus_reg_dataout_1758_port, 
      DataPath_RF_bus_reg_dataout_1759_port, 
      DataPath_RF_bus_reg_dataout_1760_port, 
      DataPath_RF_bus_reg_dataout_1761_port, 
      DataPath_RF_bus_reg_dataout_1762_port, 
      DataPath_RF_bus_reg_dataout_1763_port, 
      DataPath_RF_bus_reg_dataout_1764_port, 
      DataPath_RF_bus_reg_dataout_1765_port, 
      DataPath_RF_bus_reg_dataout_1766_port, 
      DataPath_RF_bus_reg_dataout_1767_port, 
      DataPath_RF_bus_reg_dataout_1768_port, 
      DataPath_RF_bus_reg_dataout_1769_port, 
      DataPath_RF_bus_reg_dataout_1770_port, 
      DataPath_RF_bus_reg_dataout_1771_port, 
      DataPath_RF_bus_reg_dataout_1772_port, 
      DataPath_RF_bus_reg_dataout_1773_port, 
      DataPath_RF_bus_reg_dataout_1774_port, 
      DataPath_RF_bus_reg_dataout_1775_port, 
      DataPath_RF_bus_reg_dataout_1776_port, 
      DataPath_RF_bus_reg_dataout_1777_port, 
      DataPath_RF_bus_reg_dataout_1778_port, 
      DataPath_RF_bus_reg_dataout_1779_port, 
      DataPath_RF_bus_reg_dataout_1780_port, 
      DataPath_RF_bus_reg_dataout_1781_port, 
      DataPath_RF_bus_reg_dataout_1782_port, 
      DataPath_RF_bus_reg_dataout_1783_port, 
      DataPath_RF_bus_reg_dataout_1784_port, 
      DataPath_RF_bus_reg_dataout_1785_port, 
      DataPath_RF_bus_reg_dataout_1786_port, 
      DataPath_RF_bus_reg_dataout_1787_port, 
      DataPath_RF_bus_reg_dataout_1788_port, 
      DataPath_RF_bus_reg_dataout_1789_port, 
      DataPath_RF_bus_reg_dataout_1790_port, 
      DataPath_RF_bus_reg_dataout_1791_port, 
      DataPath_RF_bus_reg_dataout_1792_port, 
      DataPath_RF_bus_reg_dataout_1793_port, 
      DataPath_RF_bus_reg_dataout_1794_port, 
      DataPath_RF_bus_reg_dataout_1795_port, 
      DataPath_RF_bus_reg_dataout_1796_port, 
      DataPath_RF_bus_reg_dataout_1797_port, 
      DataPath_RF_bus_reg_dataout_1798_port, 
      DataPath_RF_bus_reg_dataout_1799_port, 
      DataPath_RF_bus_reg_dataout_1800_port, 
      DataPath_RF_bus_reg_dataout_1801_port, 
      DataPath_RF_bus_reg_dataout_1802_port, 
      DataPath_RF_bus_reg_dataout_1803_port, 
      DataPath_RF_bus_reg_dataout_1804_port, 
      DataPath_RF_bus_reg_dataout_1805_port, 
      DataPath_RF_bus_reg_dataout_1806_port, 
      DataPath_RF_bus_reg_dataout_1807_port, 
      DataPath_RF_bus_reg_dataout_1808_port, 
      DataPath_RF_bus_reg_dataout_1809_port, 
      DataPath_RF_bus_reg_dataout_1810_port, 
      DataPath_RF_bus_reg_dataout_1811_port, 
      DataPath_RF_bus_reg_dataout_1812_port, 
      DataPath_RF_bus_reg_dataout_1813_port, 
      DataPath_RF_bus_reg_dataout_1814_port, 
      DataPath_RF_bus_reg_dataout_1815_port, 
      DataPath_RF_bus_reg_dataout_1816_port, 
      DataPath_RF_bus_reg_dataout_1817_port, 
      DataPath_RF_bus_reg_dataout_1818_port, 
      DataPath_RF_bus_reg_dataout_1819_port, 
      DataPath_RF_bus_reg_dataout_1820_port, 
      DataPath_RF_bus_reg_dataout_1821_port, 
      DataPath_RF_bus_reg_dataout_1822_port, 
      DataPath_RF_bus_reg_dataout_1823_port, 
      DataPath_RF_bus_reg_dataout_1824_port, 
      DataPath_RF_bus_reg_dataout_1825_port, 
      DataPath_RF_bus_reg_dataout_1826_port, 
      DataPath_RF_bus_reg_dataout_1827_port, 
      DataPath_RF_bus_reg_dataout_1828_port, 
      DataPath_RF_bus_reg_dataout_1829_port, 
      DataPath_RF_bus_reg_dataout_1830_port, 
      DataPath_RF_bus_reg_dataout_1831_port, 
      DataPath_RF_bus_reg_dataout_1832_port, 
      DataPath_RF_bus_reg_dataout_1833_port, 
      DataPath_RF_bus_reg_dataout_1834_port, 
      DataPath_RF_bus_reg_dataout_1835_port, 
      DataPath_RF_bus_reg_dataout_1836_port, 
      DataPath_RF_bus_reg_dataout_1837_port, 
      DataPath_RF_bus_reg_dataout_1838_port, 
      DataPath_RF_bus_reg_dataout_1839_port, 
      DataPath_RF_bus_reg_dataout_1840_port, 
      DataPath_RF_bus_reg_dataout_1841_port, 
      DataPath_RF_bus_reg_dataout_1842_port, 
      DataPath_RF_bus_reg_dataout_1843_port, 
      DataPath_RF_bus_reg_dataout_1844_port, 
      DataPath_RF_bus_reg_dataout_1845_port, 
      DataPath_RF_bus_reg_dataout_1846_port, 
      DataPath_RF_bus_reg_dataout_1847_port, 
      DataPath_RF_bus_reg_dataout_1848_port, 
      DataPath_RF_bus_reg_dataout_1849_port, 
      DataPath_RF_bus_reg_dataout_1850_port, 
      DataPath_RF_bus_reg_dataout_1851_port, 
      DataPath_RF_bus_reg_dataout_1852_port, 
      DataPath_RF_bus_reg_dataout_1853_port, 
      DataPath_RF_bus_reg_dataout_1854_port, 
      DataPath_RF_bus_reg_dataout_1855_port, 
      DataPath_RF_bus_reg_dataout_1856_port, 
      DataPath_RF_bus_reg_dataout_1857_port, 
      DataPath_RF_bus_reg_dataout_1858_port, 
      DataPath_RF_bus_reg_dataout_1859_port, 
      DataPath_RF_bus_reg_dataout_1860_port, 
      DataPath_RF_bus_reg_dataout_1861_port, 
      DataPath_RF_bus_reg_dataout_1862_port, 
      DataPath_RF_bus_reg_dataout_1863_port, 
      DataPath_RF_bus_reg_dataout_1864_port, 
      DataPath_RF_bus_reg_dataout_1865_port, 
      DataPath_RF_bus_reg_dataout_1866_port, 
      DataPath_RF_bus_reg_dataout_1867_port, 
      DataPath_RF_bus_reg_dataout_1868_port, 
      DataPath_RF_bus_reg_dataout_1869_port, 
      DataPath_RF_bus_reg_dataout_1870_port, 
      DataPath_RF_bus_reg_dataout_1871_port, 
      DataPath_RF_bus_reg_dataout_1872_port, 
      DataPath_RF_bus_reg_dataout_1873_port, 
      DataPath_RF_bus_reg_dataout_1874_port, 
      DataPath_RF_bus_reg_dataout_1875_port, 
      DataPath_RF_bus_reg_dataout_1876_port, 
      DataPath_RF_bus_reg_dataout_1877_port, 
      DataPath_RF_bus_reg_dataout_1878_port, 
      DataPath_RF_bus_reg_dataout_1879_port, 
      DataPath_RF_bus_reg_dataout_1880_port, 
      DataPath_RF_bus_reg_dataout_1881_port, 
      DataPath_RF_bus_reg_dataout_1882_port, 
      DataPath_RF_bus_reg_dataout_1883_port, 
      DataPath_RF_bus_reg_dataout_1884_port, 
      DataPath_RF_bus_reg_dataout_1885_port, 
      DataPath_RF_bus_reg_dataout_1886_port, 
      DataPath_RF_bus_reg_dataout_1887_port, 
      DataPath_RF_bus_reg_dataout_1888_port, 
      DataPath_RF_bus_reg_dataout_1889_port, 
      DataPath_RF_bus_reg_dataout_1890_port, 
      DataPath_RF_bus_reg_dataout_1891_port, 
      DataPath_RF_bus_reg_dataout_1892_port, 
      DataPath_RF_bus_reg_dataout_1893_port, 
      DataPath_RF_bus_reg_dataout_1894_port, 
      DataPath_RF_bus_reg_dataout_1895_port, 
      DataPath_RF_bus_reg_dataout_1896_port, 
      DataPath_RF_bus_reg_dataout_1897_port, 
      DataPath_RF_bus_reg_dataout_1898_port, 
      DataPath_RF_bus_reg_dataout_1899_port, 
      DataPath_RF_bus_reg_dataout_1900_port, 
      DataPath_RF_bus_reg_dataout_1901_port, 
      DataPath_RF_bus_reg_dataout_1902_port, 
      DataPath_RF_bus_reg_dataout_1903_port, 
      DataPath_RF_bus_reg_dataout_1904_port, 
      DataPath_RF_bus_reg_dataout_1905_port, 
      DataPath_RF_bus_reg_dataout_1906_port, 
      DataPath_RF_bus_reg_dataout_1907_port, 
      DataPath_RF_bus_reg_dataout_1908_port, 
      DataPath_RF_bus_reg_dataout_1909_port, 
      DataPath_RF_bus_reg_dataout_1910_port, 
      DataPath_RF_bus_reg_dataout_1911_port, 
      DataPath_RF_bus_reg_dataout_1912_port, 
      DataPath_RF_bus_reg_dataout_1913_port, 
      DataPath_RF_bus_reg_dataout_1914_port, 
      DataPath_RF_bus_reg_dataout_1915_port, 
      DataPath_RF_bus_reg_dataout_1916_port, 
      DataPath_RF_bus_reg_dataout_1917_port, 
      DataPath_RF_bus_reg_dataout_1918_port, 
      DataPath_RF_bus_reg_dataout_1919_port, 
      DataPath_RF_bus_reg_dataout_1920_port, 
      DataPath_RF_bus_reg_dataout_1921_port, 
      DataPath_RF_bus_reg_dataout_1922_port, 
      DataPath_RF_bus_reg_dataout_1923_port, 
      DataPath_RF_bus_reg_dataout_1924_port, 
      DataPath_RF_bus_reg_dataout_1925_port, 
      DataPath_RF_bus_reg_dataout_1926_port, 
      DataPath_RF_bus_reg_dataout_1927_port, 
      DataPath_RF_bus_reg_dataout_1928_port, 
      DataPath_RF_bus_reg_dataout_1929_port, 
      DataPath_RF_bus_reg_dataout_1930_port, 
      DataPath_RF_bus_reg_dataout_1931_port, 
      DataPath_RF_bus_reg_dataout_1932_port, 
      DataPath_RF_bus_reg_dataout_1933_port, 
      DataPath_RF_bus_reg_dataout_1934_port, 
      DataPath_RF_bus_reg_dataout_1935_port, 
      DataPath_RF_bus_reg_dataout_1936_port, 
      DataPath_RF_bus_reg_dataout_1937_port, 
      DataPath_RF_bus_reg_dataout_1938_port, 
      DataPath_RF_bus_reg_dataout_1939_port, 
      DataPath_RF_bus_reg_dataout_1940_port, 
      DataPath_RF_bus_reg_dataout_1941_port, 
      DataPath_RF_bus_reg_dataout_1942_port, 
      DataPath_RF_bus_reg_dataout_1943_port, 
      DataPath_RF_bus_reg_dataout_1944_port, 
      DataPath_RF_bus_reg_dataout_1945_port, 
      DataPath_RF_bus_reg_dataout_1946_port, 
      DataPath_RF_bus_reg_dataout_1947_port, 
      DataPath_RF_bus_reg_dataout_1948_port, 
      DataPath_RF_bus_reg_dataout_1949_port, 
      DataPath_RF_bus_reg_dataout_1950_port, 
      DataPath_RF_bus_reg_dataout_1951_port, 
      DataPath_RF_bus_reg_dataout_1952_port, 
      DataPath_RF_bus_reg_dataout_1953_port, 
      DataPath_RF_bus_reg_dataout_1954_port, 
      DataPath_RF_bus_reg_dataout_1955_port, 
      DataPath_RF_bus_reg_dataout_1956_port, 
      DataPath_RF_bus_reg_dataout_1957_port, 
      DataPath_RF_bus_reg_dataout_1958_port, 
      DataPath_RF_bus_reg_dataout_1959_port, 
      DataPath_RF_bus_reg_dataout_1960_port, 
      DataPath_RF_bus_reg_dataout_1961_port, 
      DataPath_RF_bus_reg_dataout_1962_port, 
      DataPath_RF_bus_reg_dataout_1963_port, 
      DataPath_RF_bus_reg_dataout_1964_port, 
      DataPath_RF_bus_reg_dataout_1965_port, 
      DataPath_RF_bus_reg_dataout_1966_port, 
      DataPath_RF_bus_reg_dataout_1967_port, 
      DataPath_RF_bus_reg_dataout_1968_port, 
      DataPath_RF_bus_reg_dataout_1969_port, 
      DataPath_RF_bus_reg_dataout_1970_port, 
      DataPath_RF_bus_reg_dataout_1971_port, 
      DataPath_RF_bus_reg_dataout_1972_port, 
      DataPath_RF_bus_reg_dataout_1973_port, 
      DataPath_RF_bus_reg_dataout_1974_port, 
      DataPath_RF_bus_reg_dataout_1975_port, 
      DataPath_RF_bus_reg_dataout_1976_port, 
      DataPath_RF_bus_reg_dataout_1977_port, 
      DataPath_RF_bus_reg_dataout_1978_port, 
      DataPath_RF_bus_reg_dataout_1979_port, 
      DataPath_RF_bus_reg_dataout_1980_port, 
      DataPath_RF_bus_reg_dataout_1981_port, 
      DataPath_RF_bus_reg_dataout_1982_port, 
      DataPath_RF_bus_reg_dataout_1983_port, 
      DataPath_RF_bus_reg_dataout_1984_port, 
      DataPath_RF_bus_reg_dataout_1985_port, 
      DataPath_RF_bus_reg_dataout_1986_port, 
      DataPath_RF_bus_reg_dataout_1987_port, 
      DataPath_RF_bus_reg_dataout_1988_port, 
      DataPath_RF_bus_reg_dataout_1989_port, 
      DataPath_RF_bus_reg_dataout_1990_port, 
      DataPath_RF_bus_reg_dataout_1991_port, 
      DataPath_RF_bus_reg_dataout_1992_port, 
      DataPath_RF_bus_reg_dataout_1993_port, 
      DataPath_RF_bus_reg_dataout_1994_port, 
      DataPath_RF_bus_reg_dataout_1995_port, 
      DataPath_RF_bus_reg_dataout_1996_port, 
      DataPath_RF_bus_reg_dataout_1997_port, 
      DataPath_RF_bus_reg_dataout_1998_port, 
      DataPath_RF_bus_reg_dataout_1999_port, 
      DataPath_RF_bus_reg_dataout_2000_port, 
      DataPath_RF_bus_reg_dataout_2001_port, 
      DataPath_RF_bus_reg_dataout_2002_port, 
      DataPath_RF_bus_reg_dataout_2003_port, 
      DataPath_RF_bus_reg_dataout_2004_port, 
      DataPath_RF_bus_reg_dataout_2005_port, 
      DataPath_RF_bus_reg_dataout_2006_port, 
      DataPath_RF_bus_reg_dataout_2007_port, 
      DataPath_RF_bus_reg_dataout_2008_port, 
      DataPath_RF_bus_reg_dataout_2009_port, 
      DataPath_RF_bus_reg_dataout_2010_port, 
      DataPath_RF_bus_reg_dataout_2011_port, 
      DataPath_RF_bus_reg_dataout_2012_port, 
      DataPath_RF_bus_reg_dataout_2013_port, 
      DataPath_RF_bus_reg_dataout_2014_port, 
      DataPath_RF_bus_reg_dataout_2015_port, 
      DataPath_RF_bus_reg_dataout_2016_port, 
      DataPath_RF_bus_reg_dataout_2017_port, 
      DataPath_RF_bus_reg_dataout_2018_port, 
      DataPath_RF_bus_reg_dataout_2019_port, 
      DataPath_RF_bus_reg_dataout_2020_port, 
      DataPath_RF_bus_reg_dataout_2021_port, 
      DataPath_RF_bus_reg_dataout_2022_port, 
      DataPath_RF_bus_reg_dataout_2023_port, 
      DataPath_RF_bus_reg_dataout_2024_port, 
      DataPath_RF_bus_reg_dataout_2025_port, 
      DataPath_RF_bus_reg_dataout_2026_port, 
      DataPath_RF_bus_reg_dataout_2027_port, 
      DataPath_RF_bus_reg_dataout_2028_port, 
      DataPath_RF_bus_reg_dataout_2029_port, 
      DataPath_RF_bus_reg_dataout_2030_port, 
      DataPath_RF_bus_reg_dataout_2031_port, 
      DataPath_RF_bus_reg_dataout_2032_port, 
      DataPath_RF_bus_reg_dataout_2033_port, 
      DataPath_RF_bus_reg_dataout_2034_port, 
      DataPath_RF_bus_reg_dataout_2035_port, 
      DataPath_RF_bus_reg_dataout_2036_port, 
      DataPath_RF_bus_reg_dataout_2037_port, 
      DataPath_RF_bus_reg_dataout_2038_port, 
      DataPath_RF_bus_reg_dataout_2039_port, 
      DataPath_RF_bus_reg_dataout_2040_port, 
      DataPath_RF_bus_reg_dataout_2041_port, 
      DataPath_RF_bus_reg_dataout_2042_port, 
      DataPath_RF_bus_reg_dataout_2043_port, 
      DataPath_RF_bus_reg_dataout_2044_port, 
      DataPath_RF_bus_reg_dataout_2045_port, 
      DataPath_RF_bus_reg_dataout_2046_port, 
      DataPath_RF_bus_reg_dataout_2047_port, 
      DataPath_RF_bus_reg_dataout_2048_port, 
      DataPath_RF_bus_reg_dataout_2049_port, 
      DataPath_RF_bus_reg_dataout_2050_port, 
      DataPath_RF_bus_reg_dataout_2051_port, 
      DataPath_RF_bus_reg_dataout_2052_port, 
      DataPath_RF_bus_reg_dataout_2053_port, 
      DataPath_RF_bus_reg_dataout_2054_port, 
      DataPath_RF_bus_reg_dataout_2055_port, 
      DataPath_RF_bus_reg_dataout_2056_port, 
      DataPath_RF_bus_reg_dataout_2057_port, 
      DataPath_RF_bus_reg_dataout_2058_port, 
      DataPath_RF_bus_reg_dataout_2059_port, 
      DataPath_RF_bus_reg_dataout_2060_port, 
      DataPath_RF_bus_reg_dataout_2061_port, 
      DataPath_RF_bus_reg_dataout_2062_port, 
      DataPath_RF_bus_reg_dataout_2063_port, 
      DataPath_RF_bus_reg_dataout_2064_port, 
      DataPath_RF_bus_reg_dataout_2065_port, 
      DataPath_RF_bus_reg_dataout_2066_port, 
      DataPath_RF_bus_reg_dataout_2067_port, 
      DataPath_RF_bus_reg_dataout_2068_port, 
      DataPath_RF_bus_reg_dataout_2069_port, 
      DataPath_RF_bus_reg_dataout_2070_port, 
      DataPath_RF_bus_reg_dataout_2071_port, 
      DataPath_RF_bus_reg_dataout_2072_port, 
      DataPath_RF_bus_reg_dataout_2073_port, 
      DataPath_RF_bus_reg_dataout_2074_port, 
      DataPath_RF_bus_reg_dataout_2075_port, 
      DataPath_RF_bus_reg_dataout_2076_port, 
      DataPath_RF_bus_reg_dataout_2077_port, 
      DataPath_RF_bus_reg_dataout_2078_port, 
      DataPath_RF_bus_reg_dataout_2079_port, 
      DataPath_RF_bus_reg_dataout_2080_port, 
      DataPath_RF_bus_reg_dataout_2081_port, 
      DataPath_RF_bus_reg_dataout_2082_port, 
      DataPath_RF_bus_reg_dataout_2083_port, 
      DataPath_RF_bus_reg_dataout_2084_port, 
      DataPath_RF_bus_reg_dataout_2085_port, 
      DataPath_RF_bus_reg_dataout_2086_port, 
      DataPath_RF_bus_reg_dataout_2087_port, 
      DataPath_RF_bus_reg_dataout_2088_port, 
      DataPath_RF_bus_reg_dataout_2089_port, 
      DataPath_RF_bus_reg_dataout_2090_port, 
      DataPath_RF_bus_reg_dataout_2091_port, 
      DataPath_RF_bus_reg_dataout_2092_port, 
      DataPath_RF_bus_reg_dataout_2093_port, 
      DataPath_RF_bus_reg_dataout_2094_port, 
      DataPath_RF_bus_reg_dataout_2095_port, 
      DataPath_RF_bus_reg_dataout_2096_port, 
      DataPath_RF_bus_reg_dataout_2097_port, 
      DataPath_RF_bus_reg_dataout_2098_port, 
      DataPath_RF_bus_reg_dataout_2099_port, 
      DataPath_RF_bus_reg_dataout_2100_port, 
      DataPath_RF_bus_reg_dataout_2101_port, 
      DataPath_RF_bus_reg_dataout_2102_port, 
      DataPath_RF_bus_reg_dataout_2103_port, 
      DataPath_RF_bus_reg_dataout_2104_port, 
      DataPath_RF_bus_reg_dataout_2105_port, 
      DataPath_RF_bus_reg_dataout_2106_port, 
      DataPath_RF_bus_reg_dataout_2107_port, 
      DataPath_RF_bus_reg_dataout_2108_port, 
      DataPath_RF_bus_reg_dataout_2109_port, 
      DataPath_RF_bus_reg_dataout_2110_port, 
      DataPath_RF_bus_reg_dataout_2111_port, 
      DataPath_RF_bus_reg_dataout_2112_port, 
      DataPath_RF_bus_reg_dataout_2113_port, 
      DataPath_RF_bus_reg_dataout_2114_port, 
      DataPath_RF_bus_reg_dataout_2115_port, 
      DataPath_RF_bus_reg_dataout_2116_port, 
      DataPath_RF_bus_reg_dataout_2117_port, 
      DataPath_RF_bus_reg_dataout_2118_port, 
      DataPath_RF_bus_reg_dataout_2119_port, 
      DataPath_RF_bus_reg_dataout_2120_port, 
      DataPath_RF_bus_reg_dataout_2121_port, 
      DataPath_RF_bus_reg_dataout_2122_port, 
      DataPath_RF_bus_reg_dataout_2123_port, 
      DataPath_RF_bus_reg_dataout_2124_port, 
      DataPath_RF_bus_reg_dataout_2125_port, 
      DataPath_RF_bus_reg_dataout_2126_port, 
      DataPath_RF_bus_reg_dataout_2127_port, 
      DataPath_RF_bus_reg_dataout_2128_port, 
      DataPath_RF_bus_reg_dataout_2129_port, 
      DataPath_RF_bus_reg_dataout_2130_port, 
      DataPath_RF_bus_reg_dataout_2131_port, 
      DataPath_RF_bus_reg_dataout_2132_port, 
      DataPath_RF_bus_reg_dataout_2133_port, 
      DataPath_RF_bus_reg_dataout_2134_port, 
      DataPath_RF_bus_reg_dataout_2135_port, 
      DataPath_RF_bus_reg_dataout_2136_port, 
      DataPath_RF_bus_reg_dataout_2137_port, 
      DataPath_RF_bus_reg_dataout_2138_port, 
      DataPath_RF_bus_reg_dataout_2139_port, 
      DataPath_RF_bus_reg_dataout_2140_port, 
      DataPath_RF_bus_reg_dataout_2141_port, 
      DataPath_RF_bus_reg_dataout_2142_port, 
      DataPath_RF_bus_reg_dataout_2143_port, 
      DataPath_RF_bus_reg_dataout_2144_port, 
      DataPath_RF_bus_reg_dataout_2145_port, 
      DataPath_RF_bus_reg_dataout_2146_port, 
      DataPath_RF_bus_reg_dataout_2147_port, 
      DataPath_RF_bus_reg_dataout_2148_port, 
      DataPath_RF_bus_reg_dataout_2149_port, 
      DataPath_RF_bus_reg_dataout_2150_port, 
      DataPath_RF_bus_reg_dataout_2151_port, 
      DataPath_RF_bus_reg_dataout_2152_port, 
      DataPath_RF_bus_reg_dataout_2153_port, 
      DataPath_RF_bus_reg_dataout_2154_port, 
      DataPath_RF_bus_reg_dataout_2155_port, 
      DataPath_RF_bus_reg_dataout_2156_port, 
      DataPath_RF_bus_reg_dataout_2157_port, 
      DataPath_RF_bus_reg_dataout_2158_port, 
      DataPath_RF_bus_reg_dataout_2159_port, 
      DataPath_RF_bus_reg_dataout_2160_port, 
      DataPath_RF_bus_reg_dataout_2161_port, 
      DataPath_RF_bus_reg_dataout_2162_port, 
      DataPath_RF_bus_reg_dataout_2163_port, 
      DataPath_RF_bus_reg_dataout_2164_port, 
      DataPath_RF_bus_reg_dataout_2165_port, 
      DataPath_RF_bus_reg_dataout_2166_port, 
      DataPath_RF_bus_reg_dataout_2167_port, 
      DataPath_RF_bus_reg_dataout_2168_port, 
      DataPath_RF_bus_reg_dataout_2169_port, 
      DataPath_RF_bus_reg_dataout_2170_port, 
      DataPath_RF_bus_reg_dataout_2171_port, 
      DataPath_RF_bus_reg_dataout_2172_port, 
      DataPath_RF_bus_reg_dataout_2173_port, 
      DataPath_RF_bus_reg_dataout_2174_port, 
      DataPath_RF_bus_reg_dataout_2175_port, 
      DataPath_RF_bus_reg_dataout_2176_port, 
      DataPath_RF_bus_reg_dataout_2177_port, 
      DataPath_RF_bus_reg_dataout_2178_port, 
      DataPath_RF_bus_reg_dataout_2179_port, 
      DataPath_RF_bus_reg_dataout_2180_port, 
      DataPath_RF_bus_reg_dataout_2181_port, 
      DataPath_RF_bus_reg_dataout_2182_port, 
      DataPath_RF_bus_reg_dataout_2183_port, 
      DataPath_RF_bus_reg_dataout_2184_port, 
      DataPath_RF_bus_reg_dataout_2185_port, 
      DataPath_RF_bus_reg_dataout_2186_port, 
      DataPath_RF_bus_reg_dataout_2187_port, 
      DataPath_RF_bus_reg_dataout_2188_port, 
      DataPath_RF_bus_reg_dataout_2189_port, 
      DataPath_RF_bus_reg_dataout_2190_port, 
      DataPath_RF_bus_reg_dataout_2191_port, 
      DataPath_RF_bus_reg_dataout_2192_port, 
      DataPath_RF_bus_reg_dataout_2193_port, 
      DataPath_RF_bus_reg_dataout_2194_port, 
      DataPath_RF_bus_reg_dataout_2195_port, 
      DataPath_RF_bus_reg_dataout_2196_port, 
      DataPath_RF_bus_reg_dataout_2197_port, 
      DataPath_RF_bus_reg_dataout_2198_port, 
      DataPath_RF_bus_reg_dataout_2199_port, 
      DataPath_RF_bus_reg_dataout_2200_port, 
      DataPath_RF_bus_reg_dataout_2201_port, 
      DataPath_RF_bus_reg_dataout_2202_port, 
      DataPath_RF_bus_reg_dataout_2203_port, 
      DataPath_RF_bus_reg_dataout_2204_port, 
      DataPath_RF_bus_reg_dataout_2205_port, 
      DataPath_RF_bus_reg_dataout_2206_port, 
      DataPath_RF_bus_reg_dataout_2207_port, 
      DataPath_RF_bus_reg_dataout_2208_port, 
      DataPath_RF_bus_reg_dataout_2209_port, 
      DataPath_RF_bus_reg_dataout_2210_port, 
      DataPath_RF_bus_reg_dataout_2211_port, 
      DataPath_RF_bus_reg_dataout_2212_port, 
      DataPath_RF_bus_reg_dataout_2213_port, 
      DataPath_RF_bus_reg_dataout_2214_port, 
      DataPath_RF_bus_reg_dataout_2215_port, 
      DataPath_RF_bus_reg_dataout_2216_port, 
      DataPath_RF_bus_reg_dataout_2217_port, 
      DataPath_RF_bus_reg_dataout_2218_port, 
      DataPath_RF_bus_reg_dataout_2219_port, 
      DataPath_RF_bus_reg_dataout_2220_port, 
      DataPath_RF_bus_reg_dataout_2221_port, 
      DataPath_RF_bus_reg_dataout_2222_port, 
      DataPath_RF_bus_reg_dataout_2223_port, 
      DataPath_RF_bus_reg_dataout_2224_port, 
      DataPath_RF_bus_reg_dataout_2225_port, 
      DataPath_RF_bus_reg_dataout_2226_port, 
      DataPath_RF_bus_reg_dataout_2227_port, 
      DataPath_RF_bus_reg_dataout_2228_port, 
      DataPath_RF_bus_reg_dataout_2229_port, 
      DataPath_RF_bus_reg_dataout_2230_port, 
      DataPath_RF_bus_reg_dataout_2231_port, 
      DataPath_RF_bus_reg_dataout_2232_port, 
      DataPath_RF_bus_reg_dataout_2233_port, 
      DataPath_RF_bus_reg_dataout_2234_port, 
      DataPath_RF_bus_reg_dataout_2235_port, 
      DataPath_RF_bus_reg_dataout_2236_port, 
      DataPath_RF_bus_reg_dataout_2237_port, 
      DataPath_RF_bus_reg_dataout_2238_port, 
      DataPath_RF_bus_reg_dataout_2239_port, 
      DataPath_RF_bus_reg_dataout_2240_port, 
      DataPath_RF_bus_reg_dataout_2241_port, 
      DataPath_RF_bus_reg_dataout_2242_port, 
      DataPath_RF_bus_reg_dataout_2243_port, 
      DataPath_RF_bus_reg_dataout_2244_port, 
      DataPath_RF_bus_reg_dataout_2245_port, 
      DataPath_RF_bus_reg_dataout_2246_port, 
      DataPath_RF_bus_reg_dataout_2247_port, 
      DataPath_RF_bus_reg_dataout_2248_port, 
      DataPath_RF_bus_reg_dataout_2249_port, 
      DataPath_RF_bus_reg_dataout_2250_port, 
      DataPath_RF_bus_reg_dataout_2251_port, 
      DataPath_RF_bus_reg_dataout_2252_port, 
      DataPath_RF_bus_reg_dataout_2253_port, 
      DataPath_RF_bus_reg_dataout_2254_port, 
      DataPath_RF_bus_reg_dataout_2255_port, 
      DataPath_RF_bus_reg_dataout_2256_port, 
      DataPath_RF_bus_reg_dataout_2257_port, 
      DataPath_RF_bus_reg_dataout_2258_port, 
      DataPath_RF_bus_reg_dataout_2259_port, 
      DataPath_RF_bus_reg_dataout_2260_port, 
      DataPath_RF_bus_reg_dataout_2261_port, 
      DataPath_RF_bus_reg_dataout_2262_port, 
      DataPath_RF_bus_reg_dataout_2263_port, 
      DataPath_RF_bus_reg_dataout_2264_port, 
      DataPath_RF_bus_reg_dataout_2265_port, 
      DataPath_RF_bus_reg_dataout_2266_port, 
      DataPath_RF_bus_reg_dataout_2267_port, 
      DataPath_RF_bus_reg_dataout_2268_port, 
      DataPath_RF_bus_reg_dataout_2269_port, 
      DataPath_RF_bus_reg_dataout_2270_port, 
      DataPath_RF_bus_reg_dataout_2271_port, 
      DataPath_RF_bus_reg_dataout_2272_port, 
      DataPath_RF_bus_reg_dataout_2273_port, 
      DataPath_RF_bus_reg_dataout_2274_port, 
      DataPath_RF_bus_reg_dataout_2275_port, 
      DataPath_RF_bus_reg_dataout_2276_port, 
      DataPath_RF_bus_reg_dataout_2277_port, 
      DataPath_RF_bus_reg_dataout_2278_port, 
      DataPath_RF_bus_reg_dataout_2279_port, 
      DataPath_RF_bus_reg_dataout_2280_port, 
      DataPath_RF_bus_reg_dataout_2281_port, 
      DataPath_RF_bus_reg_dataout_2282_port, 
      DataPath_RF_bus_reg_dataout_2283_port, 
      DataPath_RF_bus_reg_dataout_2284_port, 
      DataPath_RF_bus_reg_dataout_2285_port, 
      DataPath_RF_bus_reg_dataout_2286_port, 
      DataPath_RF_bus_reg_dataout_2287_port, 
      DataPath_RF_bus_reg_dataout_2288_port, 
      DataPath_RF_bus_reg_dataout_2289_port, 
      DataPath_RF_bus_reg_dataout_2290_port, 
      DataPath_RF_bus_reg_dataout_2291_port, 
      DataPath_RF_bus_reg_dataout_2292_port, 
      DataPath_RF_bus_reg_dataout_2293_port, 
      DataPath_RF_bus_reg_dataout_2294_port, 
      DataPath_RF_bus_reg_dataout_2295_port, 
      DataPath_RF_bus_reg_dataout_2296_port, 
      DataPath_RF_bus_reg_dataout_2297_port, 
      DataPath_RF_bus_reg_dataout_2298_port, 
      DataPath_RF_bus_reg_dataout_2299_port, 
      DataPath_RF_bus_reg_dataout_2300_port, 
      DataPath_RF_bus_reg_dataout_2301_port, 
      DataPath_RF_bus_reg_dataout_2302_port, 
      DataPath_RF_bus_reg_dataout_2303_port, 
      DataPath_RF_bus_reg_dataout_2304_port, 
      DataPath_RF_bus_reg_dataout_2305_port, 
      DataPath_RF_bus_reg_dataout_2306_port, 
      DataPath_RF_bus_reg_dataout_2307_port, 
      DataPath_RF_bus_reg_dataout_2308_port, 
      DataPath_RF_bus_reg_dataout_2309_port, 
      DataPath_RF_bus_reg_dataout_2310_port, 
      DataPath_RF_bus_reg_dataout_2311_port, 
      DataPath_RF_bus_reg_dataout_2312_port, 
      DataPath_RF_bus_reg_dataout_2313_port, 
      DataPath_RF_bus_reg_dataout_2314_port, 
      DataPath_RF_bus_reg_dataout_2315_port, 
      DataPath_RF_bus_reg_dataout_2316_port, 
      DataPath_RF_bus_reg_dataout_2317_port, 
      DataPath_RF_bus_reg_dataout_2318_port, 
      DataPath_RF_bus_reg_dataout_2319_port, 
      DataPath_RF_bus_reg_dataout_2320_port, 
      DataPath_RF_bus_reg_dataout_2321_port, 
      DataPath_RF_bus_reg_dataout_2322_port, 
      DataPath_RF_bus_reg_dataout_2323_port, 
      DataPath_RF_bus_reg_dataout_2324_port, 
      DataPath_RF_bus_reg_dataout_2325_port, 
      DataPath_RF_bus_reg_dataout_2326_port, 
      DataPath_RF_bus_reg_dataout_2327_port, 
      DataPath_RF_bus_reg_dataout_2328_port, 
      DataPath_RF_bus_reg_dataout_2329_port, 
      DataPath_RF_bus_reg_dataout_2330_port, 
      DataPath_RF_bus_reg_dataout_2331_port, 
      DataPath_RF_bus_reg_dataout_2332_port, 
      DataPath_RF_bus_reg_dataout_2333_port, 
      DataPath_RF_bus_reg_dataout_2334_port, 
      DataPath_RF_bus_reg_dataout_2335_port, 
      DataPath_RF_bus_reg_dataout_2336_port, 
      DataPath_RF_bus_reg_dataout_2337_port, 
      DataPath_RF_bus_reg_dataout_2338_port, 
      DataPath_RF_bus_reg_dataout_2339_port, 
      DataPath_RF_bus_reg_dataout_2340_port, 
      DataPath_RF_bus_reg_dataout_2341_port, 
      DataPath_RF_bus_reg_dataout_2342_port, 
      DataPath_RF_bus_reg_dataout_2343_port, 
      DataPath_RF_bus_reg_dataout_2344_port, 
      DataPath_RF_bus_reg_dataout_2345_port, 
      DataPath_RF_bus_reg_dataout_2346_port, 
      DataPath_RF_bus_reg_dataout_2347_port, 
      DataPath_RF_bus_reg_dataout_2348_port, 
      DataPath_RF_bus_reg_dataout_2349_port, 
      DataPath_RF_bus_reg_dataout_2350_port, 
      DataPath_RF_bus_reg_dataout_2351_port, 
      DataPath_RF_bus_reg_dataout_2352_port, 
      DataPath_RF_bus_reg_dataout_2353_port, 
      DataPath_RF_bus_reg_dataout_2354_port, 
      DataPath_RF_bus_reg_dataout_2355_port, 
      DataPath_RF_bus_reg_dataout_2356_port, 
      DataPath_RF_bus_reg_dataout_2357_port, 
      DataPath_RF_bus_reg_dataout_2358_port, 
      DataPath_RF_bus_reg_dataout_2359_port, 
      DataPath_RF_bus_reg_dataout_2360_port, 
      DataPath_RF_bus_reg_dataout_2361_port, 
      DataPath_RF_bus_reg_dataout_2362_port, 
      DataPath_RF_bus_reg_dataout_2363_port, 
      DataPath_RF_bus_reg_dataout_2364_port, 
      DataPath_RF_bus_reg_dataout_2365_port, 
      DataPath_RF_bus_reg_dataout_2366_port, 
      DataPath_RF_bus_reg_dataout_2367_port, 
      DataPath_RF_bus_reg_dataout_2368_port, 
      DataPath_RF_bus_reg_dataout_2369_port, 
      DataPath_RF_bus_reg_dataout_2370_port, 
      DataPath_RF_bus_reg_dataout_2371_port, 
      DataPath_RF_bus_reg_dataout_2372_port, 
      DataPath_RF_bus_reg_dataout_2373_port, 
      DataPath_RF_bus_reg_dataout_2374_port, 
      DataPath_RF_bus_reg_dataout_2375_port, 
      DataPath_RF_bus_reg_dataout_2376_port, 
      DataPath_RF_bus_reg_dataout_2377_port, 
      DataPath_RF_bus_reg_dataout_2378_port, 
      DataPath_RF_bus_reg_dataout_2379_port, 
      DataPath_RF_bus_reg_dataout_2380_port, 
      DataPath_RF_bus_reg_dataout_2381_port, 
      DataPath_RF_bus_reg_dataout_2382_port, 
      DataPath_RF_bus_reg_dataout_2383_port, 
      DataPath_RF_bus_reg_dataout_2384_port, 
      DataPath_RF_bus_reg_dataout_2385_port, 
      DataPath_RF_bus_reg_dataout_2386_port, 
      DataPath_RF_bus_reg_dataout_2387_port, 
      DataPath_RF_bus_reg_dataout_2388_port, 
      DataPath_RF_bus_reg_dataout_2389_port, 
      DataPath_RF_bus_reg_dataout_2390_port, 
      DataPath_RF_bus_reg_dataout_2391_port, 
      DataPath_RF_bus_reg_dataout_2392_port, 
      DataPath_RF_bus_reg_dataout_2393_port, 
      DataPath_RF_bus_reg_dataout_2394_port, 
      DataPath_RF_bus_reg_dataout_2395_port, 
      DataPath_RF_bus_reg_dataout_2396_port, 
      DataPath_RF_bus_reg_dataout_2397_port, 
      DataPath_RF_bus_reg_dataout_2398_port, 
      DataPath_RF_bus_reg_dataout_2399_port, 
      DataPath_RF_bus_reg_dataout_2400_port, 
      DataPath_RF_bus_reg_dataout_2401_port, 
      DataPath_RF_bus_reg_dataout_2402_port, 
      DataPath_RF_bus_reg_dataout_2403_port, 
      DataPath_RF_bus_reg_dataout_2404_port, 
      DataPath_RF_bus_reg_dataout_2405_port, 
      DataPath_RF_bus_reg_dataout_2406_port, 
      DataPath_RF_bus_reg_dataout_2407_port, 
      DataPath_RF_bus_reg_dataout_2408_port, 
      DataPath_RF_bus_reg_dataout_2409_port, 
      DataPath_RF_bus_reg_dataout_2410_port, 
      DataPath_RF_bus_reg_dataout_2411_port, 
      DataPath_RF_bus_reg_dataout_2412_port, 
      DataPath_RF_bus_reg_dataout_2413_port, 
      DataPath_RF_bus_reg_dataout_2414_port, 
      DataPath_RF_bus_reg_dataout_2415_port, 
      DataPath_RF_bus_reg_dataout_2416_port, 
      DataPath_RF_bus_reg_dataout_2417_port, 
      DataPath_RF_bus_reg_dataout_2418_port, 
      DataPath_RF_bus_reg_dataout_2419_port, 
      DataPath_RF_bus_reg_dataout_2420_port, 
      DataPath_RF_bus_reg_dataout_2421_port, 
      DataPath_RF_bus_reg_dataout_2422_port, 
      DataPath_RF_bus_reg_dataout_2423_port, 
      DataPath_RF_bus_reg_dataout_2424_port, 
      DataPath_RF_bus_reg_dataout_2425_port, 
      DataPath_RF_bus_reg_dataout_2426_port, 
      DataPath_RF_bus_reg_dataout_2427_port, 
      DataPath_RF_bus_reg_dataout_2428_port, 
      DataPath_RF_bus_reg_dataout_2429_port, 
      DataPath_RF_bus_reg_dataout_2430_port, 
      DataPath_RF_bus_reg_dataout_2431_port, 
      DataPath_RF_bus_reg_dataout_2432_port, 
      DataPath_RF_bus_reg_dataout_2433_port, 
      DataPath_RF_bus_reg_dataout_2434_port, 
      DataPath_RF_bus_reg_dataout_2435_port, 
      DataPath_RF_bus_reg_dataout_2436_port, 
      DataPath_RF_bus_reg_dataout_2437_port, 
      DataPath_RF_bus_reg_dataout_2438_port, 
      DataPath_RF_bus_reg_dataout_2439_port, 
      DataPath_RF_bus_reg_dataout_2440_port, 
      DataPath_RF_bus_reg_dataout_2441_port, 
      DataPath_RF_bus_reg_dataout_2442_port, 
      DataPath_RF_bus_reg_dataout_2443_port, 
      DataPath_RF_bus_reg_dataout_2444_port, 
      DataPath_RF_bus_reg_dataout_2445_port, 
      DataPath_RF_bus_reg_dataout_2446_port, 
      DataPath_RF_bus_reg_dataout_2447_port, 
      DataPath_RF_bus_reg_dataout_2448_port, 
      DataPath_RF_bus_reg_dataout_2449_port, 
      DataPath_RF_bus_reg_dataout_2450_port, 
      DataPath_RF_bus_reg_dataout_2451_port, 
      DataPath_RF_bus_reg_dataout_2452_port, 
      DataPath_RF_bus_reg_dataout_2453_port, 
      DataPath_RF_bus_reg_dataout_2454_port, 
      DataPath_RF_bus_reg_dataout_2455_port, 
      DataPath_RF_bus_reg_dataout_2456_port, 
      DataPath_RF_bus_reg_dataout_2457_port, 
      DataPath_RF_bus_reg_dataout_2458_port, 
      DataPath_RF_bus_reg_dataout_2459_port, 
      DataPath_RF_bus_reg_dataout_2460_port, 
      DataPath_RF_bus_reg_dataout_2461_port, 
      DataPath_RF_bus_reg_dataout_2462_port, 
      DataPath_RF_bus_reg_dataout_2463_port, 
      DataPath_RF_bus_reg_dataout_2464_port, 
      DataPath_RF_bus_reg_dataout_2465_port, 
      DataPath_RF_bus_reg_dataout_2466_port, 
      DataPath_RF_bus_reg_dataout_2467_port, 
      DataPath_RF_bus_reg_dataout_2468_port, 
      DataPath_RF_bus_reg_dataout_2469_port, 
      DataPath_RF_bus_reg_dataout_2470_port, 
      DataPath_RF_bus_reg_dataout_2471_port, 
      DataPath_RF_bus_reg_dataout_2472_port, 
      DataPath_RF_bus_reg_dataout_2473_port, 
      DataPath_RF_bus_reg_dataout_2474_port, 
      DataPath_RF_bus_reg_dataout_2475_port, 
      DataPath_RF_bus_reg_dataout_2476_port, 
      DataPath_RF_bus_reg_dataout_2477_port, 
      DataPath_RF_bus_reg_dataout_2478_port, 
      DataPath_RF_bus_reg_dataout_2479_port, 
      DataPath_RF_bus_reg_dataout_2480_port, 
      DataPath_RF_bus_reg_dataout_2481_port, 
      DataPath_RF_bus_reg_dataout_2482_port, 
      DataPath_RF_bus_reg_dataout_2483_port, 
      DataPath_RF_bus_reg_dataout_2484_port, 
      DataPath_RF_bus_reg_dataout_2485_port, 
      DataPath_RF_bus_reg_dataout_2486_port, 
      DataPath_RF_bus_reg_dataout_2487_port, 
      DataPath_RF_bus_reg_dataout_2488_port, 
      DataPath_RF_bus_reg_dataout_2489_port, 
      DataPath_RF_bus_reg_dataout_2490_port, 
      DataPath_RF_bus_reg_dataout_2491_port, 
      DataPath_RF_bus_reg_dataout_2492_port, 
      DataPath_RF_bus_reg_dataout_2493_port, 
      DataPath_RF_bus_reg_dataout_2494_port, 
      DataPath_RF_bus_reg_dataout_2495_port, 
      DataPath_RF_bus_reg_dataout_2496_port, 
      DataPath_RF_bus_reg_dataout_2497_port, 
      DataPath_RF_bus_reg_dataout_2498_port, 
      DataPath_RF_bus_reg_dataout_2499_port, 
      DataPath_RF_bus_reg_dataout_2500_port, 
      DataPath_RF_bus_reg_dataout_2501_port, 
      DataPath_RF_bus_reg_dataout_2502_port, 
      DataPath_RF_bus_reg_dataout_2503_port, 
      DataPath_RF_bus_reg_dataout_2504_port, 
      DataPath_RF_bus_reg_dataout_2505_port, 
      DataPath_RF_bus_reg_dataout_2506_port, 
      DataPath_RF_bus_reg_dataout_2507_port, 
      DataPath_RF_bus_reg_dataout_2508_port, 
      DataPath_RF_bus_reg_dataout_2509_port, 
      DataPath_RF_bus_reg_dataout_2510_port, 
      DataPath_RF_bus_reg_dataout_2511_port, 
      DataPath_RF_bus_reg_dataout_2512_port, 
      DataPath_RF_bus_reg_dataout_2513_port, 
      DataPath_RF_bus_reg_dataout_2514_port, 
      DataPath_RF_bus_reg_dataout_2515_port, 
      DataPath_RF_bus_reg_dataout_2516_port, 
      DataPath_RF_bus_reg_dataout_2517_port, 
      DataPath_RF_bus_reg_dataout_2518_port, 
      DataPath_RF_bus_reg_dataout_2519_port, 
      DataPath_RF_bus_reg_dataout_2520_port, 
      DataPath_RF_bus_reg_dataout_2521_port, 
      DataPath_RF_bus_reg_dataout_2522_port, 
      DataPath_RF_bus_reg_dataout_2523_port, 
      DataPath_RF_bus_reg_dataout_2524_port, 
      DataPath_RF_bus_reg_dataout_2525_port, 
      DataPath_RF_bus_reg_dataout_2526_port, 
      DataPath_RF_bus_reg_dataout_2527_port, 
      DataPath_RF_bus_reg_dataout_2528_port, 
      DataPath_RF_bus_reg_dataout_2529_port, 
      DataPath_RF_bus_reg_dataout_2530_port, 
      DataPath_RF_bus_reg_dataout_2531_port, 
      DataPath_RF_bus_reg_dataout_2532_port, 
      DataPath_RF_bus_reg_dataout_2533_port, 
      DataPath_RF_bus_reg_dataout_2534_port, 
      DataPath_RF_bus_reg_dataout_2535_port, 
      DataPath_RF_bus_reg_dataout_2536_port, 
      DataPath_RF_bus_reg_dataout_2537_port, 
      DataPath_RF_bus_reg_dataout_2538_port, 
      DataPath_RF_bus_reg_dataout_2539_port, 
      DataPath_RF_bus_reg_dataout_2540_port, 
      DataPath_RF_bus_reg_dataout_2541_port, 
      DataPath_RF_bus_reg_dataout_2542_port, 
      DataPath_RF_bus_reg_dataout_2543_port, 
      DataPath_RF_bus_reg_dataout_2544_port, 
      DataPath_RF_bus_reg_dataout_2545_port, 
      DataPath_RF_bus_reg_dataout_2546_port, 
      DataPath_RF_bus_reg_dataout_2547_port, 
      DataPath_RF_bus_reg_dataout_2548_port, 
      DataPath_RF_bus_reg_dataout_2549_port, 
      DataPath_RF_bus_reg_dataout_2550_port, 
      DataPath_RF_bus_reg_dataout_2551_port, 
      DataPath_RF_bus_reg_dataout_2552_port, 
      DataPath_RF_bus_reg_dataout_2553_port, 
      DataPath_RF_bus_reg_dataout_2554_port, 
      DataPath_RF_bus_reg_dataout_2555_port, 
      DataPath_RF_bus_reg_dataout_2556_port, 
      DataPath_RF_bus_reg_dataout_2557_port, 
      DataPath_RF_bus_reg_dataout_2558_port, 
      DataPath_RF_bus_reg_dataout_2559_port, DataPath_RF_c_win_0_port, 
      DataPath_RF_c_win_1_port, DataPath_RF_c_win_2_port, 
      DataPath_RF_c_win_3_port, DataPath_RF_c_win_4_port, 
      DataPath_WRF_CUhw_N145, DataPath_WRF_CUhw_curr_addr_2_port, 
      DataPath_WRF_CUhw_curr_addr_3_port, DataPath_WRF_CUhw_curr_addr_4_port, 
      DataPath_WRF_CUhw_curr_addr_5_port, DataPath_WRF_CUhw_curr_addr_6_port, 
      DataPath_WRF_CUhw_curr_addr_7_port, DataPath_WRF_CUhw_curr_addr_8_port, 
      DataPath_WRF_CUhw_curr_addr_9_port, DataPath_WRF_CUhw_curr_addr_10_port, 
      DataPath_WRF_CUhw_curr_addr_11_port, DataPath_WRF_CUhw_curr_addr_12_port,
      DataPath_WRF_CUhw_curr_addr_13_port, DataPath_WRF_CUhw_curr_addr_14_port,
      DataPath_WRF_CUhw_curr_addr_15_port, DataPath_WRF_CUhw_curr_addr_16_port,
      DataPath_WRF_CUhw_curr_addr_17_port, DataPath_WRF_CUhw_curr_addr_18_port,
      DataPath_WRF_CUhw_curr_addr_19_port, DataPath_WRF_CUhw_curr_addr_20_port,
      DataPath_WRF_CUhw_curr_addr_21_port, DataPath_WRF_CUhw_curr_addr_22_port,
      DataPath_WRF_CUhw_curr_addr_23_port, DataPath_WRF_CUhw_curr_addr_24_port,
      DataPath_WRF_CUhw_curr_addr_25_port, DataPath_WRF_CUhw_curr_addr_26_port,
      DataPath_WRF_CUhw_curr_addr_27_port, DataPath_WRF_CUhw_curr_addr_28_port,
      DataPath_WRF_CUhw_curr_addr_29_port, DataPath_WRF_CUhw_curr_addr_30_port,
      DataPath_WRF_CUhw_curr_addr_31_port, DataPath_WRF_CUhw_curr_data_0_port, 
      DataPath_WRF_CUhw_curr_data_1_port, DataPath_WRF_CUhw_curr_data_2_port, 
      DataPath_WRF_CUhw_curr_data_3_port, DataPath_WRF_CUhw_curr_data_4_port, 
      DataPath_WRF_CUhw_curr_data_5_port, DataPath_WRF_CUhw_curr_data_6_port, 
      DataPath_WRF_CUhw_curr_data_7_port, DataPath_WRF_CUhw_curr_data_8_port, 
      DataPath_WRF_CUhw_curr_data_9_port, DataPath_WRF_CUhw_curr_data_10_port, 
      DataPath_WRF_CUhw_curr_data_11_port, DataPath_WRF_CUhw_curr_data_12_port,
      DataPath_WRF_CUhw_curr_data_13_port, DataPath_WRF_CUhw_curr_data_14_port,
      DataPath_WRF_CUhw_curr_data_15_port, DataPath_WRF_CUhw_curr_data_16_port,
      DataPath_WRF_CUhw_curr_data_17_port, DataPath_WRF_CUhw_curr_data_18_port,
      DataPath_WRF_CUhw_curr_data_19_port, DataPath_WRF_CUhw_curr_data_20_port,
      DataPath_WRF_CUhw_curr_data_21_port, DataPath_WRF_CUhw_curr_data_22_port,
      DataPath_WRF_CUhw_curr_data_23_port, DataPath_WRF_CUhw_curr_data_24_port,
      DataPath_WRF_CUhw_curr_data_25_port, DataPath_WRF_CUhw_curr_data_26_port,
      DataPath_WRF_CUhw_curr_data_27_port, DataPath_WRF_CUhw_curr_data_28_port,
      DataPath_WRF_CUhw_curr_data_29_port, DataPath_WRF_CUhw_curr_data_30_port,
      DataPath_WRF_CUhw_curr_data_31_port, DataPath_ALUhw_i_Q_EXTENDED_34_port,
      DataPath_ALUhw_i_Q_EXTENDED_36_port, DataPath_ALUhw_i_Q_EXTENDED_37_port,
      DataPath_ALUhw_i_Q_EXTENDED_40_port, DataPath_ALUhw_i_Q_EXTENDED_41_port,
      DataPath_ALUhw_i_Q_EXTENDED_42_port, DataPath_ALUhw_i_Q_EXTENDED_43_port,
      DataPath_ALUhw_i_Q_EXTENDED_44_port, DataPath_ALUhw_i_Q_EXTENDED_46_port,
      DataPath_ALUhw_i_Q_EXTENDED_47_port, DataPath_ALUhw_i_Q_EXTENDED_50_port,
      DataPath_ALUhw_i_Q_EXTENDED_51_port, DataPath_ALUhw_i_Q_EXTENDED_52_port,
      DataPath_ALUhw_i_Q_EXTENDED_54_port, DataPath_ALUhw_i_Q_EXTENDED_55_port,
      DataPath_ALUhw_i_Q_EXTENDED_56_port, DataPath_ALUhw_i_Q_EXTENDED_57_port,
      DataPath_ALUhw_i_Q_EXTENDED_58_port, DataPath_ALUhw_i_Q_EXTENDED_59_port,
      DataPath_ALUhw_i_Q_EXTENDED_60_port, DataPath_ALUhw_i_Q_EXTENDED_61_port,
      DataPath_RF_RDPORT0_OUTLATCH_N35, DataPath_RF_RDPORT0_OUTLATCH_N34, 
      DataPath_RF_RDPORT0_OUTLATCH_N33, DataPath_RF_RDPORT0_OUTLATCH_N32, 
      DataPath_RF_RDPORT0_OUTLATCH_N31, DataPath_RF_RDPORT0_OUTLATCH_N30, 
      DataPath_RF_RDPORT0_OUTLATCH_N29, DataPath_RF_RDPORT0_OUTLATCH_N28, 
      DataPath_RF_RDPORT0_OUTLATCH_N27, DataPath_RF_RDPORT0_OUTLATCH_N26, 
      DataPath_RF_RDPORT0_OUTLATCH_N25, DataPath_RF_RDPORT0_OUTLATCH_N24, 
      DataPath_RF_RDPORT0_OUTLATCH_N23, DataPath_RF_RDPORT0_OUTLATCH_N22, 
      DataPath_RF_RDPORT0_OUTLATCH_N21, DataPath_RF_RDPORT0_OUTLATCH_N20, 
      DataPath_RF_RDPORT0_OUTLATCH_N19, DataPath_RF_RDPORT0_OUTLATCH_N18, 
      DataPath_RF_RDPORT0_OUTLATCH_N17, DataPath_RF_RDPORT0_OUTLATCH_N16, 
      DataPath_RF_RDPORT0_OUTLATCH_N15, DataPath_RF_RDPORT0_OUTLATCH_N14, 
      DataPath_RF_RDPORT0_OUTLATCH_N13, DataPath_RF_RDPORT0_OUTLATCH_N12, 
      DataPath_RF_RDPORT0_OUTLATCH_N11, DataPath_RF_RDPORT0_OUTLATCH_N10, 
      DataPath_RF_RDPORT0_OUTLATCH_N9, DataPath_RF_RDPORT0_OUTLATCH_N8, 
      DataPath_RF_RDPORT0_OUTLATCH_N7, DataPath_RF_RDPORT0_OUTLATCH_N6, 
      DataPath_RF_RDPORT0_OUTLATCH_N5, DataPath_RF_RDPORT0_OUTLATCH_N4, 
      DataPath_RF_RDPORT0_OUTLATCH_N3, DataPath_RF_RDPORT1_OUTLATCH_N35, 
      DataPath_RF_RDPORT1_OUTLATCH_N34, DataPath_RF_RDPORT1_OUTLATCH_N33, 
      DataPath_RF_RDPORT1_OUTLATCH_N32, DataPath_RF_RDPORT1_OUTLATCH_N31, 
      DataPath_RF_RDPORT1_OUTLATCH_N30, DataPath_RF_RDPORT1_OUTLATCH_N29, 
      DataPath_RF_RDPORT1_OUTLATCH_N28, DataPath_RF_RDPORT1_OUTLATCH_N27, 
      DataPath_RF_RDPORT1_OUTLATCH_N26, DataPath_RF_RDPORT1_OUTLATCH_N25, 
      DataPath_RF_RDPORT1_OUTLATCH_N24, DataPath_RF_RDPORT1_OUTLATCH_N23, 
      DataPath_RF_RDPORT1_OUTLATCH_N22, DataPath_RF_RDPORT1_OUTLATCH_N21, 
      DataPath_RF_RDPORT1_OUTLATCH_N20, DataPath_RF_RDPORT1_OUTLATCH_N19, 
      DataPath_RF_RDPORT1_OUTLATCH_N18, DataPath_RF_RDPORT1_OUTLATCH_N17, 
      DataPath_RF_RDPORT1_OUTLATCH_N16, DataPath_RF_RDPORT1_OUTLATCH_N15, 
      DataPath_RF_RDPORT1_OUTLATCH_N14, DataPath_RF_RDPORT1_OUTLATCH_N13, 
      DataPath_RF_RDPORT1_OUTLATCH_N12, DataPath_RF_RDPORT1_OUTLATCH_N11, 
      DataPath_RF_RDPORT1_OUTLATCH_N10, DataPath_RF_RDPORT1_OUTLATCH_N9, 
      DataPath_RF_RDPORT1_OUTLATCH_N8, DataPath_RF_RDPORT1_OUTLATCH_N7, 
      DataPath_RF_RDPORT1_OUTLATCH_N6, DataPath_RF_RDPORT1_OUTLATCH_N5, 
      DataPath_RF_RDPORT1_OUTLATCH_N4, DataPath_RF_RDPORT1_OUTLATCH_N3, 
      DataPath_RF_PUSH_ADDRGEN_N61, DataPath_RF_PUSH_ADDRGEN_N60, 
      DataPath_RF_PUSH_ADDRGEN_N59, DataPath_RF_PUSH_ADDRGEN_N58, 
      DataPath_RF_PUSH_ADDRGEN_N57, DataPath_RF_PUSH_ADDRGEN_N56, 
      DataPath_RF_PUSH_ADDRGEN_N55, DataPath_RF_PUSH_ADDRGEN_N54, 
      DataPath_RF_PUSH_ADDRGEN_N53, DataPath_RF_PUSH_ADDRGEN_N52, 
      DataPath_RF_PUSH_ADDRGEN_N51, DataPath_RF_PUSH_ADDRGEN_N50, 
      DataPath_RF_PUSH_ADDRGEN_N49, DataPath_RF_PUSH_ADDRGEN_N48, 
      DataPath_RF_PUSH_ADDRGEN_N47, DataPath_RF_PUSH_ADDRGEN_N46, 
      DataPath_RF_PUSH_ADDRGEN_curr_state_0_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, 
      DataPath_RF_PUSH_ADDRGEN_curr_addr_15_port, DataPath_RF_POP_ADDRGEN_N61, 
      DataPath_RF_POP_ADDRGEN_N60, DataPath_RF_POP_ADDRGEN_N59, 
      DataPath_RF_POP_ADDRGEN_N58, DataPath_RF_POP_ADDRGEN_N57, 
      DataPath_RF_POP_ADDRGEN_N56, DataPath_RF_POP_ADDRGEN_N55, 
      DataPath_RF_POP_ADDRGEN_N54, DataPath_RF_POP_ADDRGEN_N53, 
      DataPath_RF_POP_ADDRGEN_N52, DataPath_RF_POP_ADDRGEN_N51, 
      DataPath_RF_POP_ADDRGEN_N50, DataPath_RF_POP_ADDRGEN_N49, 
      DataPath_RF_POP_ADDRGEN_N48, DataPath_RF_POP_ADDRGEN_N47, 
      DataPath_RF_POP_ADDRGEN_N46, DataPath_RF_POP_ADDRGEN_curr_state_1_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_0_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_1_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_2_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_3_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_4_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_5_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_6_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_7_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_8_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_9_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_10_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_11_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_12_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_13_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_14_port, 
      DataPath_RF_POP_ADDRGEN_curr_addr_15_port, 
      DataPath_ALUhw_MULT_mux_out_15_30_port, 
      DataPath_ALUhw_MULT_mux_out_15_31_port, 
      DataPath_ALUhw_MULT_mux_out_14_28_port, 
      DataPath_ALUhw_MULT_mux_out_14_29_port, 
      DataPath_ALUhw_MULT_mux_out_14_30_port, 
      DataPath_ALUhw_MULT_mux_out_14_31_port, 
      DataPath_ALUhw_MULT_mux_out_13_26_port, 
      DataPath_ALUhw_MULT_mux_out_13_27_port, 
      DataPath_ALUhw_MULT_mux_out_13_28_port, 
      DataPath_ALUhw_MULT_mux_out_13_29_port, 
      DataPath_ALUhw_MULT_mux_out_13_30_port, 
      DataPath_ALUhw_MULT_mux_out_13_31_port, 
      DataPath_ALUhw_MULT_mux_out_12_24_port, 
      DataPath_ALUhw_MULT_mux_out_12_25_port, 
      DataPath_ALUhw_MULT_mux_out_12_26_port, 
      DataPath_ALUhw_MULT_mux_out_12_27_port, 
      DataPath_ALUhw_MULT_mux_out_12_28_port, 
      DataPath_ALUhw_MULT_mux_out_12_29_port, 
      DataPath_ALUhw_MULT_mux_out_12_30_port, 
      DataPath_ALUhw_MULT_mux_out_12_31_port, 
      DataPath_ALUhw_MULT_mux_out_11_22_port, 
      DataPath_ALUhw_MULT_mux_out_11_23_port, 
      DataPath_ALUhw_MULT_mux_out_11_24_port, 
      DataPath_ALUhw_MULT_mux_out_11_26_port, 
      DataPath_ALUhw_MULT_mux_out_11_27_port, 
      DataPath_ALUhw_MULT_mux_out_11_28_port, 
      DataPath_ALUhw_MULT_mux_out_11_29_port, 
      DataPath_ALUhw_MULT_mux_out_11_30_port, 
      DataPath_ALUhw_MULT_mux_out_11_31_port, 
      DataPath_ALUhw_MULT_mux_out_10_20_port, 
      DataPath_ALUhw_MULT_mux_out_10_21_port, 
      DataPath_ALUhw_MULT_mux_out_10_22_port, 
      DataPath_ALUhw_MULT_mux_out_10_23_port, 
      DataPath_ALUhw_MULT_mux_out_10_24_port, 
      DataPath_ALUhw_MULT_mux_out_10_25_port, 
      DataPath_ALUhw_MULT_mux_out_10_26_port, 
      DataPath_ALUhw_MULT_mux_out_10_27_port, 
      DataPath_ALUhw_MULT_mux_out_10_28_port, 
      DataPath_ALUhw_MULT_mux_out_10_29_port, 
      DataPath_ALUhw_MULT_mux_out_10_30_port, 
      DataPath_ALUhw_MULT_mux_out_10_31_port, 
      DataPath_ALUhw_MULT_mux_out_9_19_port, 
      DataPath_ALUhw_MULT_mux_out_9_20_port, 
      DataPath_ALUhw_MULT_mux_out_9_21_port, 
      DataPath_ALUhw_MULT_mux_out_9_22_port, 
      DataPath_ALUhw_MULT_mux_out_9_23_port, 
      DataPath_ALUhw_MULT_mux_out_9_24_port, 
      DataPath_ALUhw_MULT_mux_out_9_25_port, 
      DataPath_ALUhw_MULT_mux_out_9_26_port, 
      DataPath_ALUhw_MULT_mux_out_9_27_port, 
      DataPath_ALUhw_MULT_mux_out_9_28_port, 
      DataPath_ALUhw_MULT_mux_out_9_29_port, 
      DataPath_ALUhw_MULT_mux_out_9_30_port, 
      DataPath_ALUhw_MULT_mux_out_9_31_port, 
      DataPath_ALUhw_MULT_mux_out_8_16_port, 
      DataPath_ALUhw_MULT_mux_out_8_17_port, 
      DataPath_ALUhw_MULT_mux_out_8_18_port, 
      DataPath_ALUhw_MULT_mux_out_8_19_port, 
      DataPath_ALUhw_MULT_mux_out_8_20_port, 
      DataPath_ALUhw_MULT_mux_out_8_21_port, 
      DataPath_ALUhw_MULT_mux_out_8_22_port, 
      DataPath_ALUhw_MULT_mux_out_8_23_port, 
      DataPath_ALUhw_MULT_mux_out_8_24_port, 
      DataPath_ALUhw_MULT_mux_out_8_25_port, 
      DataPath_ALUhw_MULT_mux_out_8_26_port, 
      DataPath_ALUhw_MULT_mux_out_8_27_port, 
      DataPath_ALUhw_MULT_mux_out_8_28_port, 
      DataPath_ALUhw_MULT_mux_out_8_29_port, 
      DataPath_ALUhw_MULT_mux_out_8_30_port, 
      DataPath_ALUhw_MULT_mux_out_8_31_port, 
      DataPath_ALUhw_MULT_mux_out_7_14_port, 
      DataPath_ALUhw_MULT_mux_out_7_15_port, 
      DataPath_ALUhw_MULT_mux_out_7_16_port, 
      DataPath_ALUhw_MULT_mux_out_7_17_port, 
      DataPath_ALUhw_MULT_mux_out_7_18_port, 
      DataPath_ALUhw_MULT_mux_out_7_19_port, 
      DataPath_ALUhw_MULT_mux_out_7_20_port, 
      DataPath_ALUhw_MULT_mux_out_7_21_port, 
      DataPath_ALUhw_MULT_mux_out_7_22_port, 
      DataPath_ALUhw_MULT_mux_out_7_23_port, 
      DataPath_ALUhw_MULT_mux_out_7_24_port, 
      DataPath_ALUhw_MULT_mux_out_7_25_port, 
      DataPath_ALUhw_MULT_mux_out_7_26_port, 
      DataPath_ALUhw_MULT_mux_out_7_27_port, 
      DataPath_ALUhw_MULT_mux_out_7_28_port, 
      DataPath_ALUhw_MULT_mux_out_7_29_port, 
      DataPath_ALUhw_MULT_mux_out_7_30_port, 
      DataPath_ALUhw_MULT_mux_out_7_31_port, 
      DataPath_ALUhw_MULT_mux_out_6_12_port, 
      DataPath_ALUhw_MULT_mux_out_6_13_port, 
      DataPath_ALUhw_MULT_mux_out_6_14_port, 
      DataPath_ALUhw_MULT_mux_out_6_15_port, 
      DataPath_ALUhw_MULT_mux_out_6_16_port, 
      DataPath_ALUhw_MULT_mux_out_6_17_port, 
      DataPath_ALUhw_MULT_mux_out_6_18_port, 
      DataPath_ALUhw_MULT_mux_out_6_19_port, 
      DataPath_ALUhw_MULT_mux_out_6_20_port, 
      DataPath_ALUhw_MULT_mux_out_6_21_port, 
      DataPath_ALUhw_MULT_mux_out_6_22_port, 
      DataPath_ALUhw_MULT_mux_out_6_23_port, 
      DataPath_ALUhw_MULT_mux_out_6_25_port, 
      DataPath_ALUhw_MULT_mux_out_6_26_port, 
      DataPath_ALUhw_MULT_mux_out_6_27_port, 
      DataPath_ALUhw_MULT_mux_out_6_28_port, 
      DataPath_ALUhw_MULT_mux_out_6_29_port, 
      DataPath_ALUhw_MULT_mux_out_6_30_port, 
      DataPath_ALUhw_MULT_mux_out_6_31_port, 
      DataPath_ALUhw_MULT_mux_out_5_11_port, 
      DataPath_ALUhw_MULT_mux_out_5_12_port, 
      DataPath_ALUhw_MULT_mux_out_5_13_port, 
      DataPath_ALUhw_MULT_mux_out_5_14_port, 
      DataPath_ALUhw_MULT_mux_out_5_15_port, 
      DataPath_ALUhw_MULT_mux_out_5_16_port, 
      DataPath_ALUhw_MULT_mux_out_5_17_port, 
      DataPath_ALUhw_MULT_mux_out_5_18_port, 
      DataPath_ALUhw_MULT_mux_out_5_19_port, 
      DataPath_ALUhw_MULT_mux_out_5_20_port, 
      DataPath_ALUhw_MULT_mux_out_5_21_port, 
      DataPath_ALUhw_MULT_mux_out_5_22_port, 
      DataPath_ALUhw_MULT_mux_out_5_23_port, 
      DataPath_ALUhw_MULT_mux_out_5_24_port, 
      DataPath_ALUhw_MULT_mux_out_5_25_port, 
      DataPath_ALUhw_MULT_mux_out_5_26_port, 
      DataPath_ALUhw_MULT_mux_out_5_27_port, 
      DataPath_ALUhw_MULT_mux_out_5_28_port, 
      DataPath_ALUhw_MULT_mux_out_5_29_port, 
      DataPath_ALUhw_MULT_mux_out_5_30_port, 
      DataPath_ALUhw_MULT_mux_out_5_31_port, 
      DataPath_ALUhw_MULT_mux_out_4_9_port, 
      DataPath_ALUhw_MULT_mux_out_4_10_port, 
      DataPath_ALUhw_MULT_mux_out_4_11_port, 
      DataPath_ALUhw_MULT_mux_out_4_12_port, 
      DataPath_ALUhw_MULT_mux_out_4_13_port, 
      DataPath_ALUhw_MULT_mux_out_4_14_port, 
      DataPath_ALUhw_MULT_mux_out_4_15_port, 
      DataPath_ALUhw_MULT_mux_out_4_16_port, 
      DataPath_ALUhw_MULT_mux_out_4_17_port, 
      DataPath_ALUhw_MULT_mux_out_4_18_port, 
      DataPath_ALUhw_MULT_mux_out_4_19_port, 
      DataPath_ALUhw_MULT_mux_out_4_20_port, 
      DataPath_ALUhw_MULT_mux_out_4_21_port, 
      DataPath_ALUhw_MULT_mux_out_4_23_port, 
      DataPath_ALUhw_MULT_mux_out_4_24_port, 
      DataPath_ALUhw_MULT_mux_out_4_25_port, 
      DataPath_ALUhw_MULT_mux_out_4_26_port, 
      DataPath_ALUhw_MULT_mux_out_4_27_port, 
      DataPath_ALUhw_MULT_mux_out_4_28_port, 
      DataPath_ALUhw_MULT_mux_out_4_29_port, 
      DataPath_ALUhw_MULT_mux_out_4_30_port, 
      DataPath_ALUhw_MULT_mux_out_4_31_port, 
      DataPath_ALUhw_MULT_mux_out_3_6_port, 
      DataPath_ALUhw_MULT_mux_out_3_7_port, 
      DataPath_ALUhw_MULT_mux_out_3_8_port, 
      DataPath_ALUhw_MULT_mux_out_3_9_port, 
      DataPath_ALUhw_MULT_mux_out_3_10_port, 
      DataPath_ALUhw_MULT_mux_out_3_11_port, 
      DataPath_ALUhw_MULT_mux_out_3_12_port, 
      DataPath_ALUhw_MULT_mux_out_3_13_port, 
      DataPath_ALUhw_MULT_mux_out_3_14_port, 
      DataPath_ALUhw_MULT_mux_out_3_15_port, 
      DataPath_ALUhw_MULT_mux_out_3_16_port, 
      DataPath_ALUhw_MULT_mux_out_3_17_port, 
      DataPath_ALUhw_MULT_mux_out_3_18_port, 
      DataPath_ALUhw_MULT_mux_out_3_19_port, 
      DataPath_ALUhw_MULT_mux_out_3_20_port, 
      DataPath_ALUhw_MULT_mux_out_3_21_port, 
      DataPath_ALUhw_MULT_mux_out_3_22_port, 
      DataPath_ALUhw_MULT_mux_out_3_23_port, 
      DataPath_ALUhw_MULT_mux_out_3_24_port, 
      DataPath_ALUhw_MULT_mux_out_3_26_port, 
      DataPath_ALUhw_MULT_mux_out_3_27_port, 
      DataPath_ALUhw_MULT_mux_out_3_28_port, 
      DataPath_ALUhw_MULT_mux_out_3_29_port, 
      DataPath_ALUhw_MULT_mux_out_3_30_port, 
      DataPath_ALUhw_MULT_mux_out_3_31_port, 
      DataPath_ALUhw_MULT_mux_out_2_5_port, 
      DataPath_ALUhw_MULT_mux_out_2_6_port, 
      DataPath_ALUhw_MULT_mux_out_2_7_port, 
      DataPath_ALUhw_MULT_mux_out_2_8_port, 
      DataPath_ALUhw_MULT_mux_out_2_9_port, 
      DataPath_ALUhw_MULT_mux_out_2_10_port, 
      DataPath_ALUhw_MULT_mux_out_2_11_port, 
      DataPath_ALUhw_MULT_mux_out_2_12_port, 
      DataPath_ALUhw_MULT_mux_out_2_13_port, 
      DataPath_ALUhw_MULT_mux_out_2_14_port, 
      DataPath_ALUhw_MULT_mux_out_2_15_port, 
      DataPath_ALUhw_MULT_mux_out_2_16_port, 
      DataPath_ALUhw_MULT_mux_out_2_17_port, 
      DataPath_ALUhw_MULT_mux_out_2_18_port, 
      DataPath_ALUhw_MULT_mux_out_2_19_port, 
      DataPath_ALUhw_MULT_mux_out_2_20_port, 
      DataPath_ALUhw_MULT_mux_out_2_21_port, 
      DataPath_ALUhw_MULT_mux_out_2_22_port, 
      DataPath_ALUhw_MULT_mux_out_2_23_port, 
      DataPath_ALUhw_MULT_mux_out_2_24_port, 
      DataPath_ALUhw_MULT_mux_out_2_25_port, 
      DataPath_ALUhw_MULT_mux_out_2_26_port, 
      DataPath_ALUhw_MULT_mux_out_2_27_port, 
      DataPath_ALUhw_MULT_mux_out_2_28_port, 
      DataPath_ALUhw_MULT_mux_out_2_29_port, 
      DataPath_ALUhw_MULT_mux_out_2_30_port, 
      DataPath_ALUhw_MULT_mux_out_2_31_port, 
      DataPath_ALUhw_MULT_mux_out_1_3_port, 
      DataPath_ALUhw_MULT_mux_out_1_5_port, 
      DataPath_ALUhw_MULT_mux_out_1_8_port, 
      DataPath_ALUhw_MULT_mux_out_1_10_port, 
      DataPath_ALUhw_MULT_mux_out_1_11_port, 
      DataPath_ALUhw_MULT_mux_out_1_12_port, 
      DataPath_ALUhw_MULT_mux_out_1_13_port, 
      DataPath_ALUhw_MULT_mux_out_1_14_port, 
      DataPath_ALUhw_MULT_mux_out_1_15_port, 
      DataPath_ALUhw_MULT_mux_out_1_16_port, 
      DataPath_ALUhw_MULT_mux_out_1_17_port, 
      DataPath_ALUhw_MULT_mux_out_1_18_port, 
      DataPath_ALUhw_MULT_mux_out_1_19_port, 
      DataPath_ALUhw_MULT_mux_out_1_20_port, 
      DataPath_ALUhw_MULT_mux_out_1_21_port, 
      DataPath_ALUhw_MULT_mux_out_1_22_port, 
      DataPath_ALUhw_MULT_mux_out_1_23_port, 
      DataPath_ALUhw_MULT_mux_out_1_24_port, 
      DataPath_ALUhw_MULT_mux_out_1_25_port, 
      DataPath_ALUhw_MULT_mux_out_1_26_port, 
      DataPath_ALUhw_MULT_mux_out_1_27_port, 
      DataPath_ALUhw_MULT_mux_out_1_28_port, 
      DataPath_ALUhw_MULT_mux_out_1_29_port, 
      DataPath_ALUhw_MULT_mux_out_1_30_port, 
      DataPath_ALUhw_MULT_mux_out_1_31_port, 
      DataPath_ALUhw_MULT_mux_out_0_0_port, 
      DataPath_ALUhw_MULT_mux_out_0_4_port, 
      DataPath_ALUhw_MULT_mux_out_0_5_port, 
      DataPath_ALUhw_MULT_mux_out_0_8_port, 
      DataPath_ALUhw_MULT_mux_out_0_9_port, 
      DataPath_ALUhw_MULT_mux_out_0_12_port, 
      DataPath_ALUhw_MULT_mux_out_0_14_port, 
      DataPath_ALUhw_MULT_mux_out_0_16_port, 
      DataPath_ALUhw_MULT_mux_out_0_17_port, 
      DataPath_ALUhw_MULT_mux_out_0_22_port, 
      DataPath_ALUhw_MULT_mux_out_0_25_port, 
      DataPath_ALUhw_MULT_mux_out_0_27_port, 
      DataPath_ALUhw_MULT_mux_out_0_29_port, 
      DataPath_ALUhw_MULT_mux_out_0_31_port, C620_DATA2_4, C620_DATA2_5, 
      C620_DATA2_6, C620_DATA2_7, C620_DATA2_8, C620_DATA2_12, C620_DATA2_14, 
      C620_DATA2_15, C620_DATA2_16, C620_DATA2_17, C620_DATA2_18, C620_DATA2_21
      , C620_DATA2_23, C620_DATA2_29, C620_DATA2_30, C620_DATA2_31, n34, n36, 
      n37, n38, n39, n40, n41, n42, n43, n90, n99, n143, n159, n161, n163, n167
      , n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
      n193, n205, n206, n207, n211, n212, n213, n217, n219, n355, n356, n357, 
      n358, n359, n364, n365, n366, n367, n368, n375, n376, n403, n460, n461, 
      n465, n466, n477, n486, n492, n493, n494, n495, n496, n497, n498, n499, 
      n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, 
      n512, n513, n514, n515, n523, n525, n541, n542, n544, n546, n548, n550, 
      n552, n554, n556, n558, n560, n562, n564, n566, n568, n569, n570, n575, 
      n576, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, 
      n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, 
      n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, 
      n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, 
      n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, 
      n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, 
      n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, 
      n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, 
      n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, 
      n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, 
      n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, 
      n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, 
      n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, 
      n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, 
      n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, 
      n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, 
      n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, 
      n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, 
      n814, n815, n816, n817, n818, n819, n820, n821, n822, n824, n825, n826, 
      n838, n866, n880, n884, n886, n888, n890, n892, n894, n896, n898, n900, 
      n902, n904, n906, n908, n910, n912, n914, n918, n920, n922, n924, n926, 
      n928, n930, n932, n934, n936, n938, n940, n942, n944, n946, n948, n949, 
      n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, 
      n962, n963, n968, n971, n972, n973, n974, n975, n976, n977, n978, n979, 
      n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, 
      n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1005, 
      n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, 
      n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, 
      n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, 
      n1038, n1042, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1079, n1082, n1083, n1084, n1085, n1086, n1087, 
      n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, 
      n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, 
      n1108, n1109, n1110, n1111, n1112, n1116, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1998, n2119, n2151, 
      n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, 
      n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, 
      n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, 
      n2208, n2209, n2332, n2334, n2336, n2338, n2340, n2342, n2344, n2346, 
      n2348, n2350, n2352, n2357, n2359, n2361, n2363, n2365, n2370, n2373, 
      n2375, n2377, n2380, n2384, n2387, n2700, n2701, n2702, n2703, n2704, 
      n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, 
      n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, 
      n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, 
      n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, 
      n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, 
      n2755, n2762, n2763, n2764, n2765, n2766, n2767, n2832, n2833, n2838, 
      n2839, n2840, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, 
      n2850, n2851, n2852, n2853, n2854, n2858, n2859, n2861, n2862, n2863, 
      n2864, n2865, n2867, n2875, n2878, n2883, n2886, n3154, n3160, n3204, 
      n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, 
      n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, 
      n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, 
      n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, 
      n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, 
      n3257, n3258, n3259, n3260, n3261, n3312, n3314, n3316, n3318, n3320, 
      n3322, n3324, n3326, n3328, n3330, n3332, n3334, n3336, n3338, n3340, 
      n3342, n3344, n3346, n3348, n3350, n3352, n3354, n3356, n3358, n3360, 
      n3362, n3364, n3366, n3368, n3370, n3372, n3379, n3382, n3383, n3384, 
      n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, 
      n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, 
      n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3417, n3420, 
      n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, 
      n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, 
      n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, 
      n3455, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, 
      n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, 
      n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, 
      n3487, n3488, n3493, n3496, n3497, n3498, n3499, n3500, n3501, n3502, 
      n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, 
      n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, 
      n3523, n3524, n3525, n3526, n3531, n3534, n3535, n3536, n3537, n3538, 
      n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, 
      n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, 
      n3559, n3560, n3561, n3562, n3563, n3564, n3569, n3572, n3573, n3574, 
      n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, 
      n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, 
      n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3607, n3610, 
      n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, 
      n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, 
      n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, 
      n3645, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, 
      n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, 
      n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, 
      n3677, n3678, n3682, n3685, n3686, n3687, n3688, n3689, n3690, n3691, 
      n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, 
      n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, 
      n3712, n3713, n3714, n3715, n3719, n3722, n3723, n3724, n3725, n3726, 
      n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, 
      n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, 
      n3747, n3748, n3749, n3750, n3751, n3752, n3756, n3759, n3760, n3761, 
      n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, 
      n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, 
      n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3791, n3794, 
      n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, 
      n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, 
      n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, 
      n3826, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, 
      n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, 
      n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, 
      n3858, n3859, n3861, n3864, n3865, n3866, n3867, n3868, n3869, n3870, 
      n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, 
      n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, 
      n3891, n3892, n3893, n3894, n3896, n3900, n3902, n3904, n3906, n3908, 
      n3910, n3912, n3914, n3916, n3918, n3920, n3922, n3924, n3926, n3928, 
      n3930, n3932, n3934, n3936, n3938, n3940, n3942, n3944, n3946, n3948, 
      n3950, n3952, n3954, n3956, n3958, n3960, n3964, n3968, n3970, n3972, 
      n3974, n3976, n3978, n3980, n3982, n3984, n3986, n3988, n3990, n3992, 
      n3994, n3996, n3998, n4000, n4002, n4004, n4006, n4008, n4010, n4012, 
      n4014, n4016, n4018, n4020, n4022, n4024, n4026, n4028, n4032, n4035, 
      n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, 
      n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, 
      n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, 
      n4067, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, 
      n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, 
      n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, 
      n4099, n4100, n4102, n4105, n4106, n4107, n4108, n4109, n4110, n4111, 
      n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, 
      n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, 
      n4132, n4133, n4134, n4135, n4137, n4140, n4141, n4142, n4143, n4144, 
      n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, 
      n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, 
      n4165, n4166, n4167, n4168, n4169, n4170, n4172, n4175, n4176, n4177, 
      n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, 
      n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, 
      n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4207, n4210, 
      n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, 
      n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, 
      n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, 
      n4242, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, 
      n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, 
      n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, 
      n4274, n4275, n4277, n4280, n4281, n4282, n4283, n4284, n4285, n4286, 
      n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, 
      n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, 
      n4307, n4308, n4309, n4310, n4312, n4315, n4316, n4317, n4318, n4319, 
      n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, 
      n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, 
      n4340, n4341, n4342, n4343, n4344, n4345, n4347, n4350, n4351, n4352, 
      n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, 
      n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, 
      n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4382, n4385, 
      n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, 
      n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, 
      n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, 
      n4417, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, 
      n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, 
      n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, 
      n4449, n4450, n4452, n4455, n4456, n4457, n4458, n4459, n4460, n4461, 
      n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, 
      n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, 
      n4482, n4483, n4484, n4485, n4487, n4490, n4491, n4492, n4493, n4494, 
      n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, 
      n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, 
      n4515, n4516, n4517, n4518, n4519, n4520, n4522, n4525, n4526, n4527, 
      n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, 
      n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, 
      n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4557, n4561, 
      n4563, n4565, n4567, n4569, n4571, n4573, n4575, n4577, n4579, n4581, 
      n4583, n4585, n4587, n4589, n4591, n4593, n4595, n4597, n4599, n4601, 
      n4603, n4605, n4607, n4609, n4611, n4613, n4615, n4617, n4619, n4621, 
      n4625, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, 
      n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, 
      n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, 
      n4657, n4658, n4660, n4663, n4664, n4665, n4666, n4667, n4668, n4669, 
      n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, 
      n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, 
      n4690, n4691, n4692, n4693, n4695, n4698, n4699, n4700, n4701, n4702, 
      n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, 
      n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, 
      n4723, n4724, n4725, n4726, n4727, n4728, n4730, n4733, n4734, n4735, 
      n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, 
      n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, 
      n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4765, n4768, 
      n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, 
      n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, 
      n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, 
      n4800, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, 
      n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, 
      n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, 
      n4832, n4833, n4835, n4838, n4839, n4840, n4841, n4842, n4843, n4844, 
      n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, 
      n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, 
      n4865, n4866, n4867, n4868, n4870, n4873, n4874, n4875, n4876, n4877, 
      n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, 
      n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, 
      n4898, n4899, n4900, n4901, n4902, n4903, n4905, n4908, n4909, n4910, 
      n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, 
      n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, 
      n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4940, n4943, 
      n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, 
      n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, 
      n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, 
      n4975, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, 
      n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, 
      n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, 
      n5007, n5008, n5010, n5013, n5014, n5015, n5016, n5017, n5018, n5019, 
      n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, 
      n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, 
      n5040, n5041, n5042, n5043, n5045, n5048, n5049, n5050, n5051, n5052, 
      n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, 
      n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, 
      n5073, n5074, n5075, n5076, n5077, n5078, n5080, n5083, n5084, n5085, 
      n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, 
      n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, 
      n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5115, n5118, 
      n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, 
      n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, 
      n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, 
      n5150, n5154, n5156, n5158, n5160, n5162, n5164, n5166, n5168, n5170, 
      n5172, n5174, n5176, n5178, n5180, n5182, n5184, n5186, n5188, n5190, 
      n5192, n5194, n5196, n5198, n5200, n5202, n5204, n5206, n5208, n5210, 
      n5212, n5214, n5217, n5220, n5221, n5222, n5223, n5224, n5225, n5226, 
      n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, 
      n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, 
      n5247, n5248, n5249, n5250, n5253, n5256, n5257, n5258, n5259, n5260, 
      n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, 
      n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, 
      n5281, n5282, n5283, n5284, n5285, n5286, n5288, n5291, n5292, n5293, 
      n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, 
      n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, 
      n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5323, n5326, 
      n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, 
      n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, 
      n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, 
      n5358, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, 
      n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, 
      n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, 
      n5390, n5391, n5393, n5396, n5397, n5398, n5399, n5400, n5401, n5402, 
      n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, 
      n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, 
      n5423, n5424, n5425, n5426, n5428, n5431, n5432, n5433, n5434, n5435, 
      n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, 
      n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, 
      n5456, n5457, n5458, n5459, n5460, n5461, n5463, n5466, n5467, n5468, 
      n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, 
      n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, 
      n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5498, n5501, 
      n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, 
      n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, 
      n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, 
      n5533, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, 
      n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, 
      n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, 
      n5565, n5566, n5568, n5571, n5572, n5573, n5574, n5575, n5576, n5577, 
      n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, 
      n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, 
      n5598, n5599, n5600, n5601, n5607, n5610, n5611, n5612, n5613, n5614, 
      n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, 
      n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, 
      n5635, n5636, n5637, n5638, n5639, n5640, n5644, n5647, n5648, n5649, 
      n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, 
      n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, 
      n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5681, n5684, 
      n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, 
      n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, 
      n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, 
      n5718, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, 
      n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, 
      n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, 
      n5750, n5751, n5755, n5758, n5759, n5760, n5761, n5762, n5763, n5764, 
      n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, 
      n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, 
      n5785, n5786, n5787, n5788, n5794, n5797, n5798, n5799, n5800, n5801, 
      n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, 
      n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, 
      n5822, n5823, n5824, n5825, n5826, n5827, n5830, n5833, n5834, n5835, 
      n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, 
      n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, 
      n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5866, n5869, 
      n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, 
      n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, 
      n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, 
      n5902, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, 
      n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, 
      n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, 
      n5934, n5935, n5938, n5941, n5942, n5943, n5944, n5945, n5946, n5947, 
      n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, 
      n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, 
      n5968, n5969, n5970, n5971, n5974, n5977, n5978, n5979, n5980, n5981, 
      n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, 
      n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, 
      n6002, n6003, n6004, n6005, n6006, n6007, n6010, n6013, n6014, n6015, 
      n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, 
      n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, 
      n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6047, n6050, 
      n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, 
      n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, 
      n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, 
      n6083, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, 
      n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, 
      n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, 
      n6115, n6116, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, 
      n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6692, n6728, 
      n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6768, n6769, n6770, 
      n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, 
      n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, 
      n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, 
      n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, 
      n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, 
      n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, 
      n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, 
      n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, 
      n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, 
      n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, 
      n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, 
      n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, 
      n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, 
      n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, 
      n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, 
      n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, 
      n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, 
      n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, 
      n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, 
      n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, 
      n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, 
      n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, 
      n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, 
      n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, 
      n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, 
      n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, 
      n7031, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, 
      n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, 
      n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, 
      n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, 
      n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, 
      n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, 
      n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7116, n7117, n7118, 
      n7119, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, 
      n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, 
      n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, 
      n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, 
      n7160, n7162, n7164, n7165, n7166, intadd_1_B_2_port, intadd_1_B_1_port, 
      intadd_1_B_0_port, intadd_1_n27, intadd_1_n26, intadd_1_n23, intadd_1_n22
      , intadd_1_n21, intadd_1_n20, intadd_1_n18, intadd_1_n17, intadd_1_n16, 
      intadd_1_n15, intadd_1_n14, intadd_1_n13, intadd_1_n12, intadd_1_n6, 
      intadd_1_n3, intadd_1_n2, intadd_1_n1, intadd_0_B_3_port, 
      intadd_0_B_2_port, intadd_0_B_1_port, intadd_0_B_0_port, 
      intadd_0_SUM_1_port, intadd_0_CO, intadd_0_n23, intadd_0_n22, 
      intadd_0_n21, intadd_0_n19, intadd_0_n18, intadd_0_n17, intadd_0_n16, 
      intadd_0_n15, intadd_0_n14, intadd_0_n13, intadd_0_n12, intadd_0_n11, 
      intadd_0_n10, intadd_0_n9, intadd_0_n8, intadd_0_n7, intadd_0_n6, 
      intadd_0_n3, intadd_0_n2, intadd_0_n1, DP_OP_1091J1_126_6973_n75, 
      DP_OP_1091J1_126_6973_n72, DP_OP_1091J1_126_6973_n31, 
      DP_OP_1091J1_126_6973_n29, DP_OP_1091J1_126_6973_n28, 
      DP_OP_1091J1_126_6973_n27, DP_OP_1091J1_126_6973_n26, 
      DP_OP_1091J1_126_6973_n25, DP_OP_1091J1_126_6973_n23, 
      DP_OP_1091J1_126_6973_n22, DP_OP_1091J1_126_6973_n21, 
      DP_OP_1091J1_126_6973_n20, DP_OP_1091J1_126_6973_n19, 
      DP_OP_1091J1_126_6973_n18, DP_OP_1091J1_126_6973_n17, 
      DP_OP_1091J1_126_6973_n16, DP_OP_1091J1_126_6973_n15, 
      DP_OP_1091J1_126_6973_n14, DP_OP_1091J1_126_6973_n13, 
      DP_OP_1091J1_126_6973_n12, DP_OP_1091J1_126_6973_n11, 
      DP_OP_1091J1_126_6973_n10, DP_OP_1091J1_126_6973_n6, 
      DP_OP_751_130_6421_I2, DP_OP_751_130_6421_n1795, DP_OP_751_130_6421_n1794
      , DP_OP_751_130_6421_n1791, DP_OP_751_130_6421_n1790, 
      DP_OP_751_130_6421_n1787, DP_OP_751_130_6421_n1785, 
      DP_OP_751_130_6421_n1783, DP_OP_751_130_6421_n1782, 
      DP_OP_751_130_6421_n1777, DP_OP_751_130_6421_n1774, 
      DP_OP_751_130_6421_n1772, DP_OP_751_130_6421_n1770, 
      DP_OP_751_130_6421_n1768, DP_OP_751_130_6421_n1765, 
      DP_OP_751_130_6421_n1764, DP_OP_751_130_6421_n1762, 
      DP_OP_751_130_6421_n1760, DP_OP_751_130_6421_n1759, 
      DP_OP_751_130_6421_n1756, DP_OP_751_130_6421_n1754, 
      DP_OP_751_130_6421_n1750, DP_OP_751_130_6421_n1748, 
      DP_OP_751_130_6421_n1746, DP_OP_751_130_6421_n1745, 
      DP_OP_751_130_6421_n1743, DP_OP_751_130_6421_n1742, 
      DP_OP_751_130_6421_n1739, DP_OP_751_130_6421_n1738, 
      DP_OP_751_130_6421_n1737, DP_OP_751_130_6421_n1736, 
      DP_OP_751_130_6421_n1735, DP_OP_751_130_6421_n1734, 
      DP_OP_751_130_6421_n1733, DP_OP_751_130_6421_n1731, 
      DP_OP_751_130_6421_n1729, DP_OP_751_130_6421_n1726, 
      DP_OP_751_130_6421_n1724, DP_OP_751_130_6421_n1720, 
      DP_OP_751_130_6421_n1715, DP_OP_751_130_6421_n1714, 
      DP_OP_751_130_6421_n1713, DP_OP_751_130_6421_n1712, 
      DP_OP_751_130_6421_n1711, DP_OP_751_130_6421_n1710, 
      DP_OP_751_130_6421_n1709, DP_OP_751_130_6421_n1708, 
      DP_OP_751_130_6421_n1707, DP_OP_751_130_6421_n1706, 
      DP_OP_751_130_6421_n1705, DP_OP_751_130_6421_n1703, 
      DP_OP_751_130_6421_n1698, DP_OP_751_130_6421_n1697, 
      DP_OP_751_130_6421_n1696, DP_OP_751_130_6421_n1695, 
      DP_OP_751_130_6421_n1694, DP_OP_751_130_6421_n1692, 
      DP_OP_751_130_6421_n1691, DP_OP_751_130_6421_n1690, 
      DP_OP_751_130_6421_n1689, DP_OP_751_130_6421_n1688, 
      DP_OP_751_130_6421_n1687, DP_OP_751_130_6421_n1686, 
      DP_OP_751_130_6421_n1685, DP_OP_751_130_6421_n1684, 
      DP_OP_751_130_6421_n1683, DP_OP_751_130_6421_n1682, 
      DP_OP_751_130_6421_n1681, DP_OP_751_130_6421_n1680, 
      DP_OP_751_130_6421_n1678, DP_OP_751_130_6421_n1677, 
      DP_OP_751_130_6421_n1676, DP_OP_751_130_6421_n1675, 
      DP_OP_751_130_6421_n1674, DP_OP_751_130_6421_n1673, 
      DP_OP_751_130_6421_n1672, DP_OP_751_130_6421_n1671, 
      DP_OP_751_130_6421_n1670, DP_OP_751_130_6421_n1669, 
      DP_OP_751_130_6421_n1668, DP_OP_751_130_6421_n1667, 
      DP_OP_751_130_6421_n1666, DP_OP_751_130_6421_n1665, 
      DP_OP_751_130_6421_n1664, DP_OP_751_130_6421_n1663, 
      DP_OP_751_130_6421_n1662, DP_OP_751_130_6421_n1661, 
      DP_OP_751_130_6421_n1660, DP_OP_751_130_6421_n1659, 
      DP_OP_751_130_6421_n1658, DP_OP_751_130_6421_n1657, 
      DP_OP_751_130_6421_n1655, DP_OP_751_130_6421_n1654, 
      DP_OP_751_130_6421_n1653, DP_OP_751_130_6421_n1652, 
      DP_OP_751_130_6421_n1651, DP_OP_751_130_6421_n1649, 
      DP_OP_751_130_6421_n1647, DP_OP_751_130_6421_n1646, 
      DP_OP_751_130_6421_n1645, DP_OP_751_130_6421_n1644, 
      DP_OP_751_130_6421_n1643, DP_OP_751_130_6421_n1642, 
      DP_OP_751_130_6421_n1641, DP_OP_751_130_6421_n1640, 
      DP_OP_751_130_6421_n1639, DP_OP_751_130_6421_n1638, 
      DP_OP_751_130_6421_n1629, DP_OP_751_130_6421_n1627, 
      DP_OP_751_130_6421_n1626, DP_OP_751_130_6421_n1625, 
      DP_OP_751_130_6421_n1624, DP_OP_751_130_6421_n1623, 
      DP_OP_751_130_6421_n1622, DP_OP_751_130_6421_n1621, 
      DP_OP_751_130_6421_n1620, DP_OP_751_130_6421_n1619, 
      DP_OP_751_130_6421_n1618, DP_OP_751_130_6421_n1617, 
      DP_OP_751_130_6421_n1616, DP_OP_751_130_6421_n1615, 
      DP_OP_751_130_6421_n1614, DP_OP_751_130_6421_n1613, 
      DP_OP_751_130_6421_n1612, DP_OP_751_130_6421_n1611, 
      DP_OP_751_130_6421_n1610, DP_OP_751_130_6421_n1609, 
      DP_OP_751_130_6421_n1608, DP_OP_751_130_6421_n1607, 
      DP_OP_751_130_6421_n1606, DP_OP_751_130_6421_n1605, 
      DP_OP_751_130_6421_n1604, DP_OP_751_130_6421_n1603, 
      DP_OP_751_130_6421_n1602, DP_OP_751_130_6421_n1601, 
      DP_OP_751_130_6421_n1594, DP_OP_751_130_6421_n1593, 
      DP_OP_751_130_6421_n1592, DP_OP_751_130_6421_n1591, 
      DP_OP_751_130_6421_n1590, DP_OP_751_130_6421_n1589, 
      DP_OP_751_130_6421_n1588, DP_OP_751_130_6421_n1587, 
      DP_OP_751_130_6421_n1586, DP_OP_751_130_6421_n1585, 
      DP_OP_751_130_6421_n1584, DP_OP_751_130_6421_n1583, 
      DP_OP_751_130_6421_n1582, DP_OP_751_130_6421_n1581, 
      DP_OP_751_130_6421_n1580, DP_OP_751_130_6421_n1579, 
      DP_OP_751_130_6421_n1578, DP_OP_751_130_6421_n1577, 
      DP_OP_751_130_6421_n1576, DP_OP_751_130_6421_n1575, 
      DP_OP_751_130_6421_n1574, DP_OP_751_130_6421_n1573, 
      DP_OP_751_130_6421_n1572, DP_OP_751_130_6421_n1571, 
      DP_OP_751_130_6421_n1570, DP_OP_751_130_6421_n1569, 
      DP_OP_751_130_6421_n1567, DP_OP_751_130_6421_n1566, 
      DP_OP_751_130_6421_n1565, DP_OP_751_130_6421_n1564, 
      DP_OP_751_130_6421_n1563, DP_OP_751_130_6421_n1562, 
      DP_OP_751_130_6421_n1561, DP_OP_751_130_6421_n1559, 
      DP_OP_751_130_6421_n1558, DP_OP_751_130_6421_n1557, 
      DP_OP_751_130_6421_n1556, DP_OP_751_130_6421_n1555, 
      DP_OP_751_130_6421_n1554, DP_OP_751_130_6421_n1553, 
      DP_OP_751_130_6421_n1551, DP_OP_751_130_6421_n1550, 
      DP_OP_751_130_6421_n1549, DP_OP_751_130_6421_n1548, 
      DP_OP_751_130_6421_n1547, DP_OP_751_130_6421_n1546, 
      DP_OP_751_130_6421_n1545, DP_OP_751_130_6421_n1543, 
      DP_OP_751_130_6421_n1542, DP_OP_751_130_6421_n1541, 
      DP_OP_751_130_6421_n1540, DP_OP_751_130_6421_n1527, 
      DP_OP_751_130_6421_n1526, DP_OP_751_130_6421_n1525, 
      DP_OP_751_130_6421_n1524, DP_OP_751_130_6421_n1523, 
      DP_OP_751_130_6421_n1522, DP_OP_751_130_6421_n1521, 
      DP_OP_751_130_6421_n1520, DP_OP_751_130_6421_n1519, 
      DP_OP_751_130_6421_n1518, DP_OP_751_130_6421_n1517, 
      DP_OP_751_130_6421_n1516, DP_OP_751_130_6421_n1515, 
      DP_OP_751_130_6421_n1514, DP_OP_751_130_6421_n1513, 
      DP_OP_751_130_6421_n1512, DP_OP_751_130_6421_n1511, 
      DP_OP_751_130_6421_n1510, DP_OP_751_130_6421_n1509, 
      DP_OP_751_130_6421_n1508, DP_OP_751_130_6421_n1507, 
      DP_OP_751_130_6421_n1506, DP_OP_751_130_6421_n1505, 
      DP_OP_751_130_6421_n1504, DP_OP_751_130_6421_n1503, 
      DP_OP_751_130_6421_n1502, DP_OP_751_130_6421_n1501, 
      DP_OP_751_130_6421_n1492, DP_OP_751_130_6421_n1491, 
      DP_OP_751_130_6421_n1490, DP_OP_751_130_6421_n1489, 
      DP_OP_751_130_6421_n1488, DP_OP_751_130_6421_n1487, 
      DP_OP_751_130_6421_n1486, DP_OP_751_130_6421_n1485, 
      DP_OP_751_130_6421_n1484, DP_OP_751_130_6421_n1483, 
      DP_OP_751_130_6421_n1482, DP_OP_751_130_6421_n1481, 
      DP_OP_751_130_6421_n1480, DP_OP_751_130_6421_n1479, 
      DP_OP_751_130_6421_n1478, DP_OP_751_130_6421_n1477, 
      DP_OP_751_130_6421_n1476, DP_OP_751_130_6421_n1475, 
      DP_OP_751_130_6421_n1474, DP_OP_751_130_6421_n1473, 
      DP_OP_751_130_6421_n1472, DP_OP_751_130_6421_n1471, 
      DP_OP_751_130_6421_n1470, DP_OP_751_130_6421_n1469, 
      DP_OP_751_130_6421_n1468, DP_OP_751_130_6421_n1467, 
      DP_OP_751_130_6421_n1466, DP_OP_751_130_6421_n1465, 
      DP_OP_751_130_6421_n1464, DP_OP_751_130_6421_n1463, 
      DP_OP_751_130_6421_n1462, DP_OP_751_130_6421_n1461, 
      DP_OP_751_130_6421_n1460, DP_OP_751_130_6421_n1459, 
      DP_OP_751_130_6421_n1458, DP_OP_751_130_6421_n1457, 
      DP_OP_751_130_6421_n1456, DP_OP_751_130_6421_n1455, 
      DP_OP_751_130_6421_n1454, DP_OP_751_130_6421_n1453, 
      DP_OP_751_130_6421_n1452, DP_OP_751_130_6421_n1451, 
      DP_OP_751_130_6421_n1449, DP_OP_751_130_6421_n1448, 
      DP_OP_751_130_6421_n1447, DP_OP_751_130_6421_n1445, 
      DP_OP_751_130_6421_n1444, DP_OP_751_130_6421_n1443, 
      DP_OP_751_130_6421_n1442, DP_OP_751_130_6421_n1425, 
      DP_OP_751_130_6421_n1423, DP_OP_751_130_6421_n1422, 
      DP_OP_751_130_6421_n1421, DP_OP_751_130_6421_n1420, 
      DP_OP_751_130_6421_n1419, DP_OP_751_130_6421_n1418, 
      DP_OP_751_130_6421_n1417, DP_OP_751_130_6421_n1416, 
      DP_OP_751_130_6421_n1415, DP_OP_751_130_6421_n1414, 
      DP_OP_751_130_6421_n1413, DP_OP_751_130_6421_n1412, 
      DP_OP_751_130_6421_n1411, DP_OP_751_130_6421_n1410, 
      DP_OP_751_130_6421_n1409, DP_OP_751_130_6421_n1408, 
      DP_OP_751_130_6421_n1407, DP_OP_751_130_6421_n1406, 
      DP_OP_751_130_6421_n1405, DP_OP_751_130_6421_n1404, 
      DP_OP_751_130_6421_n1403, DP_OP_751_130_6421_n1402, 
      DP_OP_751_130_6421_n1401, DP_OP_751_130_6421_n1390, 
      DP_OP_751_130_6421_n1389, DP_OP_751_130_6421_n1388, 
      DP_OP_751_130_6421_n1387, DP_OP_751_130_6421_n1386, 
      DP_OP_751_130_6421_n1385, DP_OP_751_130_6421_n1384, 
      DP_OP_751_130_6421_n1383, DP_OP_751_130_6421_n1382, 
      DP_OP_751_130_6421_n1381, DP_OP_751_130_6421_n1380, 
      DP_OP_751_130_6421_n1379, DP_OP_751_130_6421_n1378, 
      DP_OP_751_130_6421_n1377, DP_OP_751_130_6421_n1376, 
      DP_OP_751_130_6421_n1375, DP_OP_751_130_6421_n1374, 
      DP_OP_751_130_6421_n1373, DP_OP_751_130_6421_n1372, 
      DP_OP_751_130_6421_n1371, DP_OP_751_130_6421_n1370, 
      DP_OP_751_130_6421_n1369, DP_OP_751_130_6421_n1368, 
      DP_OP_751_130_6421_n1367, DP_OP_751_130_6421_n1366, 
      DP_OP_751_130_6421_n1365, DP_OP_751_130_6421_n1364, 
      DP_OP_751_130_6421_n1363, DP_OP_751_130_6421_n1362, 
      DP_OP_751_130_6421_n1361, DP_OP_751_130_6421_n1360, 
      DP_OP_751_130_6421_n1359, DP_OP_751_130_6421_n1358, 
      DP_OP_751_130_6421_n1357, DP_OP_751_130_6421_n1356, 
      DP_OP_751_130_6421_n1355, DP_OP_751_130_6421_n1354, 
      DP_OP_751_130_6421_n1353, DP_OP_751_130_6421_n1352, 
      DP_OP_751_130_6421_n1351, DP_OP_751_130_6421_n1350, 
      DP_OP_751_130_6421_n1349, DP_OP_751_130_6421_n1348, 
      DP_OP_751_130_6421_n1347, DP_OP_751_130_6421_n1346, 
      DP_OP_751_130_6421_n1345, DP_OP_751_130_6421_n1344, 
      DP_OP_751_130_6421_n1323, DP_OP_751_130_6421_n1321, 
      DP_OP_751_130_6421_n1320, DP_OP_751_130_6421_n1319, 
      DP_OP_751_130_6421_n1318, DP_OP_751_130_6421_n1317, 
      DP_OP_751_130_6421_n1316, DP_OP_751_130_6421_n1315, 
      DP_OP_751_130_6421_n1314, DP_OP_751_130_6421_n1313, 
      DP_OP_751_130_6421_n1312, DP_OP_751_130_6421_n1311, 
      DP_OP_751_130_6421_n1310, DP_OP_751_130_6421_n1309, 
      DP_OP_751_130_6421_n1308, DP_OP_751_130_6421_n1307, 
      DP_OP_751_130_6421_n1306, DP_OP_751_130_6421_n1305, 
      DP_OP_751_130_6421_n1304, DP_OP_751_130_6421_n1303, 
      DP_OP_751_130_6421_n1302, DP_OP_751_130_6421_n1301, 
      DP_OP_751_130_6421_n1288, DP_OP_751_130_6421_n1287, 
      DP_OP_751_130_6421_n1286, DP_OP_751_130_6421_n1285, 
      DP_OP_751_130_6421_n1284, DP_OP_751_130_6421_n1283, 
      DP_OP_751_130_6421_n1282, DP_OP_751_130_6421_n1281, 
      DP_OP_751_130_6421_n1280, DP_OP_751_130_6421_n1279, 
      DP_OP_751_130_6421_n1278, DP_OP_751_130_6421_n1277, 
      DP_OP_751_130_6421_n1276, DP_OP_751_130_6421_n1275, 
      DP_OP_751_130_6421_n1274, DP_OP_751_130_6421_n1273, 
      DP_OP_751_130_6421_n1272, DP_OP_751_130_6421_n1271, 
      DP_OP_751_130_6421_n1270, DP_OP_751_130_6421_n1269, 
      DP_OP_751_130_6421_n1268, DP_OP_751_130_6421_n1267, 
      DP_OP_751_130_6421_n1266, DP_OP_751_130_6421_n1265, 
      DP_OP_751_130_6421_n1264, DP_OP_751_130_6421_n1263, 
      DP_OP_751_130_6421_n1262, DP_OP_751_130_6421_n1261, 
      DP_OP_751_130_6421_n1260, DP_OP_751_130_6421_n1259, 
      DP_OP_751_130_6421_n1258, DP_OP_751_130_6421_n1257, 
      DP_OP_751_130_6421_n1256, DP_OP_751_130_6421_n1255, 
      DP_OP_751_130_6421_n1253, DP_OP_751_130_6421_n1252, 
      DP_OP_751_130_6421_n1251, DP_OP_751_130_6421_n1250, 
      DP_OP_751_130_6421_n1249, DP_OP_751_130_6421_n1248, 
      DP_OP_751_130_6421_n1247, DP_OP_751_130_6421_n1246, 
      DP_OP_751_130_6421_n1221, DP_OP_751_130_6421_n1220, 
      DP_OP_751_130_6421_n1219, DP_OP_751_130_6421_n1218, 
      DP_OP_751_130_6421_n1217, DP_OP_751_130_6421_n1216, 
      DP_OP_751_130_6421_n1215, DP_OP_751_130_6421_n1214, 
      DP_OP_751_130_6421_n1213, DP_OP_751_130_6421_n1212, 
      DP_OP_751_130_6421_n1211, DP_OP_751_130_6421_n1210, 
      DP_OP_751_130_6421_n1209, DP_OP_751_130_6421_n1208, 
      DP_OP_751_130_6421_n1207, DP_OP_751_130_6421_n1206, 
      DP_OP_751_130_6421_n1205, DP_OP_751_130_6421_n1204, 
      DP_OP_751_130_6421_n1203, DP_OP_751_130_6421_n1202, 
      DP_OP_751_130_6421_n1201, DP_OP_751_130_6421_n1186, 
      DP_OP_751_130_6421_n1185, DP_OP_751_130_6421_n1184, 
      DP_OP_751_130_6421_n1183, DP_OP_751_130_6421_n1182, 
      DP_OP_751_130_6421_n1181, DP_OP_751_130_6421_n1180, 
      DP_OP_751_130_6421_n1179, DP_OP_751_130_6421_n1178, 
      DP_OP_751_130_6421_n1177, DP_OP_751_130_6421_n1176, 
      DP_OP_751_130_6421_n1175, DP_OP_751_130_6421_n1174, 
      DP_OP_751_130_6421_n1173, DP_OP_751_130_6421_n1172, 
      DP_OP_751_130_6421_n1171, DP_OP_751_130_6421_n1170, 
      DP_OP_751_130_6421_n1169, DP_OP_751_130_6421_n1168, 
      DP_OP_751_130_6421_n1167, DP_OP_751_130_6421_n1166, 
      DP_OP_751_130_6421_n1165, DP_OP_751_130_6421_n1164, 
      DP_OP_751_130_6421_n1163, DP_OP_751_130_6421_n1162, 
      DP_OP_751_130_6421_n1161, DP_OP_751_130_6421_n1160, 
      DP_OP_751_130_6421_n1159, DP_OP_751_130_6421_n1158, 
      DP_OP_751_130_6421_n1157, DP_OP_751_130_6421_n1156, 
      DP_OP_751_130_6421_n1155, DP_OP_751_130_6421_n1154, 
      DP_OP_751_130_6421_n1153, DP_OP_751_130_6421_n1152, 
      DP_OP_751_130_6421_n1151, DP_OP_751_130_6421_n1150, 
      DP_OP_751_130_6421_n1149, DP_OP_751_130_6421_n1148, 
      DP_OP_751_130_6421_n1119, DP_OP_751_130_6421_n1118, 
      DP_OP_751_130_6421_n1117, DP_OP_751_130_6421_n1116, 
      DP_OP_751_130_6421_n1115, DP_OP_751_130_6421_n1114, 
      DP_OP_751_130_6421_n1113, DP_OP_751_130_6421_n1112, 
      DP_OP_751_130_6421_n1111, DP_OP_751_130_6421_n1110, 
      DP_OP_751_130_6421_n1109, DP_OP_751_130_6421_n1108, 
      DP_OP_751_130_6421_n1107, DP_OP_751_130_6421_n1106, 
      DP_OP_751_130_6421_n1105, DP_OP_751_130_6421_n1104, 
      DP_OP_751_130_6421_n1103, DP_OP_751_130_6421_n1102, 
      DP_OP_751_130_6421_n1101, DP_OP_751_130_6421_n1084, 
      DP_OP_751_130_6421_n1083, DP_OP_751_130_6421_n1082, 
      DP_OP_751_130_6421_n1081, DP_OP_751_130_6421_n1080, 
      DP_OP_751_130_6421_n1079, DP_OP_751_130_6421_n1078, 
      DP_OP_751_130_6421_n1077, DP_OP_751_130_6421_n1076, 
      DP_OP_751_130_6421_n1075, DP_OP_751_130_6421_n1074, 
      DP_OP_751_130_6421_n1073, DP_OP_751_130_6421_n1072, 
      DP_OP_751_130_6421_n1071, DP_OP_751_130_6421_n1070, 
      DP_OP_751_130_6421_n1069, DP_OP_751_130_6421_n1068, 
      DP_OP_751_130_6421_n1067, DP_OP_751_130_6421_n1066, 
      DP_OP_751_130_6421_n1065, DP_OP_751_130_6421_n1064, 
      DP_OP_751_130_6421_n1063, DP_OP_751_130_6421_n1062, 
      DP_OP_751_130_6421_n1061, DP_OP_751_130_6421_n1060, 
      DP_OP_751_130_6421_n1059, DP_OP_751_130_6421_n1058, 
      DP_OP_751_130_6421_n1057, DP_OP_751_130_6421_n1056, 
      DP_OP_751_130_6421_n1055, DP_OP_751_130_6421_n1054, 
      DP_OP_751_130_6421_n1053, DP_OP_751_130_6421_n1052, 
      DP_OP_751_130_6421_n1051, DP_OP_751_130_6421_n1050, 
      DP_OP_751_130_6421_n1017, DP_OP_751_130_6421_n1016, 
      DP_OP_751_130_6421_n1015, DP_OP_751_130_6421_n1014, 
      DP_OP_751_130_6421_n1013, DP_OP_751_130_6421_n1012, 
      DP_OP_751_130_6421_n1011, DP_OP_751_130_6421_n1010, 
      DP_OP_751_130_6421_n1009, DP_OP_751_130_6421_n1008, 
      DP_OP_751_130_6421_n1007, DP_OP_751_130_6421_n1006, 
      DP_OP_751_130_6421_n1005, DP_OP_751_130_6421_n1004, 
      DP_OP_751_130_6421_n1003, DP_OP_751_130_6421_n1002, 
      DP_OP_751_130_6421_n1001, DP_OP_751_130_6421_n982, 
      DP_OP_751_130_6421_n981, DP_OP_751_130_6421_n980, DP_OP_751_130_6421_n979
      , DP_OP_751_130_6421_n978, DP_OP_751_130_6421_n977, 
      DP_OP_751_130_6421_n976, DP_OP_751_130_6421_n975, DP_OP_751_130_6421_n974
      , DP_OP_751_130_6421_n973, DP_OP_751_130_6421_n972, 
      DP_OP_751_130_6421_n971, DP_OP_751_130_6421_n970, DP_OP_751_130_6421_n969
      , DP_OP_751_130_6421_n968, DP_OP_751_130_6421_n967, 
      DP_OP_751_130_6421_n966, DP_OP_751_130_6421_n965, DP_OP_751_130_6421_n964
      , DP_OP_751_130_6421_n963, DP_OP_751_130_6421_n962, 
      DP_OP_751_130_6421_n961, DP_OP_751_130_6421_n960, DP_OP_751_130_6421_n959
      , DP_OP_751_130_6421_n958, DP_OP_751_130_6421_n957, 
      DP_OP_751_130_6421_n956, DP_OP_751_130_6421_n955, DP_OP_751_130_6421_n954
      , DP_OP_751_130_6421_n953, DP_OP_751_130_6421_n952, 
      DP_OP_751_130_6421_n915, DP_OP_751_130_6421_n913, DP_OP_751_130_6421_n912
      , DP_OP_751_130_6421_n911, DP_OP_751_130_6421_n910, 
      DP_OP_751_130_6421_n909, DP_OP_751_130_6421_n908, DP_OP_751_130_6421_n907
      , DP_OP_751_130_6421_n906, DP_OP_751_130_6421_n905, 
      DP_OP_751_130_6421_n904, DP_OP_751_130_6421_n903, DP_OP_751_130_6421_n902
      , DP_OP_751_130_6421_n901, DP_OP_751_130_6421_n880, 
      DP_OP_751_130_6421_n879, DP_OP_751_130_6421_n878, DP_OP_751_130_6421_n877
      , DP_OP_751_130_6421_n876, DP_OP_751_130_6421_n875, 
      DP_OP_751_130_6421_n874, DP_OP_751_130_6421_n873, DP_OP_751_130_6421_n872
      , DP_OP_751_130_6421_n871, DP_OP_751_130_6421_n870, 
      DP_OP_751_130_6421_n869, DP_OP_751_130_6421_n868, DP_OP_751_130_6421_n867
      , DP_OP_751_130_6421_n866, DP_OP_751_130_6421_n865, 
      DP_OP_751_130_6421_n864, DP_OP_751_130_6421_n863, DP_OP_751_130_6421_n862
      , DP_OP_751_130_6421_n861, DP_OP_751_130_6421_n860, 
      DP_OP_751_130_6421_n859, DP_OP_751_130_6421_n858, DP_OP_751_130_6421_n857
      , DP_OP_751_130_6421_n856, DP_OP_751_130_6421_n855, 
      DP_OP_751_130_6421_n854, DP_OP_751_130_6421_n813, DP_OP_751_130_6421_n812
      , DP_OP_751_130_6421_n811, DP_OP_751_130_6421_n810, 
      DP_OP_751_130_6421_n809, DP_OP_751_130_6421_n808, DP_OP_751_130_6421_n807
      , DP_OP_751_130_6421_n806, DP_OP_751_130_6421_n805, 
      DP_OP_751_130_6421_n804, DP_OP_751_130_6421_n803, DP_OP_751_130_6421_n802
      , DP_OP_751_130_6421_n801, DP_OP_751_130_6421_n778, 
      DP_OP_751_130_6421_n777, DP_OP_751_130_6421_n776, DP_OP_751_130_6421_n775
      , DP_OP_751_130_6421_n774, DP_OP_751_130_6421_n773, 
      DP_OP_751_130_6421_n772, DP_OP_751_130_6421_n771, DP_OP_751_130_6421_n770
      , DP_OP_751_130_6421_n769, DP_OP_751_130_6421_n768, 
      DP_OP_751_130_6421_n767, DP_OP_751_130_6421_n766, DP_OP_751_130_6421_n765
      , DP_OP_751_130_6421_n764, DP_OP_751_130_6421_n763, 
      DP_OP_751_130_6421_n762, DP_OP_751_130_6421_n761, DP_OP_751_130_6421_n760
      , DP_OP_751_130_6421_n759, DP_OP_751_130_6421_n758, 
      DP_OP_751_130_6421_n757, DP_OP_751_130_6421_n756, DP_OP_751_130_6421_n711
      , DP_OP_751_130_6421_n710, DP_OP_751_130_6421_n709, 
      DP_OP_751_130_6421_n708, DP_OP_751_130_6421_n707, DP_OP_751_130_6421_n706
      , DP_OP_751_130_6421_n705, DP_OP_751_130_6421_n704, 
      DP_OP_751_130_6421_n703, DP_OP_751_130_6421_n702, DP_OP_751_130_6421_n701
      , DP_OP_751_130_6421_n676, DP_OP_751_130_6421_n675, 
      DP_OP_751_130_6421_n674, DP_OP_751_130_6421_n673, DP_OP_751_130_6421_n672
      , DP_OP_751_130_6421_n671, DP_OP_751_130_6421_n670, 
      DP_OP_751_130_6421_n669, DP_OP_751_130_6421_n668, DP_OP_751_130_6421_n667
      , DP_OP_751_130_6421_n666, DP_OP_751_130_6421_n665, 
      DP_OP_751_130_6421_n664, DP_OP_751_130_6421_n663, DP_OP_751_130_6421_n662
      , DP_OP_751_130_6421_n661, DP_OP_751_130_6421_n660, 
      DP_OP_751_130_6421_n659, DP_OP_751_130_6421_n658, DP_OP_751_130_6421_n609
      , DP_OP_751_130_6421_n608, DP_OP_751_130_6421_n607, 
      DP_OP_751_130_6421_n606, DP_OP_751_130_6421_n605, DP_OP_751_130_6421_n604
      , DP_OP_751_130_6421_n603, DP_OP_751_130_6421_n602, 
      DP_OP_751_130_6421_n601, DP_OP_751_130_6421_n574, DP_OP_751_130_6421_n573
      , DP_OP_751_130_6421_n572, DP_OP_751_130_6421_n571, 
      DP_OP_751_130_6421_n570, DP_OP_751_130_6421_n569, DP_OP_751_130_6421_n568
      , DP_OP_751_130_6421_n567, DP_OP_751_130_6421_n566, 
      DP_OP_751_130_6421_n565, DP_OP_751_130_6421_n564, DP_OP_751_130_6421_n563
      , DP_OP_751_130_6421_n562, DP_OP_751_130_6421_n561, 
      DP_OP_751_130_6421_n560, DP_OP_751_130_6421_n507, DP_OP_751_130_6421_n506
      , DP_OP_751_130_6421_n505, DP_OP_751_130_6421_n504, 
      DP_OP_751_130_6421_n503, DP_OP_751_130_6421_n502, DP_OP_751_130_6421_n501
      , DP_OP_751_130_6421_n472, DP_OP_751_130_6421_n471, 
      DP_OP_751_130_6421_n470, DP_OP_751_130_6421_n469, DP_OP_751_130_6421_n468
      , DP_OP_751_130_6421_n467, DP_OP_751_130_6421_n466, 
      DP_OP_751_130_6421_n465, DP_OP_751_130_6421_n464, DP_OP_751_130_6421_n463
      , DP_OP_751_130_6421_n462, DP_OP_751_130_6421_n405, 
      DP_OP_751_130_6421_n404, DP_OP_751_130_6421_n403, DP_OP_751_130_6421_n402
      , DP_OP_751_130_6421_n401, DP_OP_751_130_6421_n370, 
      DP_OP_751_130_6421_n369, DP_OP_751_130_6421_n368, DP_OP_751_130_6421_n367
      , DP_OP_751_130_6421_n366, DP_OP_751_130_6421_n365, 
      DP_OP_751_130_6421_n303, DP_OP_751_130_6421_n302, DP_OP_751_130_6421_n301
      , DP_OP_751_130_6421_n268, DP_OP_751_130_6421_n267, 
      DP_OP_751_130_6421_n193, DP_OP_751_130_6421_n190, DP_OP_751_130_6421_n183
      , DP_OP_751_130_6421_n181, DP_OP_751_130_6421_n179, 
      DP_OP_751_130_6421_n174, DP_OP_751_130_6421_n172, DP_OP_751_130_6421_n170
      , DP_OP_751_130_6421_n167, DP_OP_751_130_6421_n166, 
      DP_OP_751_130_6421_n165, DP_OP_751_130_6421_n163, DP_OP_751_130_6421_n162
      , DP_OP_751_130_6421_n161, DP_OP_751_130_6421_n160, 
      DP_OP_751_130_6421_n159, DP_OP_751_130_6421_n154, DP_OP_751_130_6421_n153
      , DP_OP_751_130_6421_n151, DP_OP_751_130_6421_n149, 
      DP_OP_751_130_6421_n148, DP_OP_751_130_6421_n147, DP_OP_751_130_6421_n146
      , DP_OP_751_130_6421_n145, DP_OP_751_130_6421_n143, 
      DP_OP_751_130_6421_n141, DP_OP_751_130_6421_n140, DP_OP_751_130_6421_n139
      , DP_OP_751_130_6421_n138, DP_OP_751_130_6421_n137, 
      DP_OP_751_130_6421_n132, DP_OP_751_130_6421_n131, DP_OP_751_130_6421_n129
      , DP_OP_751_130_6421_n127, DP_OP_751_130_6421_n126, 
      DP_OP_751_130_6421_n125, DP_OP_751_130_6421_n124, DP_OP_751_130_6421_n123
      , DP_OP_751_130_6421_n119, DP_OP_751_130_6421_n118, 
      DP_OP_751_130_6421_n117, DP_OP_751_130_6421_n116, DP_OP_751_130_6421_n115
      , DP_OP_751_130_6421_n113, DP_OP_751_130_6421_n111, 
      DP_OP_751_130_6421_n110, DP_OP_751_130_6421_n109, DP_OP_751_130_6421_n106
      , DP_OP_751_130_6421_n105, DP_OP_751_130_6421_n103, 
      DP_OP_751_130_6421_n99, DP_OP_751_130_6421_n98, DP_OP_751_130_6421_n97, 
      DP_OP_751_130_6421_n96, DP_OP_751_130_6421_n95, DP_OP_751_130_6421_n91, 
      DP_OP_751_130_6421_n90, DP_OP_751_130_6421_n89, DP_OP_751_130_6421_n88, 
      DP_OP_751_130_6421_n83, DP_OP_751_130_6421_n82, DP_OP_751_130_6421_n81, 
      DP_OP_751_130_6421_n80, DP_OP_751_130_6421_n79, DP_OP_751_130_6421_n74, 
      DP_OP_751_130_6421_n73, DP_OP_751_130_6421_n68, DP_OP_751_130_6421_n67, 
      DP_OP_751_130_6421_n66, DP_OP_751_130_6421_n64, DP_OP_751_130_6421_n63, 
      DP_OP_751_130_6421_n26, DP_OP_751_130_6421_n24, DP_OP_751_130_6421_n23, 
      DP_OP_751_130_6421_n20, DP_OP_751_130_6421_n19, DP_OP_751_130_6421_n18, 
      DP_OP_751_130_6421_n17, DP_OP_751_130_6421_n16, DP_OP_751_130_6421_n14, 
      DP_OP_751_130_6421_n13, DP_OP_751_130_6421_n10, DP_OP_751_130_6421_n9, 
      DP_OP_751_130_6421_n8, DP_OP_751_130_6421_n6, DP_OP_751_130_6421_n5, 
      DP_OP_751_130_6421_n4, n7187, n7188, n7189, n7190, n7191, n7192, n7193, 
      n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, 
      n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, 
      n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, 
      n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, 
      n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, 
      n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, 
      n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, 
      n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, 
      n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, 
      n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, 
      n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, 
      n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, 
      n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, 
      n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, 
      n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, 
      n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, 
      n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, 
      n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, 
      n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, 
      n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, 
      n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, 
      n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, 
      n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, 
      n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, 
      n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, 
      n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, 
      n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, 
      n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, 
      n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, 
      n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, 
      n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, 
      n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, 
      n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, 
      n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, 
      n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, 
      n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, 
      n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, 
      n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, 
      n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, 
      n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, 
      n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, 
      n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, 
      n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, 
      n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, 
      n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, 
      n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, 
      n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, 
      n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, 
      n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, 
      n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, 
      n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, 
      n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, 
      n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, 
      n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, 
      n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, 
      n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, 
      n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, 
      n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, 
      n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, 
      n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, 
      n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, 
      n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, 
      n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, 
      n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, 
      n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, 
      n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, 
      n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, 
      n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, 
      n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, 
      n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, 
      n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, 
      n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, 
      n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, 
      n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, 
      n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, 
      n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, 
      n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, 
      n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, 
      n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, 
      n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, 
      n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, 
      n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, 
      n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, 
      n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, 
      n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, 
      n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, 
      n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, 
      n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, 
      n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, 
      n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, 
      n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, 
      n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, 
      n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, 
      n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, 
      n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, 
      n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, 
      n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, 
      n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, 
      n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, 
      n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, 
      n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, 
      n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, 
      n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, 
      n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, 
      n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, 
      n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, 
      n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, 
      n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, 
      n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, 
      n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, 
      n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, 
      n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, 
      n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, 
      n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, 
      n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, 
      n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, 
      n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, 
      n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, 
      n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, 
      n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, 
      n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, 
      n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, 
      n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, 
      n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, 
      n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, 
      n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, 
      n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, 
      n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, 
      n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, 
      n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, 
      n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, 
      n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, 
      n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, 
      n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, 
      n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, 
      n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, 
      n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, 
      n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, 
      n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, 
      n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, 
      n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, 
      n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, 
      n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, 
      n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, 
      n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, 
      n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, 
      n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, 
      n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, 
      n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, 
      n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, 
      n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, 
      n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, 
      n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, 
      n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, 
      n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, 
      n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, 
      n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, 
      n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, 
      n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, 
      n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, 
      n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, 
      n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, 
      n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, 
      n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, 
      n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, 
      n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, 
      n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, 
      n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, 
      n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, 
      n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, 
      n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, 
      n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, 
      n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, 
      n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, 
      n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, 
      n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, 
      n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, 
      n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, 
      n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, 
      n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, 
      n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, 
      n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, 
      n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, 
      n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, 
      n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, 
      n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, 
      n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, 
      n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, 
      n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, 
      n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, 
      n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, 
      n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, 
      n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, 
      n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, 
      n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, 
      n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, 
      n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, 
      n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, 
      n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, 
      n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, 
      n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, 
      n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, 
      n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, 
      n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, 
      n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, 
      n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, 
      n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, 
      n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, 
      n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, 
      n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, 
      n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, 
      n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, 
      n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, 
      n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, 
      n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, 
      n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, 
      n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, 
      n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, 
      n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, 
      n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, 
      n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, 
      n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, 
      n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, 
      n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, 
      n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, 
      n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, 
      n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, 
      n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, 
      n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, 
      n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, 
      n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, 
      n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, 
      n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, 
      n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, 
      n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, 
      n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, 
      n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, 
      n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, 
      n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, 
      n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, 
      n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, 
      n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, 
      n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, 
      n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, 
      n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, 
      n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, 
      n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, 
      n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, 
      n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, 
      n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, 
      n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, 
      n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, 
      n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, 
      n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, 
      n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, 
      n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, 
      n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, 
      n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, 
      n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, 
      n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, 
      n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, 
      n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, 
      n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, 
      n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, 
      n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, 
      n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, 
      n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, 
      n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, 
      n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, 
      n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, 
      n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, 
      n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, 
      n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, 
      n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, 
      n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, 
      n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, 
      n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, 
      n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, 
      n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, 
      n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, 
      n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
      n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, 
      n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, 
      n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, 
      n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, 
      n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, 
      n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, 
      n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, 
      n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, 
      n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, 
      n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, 
      n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, 
      n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, 
      n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, 
      n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, 
      n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, 
      n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, 
      n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, 
      n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, 
      n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174, 
      n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183, 
      n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, 
      n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201, 
      n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210, 
      n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, 
      n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228, 
      n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237, 
      n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246, 
      n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255, 
      n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264, 
      n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273, 
      n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282, 
      n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291, 
      n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300, 
      n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309, 
      n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318, 
      n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327, 
      n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336, 
      n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, 
      n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354, 
      n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363, 
      n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372, 
      n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381, 
      n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390, 
      n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399, 
      n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, 
      n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, 
      n10418, n10419, n10420, n10421, n10422, n10423, DRAMRF_ADDRESS_0_port, 
      n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433, 
      n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442, 
      n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451, 
      n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460, 
      n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469, 
      n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478, 
      n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487, 
      n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496, 
      n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505, 
      n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514, 
      n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523, 
      n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532, 
      n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541, 
      n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550, 
      n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559, 
      n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568, 
      n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577, 
      n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586, 
      n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595, 
      n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604, 
      n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613, 
      n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622, 
      n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631, 
      n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640, 
      n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649, 
      n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658, 
      n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667, 
      n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676, 
      n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685, 
      n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694, 
      n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703, 
      n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712, 
      n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721, 
      n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730, 
      n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739, 
      n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748, 
      n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757, 
      n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766, 
      n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, 
      n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, 
      n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, 
      n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802, 
      n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811, 
      n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820, 
      n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829, 
      n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838, 
      n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847, 
      n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856, 
      n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865, 
      n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874, 
      n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883, 
      n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892, 
      n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901, 
      n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910, 
      n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919, 
      n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928, 
      n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937, 
      n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946, 
      n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955, 
      n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964, 
      n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973, 
      n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982, 
      n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991, 
      n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000, 
      n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009, 
      n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018, 
      n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027, 
      n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036, 
      n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045, 
      n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054, 
      n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063, 
      n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072, 
      n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081, 
      n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090, 
      n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099, 
      n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108, 
      n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117, 
      n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126, 
      n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135, 
      n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144, 
      n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153, 
      n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162, 
      n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171, 
      n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180, 
      n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189, 
      n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198, 
      n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207, 
      n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216, 
      n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225, 
      n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234, 
      n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243, 
      n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252, 
      n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261, 
      n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270, 
      n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279, 
      n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288, 
      n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297, 
      n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306, 
      n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315, 
      n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324, 
      n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333, 
      n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342, 
      n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351, 
      n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360, 
      n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369, 
      n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378, 
      n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387, 
      n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396, 
      n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, 
      n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, 
      n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, 
      n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432, 
      n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441, 
      n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450, 
      n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459, 
      n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468, 
      n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477, 
      n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486, 
      n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495, 
      n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504, 
      n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513, 
      n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522, 
      n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, 
      n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540, 
      n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549, 
      n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558, 
      n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567, 
      n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576, 
      n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585, 
      n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594, 
      n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603, 
      n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612, 
      n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621, 
      n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630, 
      n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639, 
      n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648, 
      n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657, 
      n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666, 
      n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675, 
      n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684, 
      n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693, 
      n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, 
      n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, 
      n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, 
      n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, 
      n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, 
      n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, 
      n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, 
      n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, 
      n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, 
      n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, 
      n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, 
      n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, 
      n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810, 
      n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819, 
      n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828, 
      n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837, 
      n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846, 
      n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855, 
      n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, 
      n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, 
      n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, 
      n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, 
      n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, 
      n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909, 
      n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918, 
      n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927, 
      n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936, 
      n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945, 
      n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954, 
      n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963, 
      n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972, 
      n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981, 
      n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990, 
      n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999, 
      n12000, n12001, n12002, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, 
      n_1071, n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, 
      n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, 
      n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, 
      n_1098, n_1099, n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, 
      n_1107, n_1108, n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, 
      n_1116, n_1117, n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, 
      n_1125, n_1126, n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, 
      n_1134, n_1135, n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, 
      n_1143, n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, 
      n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, 
      n_1161, n_1162, n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, 
      n_1170, n_1171, n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, 
      n_1179, n_1180, n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, 
      n_1188, n_1189, n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, 
      n_1197, n_1198, n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, 
      n_1206, n_1207, n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, 
      n_1215, n_1216, n_1217, n_1218, n_1219, n_1220, n_1221, n_1222, n_1223, 
      n_1224, n_1225, n_1226, n_1227, n_1228, n_1229, n_1230, n_1231, n_1232, 
      n_1233, n_1234, n_1235, n_1236, n_1237, n_1238, n_1239, n_1240, n_1241, 
      n_1242, n_1243, n_1244, n_1245, n_1246, n_1247, n_1248, n_1249, n_1250, 
      n_1251, n_1252, n_1253, n_1254, n_1255, n_1256, n_1257, n_1258, n_1259, 
      n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, 
      n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, 
      n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, 
      n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, 
      n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, 
      n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, 
      n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, 
      n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, 
      n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, 
      n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, 
      n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357, n_1358, 
      n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365, n_1366, n_1367, 
      n_1368, n_1369, n_1370, n_1371, n_1372, n_1373, n_1374, n_1375, n_1376, 
      n_1377, n_1378, n_1379, n_1380, n_1381, n_1382, n_1383, n_1384, n_1385, 
      n_1386, n_1387, n_1388, n_1389, n_1390, n_1391, n_1392, n_1393, n_1394, 
      n_1395, n_1396, n_1397, n_1398, n_1399, n_1400, n_1401, n_1402, n_1403, 
      n_1404, n_1405, n_1406, n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, 
      n_1413, n_1414, n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, 
      n_1422, n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1429, n_1430, 
      n_1431, n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1439, 
      n_1440, n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448, 
      n_1449, n_1450, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457, 
      n_1458, n_1459, n_1460, n_1461, n_1462, n_1463, n_1464, n_1465, n_1466, 
      n_1467, n_1468, n_1469, n_1470, n_1471, n_1472, n_1473, n_1474, n_1475, 
      n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483, n_1484, 
      n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492, n_1493, 
      n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501, n_1502, 
      n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510, n_1511, 
      n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519, n_1520, 
      n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528, n_1529, 
      n_1530, n_1531, n_1532, n_1533, n_1534, n_1535, n_1536, n_1537, n_1538, 
      n_1539, n_1540, n_1541, n_1542, n_1543, n_1544, n_1545, n_1546, n_1547, 
      n_1548, n_1549, n_1550, n_1551, n_1552, n_1553, n_1554, n_1555, n_1556, 
      n_1557, n_1558, n_1559, n_1560, n_1561, n_1562, n_1563, n_1564, n_1565, 
      n_1566, n_1567, n_1568, n_1569, n_1570, n_1571, n_1572, n_1573, n_1574, 
      n_1575, n_1576, n_1577, n_1578, n_1579, n_1580, n_1581, n_1582, n_1583, 
      n_1584, n_1585, n_1586, n_1587, n_1588, n_1589, n_1590, n_1591, n_1592, 
      n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599, n_1600, n_1601, 
      n_1602, n_1603, n_1604, n_1605, n_1606, n_1607, n_1608, n_1609, n_1610, 
      n_1611, n_1612, n_1613, n_1614, n_1615, n_1616, n_1617, n_1618, n_1619, 
      n_1620, n_1621, n_1622, n_1623, n_1624, n_1625, n_1626, n_1627, n_1628, 
      n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, 
      n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, 
      n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, 
      n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, 
      n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, 
      n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, 
      n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, 
      n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, 
      n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, 
      n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, 
      n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, 
      n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, 
      n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, 
      n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, 
      n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, 
      n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, 
      n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, 
      n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, 
      n_1791, n_1792, n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, 
      n_1800, n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808, 
      n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816, n_1817, 
      n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824, n_1825, n_1826, 
      n_1827, n_1828, n_1829, n_1830, n_1831, n_1832, n_1833, n_1834, n_1835, 
      n_1836, n_1837, n_1838, n_1839, n_1840, n_1841, n_1842, n_1843, n_1844, 
      n_1845, n_1846, n_1847, n_1848, n_1849, n_1850, n_1851, n_1852, n_1853, 
      n_1854, n_1855, n_1856, n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, 
      n_1863, n_1864, n_1865, n_1866, n_1867, n_1868, n_1869, n_1870, n_1871, 
      n_1872, n_1873, n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, 
      n_1881, n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889, 
      n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897, n_1898, 
      n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905, n_1906, n_1907, 
      n_1908, n_1909, n_1910, n_1911, n_1912, n_1913, n_1914, n_1915, n_1916, 
      n_1917, n_1918, n_1919, n_1920, n_1921, n_1922, n_1923, n_1924, n_1925, 
      n_1926, n_1927, n_1928, n_1929, n_1930, n_1931, n_1932, n_1933, n_1934, 
      n_1935, n_1936, n_1937, n_1938, n_1939, n_1940, n_1941, n_1942, n_1943, 
      n_1944, n_1945, n_1946, n_1947, n_1948, n_1949, n_1950, n_1951, n_1952, 
      n_1953, n_1954, n_1955, n_1956, n_1957, n_1958, n_1959, n_1960, n_1961, 
      n_1962, n_1963, n_1964, n_1965, n_1966, n_1967, n_1968, n_1969, n_1970, 
      n_1971, n_1972, n_1973, n_1974, n_1975, n_1976, n_1977, n_1978, n_1979, 
      n_1980, n_1981, n_1982, n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, 
      n_1989, n_1990, n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, 
      n_1998, n_1999, n_2000, n_2001, n_2002, n_2003, n_2004, n_2005, n_2006, 
      n_2007, n_2008, n_2009, n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, 
      n_2016, n_2017, n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, 
      n_2025, n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033, 
      n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041, n_2042, 
      n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2049, n_2050, n_2051, 
      n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058, n_2059, n_2060, 
      n_2061, n_2062, n_2063, n_2064, n_2065, n_2066, n_2067, n_2068, n_2069, 
      n_2070, n_2071, n_2072, n_2073, n_2074, n_2075, n_2076, n_2077, n_2078, 
      n_2079, n_2080, n_2081, n_2082, n_2083, n_2084, n_2085, n_2086, n_2087, 
      n_2088, n_2089, n_2090, n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, 
      n_2097, n_2098, n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, 
      n_2106, n_2107, n_2108, n_2109, n_2110, n_2111, n_2112, n_2113, n_2114, 
      n_2115, n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123, 
      n_2124, n_2125, n_2126, n_2127, n_2128, n_2129, n_2130, n_2131, n_2132, 
      n_2133, n_2134, n_2135, n_2136, n_2137, n_2138, n_2139, n_2140, n_2141, 
      n_2142, n_2143, n_2144, n_2145, n_2146, n_2147, n_2148, n_2149, n_2150, 
      n_2151, n_2152, n_2153, n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, 
      n_2160, n_2161, n_2162, n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, 
      n_2169, n_2170, n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, 
      n_2178, n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186, 
      n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194, n_2195, 
      n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202, n_2203, n_2204, 
      n_2205, n_2206, n_2207, n_2208, n_2209, n_2210, n_2211, n_2212, n_2213, 
      n_2214, n_2215, n_2216, n_2217, n_2218, n_2219, n_2220, n_2221, n_2222, 
      n_2223, n_2224, n_2225, n_2226, n_2227, n_2228, n_2229, n_2230, n_2231, 
      n_2232, n_2233, n_2234, n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, 
      n_2241, n_2242, n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, 
      n_2250, n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258, 
      n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266, n_2267, 
      n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274, n_2275, n_2276, 
      n_2277, n_2278, n_2279, n_2280, n_2281, n_2282, n_2283, n_2284, n_2285, 
      n_2286, n_2287, n_2288, n_2289, n_2290, n_2291, n_2292, n_2293, n_2294, 
      n_2295, n_2296, n_2297, n_2298, n_2299, n_2300, n_2301, n_2302, n_2303, 
      n_2304, n_2305, n_2306, n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, 
      n_2313, n_2314, n_2315, n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, 
      n_2322, n_2323, n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, 
      n_2331, n_2332, n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, 
      n_2340, n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348, 
      n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356, n_2357, 
      n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364, n_2365, n_2366, 
      n_2367, n_2368, n_2369, n_2370, n_2371, n_2372, n_2373, n_2374, n_2375, 
      n_2376, n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384, 
      n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392, n_2393, 
      n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400, n_2401, n_2402, 
      n_2403, n_2404, n_2405, n_2406, n_2407, n_2408, n_2409, n_2410, n_2411, 
      n_2412, n_2413, n_2414, n_2415, n_2416, n_2417, n_2418, n_2419, n_2420, 
      n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427, n_2428, n_2429, 
      n_2430, n_2431, n_2432, n_2433, n_2434, n_2435, n_2436, n_2437, n_2438, 
      n_2439, n_2440, n_2441, n_2442, n_2443, n_2444, n_2445, n_2446, n_2447, 
      n_2448, n_2449, n_2450, n_2451, n_2452, n_2453, n_2454, n_2455, n_2456, 
      n_2457, n_2458, n_2459, n_2460, n_2461, n_2462, n_2463, n_2464, n_2465, 
      n_2466, n_2467, n_2468, n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, 
      n_2475, n_2476, n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, 
      n_2484, n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492, 
      n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500, n_2501, 
      n_2502, n_2503, n_2504, n_2505, n_2506, n_2507, n_2508, n_2509, n_2510, 
      n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518, n_2519, 
      n_2520, n_2521, n_2522, n_2523, n_2524, n_2525, n_2526, n_2527, n_2528, 
      n_2529, n_2530, n_2531, n_2532, n_2533, n_2534, n_2535, n_2536, n_2537, 
      n_2538, n_2539, n_2540, n_2541, n_2542, n_2543, n_2544, n_2545, n_2546, 
      n_2547, n_2548, n_2549, n_2550, n_2551, n_2552, n_2553, n_2554, n_2555, 
      n_2556, n_2557, n_2558, n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, 
      n_2565, n_2566, n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, 
      n_2574, n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582, 
      n_2583, n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591, 
      n_2592, n_2593, n_2594, n_2595, n_2596, n_2597, n_2598, n_2599, n_2600, 
      n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608, n_2609, 
      n_2610, n_2611, n_2612, n_2613, n_2614, n_2615, n_2616, n_2617, n_2618, 
      n_2619, n_2620, n_2621, n_2622, n_2623, n_2624, n_2625, n_2626, n_2627, 
      n_2628, n_2629, n_2630, n_2631, n_2632, n_2633, n_2634, n_2635, n_2636, 
      n_2637, n_2638, n_2639, n_2640, n_2641, n_2642, n_2643, n_2644, n_2645, 
      n_2646, n_2647, n_2648, n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, 
      n_2655, n_2656, n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, 
      n_2664, n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672, 
      n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680, n_2681, 
      n_2682, n_2683, n_2684, n_2685, n_2686, n_2687, n_2688, n_2689, n_2690, 
      n_2691, n_2692, n_2693, n_2694, n_2695, n_2696, n_2697, n_2698, n_2699, 
      n_2700, n_2701, n_2702, n_2703, n_2704, n_2705, n_2706, n_2707, n_2708, 
      n_2709, n_2710, n_2711, n_2712, n_2713, n_2714, n_2715, n_2716, n_2717, 
      n_2718, n_2719, n_2720, n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, 
      n_2727, n_2728, n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, 
      n_2736, n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744, 
      n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752, n_2753, 
      n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760, n_2761, n_2762, 
      n_2763, n_2764, n_2765, n_2766, n_2767, n_2768, n_2769, n_2770, n_2771, 
      n_2772, n_2773, n_2774, n_2775, n_2776, n_2777, n_2778, n_2779, n_2780, 
      n_2781, n_2782, n_2783, n_2784, n_2785, n_2786, n_2787, n_2788, n_2789, 
      n_2790, n_2791, n_2792, n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, 
      n_2799, n_2800, n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, 
      n_2808, n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816, 
      n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, n_2823, n_2824, n_2825, 
      n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832, n_2833, n_2834, 
      n_2835, n_2836, n_2837, n_2838, n_2839, n_2840, n_2841, n_2842, n_2843, 
      n_2844, n_2845, n_2846, n_2847, n_2848, n_2849, n_2850, n_2851, n_2852, 
      n_2853, n_2854, n_2855, n_2856, n_2857, n_2858, n_2859, n_2860, n_2861, 
      n_2862, n_2863, n_2864, n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, 
      n_2871, n_2872, n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, 
      n_2880, n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888, 
      n_2889, n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896, n_2897, 
      n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904, n_2905, n_2906, 
      n_2907, n_2908, n_2909, n_2910, n_2911, n_2912, n_2913, n_2914, n_2915, 
      n_2916, n_2917, n_2918, n_2919, n_2920, n_2921, n_2922, n_2923, n_2924, 
      n_2925, n_2926, n_2927, n_2928, n_2929, n_2930, n_2931, n_2932, n_2933, 
      n_2934, n_2935, n_2936, n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, 
      n_2943, n_2944, n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, 
      n_2952, n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960, 
      n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967, n_2968, n_2969, 
      n_2970, n_2971, n_2972, n_2973, n_2974, n_2975, n_2976, n_2977, n_2978, 
      n_2979, n_2980, n_2981, n_2982, n_2983, n_2984, n_2985, n_2986, n_2987, 
      n_2988, n_2989, n_2990, n_2991, n_2992, n_2993, n_2994, n_2995, n_2996, 
      n_2997, n_2998, n_2999, n_3000, n_3001, n_3002, n_3003, n_3004, n_3005, 
      n_3006, n_3007, n_3008, n_3009, n_3010, n_3011, n_3012, n_3013, n_3014, 
      n_3015, n_3016, n_3017, n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, 
      n_3024, n_3025, n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, 
      n_3033, n_3034, n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041, 
      n_3042, n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050, 
      n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058, n_3059, 
      n_3060, n_3061, n_3062, n_3063, n_3064, n_3065, n_3066, n_3067, n_3068, 
      n_3069, n_3070, n_3071, n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, 
      n_3078, n_3079, n_3080, n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, 
      n_3087, n_3088, n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095, 
      n_3096, n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, n_3103, n_3104, 
      n_3105, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111, n_3112, n_3113, 
      n_3114, n_3115, n_3116, n_3117, n_3118, n_3119, n_3120, n_3121, n_3122, 
      n_3123, n_3124, n_3125, n_3126, n_3127, n_3128, n_3129, n_3130, n_3131, 
      n_3132, n_3133, n_3134, n_3135, n_3136, n_3137, n_3138, n_3139, n_3140, 
      n_3141, n_3142, n_3143, n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, 
      n_3150, n_3151, n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, 
      n_3159, n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167, 
      n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175, n_3176, 
      n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183, n_3184, n_3185, 
      n_3186, n_3187, n_3188, n_3189, n_3190, n_3191, n_3192, n_3193, n_3194, 
      n_3195, n_3196, n_3197, n_3198, n_3199, n_3200, n_3201, n_3202, n_3203, 
      n_3204, n_3205, n_3206, n_3207, n_3208, n_3209, n_3210, n_3211, n_3212, 
      n_3213, n_3214, n_3215, n_3216, n_3217, n_3218, n_3219, n_3220, n_3221, 
      n_3222, n_3223, n_3224, n_3225, n_3226, n_3227, n_3228, n_3229, n_3230, 
      n_3231, n_3232, n_3233, n_3234, n_3235, n_3236, n_3237, n_3238, n_3239, 
      n_3240, n_3241, n_3242, n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, 
      n_3249, n_3250, n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, 
      n_3258, n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, n_3266, 
      n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, n_3274, n_3275, 
      n_3276, n_3277, n_3278, n_3279, n_3280, n_3281, n_3282, n_3283, n_3284, 
      n_3285, n_3286, n_3287, n_3288, n_3289, n_3290, n_3291, n_3292, n_3293, 
      n_3294, n_3295, n_3296, n_3297, n_3298, n_3299, n_3300, n_3301, n_3302, 
      n_3303, n_3304, n_3305, n_3306, n_3307, n_3308, n_3309, n_3310, n_3311, 
      n_3312, n_3313, n_3314, n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, 
      n_3321, n_3322, n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, 
      n_3330, n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338, 
      n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346, n_3347, 
      n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354, n_3355, n_3356, 
      n_3357, n_3358, n_3359, n_3360, n_3361, n_3362, n_3363, n_3364, n_3365, 
      n_3366, n_3367, n_3368, n_3369, n_3370, n_3371, n_3372, n_3373, n_3374, 
      n_3375, n_3376, n_3377, n_3378, n_3379, n_3380, n_3381, n_3382, n_3383, 
      n_3384, n_3385, n_3386, n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, 
      n_3393, n_3394, n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, 
      n_3402, n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410, 
      n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, n_3418, n_3419, 
      n_3420, n_3421, n_3422, n_3423, n_3424, n_3425, n_3426, n_3427, n_3428, 
      n_3429, n_3430, n_3431, n_3432, n_3433, n_3434, n_3435, n_3436, n_3437, 
      n_3438, n_3439, n_3440, n_3441, n_3442, n_3443, n_3444, n_3445, n_3446, 
      n_3447, n_3448, n_3449, n_3450, n_3451, n_3452, n_3453, n_3454, n_3455, 
      n_3456, n_3457, n_3458, n_3459, n_3460, n_3461, n_3462, n_3463, n_3464, 
      n_3465, n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473, 
      n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, n_3481, n_3482, 
      n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489, n_3490, n_3491, 
      n_3492, n_3493, n_3494, n_3495, n_3496, n_3497, n_3498, n_3499, n_3500, 
      n_3501, n_3502, n_3503, n_3504, n_3505, n_3506, n_3507, n_3508, n_3509, 
      n_3510, n_3511, n_3512, n_3513, n_3514, n_3515, n_3516, n_3517, n_3518, 
      n_3519, n_3520, n_3521, n_3522, n_3523, n_3524, n_3525, n_3526, n_3527, 
      n_3528, n_3529, n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, 
      n_3537, n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545, 
      n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553, n_3554, 
      n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561, n_3562, n_3563, 
      n_3564, n_3565, n_3566, n_3567, n_3568, n_3569, n_3570, n_3571, n_3572, 
      n_3573, n_3574, n_3575, n_3576, n_3577, n_3578, n_3579, n_3580, n_3581, 
      n_3582, n_3583, n_3584, n_3585, n_3586, n_3587, n_3588, n_3589, n_3590, 
      n_3591, n_3592, n_3593, n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, 
      n_3600, n_3601, n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, 
      n_3609, n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617, 
      n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625, n_3626, 
      n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633, n_3634, n_3635, 
      n_3636, n_3637, n_3638, n_3639, n_3640, n_3641, n_3642, n_3643, n_3644, 
      n_3645, n_3646, n_3647, n_3648, n_3649, n_3650, n_3651, n_3652, n_3653, 
      n_3654, n_3655, n_3656, n_3657, n_3658, n_3659, n_3660, n_3661, n_3662, 
      n_3663, n_3664, n_3665, n_3666, n_3667, n_3668, n_3669, n_3670, n_3671, 
      n_3672, n_3673, n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, 
      n_3681, n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689, 
      n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697, n_3698, 
      n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705, n_3706, n_3707, 
      n_3708, n_3709, n_3710, n_3711, n_3712, n_3713, n_3714, n_3715, n_3716, 
      n_3717, n_3718, n_3719, n_3720, n_3721, n_3722, n_3723, n_3724, n_3725, 
      n_3726, n_3727, n_3728, n_3729, n_3730, n_3731, n_3732, n_3733, n_3734, 
      n_3735, n_3736, n_3737, n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, 
      n_3744, n_3745, n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, 
      n_3753, n_3754, n_3755, n_3756, n_3757, n_3758, n_3759, n_3760, n_3761, 
      n_3762, n_3763, n_3764, n_3765, n_3766, n_3767, n_3768, n_3769, n_3770, 
      n_3771, n_3772, n_3773, n_3774, n_3775, n_3776, n_3777, n_3778, n_3779, 
      n_3780, n_3781, n_3782, n_3783, n_3784, n_3785, n_3786, n_3787, n_3788, 
      n_3789, n_3790, n_3791, n_3792, n_3793, n_3794, n_3795, n_3796, n_3797, 
      n_3798, n_3799, n_3800, n_3801, n_3802, n_3803, n_3804, n_3805, n_3806, 
      n_3807, n_3808, n_3809, n_3810, n_3811, n_3812, n_3813, n_3814, n_3815, 
      n_3816, n_3817, n_3818, n_3819, n_3820, n_3821, n_3822, n_3823, n_3824, 
      n_3825, n_3826, n_3827, n_3828, n_3829, n_3830, n_3831, n_3832, n_3833, 
      n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841, n_3842, 
      n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849, n_3850, n_3851, 
      n_3852, n_3853, n_3854, n_3855, n_3856, n_3857, n_3858, n_3859, n_3860, 
      n_3861, n_3862, n_3863, n_3864, n_3865, n_3866, n_3867, n_3868, n_3869, 
      n_3870, n_3871, n_3872, n_3873, n_3874, n_3875, n_3876, n_3877, n_3878, 
      n_3879, n_3880, n_3881, n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, 
      n_3888, n_3889, n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896, 
      n_3897, n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904, n_3905, 
      n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, n_3913, n_3914, 
      n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921, n_3922, n_3923, 
      n_3924, n_3925, n_3926, n_3927, n_3928, n_3929, n_3930, n_3931, n_3932, 
      n_3933, n_3934, n_3935, n_3936, n_3937, n_3938, n_3939, n_3940, n_3941, 
      n_3942, n_3943, n_3944, n_3945, n_3946, n_3947, n_3948, n_3949, n_3950, 
      n_3951, n_3952, n_3953, n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, 
      n_3960, n_3961, n_3962, n_3963, n_3964, n_3965, n_3966, n_3967, n_3968, 
      n_3969, n_3970, n_3971, n_3972, n_3973, n_3974, n_3975 : std_logic;

begin
   IRAM_ADDRESS <= ( IRAM_ADDRESS_31_port, IRAM_ADDRESS_30_port, 
      IRAM_ADDRESS_29_port, IRAM_ADDRESS_28_port, IRAM_ADDRESS_27_port, 
      IRAM_ADDRESS_26_port, IRAM_ADDRESS_25_port, IRAM_ADDRESS_24_port, 
      IRAM_ADDRESS_23_port, IRAM_ADDRESS_22_port, IRAM_ADDRESS_21_port, 
      IRAM_ADDRESS_20_port, IRAM_ADDRESS_19_port, IRAM_ADDRESS_18_port, 
      IRAM_ADDRESS_17_port, IRAM_ADDRESS_16_port, IRAM_ADDRESS_15_port, 
      IRAM_ADDRESS_14_port, IRAM_ADDRESS_13_port, IRAM_ADDRESS_12_port, 
      IRAM_ADDRESS_11_port, IRAM_ADDRESS_10_port, IRAM_ADDRESS_9_port, 
      IRAM_ADDRESS_8_port, IRAM_ADDRESS_7_port, IRAM_ADDRESS_6_port, 
      IRAM_ADDRESS_5_port, IRAM_ADDRESS_4_port, IRAM_ADDRESS_3_port, 
      IRAM_ADDRESS_2_port, IRAM_ADDRESS_1_port, IRAM_ADDRESS_0_port );
   DRAM_ADDRESS <= ( DRAM_ADDRESS_31_port, DRAM_ADDRESS_30_port, 
      DRAM_ADDRESS_29_port, DRAM_ADDRESS_28_port, DRAM_ADDRESS_27_port, 
      DRAM_ADDRESS_26_port, DRAM_ADDRESS_25_port, DRAM_ADDRESS_24_port, 
      DRAM_ADDRESS_23_port, DRAM_ADDRESS_22_port, DRAM_ADDRESS_21_port, 
      DRAM_ADDRESS_20_port, DRAM_ADDRESS_19_port, DRAM_ADDRESS_18_port, 
      DRAM_ADDRESS_17_port, DRAM_ADDRESS_16_port, DRAM_ADDRESS_15_port, 
      DRAM_ADDRESS_14_port, DRAM_ADDRESS_13_port, DRAM_ADDRESS_12_port, 
      DRAM_ADDRESS_11_port, DRAM_ADDRESS_10_port, DRAM_ADDRESS_9_port, 
      DRAM_ADDRESS_8_port, DRAM_ADDRESS_7_port, DRAM_ADDRESS_6_port, 
      DRAM_ADDRESS_5_port, DRAM_ADDRESS_4_port, DRAM_ADDRESS_3_port, 
      DRAM_ADDRESS_2_port, DRAM_ADDRESS_1_port, DRAM_ADDRESS_0_port );
   DRAM_DATA_OUT <= ( DRAM_DATA_OUT_31_port, DRAM_DATA_OUT_30_port, 
      DRAM_DATA_OUT_29_port, DRAM_DATA_OUT_28_port, DRAM_DATA_OUT_27_port, 
      DRAM_DATA_OUT_26_port, DRAM_DATA_OUT_25_port, DRAM_DATA_OUT_24_port, 
      DRAM_DATA_OUT_23_port, DRAM_DATA_OUT_22_port, DRAM_DATA_OUT_21_port, 
      DRAM_DATA_OUT_20_port, DRAM_DATA_OUT_19_port, DRAM_DATA_OUT_18_port, 
      DRAM_DATA_OUT_17_port, DRAM_DATA_OUT_16_port, DRAM_DATA_OUT_15_port, 
      DRAM_DATA_OUT_14_port, DRAM_DATA_OUT_13_port, DRAM_DATA_OUT_12_port, 
      DRAM_DATA_OUT_11_port, DRAM_DATA_OUT_10_port, DRAM_DATA_OUT_9_port, 
      DRAM_DATA_OUT_8_port, DRAM_DATA_OUT_7_port, DRAM_DATA_OUT_6_port, 
      DRAM_DATA_OUT_5_port, DRAM_DATA_OUT_4_port, DRAM_DATA_OUT_3_port, 
      DRAM_DATA_OUT_2_port, DRAM_DATA_OUT_1_port, DRAM_DATA_OUT_0_port );
   DATA_SIZE <= ( DATA_SIZE_1_port, DATA_SIZE_0_port );
   DRAMRF_ADDRESS <= ( DRAMRF_ADDRESS_31_port, DRAMRF_ADDRESS_30_port, 
      DRAMRF_ADDRESS_29_port, DRAMRF_ADDRESS_28_port, DRAMRF_ADDRESS_27_port, 
      DRAMRF_ADDRESS_26_port, DRAMRF_ADDRESS_25_port, DRAMRF_ADDRESS_24_port, 
      DRAMRF_ADDRESS_23_port, DRAMRF_ADDRESS_22_port, DRAMRF_ADDRESS_21_port, 
      DRAMRF_ADDRESS_20_port, DRAMRF_ADDRESS_19_port, DRAMRF_ADDRESS_18_port, 
      DRAMRF_ADDRESS_17_port, DRAMRF_ADDRESS_16_port, DRAMRF_ADDRESS_15_port, 
      DRAMRF_ADDRESS_14_port, DRAMRF_ADDRESS_13_port, DRAMRF_ADDRESS_12_port, 
      DRAMRF_ADDRESS_11_port, DRAMRF_ADDRESS_10_port, DRAMRF_ADDRESS_9_port, 
      DRAMRF_ADDRESS_8_port, DRAMRF_ADDRESS_7_port, DRAMRF_ADDRESS_6_port, 
      DRAMRF_ADDRESS_5_port, DRAMRF_ADDRESS_4_port, DRAMRF_ADDRESS_3_port, 
      DRAMRF_ADDRESS_2_port, DRAMRF_ADDRESS_1_port, DRAMRF_ADDRESS_0_port );
   DATA_SIZE_RF <= ( DataPath_RF_bus_complete_win_data_0_port, 
      DataPath_RF_bus_complete_win_data_0_port );
   
   DECODEhw_HAZARD_CTRL : hazard_table_N_REGS_LOG5 port map( CLK => CLK, RST =>
                           RST, WR1 => DECODEhw_i_WR1, WR2 => i_WF, ADD_WR1(4) 
                           => i_ADD_WS1_4_port, ADD_WR1(3) => i_ADD_WS1_3_port,
                           ADD_WR1(2) => i_ADD_WS1_2_port, ADD_WR1(1) => 
                           i_ADD_WS1_1_port, ADD_WR1(0) => i_ADD_WS1_0_port, 
                           ADD_WR2(4) => i_ADD_WB_4_port, ADD_WR2(3) => 
                           i_ADD_WB_3_port, ADD_WR2(2) => i_ADD_WB_2_port, 
                           ADD_WR2(1) => i_ADD_WB_1_port, ADD_WR2(0) => 
                           i_ADD_WB_0_port, ADD_CHECK1(4) => i_ADD_RS1_4_port, 
                           ADD_CHECK1(3) => i_ADD_RS1_3_port, ADD_CHECK1(2) => 
                           i_ADD_RS1_2_port, ADD_CHECK1(1) => i_ADD_RS1_1_port,
                           ADD_CHECK1(0) => i_ADD_RS1_0_port, ADD_CHECK2(4) => 
                           i_ADD_RS2_4_port, ADD_CHECK2(3) => i_ADD_RS2_3_port,
                           ADD_CHECK2(2) => i_ADD_RS2_2_port, ADD_CHECK2(1) => 
                           i_ADD_RS2_1_port, ADD_CHECK2(0) => i_ADD_RS2_0_port,
                           BUSY => i_HAZARD_SIG_CU, BUSY_WINDOW => 
                           i_BUSY_WINDOW);
   DataPath_RF_SELBLOCK_INLOC : in_loc_selblock_NBIT_DATA32_N8_F5 port map( 
                           regs(2559) => DataPath_RF_bus_reg_dataout_2559_port,
                           regs(2558) => DataPath_RF_bus_reg_dataout_2558_port,
                           regs(2557) => DataPath_RF_bus_reg_dataout_2557_port,
                           regs(2556) => DataPath_RF_bus_reg_dataout_2556_port,
                           regs(2555) => DataPath_RF_bus_reg_dataout_2555_port,
                           regs(2554) => DataPath_RF_bus_reg_dataout_2554_port,
                           regs(2553) => DataPath_RF_bus_reg_dataout_2553_port,
                           regs(2552) => DataPath_RF_bus_reg_dataout_2552_port,
                           regs(2551) => DataPath_RF_bus_reg_dataout_2551_port,
                           regs(2550) => DataPath_RF_bus_reg_dataout_2550_port,
                           regs(2549) => DataPath_RF_bus_reg_dataout_2549_port,
                           regs(2548) => DataPath_RF_bus_reg_dataout_2548_port,
                           regs(2547) => DataPath_RF_bus_reg_dataout_2547_port,
                           regs(2546) => DataPath_RF_bus_reg_dataout_2546_port,
                           regs(2545) => DataPath_RF_bus_reg_dataout_2545_port,
                           regs(2544) => DataPath_RF_bus_reg_dataout_2544_port,
                           regs(2543) => DataPath_RF_bus_reg_dataout_2543_port,
                           regs(2542) => DataPath_RF_bus_reg_dataout_2542_port,
                           regs(2541) => DataPath_RF_bus_reg_dataout_2541_port,
                           regs(2540) => DataPath_RF_bus_reg_dataout_2540_port,
                           regs(2539) => DataPath_RF_bus_reg_dataout_2539_port,
                           regs(2538) => DataPath_RF_bus_reg_dataout_2538_port,
                           regs(2537) => DataPath_RF_bus_reg_dataout_2537_port,
                           regs(2536) => DataPath_RF_bus_reg_dataout_2536_port,
                           regs(2535) => DataPath_RF_bus_reg_dataout_2535_port,
                           regs(2534) => DataPath_RF_bus_reg_dataout_2534_port,
                           regs(2533) => DataPath_RF_bus_reg_dataout_2533_port,
                           regs(2532) => DataPath_RF_bus_reg_dataout_2532_port,
                           regs(2531) => DataPath_RF_bus_reg_dataout_2531_port,
                           regs(2530) => DataPath_RF_bus_reg_dataout_2530_port,
                           regs(2529) => DataPath_RF_bus_reg_dataout_2529_port,
                           regs(2528) => DataPath_RF_bus_reg_dataout_2528_port,
                           regs(2527) => DataPath_RF_bus_reg_dataout_2527_port,
                           regs(2526) => DataPath_RF_bus_reg_dataout_2526_port,
                           regs(2525) => DataPath_RF_bus_reg_dataout_2525_port,
                           regs(2524) => DataPath_RF_bus_reg_dataout_2524_port,
                           regs(2523) => DataPath_RF_bus_reg_dataout_2523_port,
                           regs(2522) => DataPath_RF_bus_reg_dataout_2522_port,
                           regs(2521) => DataPath_RF_bus_reg_dataout_2521_port,
                           regs(2520) => DataPath_RF_bus_reg_dataout_2520_port,
                           regs(2519) => DataPath_RF_bus_reg_dataout_2519_port,
                           regs(2518) => DataPath_RF_bus_reg_dataout_2518_port,
                           regs(2517) => DataPath_RF_bus_reg_dataout_2517_port,
                           regs(2516) => DataPath_RF_bus_reg_dataout_2516_port,
                           regs(2515) => DataPath_RF_bus_reg_dataout_2515_port,
                           regs(2514) => DataPath_RF_bus_reg_dataout_2514_port,
                           regs(2513) => DataPath_RF_bus_reg_dataout_2513_port,
                           regs(2512) => DataPath_RF_bus_reg_dataout_2512_port,
                           regs(2511) => DataPath_RF_bus_reg_dataout_2511_port,
                           regs(2510) => DataPath_RF_bus_reg_dataout_2510_port,
                           regs(2509) => DataPath_RF_bus_reg_dataout_2509_port,
                           regs(2508) => DataPath_RF_bus_reg_dataout_2508_port,
                           regs(2507) => DataPath_RF_bus_reg_dataout_2507_port,
                           regs(2506) => DataPath_RF_bus_reg_dataout_2506_port,
                           regs(2505) => DataPath_RF_bus_reg_dataout_2505_port,
                           regs(2504) => DataPath_RF_bus_reg_dataout_2504_port,
                           regs(2503) => DataPath_RF_bus_reg_dataout_2503_port,
                           regs(2502) => DataPath_RF_bus_reg_dataout_2502_port,
                           regs(2501) => DataPath_RF_bus_reg_dataout_2501_port,
                           regs(2500) => DataPath_RF_bus_reg_dataout_2500_port,
                           regs(2499) => DataPath_RF_bus_reg_dataout_2499_port,
                           regs(2498) => DataPath_RF_bus_reg_dataout_2498_port,
                           regs(2497) => DataPath_RF_bus_reg_dataout_2497_port,
                           regs(2496) => DataPath_RF_bus_reg_dataout_2496_port,
                           regs(2495) => DataPath_RF_bus_reg_dataout_2495_port,
                           regs(2494) => DataPath_RF_bus_reg_dataout_2494_port,
                           regs(2493) => DataPath_RF_bus_reg_dataout_2493_port,
                           regs(2492) => DataPath_RF_bus_reg_dataout_2492_port,
                           regs(2491) => DataPath_RF_bus_reg_dataout_2491_port,
                           regs(2490) => DataPath_RF_bus_reg_dataout_2490_port,
                           regs(2489) => DataPath_RF_bus_reg_dataout_2489_port,
                           regs(2488) => DataPath_RF_bus_reg_dataout_2488_port,
                           regs(2487) => DataPath_RF_bus_reg_dataout_2487_port,
                           regs(2486) => DataPath_RF_bus_reg_dataout_2486_port,
                           regs(2485) => DataPath_RF_bus_reg_dataout_2485_port,
                           regs(2484) => DataPath_RF_bus_reg_dataout_2484_port,
                           regs(2483) => DataPath_RF_bus_reg_dataout_2483_port,
                           regs(2482) => DataPath_RF_bus_reg_dataout_2482_port,
                           regs(2481) => DataPath_RF_bus_reg_dataout_2481_port,
                           regs(2480) => DataPath_RF_bus_reg_dataout_2480_port,
                           regs(2479) => DataPath_RF_bus_reg_dataout_2479_port,
                           regs(2478) => DataPath_RF_bus_reg_dataout_2478_port,
                           regs(2477) => DataPath_RF_bus_reg_dataout_2477_port,
                           regs(2476) => DataPath_RF_bus_reg_dataout_2476_port,
                           regs(2475) => DataPath_RF_bus_reg_dataout_2475_port,
                           regs(2474) => DataPath_RF_bus_reg_dataout_2474_port,
                           regs(2473) => DataPath_RF_bus_reg_dataout_2473_port,
                           regs(2472) => DataPath_RF_bus_reg_dataout_2472_port,
                           regs(2471) => DataPath_RF_bus_reg_dataout_2471_port,
                           regs(2470) => DataPath_RF_bus_reg_dataout_2470_port,
                           regs(2469) => DataPath_RF_bus_reg_dataout_2469_port,
                           regs(2468) => DataPath_RF_bus_reg_dataout_2468_port,
                           regs(2467) => DataPath_RF_bus_reg_dataout_2467_port,
                           regs(2466) => DataPath_RF_bus_reg_dataout_2466_port,
                           regs(2465) => DataPath_RF_bus_reg_dataout_2465_port,
                           regs(2464) => DataPath_RF_bus_reg_dataout_2464_port,
                           regs(2463) => DataPath_RF_bus_reg_dataout_2463_port,
                           regs(2462) => DataPath_RF_bus_reg_dataout_2462_port,
                           regs(2461) => DataPath_RF_bus_reg_dataout_2461_port,
                           regs(2460) => DataPath_RF_bus_reg_dataout_2460_port,
                           regs(2459) => DataPath_RF_bus_reg_dataout_2459_port,
                           regs(2458) => DataPath_RF_bus_reg_dataout_2458_port,
                           regs(2457) => DataPath_RF_bus_reg_dataout_2457_port,
                           regs(2456) => DataPath_RF_bus_reg_dataout_2456_port,
                           regs(2455) => DataPath_RF_bus_reg_dataout_2455_port,
                           regs(2454) => DataPath_RF_bus_reg_dataout_2454_port,
                           regs(2453) => DataPath_RF_bus_reg_dataout_2453_port,
                           regs(2452) => DataPath_RF_bus_reg_dataout_2452_port,
                           regs(2451) => DataPath_RF_bus_reg_dataout_2451_port,
                           regs(2450) => DataPath_RF_bus_reg_dataout_2450_port,
                           regs(2449) => DataPath_RF_bus_reg_dataout_2449_port,
                           regs(2448) => DataPath_RF_bus_reg_dataout_2448_port,
                           regs(2447) => DataPath_RF_bus_reg_dataout_2447_port,
                           regs(2446) => DataPath_RF_bus_reg_dataout_2446_port,
                           regs(2445) => DataPath_RF_bus_reg_dataout_2445_port,
                           regs(2444) => DataPath_RF_bus_reg_dataout_2444_port,
                           regs(2443) => DataPath_RF_bus_reg_dataout_2443_port,
                           regs(2442) => DataPath_RF_bus_reg_dataout_2442_port,
                           regs(2441) => DataPath_RF_bus_reg_dataout_2441_port,
                           regs(2440) => DataPath_RF_bus_reg_dataout_2440_port,
                           regs(2439) => DataPath_RF_bus_reg_dataout_2439_port,
                           regs(2438) => DataPath_RF_bus_reg_dataout_2438_port,
                           regs(2437) => DataPath_RF_bus_reg_dataout_2437_port,
                           regs(2436) => DataPath_RF_bus_reg_dataout_2436_port,
                           regs(2435) => DataPath_RF_bus_reg_dataout_2435_port,
                           regs(2434) => DataPath_RF_bus_reg_dataout_2434_port,
                           regs(2433) => DataPath_RF_bus_reg_dataout_2433_port,
                           regs(2432) => DataPath_RF_bus_reg_dataout_2432_port,
                           regs(2431) => DataPath_RF_bus_reg_dataout_2431_port,
                           regs(2430) => DataPath_RF_bus_reg_dataout_2430_port,
                           regs(2429) => DataPath_RF_bus_reg_dataout_2429_port,
                           regs(2428) => DataPath_RF_bus_reg_dataout_2428_port,
                           regs(2427) => DataPath_RF_bus_reg_dataout_2427_port,
                           regs(2426) => DataPath_RF_bus_reg_dataout_2426_port,
                           regs(2425) => DataPath_RF_bus_reg_dataout_2425_port,
                           regs(2424) => DataPath_RF_bus_reg_dataout_2424_port,
                           regs(2423) => DataPath_RF_bus_reg_dataout_2423_port,
                           regs(2422) => DataPath_RF_bus_reg_dataout_2422_port,
                           regs(2421) => DataPath_RF_bus_reg_dataout_2421_port,
                           regs(2420) => DataPath_RF_bus_reg_dataout_2420_port,
                           regs(2419) => DataPath_RF_bus_reg_dataout_2419_port,
                           regs(2418) => DataPath_RF_bus_reg_dataout_2418_port,
                           regs(2417) => DataPath_RF_bus_reg_dataout_2417_port,
                           regs(2416) => DataPath_RF_bus_reg_dataout_2416_port,
                           regs(2415) => DataPath_RF_bus_reg_dataout_2415_port,
                           regs(2414) => DataPath_RF_bus_reg_dataout_2414_port,
                           regs(2413) => DataPath_RF_bus_reg_dataout_2413_port,
                           regs(2412) => DataPath_RF_bus_reg_dataout_2412_port,
                           regs(2411) => DataPath_RF_bus_reg_dataout_2411_port,
                           regs(2410) => DataPath_RF_bus_reg_dataout_2410_port,
                           regs(2409) => DataPath_RF_bus_reg_dataout_2409_port,
                           regs(2408) => DataPath_RF_bus_reg_dataout_2408_port,
                           regs(2407) => DataPath_RF_bus_reg_dataout_2407_port,
                           regs(2406) => DataPath_RF_bus_reg_dataout_2406_port,
                           regs(2405) => DataPath_RF_bus_reg_dataout_2405_port,
                           regs(2404) => DataPath_RF_bus_reg_dataout_2404_port,
                           regs(2403) => DataPath_RF_bus_reg_dataout_2403_port,
                           regs(2402) => DataPath_RF_bus_reg_dataout_2402_port,
                           regs(2401) => DataPath_RF_bus_reg_dataout_2401_port,
                           regs(2400) => DataPath_RF_bus_reg_dataout_2400_port,
                           regs(2399) => DataPath_RF_bus_reg_dataout_2399_port,
                           regs(2398) => DataPath_RF_bus_reg_dataout_2398_port,
                           regs(2397) => DataPath_RF_bus_reg_dataout_2397_port,
                           regs(2396) => DataPath_RF_bus_reg_dataout_2396_port,
                           regs(2395) => DataPath_RF_bus_reg_dataout_2395_port,
                           regs(2394) => DataPath_RF_bus_reg_dataout_2394_port,
                           regs(2393) => DataPath_RF_bus_reg_dataout_2393_port,
                           regs(2392) => DataPath_RF_bus_reg_dataout_2392_port,
                           regs(2391) => DataPath_RF_bus_reg_dataout_2391_port,
                           regs(2390) => DataPath_RF_bus_reg_dataout_2390_port,
                           regs(2389) => DataPath_RF_bus_reg_dataout_2389_port,
                           regs(2388) => DataPath_RF_bus_reg_dataout_2388_port,
                           regs(2387) => DataPath_RF_bus_reg_dataout_2387_port,
                           regs(2386) => DataPath_RF_bus_reg_dataout_2386_port,
                           regs(2385) => DataPath_RF_bus_reg_dataout_2385_port,
                           regs(2384) => DataPath_RF_bus_reg_dataout_2384_port,
                           regs(2383) => DataPath_RF_bus_reg_dataout_2383_port,
                           regs(2382) => DataPath_RF_bus_reg_dataout_2382_port,
                           regs(2381) => DataPath_RF_bus_reg_dataout_2381_port,
                           regs(2380) => DataPath_RF_bus_reg_dataout_2380_port,
                           regs(2379) => DataPath_RF_bus_reg_dataout_2379_port,
                           regs(2378) => DataPath_RF_bus_reg_dataout_2378_port,
                           regs(2377) => DataPath_RF_bus_reg_dataout_2377_port,
                           regs(2376) => DataPath_RF_bus_reg_dataout_2376_port,
                           regs(2375) => DataPath_RF_bus_reg_dataout_2375_port,
                           regs(2374) => DataPath_RF_bus_reg_dataout_2374_port,
                           regs(2373) => DataPath_RF_bus_reg_dataout_2373_port,
                           regs(2372) => DataPath_RF_bus_reg_dataout_2372_port,
                           regs(2371) => DataPath_RF_bus_reg_dataout_2371_port,
                           regs(2370) => DataPath_RF_bus_reg_dataout_2370_port,
                           regs(2369) => DataPath_RF_bus_reg_dataout_2369_port,
                           regs(2368) => DataPath_RF_bus_reg_dataout_2368_port,
                           regs(2367) => DataPath_RF_bus_reg_dataout_2367_port,
                           regs(2366) => DataPath_RF_bus_reg_dataout_2366_port,
                           regs(2365) => DataPath_RF_bus_reg_dataout_2365_port,
                           regs(2364) => DataPath_RF_bus_reg_dataout_2364_port,
                           regs(2363) => DataPath_RF_bus_reg_dataout_2363_port,
                           regs(2362) => DataPath_RF_bus_reg_dataout_2362_port,
                           regs(2361) => DataPath_RF_bus_reg_dataout_2361_port,
                           regs(2360) => DataPath_RF_bus_reg_dataout_2360_port,
                           regs(2359) => DataPath_RF_bus_reg_dataout_2359_port,
                           regs(2358) => DataPath_RF_bus_reg_dataout_2358_port,
                           regs(2357) => DataPath_RF_bus_reg_dataout_2357_port,
                           regs(2356) => DataPath_RF_bus_reg_dataout_2356_port,
                           regs(2355) => DataPath_RF_bus_reg_dataout_2355_port,
                           regs(2354) => DataPath_RF_bus_reg_dataout_2354_port,
                           regs(2353) => DataPath_RF_bus_reg_dataout_2353_port,
                           regs(2352) => DataPath_RF_bus_reg_dataout_2352_port,
                           regs(2351) => DataPath_RF_bus_reg_dataout_2351_port,
                           regs(2350) => DataPath_RF_bus_reg_dataout_2350_port,
                           regs(2349) => DataPath_RF_bus_reg_dataout_2349_port,
                           regs(2348) => DataPath_RF_bus_reg_dataout_2348_port,
                           regs(2347) => DataPath_RF_bus_reg_dataout_2347_port,
                           regs(2346) => DataPath_RF_bus_reg_dataout_2346_port,
                           regs(2345) => DataPath_RF_bus_reg_dataout_2345_port,
                           regs(2344) => DataPath_RF_bus_reg_dataout_2344_port,
                           regs(2343) => DataPath_RF_bus_reg_dataout_2343_port,
                           regs(2342) => DataPath_RF_bus_reg_dataout_2342_port,
                           regs(2341) => DataPath_RF_bus_reg_dataout_2341_port,
                           regs(2340) => DataPath_RF_bus_reg_dataout_2340_port,
                           regs(2339) => DataPath_RF_bus_reg_dataout_2339_port,
                           regs(2338) => DataPath_RF_bus_reg_dataout_2338_port,
                           regs(2337) => DataPath_RF_bus_reg_dataout_2337_port,
                           regs(2336) => DataPath_RF_bus_reg_dataout_2336_port,
                           regs(2335) => DataPath_RF_bus_reg_dataout_2335_port,
                           regs(2334) => DataPath_RF_bus_reg_dataout_2334_port,
                           regs(2333) => DataPath_RF_bus_reg_dataout_2333_port,
                           regs(2332) => DataPath_RF_bus_reg_dataout_2332_port,
                           regs(2331) => DataPath_RF_bus_reg_dataout_2331_port,
                           regs(2330) => DataPath_RF_bus_reg_dataout_2330_port,
                           regs(2329) => DataPath_RF_bus_reg_dataout_2329_port,
                           regs(2328) => DataPath_RF_bus_reg_dataout_2328_port,
                           regs(2327) => DataPath_RF_bus_reg_dataout_2327_port,
                           regs(2326) => DataPath_RF_bus_reg_dataout_2326_port,
                           regs(2325) => DataPath_RF_bus_reg_dataout_2325_port,
                           regs(2324) => DataPath_RF_bus_reg_dataout_2324_port,
                           regs(2323) => DataPath_RF_bus_reg_dataout_2323_port,
                           regs(2322) => DataPath_RF_bus_reg_dataout_2322_port,
                           regs(2321) => DataPath_RF_bus_reg_dataout_2321_port,
                           regs(2320) => DataPath_RF_bus_reg_dataout_2320_port,
                           regs(2319) => DataPath_RF_bus_reg_dataout_2319_port,
                           regs(2318) => DataPath_RF_bus_reg_dataout_2318_port,
                           regs(2317) => DataPath_RF_bus_reg_dataout_2317_port,
                           regs(2316) => DataPath_RF_bus_reg_dataout_2316_port,
                           regs(2315) => DataPath_RF_bus_reg_dataout_2315_port,
                           regs(2314) => DataPath_RF_bus_reg_dataout_2314_port,
                           regs(2313) => DataPath_RF_bus_reg_dataout_2313_port,
                           regs(2312) => DataPath_RF_bus_reg_dataout_2312_port,
                           regs(2311) => DataPath_RF_bus_reg_dataout_2311_port,
                           regs(2310) => DataPath_RF_bus_reg_dataout_2310_port,
                           regs(2309) => DataPath_RF_bus_reg_dataout_2309_port,
                           regs(2308) => DataPath_RF_bus_reg_dataout_2308_port,
                           regs(2307) => DataPath_RF_bus_reg_dataout_2307_port,
                           regs(2306) => DataPath_RF_bus_reg_dataout_2306_port,
                           regs(2305) => DataPath_RF_bus_reg_dataout_2305_port,
                           regs(2304) => DataPath_RF_bus_reg_dataout_2304_port,
                           regs(2303) => DataPath_RF_bus_reg_dataout_2303_port,
                           regs(2302) => DataPath_RF_bus_reg_dataout_2302_port,
                           regs(2301) => DataPath_RF_bus_reg_dataout_2301_port,
                           regs(2300) => DataPath_RF_bus_reg_dataout_2300_port,
                           regs(2299) => DataPath_RF_bus_reg_dataout_2299_port,
                           regs(2298) => DataPath_RF_bus_reg_dataout_2298_port,
                           regs(2297) => DataPath_RF_bus_reg_dataout_2297_port,
                           regs(2296) => DataPath_RF_bus_reg_dataout_2296_port,
                           regs(2295) => DataPath_RF_bus_reg_dataout_2295_port,
                           regs(2294) => DataPath_RF_bus_reg_dataout_2294_port,
                           regs(2293) => DataPath_RF_bus_reg_dataout_2293_port,
                           regs(2292) => DataPath_RF_bus_reg_dataout_2292_port,
                           regs(2291) => DataPath_RF_bus_reg_dataout_2291_port,
                           regs(2290) => DataPath_RF_bus_reg_dataout_2290_port,
                           regs(2289) => DataPath_RF_bus_reg_dataout_2289_port,
                           regs(2288) => DataPath_RF_bus_reg_dataout_2288_port,
                           regs(2287) => DataPath_RF_bus_reg_dataout_2287_port,
                           regs(2286) => DataPath_RF_bus_reg_dataout_2286_port,
                           regs(2285) => DataPath_RF_bus_reg_dataout_2285_port,
                           regs(2284) => DataPath_RF_bus_reg_dataout_2284_port,
                           regs(2283) => DataPath_RF_bus_reg_dataout_2283_port,
                           regs(2282) => DataPath_RF_bus_reg_dataout_2282_port,
                           regs(2281) => DataPath_RF_bus_reg_dataout_2281_port,
                           regs(2280) => DataPath_RF_bus_reg_dataout_2280_port,
                           regs(2279) => DataPath_RF_bus_reg_dataout_2279_port,
                           regs(2278) => DataPath_RF_bus_reg_dataout_2278_port,
                           regs(2277) => DataPath_RF_bus_reg_dataout_2277_port,
                           regs(2276) => DataPath_RF_bus_reg_dataout_2276_port,
                           regs(2275) => DataPath_RF_bus_reg_dataout_2275_port,
                           regs(2274) => DataPath_RF_bus_reg_dataout_2274_port,
                           regs(2273) => DataPath_RF_bus_reg_dataout_2273_port,
                           regs(2272) => DataPath_RF_bus_reg_dataout_2272_port,
                           regs(2271) => DataPath_RF_bus_reg_dataout_2271_port,
                           regs(2270) => DataPath_RF_bus_reg_dataout_2270_port,
                           regs(2269) => DataPath_RF_bus_reg_dataout_2269_port,
                           regs(2268) => DataPath_RF_bus_reg_dataout_2268_port,
                           regs(2267) => DataPath_RF_bus_reg_dataout_2267_port,
                           regs(2266) => DataPath_RF_bus_reg_dataout_2266_port,
                           regs(2265) => DataPath_RF_bus_reg_dataout_2265_port,
                           regs(2264) => DataPath_RF_bus_reg_dataout_2264_port,
                           regs(2263) => DataPath_RF_bus_reg_dataout_2263_port,
                           regs(2262) => DataPath_RF_bus_reg_dataout_2262_port,
                           regs(2261) => DataPath_RF_bus_reg_dataout_2261_port,
                           regs(2260) => DataPath_RF_bus_reg_dataout_2260_port,
                           regs(2259) => DataPath_RF_bus_reg_dataout_2259_port,
                           regs(2258) => DataPath_RF_bus_reg_dataout_2258_port,
                           regs(2257) => DataPath_RF_bus_reg_dataout_2257_port,
                           regs(2256) => DataPath_RF_bus_reg_dataout_2256_port,
                           regs(2255) => DataPath_RF_bus_reg_dataout_2255_port,
                           regs(2254) => DataPath_RF_bus_reg_dataout_2254_port,
                           regs(2253) => DataPath_RF_bus_reg_dataout_2253_port,
                           regs(2252) => DataPath_RF_bus_reg_dataout_2252_port,
                           regs(2251) => DataPath_RF_bus_reg_dataout_2251_port,
                           regs(2250) => DataPath_RF_bus_reg_dataout_2250_port,
                           regs(2249) => DataPath_RF_bus_reg_dataout_2249_port,
                           regs(2248) => DataPath_RF_bus_reg_dataout_2248_port,
                           regs(2247) => DataPath_RF_bus_reg_dataout_2247_port,
                           regs(2246) => DataPath_RF_bus_reg_dataout_2246_port,
                           regs(2245) => DataPath_RF_bus_reg_dataout_2245_port,
                           regs(2244) => DataPath_RF_bus_reg_dataout_2244_port,
                           regs(2243) => DataPath_RF_bus_reg_dataout_2243_port,
                           regs(2242) => DataPath_RF_bus_reg_dataout_2242_port,
                           regs(2241) => DataPath_RF_bus_reg_dataout_2241_port,
                           regs(2240) => DataPath_RF_bus_reg_dataout_2240_port,
                           regs(2239) => DataPath_RF_bus_reg_dataout_2239_port,
                           regs(2238) => DataPath_RF_bus_reg_dataout_2238_port,
                           regs(2237) => DataPath_RF_bus_reg_dataout_2237_port,
                           regs(2236) => DataPath_RF_bus_reg_dataout_2236_port,
                           regs(2235) => DataPath_RF_bus_reg_dataout_2235_port,
                           regs(2234) => DataPath_RF_bus_reg_dataout_2234_port,
                           regs(2233) => DataPath_RF_bus_reg_dataout_2233_port,
                           regs(2232) => DataPath_RF_bus_reg_dataout_2232_port,
                           regs(2231) => DataPath_RF_bus_reg_dataout_2231_port,
                           regs(2230) => DataPath_RF_bus_reg_dataout_2230_port,
                           regs(2229) => DataPath_RF_bus_reg_dataout_2229_port,
                           regs(2228) => DataPath_RF_bus_reg_dataout_2228_port,
                           regs(2227) => DataPath_RF_bus_reg_dataout_2227_port,
                           regs(2226) => DataPath_RF_bus_reg_dataout_2226_port,
                           regs(2225) => DataPath_RF_bus_reg_dataout_2225_port,
                           regs(2224) => DataPath_RF_bus_reg_dataout_2224_port,
                           regs(2223) => DataPath_RF_bus_reg_dataout_2223_port,
                           regs(2222) => DataPath_RF_bus_reg_dataout_2222_port,
                           regs(2221) => DataPath_RF_bus_reg_dataout_2221_port,
                           regs(2220) => DataPath_RF_bus_reg_dataout_2220_port,
                           regs(2219) => DataPath_RF_bus_reg_dataout_2219_port,
                           regs(2218) => DataPath_RF_bus_reg_dataout_2218_port,
                           regs(2217) => DataPath_RF_bus_reg_dataout_2217_port,
                           regs(2216) => DataPath_RF_bus_reg_dataout_2216_port,
                           regs(2215) => DataPath_RF_bus_reg_dataout_2215_port,
                           regs(2214) => DataPath_RF_bus_reg_dataout_2214_port,
                           regs(2213) => DataPath_RF_bus_reg_dataout_2213_port,
                           regs(2212) => DataPath_RF_bus_reg_dataout_2212_port,
                           regs(2211) => DataPath_RF_bus_reg_dataout_2211_port,
                           regs(2210) => DataPath_RF_bus_reg_dataout_2210_port,
                           regs(2209) => DataPath_RF_bus_reg_dataout_2209_port,
                           regs(2208) => DataPath_RF_bus_reg_dataout_2208_port,
                           regs(2207) => DataPath_RF_bus_reg_dataout_2207_port,
                           regs(2206) => DataPath_RF_bus_reg_dataout_2206_port,
                           regs(2205) => DataPath_RF_bus_reg_dataout_2205_port,
                           regs(2204) => DataPath_RF_bus_reg_dataout_2204_port,
                           regs(2203) => DataPath_RF_bus_reg_dataout_2203_port,
                           regs(2202) => DataPath_RF_bus_reg_dataout_2202_port,
                           regs(2201) => DataPath_RF_bus_reg_dataout_2201_port,
                           regs(2200) => DataPath_RF_bus_reg_dataout_2200_port,
                           regs(2199) => DataPath_RF_bus_reg_dataout_2199_port,
                           regs(2198) => DataPath_RF_bus_reg_dataout_2198_port,
                           regs(2197) => DataPath_RF_bus_reg_dataout_2197_port,
                           regs(2196) => DataPath_RF_bus_reg_dataout_2196_port,
                           regs(2195) => DataPath_RF_bus_reg_dataout_2195_port,
                           regs(2194) => DataPath_RF_bus_reg_dataout_2194_port,
                           regs(2193) => DataPath_RF_bus_reg_dataout_2193_port,
                           regs(2192) => DataPath_RF_bus_reg_dataout_2192_port,
                           regs(2191) => DataPath_RF_bus_reg_dataout_2191_port,
                           regs(2190) => DataPath_RF_bus_reg_dataout_2190_port,
                           regs(2189) => DataPath_RF_bus_reg_dataout_2189_port,
                           regs(2188) => DataPath_RF_bus_reg_dataout_2188_port,
                           regs(2187) => DataPath_RF_bus_reg_dataout_2187_port,
                           regs(2186) => DataPath_RF_bus_reg_dataout_2186_port,
                           regs(2185) => DataPath_RF_bus_reg_dataout_2185_port,
                           regs(2184) => DataPath_RF_bus_reg_dataout_2184_port,
                           regs(2183) => DataPath_RF_bus_reg_dataout_2183_port,
                           regs(2182) => DataPath_RF_bus_reg_dataout_2182_port,
                           regs(2181) => DataPath_RF_bus_reg_dataout_2181_port,
                           regs(2180) => DataPath_RF_bus_reg_dataout_2180_port,
                           regs(2179) => DataPath_RF_bus_reg_dataout_2179_port,
                           regs(2178) => DataPath_RF_bus_reg_dataout_2178_port,
                           regs(2177) => DataPath_RF_bus_reg_dataout_2177_port,
                           regs(2176) => DataPath_RF_bus_reg_dataout_2176_port,
                           regs(2175) => DataPath_RF_bus_reg_dataout_2175_port,
                           regs(2174) => DataPath_RF_bus_reg_dataout_2174_port,
                           regs(2173) => DataPath_RF_bus_reg_dataout_2173_port,
                           regs(2172) => DataPath_RF_bus_reg_dataout_2172_port,
                           regs(2171) => DataPath_RF_bus_reg_dataout_2171_port,
                           regs(2170) => DataPath_RF_bus_reg_dataout_2170_port,
                           regs(2169) => DataPath_RF_bus_reg_dataout_2169_port,
                           regs(2168) => DataPath_RF_bus_reg_dataout_2168_port,
                           regs(2167) => DataPath_RF_bus_reg_dataout_2167_port,
                           regs(2166) => DataPath_RF_bus_reg_dataout_2166_port,
                           regs(2165) => DataPath_RF_bus_reg_dataout_2165_port,
                           regs(2164) => DataPath_RF_bus_reg_dataout_2164_port,
                           regs(2163) => DataPath_RF_bus_reg_dataout_2163_port,
                           regs(2162) => DataPath_RF_bus_reg_dataout_2162_port,
                           regs(2161) => DataPath_RF_bus_reg_dataout_2161_port,
                           regs(2160) => DataPath_RF_bus_reg_dataout_2160_port,
                           regs(2159) => DataPath_RF_bus_reg_dataout_2159_port,
                           regs(2158) => DataPath_RF_bus_reg_dataout_2158_port,
                           regs(2157) => DataPath_RF_bus_reg_dataout_2157_port,
                           regs(2156) => DataPath_RF_bus_reg_dataout_2156_port,
                           regs(2155) => DataPath_RF_bus_reg_dataout_2155_port,
                           regs(2154) => DataPath_RF_bus_reg_dataout_2154_port,
                           regs(2153) => DataPath_RF_bus_reg_dataout_2153_port,
                           regs(2152) => DataPath_RF_bus_reg_dataout_2152_port,
                           regs(2151) => DataPath_RF_bus_reg_dataout_2151_port,
                           regs(2150) => DataPath_RF_bus_reg_dataout_2150_port,
                           regs(2149) => DataPath_RF_bus_reg_dataout_2149_port,
                           regs(2148) => DataPath_RF_bus_reg_dataout_2148_port,
                           regs(2147) => DataPath_RF_bus_reg_dataout_2147_port,
                           regs(2146) => DataPath_RF_bus_reg_dataout_2146_port,
                           regs(2145) => DataPath_RF_bus_reg_dataout_2145_port,
                           regs(2144) => DataPath_RF_bus_reg_dataout_2144_port,
                           regs(2143) => DataPath_RF_bus_reg_dataout_2143_port,
                           regs(2142) => DataPath_RF_bus_reg_dataout_2142_port,
                           regs(2141) => DataPath_RF_bus_reg_dataout_2141_port,
                           regs(2140) => DataPath_RF_bus_reg_dataout_2140_port,
                           regs(2139) => DataPath_RF_bus_reg_dataout_2139_port,
                           regs(2138) => DataPath_RF_bus_reg_dataout_2138_port,
                           regs(2137) => DataPath_RF_bus_reg_dataout_2137_port,
                           regs(2136) => DataPath_RF_bus_reg_dataout_2136_port,
                           regs(2135) => DataPath_RF_bus_reg_dataout_2135_port,
                           regs(2134) => DataPath_RF_bus_reg_dataout_2134_port,
                           regs(2133) => DataPath_RF_bus_reg_dataout_2133_port,
                           regs(2132) => DataPath_RF_bus_reg_dataout_2132_port,
                           regs(2131) => DataPath_RF_bus_reg_dataout_2131_port,
                           regs(2130) => DataPath_RF_bus_reg_dataout_2130_port,
                           regs(2129) => DataPath_RF_bus_reg_dataout_2129_port,
                           regs(2128) => DataPath_RF_bus_reg_dataout_2128_port,
                           regs(2127) => DataPath_RF_bus_reg_dataout_2127_port,
                           regs(2126) => DataPath_RF_bus_reg_dataout_2126_port,
                           regs(2125) => DataPath_RF_bus_reg_dataout_2125_port,
                           regs(2124) => DataPath_RF_bus_reg_dataout_2124_port,
                           regs(2123) => DataPath_RF_bus_reg_dataout_2123_port,
                           regs(2122) => DataPath_RF_bus_reg_dataout_2122_port,
                           regs(2121) => DataPath_RF_bus_reg_dataout_2121_port,
                           regs(2120) => DataPath_RF_bus_reg_dataout_2120_port,
                           regs(2119) => DataPath_RF_bus_reg_dataout_2119_port,
                           regs(2118) => DataPath_RF_bus_reg_dataout_2118_port,
                           regs(2117) => DataPath_RF_bus_reg_dataout_2117_port,
                           regs(2116) => DataPath_RF_bus_reg_dataout_2116_port,
                           regs(2115) => DataPath_RF_bus_reg_dataout_2115_port,
                           regs(2114) => DataPath_RF_bus_reg_dataout_2114_port,
                           regs(2113) => DataPath_RF_bus_reg_dataout_2113_port,
                           regs(2112) => DataPath_RF_bus_reg_dataout_2112_port,
                           regs(2111) => DataPath_RF_bus_reg_dataout_2111_port,
                           regs(2110) => DataPath_RF_bus_reg_dataout_2110_port,
                           regs(2109) => DataPath_RF_bus_reg_dataout_2109_port,
                           regs(2108) => DataPath_RF_bus_reg_dataout_2108_port,
                           regs(2107) => DataPath_RF_bus_reg_dataout_2107_port,
                           regs(2106) => DataPath_RF_bus_reg_dataout_2106_port,
                           regs(2105) => DataPath_RF_bus_reg_dataout_2105_port,
                           regs(2104) => DataPath_RF_bus_reg_dataout_2104_port,
                           regs(2103) => DataPath_RF_bus_reg_dataout_2103_port,
                           regs(2102) => DataPath_RF_bus_reg_dataout_2102_port,
                           regs(2101) => DataPath_RF_bus_reg_dataout_2101_port,
                           regs(2100) => DataPath_RF_bus_reg_dataout_2100_port,
                           regs(2099) => DataPath_RF_bus_reg_dataout_2099_port,
                           regs(2098) => DataPath_RF_bus_reg_dataout_2098_port,
                           regs(2097) => DataPath_RF_bus_reg_dataout_2097_port,
                           regs(2096) => DataPath_RF_bus_reg_dataout_2096_port,
                           regs(2095) => DataPath_RF_bus_reg_dataout_2095_port,
                           regs(2094) => DataPath_RF_bus_reg_dataout_2094_port,
                           regs(2093) => DataPath_RF_bus_reg_dataout_2093_port,
                           regs(2092) => DataPath_RF_bus_reg_dataout_2092_port,
                           regs(2091) => DataPath_RF_bus_reg_dataout_2091_port,
                           regs(2090) => DataPath_RF_bus_reg_dataout_2090_port,
                           regs(2089) => DataPath_RF_bus_reg_dataout_2089_port,
                           regs(2088) => DataPath_RF_bus_reg_dataout_2088_port,
                           regs(2087) => DataPath_RF_bus_reg_dataout_2087_port,
                           regs(2086) => DataPath_RF_bus_reg_dataout_2086_port,
                           regs(2085) => DataPath_RF_bus_reg_dataout_2085_port,
                           regs(2084) => DataPath_RF_bus_reg_dataout_2084_port,
                           regs(2083) => DataPath_RF_bus_reg_dataout_2083_port,
                           regs(2082) => DataPath_RF_bus_reg_dataout_2082_port,
                           regs(2081) => DataPath_RF_bus_reg_dataout_2081_port,
                           regs(2080) => DataPath_RF_bus_reg_dataout_2080_port,
                           regs(2079) => DataPath_RF_bus_reg_dataout_2079_port,
                           regs(2078) => DataPath_RF_bus_reg_dataout_2078_port,
                           regs(2077) => DataPath_RF_bus_reg_dataout_2077_port,
                           regs(2076) => DataPath_RF_bus_reg_dataout_2076_port,
                           regs(2075) => DataPath_RF_bus_reg_dataout_2075_port,
                           regs(2074) => DataPath_RF_bus_reg_dataout_2074_port,
                           regs(2073) => DataPath_RF_bus_reg_dataout_2073_port,
                           regs(2072) => DataPath_RF_bus_reg_dataout_2072_port,
                           regs(2071) => DataPath_RF_bus_reg_dataout_2071_port,
                           regs(2070) => DataPath_RF_bus_reg_dataout_2070_port,
                           regs(2069) => DataPath_RF_bus_reg_dataout_2069_port,
                           regs(2068) => DataPath_RF_bus_reg_dataout_2068_port,
                           regs(2067) => DataPath_RF_bus_reg_dataout_2067_port,
                           regs(2066) => DataPath_RF_bus_reg_dataout_2066_port,
                           regs(2065) => DataPath_RF_bus_reg_dataout_2065_port,
                           regs(2064) => DataPath_RF_bus_reg_dataout_2064_port,
                           regs(2063) => DataPath_RF_bus_reg_dataout_2063_port,
                           regs(2062) => DataPath_RF_bus_reg_dataout_2062_port,
                           regs(2061) => DataPath_RF_bus_reg_dataout_2061_port,
                           regs(2060) => DataPath_RF_bus_reg_dataout_2060_port,
                           regs(2059) => DataPath_RF_bus_reg_dataout_2059_port,
                           regs(2058) => DataPath_RF_bus_reg_dataout_2058_port,
                           regs(2057) => DataPath_RF_bus_reg_dataout_2057_port,
                           regs(2056) => DataPath_RF_bus_reg_dataout_2056_port,
                           regs(2055) => DataPath_RF_bus_reg_dataout_2055_port,
                           regs(2054) => DataPath_RF_bus_reg_dataout_2054_port,
                           regs(2053) => DataPath_RF_bus_reg_dataout_2053_port,
                           regs(2052) => DataPath_RF_bus_reg_dataout_2052_port,
                           regs(2051) => DataPath_RF_bus_reg_dataout_2051_port,
                           regs(2050) => DataPath_RF_bus_reg_dataout_2050_port,
                           regs(2049) => DataPath_RF_bus_reg_dataout_2049_port,
                           regs(2048) => DataPath_RF_bus_reg_dataout_2048_port,
                           regs(2047) => DataPath_RF_bus_reg_dataout_2047_port,
                           regs(2046) => DataPath_RF_bus_reg_dataout_2046_port,
                           regs(2045) => DataPath_RF_bus_reg_dataout_2045_port,
                           regs(2044) => DataPath_RF_bus_reg_dataout_2044_port,
                           regs(2043) => DataPath_RF_bus_reg_dataout_2043_port,
                           regs(2042) => DataPath_RF_bus_reg_dataout_2042_port,
                           regs(2041) => DataPath_RF_bus_reg_dataout_2041_port,
                           regs(2040) => DataPath_RF_bus_reg_dataout_2040_port,
                           regs(2039) => DataPath_RF_bus_reg_dataout_2039_port,
                           regs(2038) => DataPath_RF_bus_reg_dataout_2038_port,
                           regs(2037) => DataPath_RF_bus_reg_dataout_2037_port,
                           regs(2036) => DataPath_RF_bus_reg_dataout_2036_port,
                           regs(2035) => DataPath_RF_bus_reg_dataout_2035_port,
                           regs(2034) => DataPath_RF_bus_reg_dataout_2034_port,
                           regs(2033) => DataPath_RF_bus_reg_dataout_2033_port,
                           regs(2032) => DataPath_RF_bus_reg_dataout_2032_port,
                           regs(2031) => DataPath_RF_bus_reg_dataout_2031_port,
                           regs(2030) => DataPath_RF_bus_reg_dataout_2030_port,
                           regs(2029) => DataPath_RF_bus_reg_dataout_2029_port,
                           regs(2028) => DataPath_RF_bus_reg_dataout_2028_port,
                           regs(2027) => DataPath_RF_bus_reg_dataout_2027_port,
                           regs(2026) => DataPath_RF_bus_reg_dataout_2026_port,
                           regs(2025) => DataPath_RF_bus_reg_dataout_2025_port,
                           regs(2024) => DataPath_RF_bus_reg_dataout_2024_port,
                           regs(2023) => DataPath_RF_bus_reg_dataout_2023_port,
                           regs(2022) => DataPath_RF_bus_reg_dataout_2022_port,
                           regs(2021) => DataPath_RF_bus_reg_dataout_2021_port,
                           regs(2020) => DataPath_RF_bus_reg_dataout_2020_port,
                           regs(2019) => DataPath_RF_bus_reg_dataout_2019_port,
                           regs(2018) => DataPath_RF_bus_reg_dataout_2018_port,
                           regs(2017) => DataPath_RF_bus_reg_dataout_2017_port,
                           regs(2016) => DataPath_RF_bus_reg_dataout_2016_port,
                           regs(2015) => DataPath_RF_bus_reg_dataout_2015_port,
                           regs(2014) => DataPath_RF_bus_reg_dataout_2014_port,
                           regs(2013) => DataPath_RF_bus_reg_dataout_2013_port,
                           regs(2012) => DataPath_RF_bus_reg_dataout_2012_port,
                           regs(2011) => DataPath_RF_bus_reg_dataout_2011_port,
                           regs(2010) => DataPath_RF_bus_reg_dataout_2010_port,
                           regs(2009) => DataPath_RF_bus_reg_dataout_2009_port,
                           regs(2008) => DataPath_RF_bus_reg_dataout_2008_port,
                           regs(2007) => DataPath_RF_bus_reg_dataout_2007_port,
                           regs(2006) => DataPath_RF_bus_reg_dataout_2006_port,
                           regs(2005) => DataPath_RF_bus_reg_dataout_2005_port,
                           regs(2004) => DataPath_RF_bus_reg_dataout_2004_port,
                           regs(2003) => DataPath_RF_bus_reg_dataout_2003_port,
                           regs(2002) => DataPath_RF_bus_reg_dataout_2002_port,
                           regs(2001) => DataPath_RF_bus_reg_dataout_2001_port,
                           regs(2000) => DataPath_RF_bus_reg_dataout_2000_port,
                           regs(1999) => DataPath_RF_bus_reg_dataout_1999_port,
                           regs(1998) => DataPath_RF_bus_reg_dataout_1998_port,
                           regs(1997) => DataPath_RF_bus_reg_dataout_1997_port,
                           regs(1996) => DataPath_RF_bus_reg_dataout_1996_port,
                           regs(1995) => DataPath_RF_bus_reg_dataout_1995_port,
                           regs(1994) => DataPath_RF_bus_reg_dataout_1994_port,
                           regs(1993) => DataPath_RF_bus_reg_dataout_1993_port,
                           regs(1992) => DataPath_RF_bus_reg_dataout_1992_port,
                           regs(1991) => DataPath_RF_bus_reg_dataout_1991_port,
                           regs(1990) => DataPath_RF_bus_reg_dataout_1990_port,
                           regs(1989) => DataPath_RF_bus_reg_dataout_1989_port,
                           regs(1988) => DataPath_RF_bus_reg_dataout_1988_port,
                           regs(1987) => DataPath_RF_bus_reg_dataout_1987_port,
                           regs(1986) => DataPath_RF_bus_reg_dataout_1986_port,
                           regs(1985) => DataPath_RF_bus_reg_dataout_1985_port,
                           regs(1984) => DataPath_RF_bus_reg_dataout_1984_port,
                           regs(1983) => DataPath_RF_bus_reg_dataout_1983_port,
                           regs(1982) => DataPath_RF_bus_reg_dataout_1982_port,
                           regs(1981) => DataPath_RF_bus_reg_dataout_1981_port,
                           regs(1980) => DataPath_RF_bus_reg_dataout_1980_port,
                           regs(1979) => DataPath_RF_bus_reg_dataout_1979_port,
                           regs(1978) => DataPath_RF_bus_reg_dataout_1978_port,
                           regs(1977) => DataPath_RF_bus_reg_dataout_1977_port,
                           regs(1976) => DataPath_RF_bus_reg_dataout_1976_port,
                           regs(1975) => DataPath_RF_bus_reg_dataout_1975_port,
                           regs(1974) => DataPath_RF_bus_reg_dataout_1974_port,
                           regs(1973) => DataPath_RF_bus_reg_dataout_1973_port,
                           regs(1972) => DataPath_RF_bus_reg_dataout_1972_port,
                           regs(1971) => DataPath_RF_bus_reg_dataout_1971_port,
                           regs(1970) => DataPath_RF_bus_reg_dataout_1970_port,
                           regs(1969) => DataPath_RF_bus_reg_dataout_1969_port,
                           regs(1968) => DataPath_RF_bus_reg_dataout_1968_port,
                           regs(1967) => DataPath_RF_bus_reg_dataout_1967_port,
                           regs(1966) => DataPath_RF_bus_reg_dataout_1966_port,
                           regs(1965) => DataPath_RF_bus_reg_dataout_1965_port,
                           regs(1964) => DataPath_RF_bus_reg_dataout_1964_port,
                           regs(1963) => DataPath_RF_bus_reg_dataout_1963_port,
                           regs(1962) => DataPath_RF_bus_reg_dataout_1962_port,
                           regs(1961) => DataPath_RF_bus_reg_dataout_1961_port,
                           regs(1960) => DataPath_RF_bus_reg_dataout_1960_port,
                           regs(1959) => DataPath_RF_bus_reg_dataout_1959_port,
                           regs(1958) => DataPath_RF_bus_reg_dataout_1958_port,
                           regs(1957) => DataPath_RF_bus_reg_dataout_1957_port,
                           regs(1956) => DataPath_RF_bus_reg_dataout_1956_port,
                           regs(1955) => DataPath_RF_bus_reg_dataout_1955_port,
                           regs(1954) => DataPath_RF_bus_reg_dataout_1954_port,
                           regs(1953) => DataPath_RF_bus_reg_dataout_1953_port,
                           regs(1952) => DataPath_RF_bus_reg_dataout_1952_port,
                           regs(1951) => DataPath_RF_bus_reg_dataout_1951_port,
                           regs(1950) => DataPath_RF_bus_reg_dataout_1950_port,
                           regs(1949) => DataPath_RF_bus_reg_dataout_1949_port,
                           regs(1948) => DataPath_RF_bus_reg_dataout_1948_port,
                           regs(1947) => DataPath_RF_bus_reg_dataout_1947_port,
                           regs(1946) => DataPath_RF_bus_reg_dataout_1946_port,
                           regs(1945) => DataPath_RF_bus_reg_dataout_1945_port,
                           regs(1944) => DataPath_RF_bus_reg_dataout_1944_port,
                           regs(1943) => DataPath_RF_bus_reg_dataout_1943_port,
                           regs(1942) => DataPath_RF_bus_reg_dataout_1942_port,
                           regs(1941) => DataPath_RF_bus_reg_dataout_1941_port,
                           regs(1940) => DataPath_RF_bus_reg_dataout_1940_port,
                           regs(1939) => DataPath_RF_bus_reg_dataout_1939_port,
                           regs(1938) => DataPath_RF_bus_reg_dataout_1938_port,
                           regs(1937) => DataPath_RF_bus_reg_dataout_1937_port,
                           regs(1936) => DataPath_RF_bus_reg_dataout_1936_port,
                           regs(1935) => DataPath_RF_bus_reg_dataout_1935_port,
                           regs(1934) => DataPath_RF_bus_reg_dataout_1934_port,
                           regs(1933) => DataPath_RF_bus_reg_dataout_1933_port,
                           regs(1932) => DataPath_RF_bus_reg_dataout_1932_port,
                           regs(1931) => DataPath_RF_bus_reg_dataout_1931_port,
                           regs(1930) => DataPath_RF_bus_reg_dataout_1930_port,
                           regs(1929) => DataPath_RF_bus_reg_dataout_1929_port,
                           regs(1928) => DataPath_RF_bus_reg_dataout_1928_port,
                           regs(1927) => DataPath_RF_bus_reg_dataout_1927_port,
                           regs(1926) => DataPath_RF_bus_reg_dataout_1926_port,
                           regs(1925) => DataPath_RF_bus_reg_dataout_1925_port,
                           regs(1924) => DataPath_RF_bus_reg_dataout_1924_port,
                           regs(1923) => DataPath_RF_bus_reg_dataout_1923_port,
                           regs(1922) => DataPath_RF_bus_reg_dataout_1922_port,
                           regs(1921) => DataPath_RF_bus_reg_dataout_1921_port,
                           regs(1920) => DataPath_RF_bus_reg_dataout_1920_port,
                           regs(1919) => DataPath_RF_bus_reg_dataout_1919_port,
                           regs(1918) => DataPath_RF_bus_reg_dataout_1918_port,
                           regs(1917) => DataPath_RF_bus_reg_dataout_1917_port,
                           regs(1916) => DataPath_RF_bus_reg_dataout_1916_port,
                           regs(1915) => DataPath_RF_bus_reg_dataout_1915_port,
                           regs(1914) => DataPath_RF_bus_reg_dataout_1914_port,
                           regs(1913) => DataPath_RF_bus_reg_dataout_1913_port,
                           regs(1912) => DataPath_RF_bus_reg_dataout_1912_port,
                           regs(1911) => DataPath_RF_bus_reg_dataout_1911_port,
                           regs(1910) => DataPath_RF_bus_reg_dataout_1910_port,
                           regs(1909) => DataPath_RF_bus_reg_dataout_1909_port,
                           regs(1908) => DataPath_RF_bus_reg_dataout_1908_port,
                           regs(1907) => DataPath_RF_bus_reg_dataout_1907_port,
                           regs(1906) => DataPath_RF_bus_reg_dataout_1906_port,
                           regs(1905) => DataPath_RF_bus_reg_dataout_1905_port,
                           regs(1904) => DataPath_RF_bus_reg_dataout_1904_port,
                           regs(1903) => DataPath_RF_bus_reg_dataout_1903_port,
                           regs(1902) => DataPath_RF_bus_reg_dataout_1902_port,
                           regs(1901) => DataPath_RF_bus_reg_dataout_1901_port,
                           regs(1900) => DataPath_RF_bus_reg_dataout_1900_port,
                           regs(1899) => DataPath_RF_bus_reg_dataout_1899_port,
                           regs(1898) => DataPath_RF_bus_reg_dataout_1898_port,
                           regs(1897) => DataPath_RF_bus_reg_dataout_1897_port,
                           regs(1896) => DataPath_RF_bus_reg_dataout_1896_port,
                           regs(1895) => DataPath_RF_bus_reg_dataout_1895_port,
                           regs(1894) => DataPath_RF_bus_reg_dataout_1894_port,
                           regs(1893) => DataPath_RF_bus_reg_dataout_1893_port,
                           regs(1892) => DataPath_RF_bus_reg_dataout_1892_port,
                           regs(1891) => DataPath_RF_bus_reg_dataout_1891_port,
                           regs(1890) => DataPath_RF_bus_reg_dataout_1890_port,
                           regs(1889) => DataPath_RF_bus_reg_dataout_1889_port,
                           regs(1888) => DataPath_RF_bus_reg_dataout_1888_port,
                           regs(1887) => DataPath_RF_bus_reg_dataout_1887_port,
                           regs(1886) => DataPath_RF_bus_reg_dataout_1886_port,
                           regs(1885) => DataPath_RF_bus_reg_dataout_1885_port,
                           regs(1884) => DataPath_RF_bus_reg_dataout_1884_port,
                           regs(1883) => DataPath_RF_bus_reg_dataout_1883_port,
                           regs(1882) => DataPath_RF_bus_reg_dataout_1882_port,
                           regs(1881) => DataPath_RF_bus_reg_dataout_1881_port,
                           regs(1880) => DataPath_RF_bus_reg_dataout_1880_port,
                           regs(1879) => DataPath_RF_bus_reg_dataout_1879_port,
                           regs(1878) => DataPath_RF_bus_reg_dataout_1878_port,
                           regs(1877) => DataPath_RF_bus_reg_dataout_1877_port,
                           regs(1876) => DataPath_RF_bus_reg_dataout_1876_port,
                           regs(1875) => DataPath_RF_bus_reg_dataout_1875_port,
                           regs(1874) => DataPath_RF_bus_reg_dataout_1874_port,
                           regs(1873) => DataPath_RF_bus_reg_dataout_1873_port,
                           regs(1872) => DataPath_RF_bus_reg_dataout_1872_port,
                           regs(1871) => DataPath_RF_bus_reg_dataout_1871_port,
                           regs(1870) => DataPath_RF_bus_reg_dataout_1870_port,
                           regs(1869) => DataPath_RF_bus_reg_dataout_1869_port,
                           regs(1868) => DataPath_RF_bus_reg_dataout_1868_port,
                           regs(1867) => DataPath_RF_bus_reg_dataout_1867_port,
                           regs(1866) => DataPath_RF_bus_reg_dataout_1866_port,
                           regs(1865) => DataPath_RF_bus_reg_dataout_1865_port,
                           regs(1864) => DataPath_RF_bus_reg_dataout_1864_port,
                           regs(1863) => DataPath_RF_bus_reg_dataout_1863_port,
                           regs(1862) => DataPath_RF_bus_reg_dataout_1862_port,
                           regs(1861) => DataPath_RF_bus_reg_dataout_1861_port,
                           regs(1860) => DataPath_RF_bus_reg_dataout_1860_port,
                           regs(1859) => DataPath_RF_bus_reg_dataout_1859_port,
                           regs(1858) => DataPath_RF_bus_reg_dataout_1858_port,
                           regs(1857) => DataPath_RF_bus_reg_dataout_1857_port,
                           regs(1856) => DataPath_RF_bus_reg_dataout_1856_port,
                           regs(1855) => DataPath_RF_bus_reg_dataout_1855_port,
                           regs(1854) => DataPath_RF_bus_reg_dataout_1854_port,
                           regs(1853) => DataPath_RF_bus_reg_dataout_1853_port,
                           regs(1852) => DataPath_RF_bus_reg_dataout_1852_port,
                           regs(1851) => DataPath_RF_bus_reg_dataout_1851_port,
                           regs(1850) => DataPath_RF_bus_reg_dataout_1850_port,
                           regs(1849) => DataPath_RF_bus_reg_dataout_1849_port,
                           regs(1848) => DataPath_RF_bus_reg_dataout_1848_port,
                           regs(1847) => DataPath_RF_bus_reg_dataout_1847_port,
                           regs(1846) => DataPath_RF_bus_reg_dataout_1846_port,
                           regs(1845) => DataPath_RF_bus_reg_dataout_1845_port,
                           regs(1844) => DataPath_RF_bus_reg_dataout_1844_port,
                           regs(1843) => DataPath_RF_bus_reg_dataout_1843_port,
                           regs(1842) => DataPath_RF_bus_reg_dataout_1842_port,
                           regs(1841) => DataPath_RF_bus_reg_dataout_1841_port,
                           regs(1840) => DataPath_RF_bus_reg_dataout_1840_port,
                           regs(1839) => DataPath_RF_bus_reg_dataout_1839_port,
                           regs(1838) => DataPath_RF_bus_reg_dataout_1838_port,
                           regs(1837) => DataPath_RF_bus_reg_dataout_1837_port,
                           regs(1836) => DataPath_RF_bus_reg_dataout_1836_port,
                           regs(1835) => DataPath_RF_bus_reg_dataout_1835_port,
                           regs(1834) => DataPath_RF_bus_reg_dataout_1834_port,
                           regs(1833) => DataPath_RF_bus_reg_dataout_1833_port,
                           regs(1832) => DataPath_RF_bus_reg_dataout_1832_port,
                           regs(1831) => DataPath_RF_bus_reg_dataout_1831_port,
                           regs(1830) => DataPath_RF_bus_reg_dataout_1830_port,
                           regs(1829) => DataPath_RF_bus_reg_dataout_1829_port,
                           regs(1828) => DataPath_RF_bus_reg_dataout_1828_port,
                           regs(1827) => DataPath_RF_bus_reg_dataout_1827_port,
                           regs(1826) => DataPath_RF_bus_reg_dataout_1826_port,
                           regs(1825) => DataPath_RF_bus_reg_dataout_1825_port,
                           regs(1824) => DataPath_RF_bus_reg_dataout_1824_port,
                           regs(1823) => DataPath_RF_bus_reg_dataout_1823_port,
                           regs(1822) => DataPath_RF_bus_reg_dataout_1822_port,
                           regs(1821) => DataPath_RF_bus_reg_dataout_1821_port,
                           regs(1820) => DataPath_RF_bus_reg_dataout_1820_port,
                           regs(1819) => DataPath_RF_bus_reg_dataout_1819_port,
                           regs(1818) => DataPath_RF_bus_reg_dataout_1818_port,
                           regs(1817) => DataPath_RF_bus_reg_dataout_1817_port,
                           regs(1816) => DataPath_RF_bus_reg_dataout_1816_port,
                           regs(1815) => DataPath_RF_bus_reg_dataout_1815_port,
                           regs(1814) => DataPath_RF_bus_reg_dataout_1814_port,
                           regs(1813) => DataPath_RF_bus_reg_dataout_1813_port,
                           regs(1812) => DataPath_RF_bus_reg_dataout_1812_port,
                           regs(1811) => DataPath_RF_bus_reg_dataout_1811_port,
                           regs(1810) => DataPath_RF_bus_reg_dataout_1810_port,
                           regs(1809) => DataPath_RF_bus_reg_dataout_1809_port,
                           regs(1808) => DataPath_RF_bus_reg_dataout_1808_port,
                           regs(1807) => DataPath_RF_bus_reg_dataout_1807_port,
                           regs(1806) => DataPath_RF_bus_reg_dataout_1806_port,
                           regs(1805) => DataPath_RF_bus_reg_dataout_1805_port,
                           regs(1804) => DataPath_RF_bus_reg_dataout_1804_port,
                           regs(1803) => DataPath_RF_bus_reg_dataout_1803_port,
                           regs(1802) => DataPath_RF_bus_reg_dataout_1802_port,
                           regs(1801) => DataPath_RF_bus_reg_dataout_1801_port,
                           regs(1800) => DataPath_RF_bus_reg_dataout_1800_port,
                           regs(1799) => DataPath_RF_bus_reg_dataout_1799_port,
                           regs(1798) => DataPath_RF_bus_reg_dataout_1798_port,
                           regs(1797) => DataPath_RF_bus_reg_dataout_1797_port,
                           regs(1796) => DataPath_RF_bus_reg_dataout_1796_port,
                           regs(1795) => DataPath_RF_bus_reg_dataout_1795_port,
                           regs(1794) => DataPath_RF_bus_reg_dataout_1794_port,
                           regs(1793) => DataPath_RF_bus_reg_dataout_1793_port,
                           regs(1792) => DataPath_RF_bus_reg_dataout_1792_port,
                           regs(1791) => DataPath_RF_bus_reg_dataout_1791_port,
                           regs(1790) => DataPath_RF_bus_reg_dataout_1790_port,
                           regs(1789) => DataPath_RF_bus_reg_dataout_1789_port,
                           regs(1788) => DataPath_RF_bus_reg_dataout_1788_port,
                           regs(1787) => DataPath_RF_bus_reg_dataout_1787_port,
                           regs(1786) => DataPath_RF_bus_reg_dataout_1786_port,
                           regs(1785) => DataPath_RF_bus_reg_dataout_1785_port,
                           regs(1784) => DataPath_RF_bus_reg_dataout_1784_port,
                           regs(1783) => DataPath_RF_bus_reg_dataout_1783_port,
                           regs(1782) => DataPath_RF_bus_reg_dataout_1782_port,
                           regs(1781) => DataPath_RF_bus_reg_dataout_1781_port,
                           regs(1780) => DataPath_RF_bus_reg_dataout_1780_port,
                           regs(1779) => DataPath_RF_bus_reg_dataout_1779_port,
                           regs(1778) => DataPath_RF_bus_reg_dataout_1778_port,
                           regs(1777) => DataPath_RF_bus_reg_dataout_1777_port,
                           regs(1776) => DataPath_RF_bus_reg_dataout_1776_port,
                           regs(1775) => DataPath_RF_bus_reg_dataout_1775_port,
                           regs(1774) => DataPath_RF_bus_reg_dataout_1774_port,
                           regs(1773) => DataPath_RF_bus_reg_dataout_1773_port,
                           regs(1772) => DataPath_RF_bus_reg_dataout_1772_port,
                           regs(1771) => DataPath_RF_bus_reg_dataout_1771_port,
                           regs(1770) => DataPath_RF_bus_reg_dataout_1770_port,
                           regs(1769) => DataPath_RF_bus_reg_dataout_1769_port,
                           regs(1768) => DataPath_RF_bus_reg_dataout_1768_port,
                           regs(1767) => DataPath_RF_bus_reg_dataout_1767_port,
                           regs(1766) => DataPath_RF_bus_reg_dataout_1766_port,
                           regs(1765) => DataPath_RF_bus_reg_dataout_1765_port,
                           regs(1764) => DataPath_RF_bus_reg_dataout_1764_port,
                           regs(1763) => DataPath_RF_bus_reg_dataout_1763_port,
                           regs(1762) => DataPath_RF_bus_reg_dataout_1762_port,
                           regs(1761) => DataPath_RF_bus_reg_dataout_1761_port,
                           regs(1760) => DataPath_RF_bus_reg_dataout_1760_port,
                           regs(1759) => DataPath_RF_bus_reg_dataout_1759_port,
                           regs(1758) => DataPath_RF_bus_reg_dataout_1758_port,
                           regs(1757) => DataPath_RF_bus_reg_dataout_1757_port,
                           regs(1756) => DataPath_RF_bus_reg_dataout_1756_port,
                           regs(1755) => DataPath_RF_bus_reg_dataout_1755_port,
                           regs(1754) => DataPath_RF_bus_reg_dataout_1754_port,
                           regs(1753) => DataPath_RF_bus_reg_dataout_1753_port,
                           regs(1752) => DataPath_RF_bus_reg_dataout_1752_port,
                           regs(1751) => DataPath_RF_bus_reg_dataout_1751_port,
                           regs(1750) => DataPath_RF_bus_reg_dataout_1750_port,
                           regs(1749) => DataPath_RF_bus_reg_dataout_1749_port,
                           regs(1748) => DataPath_RF_bus_reg_dataout_1748_port,
                           regs(1747) => DataPath_RF_bus_reg_dataout_1747_port,
                           regs(1746) => DataPath_RF_bus_reg_dataout_1746_port,
                           regs(1745) => DataPath_RF_bus_reg_dataout_1745_port,
                           regs(1744) => DataPath_RF_bus_reg_dataout_1744_port,
                           regs(1743) => DataPath_RF_bus_reg_dataout_1743_port,
                           regs(1742) => DataPath_RF_bus_reg_dataout_1742_port,
                           regs(1741) => DataPath_RF_bus_reg_dataout_1741_port,
                           regs(1740) => DataPath_RF_bus_reg_dataout_1740_port,
                           regs(1739) => DataPath_RF_bus_reg_dataout_1739_port,
                           regs(1738) => DataPath_RF_bus_reg_dataout_1738_port,
                           regs(1737) => DataPath_RF_bus_reg_dataout_1737_port,
                           regs(1736) => DataPath_RF_bus_reg_dataout_1736_port,
                           regs(1735) => DataPath_RF_bus_reg_dataout_1735_port,
                           regs(1734) => DataPath_RF_bus_reg_dataout_1734_port,
                           regs(1733) => DataPath_RF_bus_reg_dataout_1733_port,
                           regs(1732) => DataPath_RF_bus_reg_dataout_1732_port,
                           regs(1731) => DataPath_RF_bus_reg_dataout_1731_port,
                           regs(1730) => DataPath_RF_bus_reg_dataout_1730_port,
                           regs(1729) => DataPath_RF_bus_reg_dataout_1729_port,
                           regs(1728) => DataPath_RF_bus_reg_dataout_1728_port,
                           regs(1727) => DataPath_RF_bus_reg_dataout_1727_port,
                           regs(1726) => DataPath_RF_bus_reg_dataout_1726_port,
                           regs(1725) => DataPath_RF_bus_reg_dataout_1725_port,
                           regs(1724) => DataPath_RF_bus_reg_dataout_1724_port,
                           regs(1723) => DataPath_RF_bus_reg_dataout_1723_port,
                           regs(1722) => DataPath_RF_bus_reg_dataout_1722_port,
                           regs(1721) => DataPath_RF_bus_reg_dataout_1721_port,
                           regs(1720) => DataPath_RF_bus_reg_dataout_1720_port,
                           regs(1719) => DataPath_RF_bus_reg_dataout_1719_port,
                           regs(1718) => DataPath_RF_bus_reg_dataout_1718_port,
                           regs(1717) => DataPath_RF_bus_reg_dataout_1717_port,
                           regs(1716) => DataPath_RF_bus_reg_dataout_1716_port,
                           regs(1715) => DataPath_RF_bus_reg_dataout_1715_port,
                           regs(1714) => DataPath_RF_bus_reg_dataout_1714_port,
                           regs(1713) => DataPath_RF_bus_reg_dataout_1713_port,
                           regs(1712) => DataPath_RF_bus_reg_dataout_1712_port,
                           regs(1711) => DataPath_RF_bus_reg_dataout_1711_port,
                           regs(1710) => DataPath_RF_bus_reg_dataout_1710_port,
                           regs(1709) => DataPath_RF_bus_reg_dataout_1709_port,
                           regs(1708) => DataPath_RF_bus_reg_dataout_1708_port,
                           regs(1707) => DataPath_RF_bus_reg_dataout_1707_port,
                           regs(1706) => DataPath_RF_bus_reg_dataout_1706_port,
                           regs(1705) => DataPath_RF_bus_reg_dataout_1705_port,
                           regs(1704) => DataPath_RF_bus_reg_dataout_1704_port,
                           regs(1703) => DataPath_RF_bus_reg_dataout_1703_port,
                           regs(1702) => DataPath_RF_bus_reg_dataout_1702_port,
                           regs(1701) => DataPath_RF_bus_reg_dataout_1701_port,
                           regs(1700) => DataPath_RF_bus_reg_dataout_1700_port,
                           regs(1699) => DataPath_RF_bus_reg_dataout_1699_port,
                           regs(1698) => DataPath_RF_bus_reg_dataout_1698_port,
                           regs(1697) => DataPath_RF_bus_reg_dataout_1697_port,
                           regs(1696) => DataPath_RF_bus_reg_dataout_1696_port,
                           regs(1695) => DataPath_RF_bus_reg_dataout_1695_port,
                           regs(1694) => DataPath_RF_bus_reg_dataout_1694_port,
                           regs(1693) => DataPath_RF_bus_reg_dataout_1693_port,
                           regs(1692) => DataPath_RF_bus_reg_dataout_1692_port,
                           regs(1691) => DataPath_RF_bus_reg_dataout_1691_port,
                           regs(1690) => DataPath_RF_bus_reg_dataout_1690_port,
                           regs(1689) => DataPath_RF_bus_reg_dataout_1689_port,
                           regs(1688) => DataPath_RF_bus_reg_dataout_1688_port,
                           regs(1687) => DataPath_RF_bus_reg_dataout_1687_port,
                           regs(1686) => DataPath_RF_bus_reg_dataout_1686_port,
                           regs(1685) => DataPath_RF_bus_reg_dataout_1685_port,
                           regs(1684) => DataPath_RF_bus_reg_dataout_1684_port,
                           regs(1683) => DataPath_RF_bus_reg_dataout_1683_port,
                           regs(1682) => DataPath_RF_bus_reg_dataout_1682_port,
                           regs(1681) => DataPath_RF_bus_reg_dataout_1681_port,
                           regs(1680) => DataPath_RF_bus_reg_dataout_1680_port,
                           regs(1679) => DataPath_RF_bus_reg_dataout_1679_port,
                           regs(1678) => DataPath_RF_bus_reg_dataout_1678_port,
                           regs(1677) => DataPath_RF_bus_reg_dataout_1677_port,
                           regs(1676) => DataPath_RF_bus_reg_dataout_1676_port,
                           regs(1675) => DataPath_RF_bus_reg_dataout_1675_port,
                           regs(1674) => DataPath_RF_bus_reg_dataout_1674_port,
                           regs(1673) => DataPath_RF_bus_reg_dataout_1673_port,
                           regs(1672) => DataPath_RF_bus_reg_dataout_1672_port,
                           regs(1671) => DataPath_RF_bus_reg_dataout_1671_port,
                           regs(1670) => DataPath_RF_bus_reg_dataout_1670_port,
                           regs(1669) => DataPath_RF_bus_reg_dataout_1669_port,
                           regs(1668) => DataPath_RF_bus_reg_dataout_1668_port,
                           regs(1667) => DataPath_RF_bus_reg_dataout_1667_port,
                           regs(1666) => DataPath_RF_bus_reg_dataout_1666_port,
                           regs(1665) => DataPath_RF_bus_reg_dataout_1665_port,
                           regs(1664) => DataPath_RF_bus_reg_dataout_1664_port,
                           regs(1663) => DataPath_RF_bus_reg_dataout_1663_port,
                           regs(1662) => DataPath_RF_bus_reg_dataout_1662_port,
                           regs(1661) => DataPath_RF_bus_reg_dataout_1661_port,
                           regs(1660) => DataPath_RF_bus_reg_dataout_1660_port,
                           regs(1659) => DataPath_RF_bus_reg_dataout_1659_port,
                           regs(1658) => DataPath_RF_bus_reg_dataout_1658_port,
                           regs(1657) => DataPath_RF_bus_reg_dataout_1657_port,
                           regs(1656) => DataPath_RF_bus_reg_dataout_1656_port,
                           regs(1655) => DataPath_RF_bus_reg_dataout_1655_port,
                           regs(1654) => DataPath_RF_bus_reg_dataout_1654_port,
                           regs(1653) => DataPath_RF_bus_reg_dataout_1653_port,
                           regs(1652) => DataPath_RF_bus_reg_dataout_1652_port,
                           regs(1651) => DataPath_RF_bus_reg_dataout_1651_port,
                           regs(1650) => DataPath_RF_bus_reg_dataout_1650_port,
                           regs(1649) => DataPath_RF_bus_reg_dataout_1649_port,
                           regs(1648) => DataPath_RF_bus_reg_dataout_1648_port,
                           regs(1647) => DataPath_RF_bus_reg_dataout_1647_port,
                           regs(1646) => DataPath_RF_bus_reg_dataout_1646_port,
                           regs(1645) => DataPath_RF_bus_reg_dataout_1645_port,
                           regs(1644) => DataPath_RF_bus_reg_dataout_1644_port,
                           regs(1643) => DataPath_RF_bus_reg_dataout_1643_port,
                           regs(1642) => DataPath_RF_bus_reg_dataout_1642_port,
                           regs(1641) => DataPath_RF_bus_reg_dataout_1641_port,
                           regs(1640) => DataPath_RF_bus_reg_dataout_1640_port,
                           regs(1639) => DataPath_RF_bus_reg_dataout_1639_port,
                           regs(1638) => DataPath_RF_bus_reg_dataout_1638_port,
                           regs(1637) => DataPath_RF_bus_reg_dataout_1637_port,
                           regs(1636) => DataPath_RF_bus_reg_dataout_1636_port,
                           regs(1635) => DataPath_RF_bus_reg_dataout_1635_port,
                           regs(1634) => DataPath_RF_bus_reg_dataout_1634_port,
                           regs(1633) => DataPath_RF_bus_reg_dataout_1633_port,
                           regs(1632) => DataPath_RF_bus_reg_dataout_1632_port,
                           regs(1631) => DataPath_RF_bus_reg_dataout_1631_port,
                           regs(1630) => DataPath_RF_bus_reg_dataout_1630_port,
                           regs(1629) => DataPath_RF_bus_reg_dataout_1629_port,
                           regs(1628) => DataPath_RF_bus_reg_dataout_1628_port,
                           regs(1627) => DataPath_RF_bus_reg_dataout_1627_port,
                           regs(1626) => DataPath_RF_bus_reg_dataout_1626_port,
                           regs(1625) => DataPath_RF_bus_reg_dataout_1625_port,
                           regs(1624) => DataPath_RF_bus_reg_dataout_1624_port,
                           regs(1623) => DataPath_RF_bus_reg_dataout_1623_port,
                           regs(1622) => DataPath_RF_bus_reg_dataout_1622_port,
                           regs(1621) => DataPath_RF_bus_reg_dataout_1621_port,
                           regs(1620) => DataPath_RF_bus_reg_dataout_1620_port,
                           regs(1619) => DataPath_RF_bus_reg_dataout_1619_port,
                           regs(1618) => DataPath_RF_bus_reg_dataout_1618_port,
                           regs(1617) => DataPath_RF_bus_reg_dataout_1617_port,
                           regs(1616) => DataPath_RF_bus_reg_dataout_1616_port,
                           regs(1615) => DataPath_RF_bus_reg_dataout_1615_port,
                           regs(1614) => DataPath_RF_bus_reg_dataout_1614_port,
                           regs(1613) => DataPath_RF_bus_reg_dataout_1613_port,
                           regs(1612) => DataPath_RF_bus_reg_dataout_1612_port,
                           regs(1611) => DataPath_RF_bus_reg_dataout_1611_port,
                           regs(1610) => DataPath_RF_bus_reg_dataout_1610_port,
                           regs(1609) => DataPath_RF_bus_reg_dataout_1609_port,
                           regs(1608) => DataPath_RF_bus_reg_dataout_1608_port,
                           regs(1607) => DataPath_RF_bus_reg_dataout_1607_port,
                           regs(1606) => DataPath_RF_bus_reg_dataout_1606_port,
                           regs(1605) => DataPath_RF_bus_reg_dataout_1605_port,
                           regs(1604) => DataPath_RF_bus_reg_dataout_1604_port,
                           regs(1603) => DataPath_RF_bus_reg_dataout_1603_port,
                           regs(1602) => DataPath_RF_bus_reg_dataout_1602_port,
                           regs(1601) => DataPath_RF_bus_reg_dataout_1601_port,
                           regs(1600) => DataPath_RF_bus_reg_dataout_1600_port,
                           regs(1599) => DataPath_RF_bus_reg_dataout_1599_port,
                           regs(1598) => DataPath_RF_bus_reg_dataout_1598_port,
                           regs(1597) => DataPath_RF_bus_reg_dataout_1597_port,
                           regs(1596) => DataPath_RF_bus_reg_dataout_1596_port,
                           regs(1595) => DataPath_RF_bus_reg_dataout_1595_port,
                           regs(1594) => DataPath_RF_bus_reg_dataout_1594_port,
                           regs(1593) => DataPath_RF_bus_reg_dataout_1593_port,
                           regs(1592) => DataPath_RF_bus_reg_dataout_1592_port,
                           regs(1591) => DataPath_RF_bus_reg_dataout_1591_port,
                           regs(1590) => DataPath_RF_bus_reg_dataout_1590_port,
                           regs(1589) => DataPath_RF_bus_reg_dataout_1589_port,
                           regs(1588) => DataPath_RF_bus_reg_dataout_1588_port,
                           regs(1587) => DataPath_RF_bus_reg_dataout_1587_port,
                           regs(1586) => DataPath_RF_bus_reg_dataout_1586_port,
                           regs(1585) => DataPath_RF_bus_reg_dataout_1585_port,
                           regs(1584) => DataPath_RF_bus_reg_dataout_1584_port,
                           regs(1583) => DataPath_RF_bus_reg_dataout_1583_port,
                           regs(1582) => DataPath_RF_bus_reg_dataout_1582_port,
                           regs(1581) => DataPath_RF_bus_reg_dataout_1581_port,
                           regs(1580) => DataPath_RF_bus_reg_dataout_1580_port,
                           regs(1579) => DataPath_RF_bus_reg_dataout_1579_port,
                           regs(1578) => DataPath_RF_bus_reg_dataout_1578_port,
                           regs(1577) => DataPath_RF_bus_reg_dataout_1577_port,
                           regs(1576) => DataPath_RF_bus_reg_dataout_1576_port,
                           regs(1575) => DataPath_RF_bus_reg_dataout_1575_port,
                           regs(1574) => DataPath_RF_bus_reg_dataout_1574_port,
                           regs(1573) => DataPath_RF_bus_reg_dataout_1573_port,
                           regs(1572) => DataPath_RF_bus_reg_dataout_1572_port,
                           regs(1571) => DataPath_RF_bus_reg_dataout_1571_port,
                           regs(1570) => DataPath_RF_bus_reg_dataout_1570_port,
                           regs(1569) => DataPath_RF_bus_reg_dataout_1569_port,
                           regs(1568) => DataPath_RF_bus_reg_dataout_1568_port,
                           regs(1567) => DataPath_RF_bus_reg_dataout_1567_port,
                           regs(1566) => DataPath_RF_bus_reg_dataout_1566_port,
                           regs(1565) => DataPath_RF_bus_reg_dataout_1565_port,
                           regs(1564) => DataPath_RF_bus_reg_dataout_1564_port,
                           regs(1563) => DataPath_RF_bus_reg_dataout_1563_port,
                           regs(1562) => DataPath_RF_bus_reg_dataout_1562_port,
                           regs(1561) => DataPath_RF_bus_reg_dataout_1561_port,
                           regs(1560) => DataPath_RF_bus_reg_dataout_1560_port,
                           regs(1559) => DataPath_RF_bus_reg_dataout_1559_port,
                           regs(1558) => DataPath_RF_bus_reg_dataout_1558_port,
                           regs(1557) => DataPath_RF_bus_reg_dataout_1557_port,
                           regs(1556) => DataPath_RF_bus_reg_dataout_1556_port,
                           regs(1555) => DataPath_RF_bus_reg_dataout_1555_port,
                           regs(1554) => DataPath_RF_bus_reg_dataout_1554_port,
                           regs(1553) => DataPath_RF_bus_reg_dataout_1553_port,
                           regs(1552) => DataPath_RF_bus_reg_dataout_1552_port,
                           regs(1551) => DataPath_RF_bus_reg_dataout_1551_port,
                           regs(1550) => DataPath_RF_bus_reg_dataout_1550_port,
                           regs(1549) => DataPath_RF_bus_reg_dataout_1549_port,
                           regs(1548) => DataPath_RF_bus_reg_dataout_1548_port,
                           regs(1547) => DataPath_RF_bus_reg_dataout_1547_port,
                           regs(1546) => DataPath_RF_bus_reg_dataout_1546_port,
                           regs(1545) => DataPath_RF_bus_reg_dataout_1545_port,
                           regs(1544) => DataPath_RF_bus_reg_dataout_1544_port,
                           regs(1543) => DataPath_RF_bus_reg_dataout_1543_port,
                           regs(1542) => DataPath_RF_bus_reg_dataout_1542_port,
                           regs(1541) => DataPath_RF_bus_reg_dataout_1541_port,
                           regs(1540) => DataPath_RF_bus_reg_dataout_1540_port,
                           regs(1539) => DataPath_RF_bus_reg_dataout_1539_port,
                           regs(1538) => DataPath_RF_bus_reg_dataout_1538_port,
                           regs(1537) => DataPath_RF_bus_reg_dataout_1537_port,
                           regs(1536) => DataPath_RF_bus_reg_dataout_1536_port,
                           regs(1535) => DataPath_RF_bus_reg_dataout_1535_port,
                           regs(1534) => DataPath_RF_bus_reg_dataout_1534_port,
                           regs(1533) => DataPath_RF_bus_reg_dataout_1533_port,
                           regs(1532) => DataPath_RF_bus_reg_dataout_1532_port,
                           regs(1531) => DataPath_RF_bus_reg_dataout_1531_port,
                           regs(1530) => DataPath_RF_bus_reg_dataout_1530_port,
                           regs(1529) => DataPath_RF_bus_reg_dataout_1529_port,
                           regs(1528) => DataPath_RF_bus_reg_dataout_1528_port,
                           regs(1527) => DataPath_RF_bus_reg_dataout_1527_port,
                           regs(1526) => DataPath_RF_bus_reg_dataout_1526_port,
                           regs(1525) => DataPath_RF_bus_reg_dataout_1525_port,
                           regs(1524) => DataPath_RF_bus_reg_dataout_1524_port,
                           regs(1523) => DataPath_RF_bus_reg_dataout_1523_port,
                           regs(1522) => DataPath_RF_bus_reg_dataout_1522_port,
                           regs(1521) => DataPath_RF_bus_reg_dataout_1521_port,
                           regs(1520) => DataPath_RF_bus_reg_dataout_1520_port,
                           regs(1519) => DataPath_RF_bus_reg_dataout_1519_port,
                           regs(1518) => DataPath_RF_bus_reg_dataout_1518_port,
                           regs(1517) => DataPath_RF_bus_reg_dataout_1517_port,
                           regs(1516) => DataPath_RF_bus_reg_dataout_1516_port,
                           regs(1515) => DataPath_RF_bus_reg_dataout_1515_port,
                           regs(1514) => DataPath_RF_bus_reg_dataout_1514_port,
                           regs(1513) => DataPath_RF_bus_reg_dataout_1513_port,
                           regs(1512) => DataPath_RF_bus_reg_dataout_1512_port,
                           regs(1511) => DataPath_RF_bus_reg_dataout_1511_port,
                           regs(1510) => DataPath_RF_bus_reg_dataout_1510_port,
                           regs(1509) => DataPath_RF_bus_reg_dataout_1509_port,
                           regs(1508) => DataPath_RF_bus_reg_dataout_1508_port,
                           regs(1507) => DataPath_RF_bus_reg_dataout_1507_port,
                           regs(1506) => DataPath_RF_bus_reg_dataout_1506_port,
                           regs(1505) => DataPath_RF_bus_reg_dataout_1505_port,
                           regs(1504) => DataPath_RF_bus_reg_dataout_1504_port,
                           regs(1503) => DataPath_RF_bus_reg_dataout_1503_port,
                           regs(1502) => DataPath_RF_bus_reg_dataout_1502_port,
                           regs(1501) => DataPath_RF_bus_reg_dataout_1501_port,
                           regs(1500) => DataPath_RF_bus_reg_dataout_1500_port,
                           regs(1499) => DataPath_RF_bus_reg_dataout_1499_port,
                           regs(1498) => DataPath_RF_bus_reg_dataout_1498_port,
                           regs(1497) => DataPath_RF_bus_reg_dataout_1497_port,
                           regs(1496) => DataPath_RF_bus_reg_dataout_1496_port,
                           regs(1495) => DataPath_RF_bus_reg_dataout_1495_port,
                           regs(1494) => DataPath_RF_bus_reg_dataout_1494_port,
                           regs(1493) => DataPath_RF_bus_reg_dataout_1493_port,
                           regs(1492) => DataPath_RF_bus_reg_dataout_1492_port,
                           regs(1491) => DataPath_RF_bus_reg_dataout_1491_port,
                           regs(1490) => DataPath_RF_bus_reg_dataout_1490_port,
                           regs(1489) => DataPath_RF_bus_reg_dataout_1489_port,
                           regs(1488) => DataPath_RF_bus_reg_dataout_1488_port,
                           regs(1487) => DataPath_RF_bus_reg_dataout_1487_port,
                           regs(1486) => DataPath_RF_bus_reg_dataout_1486_port,
                           regs(1485) => DataPath_RF_bus_reg_dataout_1485_port,
                           regs(1484) => DataPath_RF_bus_reg_dataout_1484_port,
                           regs(1483) => DataPath_RF_bus_reg_dataout_1483_port,
                           regs(1482) => DataPath_RF_bus_reg_dataout_1482_port,
                           regs(1481) => DataPath_RF_bus_reg_dataout_1481_port,
                           regs(1480) => DataPath_RF_bus_reg_dataout_1480_port,
                           regs(1479) => DataPath_RF_bus_reg_dataout_1479_port,
                           regs(1478) => DataPath_RF_bus_reg_dataout_1478_port,
                           regs(1477) => DataPath_RF_bus_reg_dataout_1477_port,
                           regs(1476) => DataPath_RF_bus_reg_dataout_1476_port,
                           regs(1475) => DataPath_RF_bus_reg_dataout_1475_port,
                           regs(1474) => DataPath_RF_bus_reg_dataout_1474_port,
                           regs(1473) => DataPath_RF_bus_reg_dataout_1473_port,
                           regs(1472) => DataPath_RF_bus_reg_dataout_1472_port,
                           regs(1471) => DataPath_RF_bus_reg_dataout_1471_port,
                           regs(1470) => DataPath_RF_bus_reg_dataout_1470_port,
                           regs(1469) => DataPath_RF_bus_reg_dataout_1469_port,
                           regs(1468) => DataPath_RF_bus_reg_dataout_1468_port,
                           regs(1467) => DataPath_RF_bus_reg_dataout_1467_port,
                           regs(1466) => DataPath_RF_bus_reg_dataout_1466_port,
                           regs(1465) => DataPath_RF_bus_reg_dataout_1465_port,
                           regs(1464) => DataPath_RF_bus_reg_dataout_1464_port,
                           regs(1463) => DataPath_RF_bus_reg_dataout_1463_port,
                           regs(1462) => DataPath_RF_bus_reg_dataout_1462_port,
                           regs(1461) => DataPath_RF_bus_reg_dataout_1461_port,
                           regs(1460) => DataPath_RF_bus_reg_dataout_1460_port,
                           regs(1459) => DataPath_RF_bus_reg_dataout_1459_port,
                           regs(1458) => DataPath_RF_bus_reg_dataout_1458_port,
                           regs(1457) => DataPath_RF_bus_reg_dataout_1457_port,
                           regs(1456) => DataPath_RF_bus_reg_dataout_1456_port,
                           regs(1455) => DataPath_RF_bus_reg_dataout_1455_port,
                           regs(1454) => DataPath_RF_bus_reg_dataout_1454_port,
                           regs(1453) => DataPath_RF_bus_reg_dataout_1453_port,
                           regs(1452) => DataPath_RF_bus_reg_dataout_1452_port,
                           regs(1451) => DataPath_RF_bus_reg_dataout_1451_port,
                           regs(1450) => DataPath_RF_bus_reg_dataout_1450_port,
                           regs(1449) => DataPath_RF_bus_reg_dataout_1449_port,
                           regs(1448) => DataPath_RF_bus_reg_dataout_1448_port,
                           regs(1447) => DataPath_RF_bus_reg_dataout_1447_port,
                           regs(1446) => DataPath_RF_bus_reg_dataout_1446_port,
                           regs(1445) => DataPath_RF_bus_reg_dataout_1445_port,
                           regs(1444) => DataPath_RF_bus_reg_dataout_1444_port,
                           regs(1443) => DataPath_RF_bus_reg_dataout_1443_port,
                           regs(1442) => DataPath_RF_bus_reg_dataout_1442_port,
                           regs(1441) => DataPath_RF_bus_reg_dataout_1441_port,
                           regs(1440) => DataPath_RF_bus_reg_dataout_1440_port,
                           regs(1439) => DataPath_RF_bus_reg_dataout_1439_port,
                           regs(1438) => DataPath_RF_bus_reg_dataout_1438_port,
                           regs(1437) => DataPath_RF_bus_reg_dataout_1437_port,
                           regs(1436) => DataPath_RF_bus_reg_dataout_1436_port,
                           regs(1435) => DataPath_RF_bus_reg_dataout_1435_port,
                           regs(1434) => DataPath_RF_bus_reg_dataout_1434_port,
                           regs(1433) => DataPath_RF_bus_reg_dataout_1433_port,
                           regs(1432) => DataPath_RF_bus_reg_dataout_1432_port,
                           regs(1431) => DataPath_RF_bus_reg_dataout_1431_port,
                           regs(1430) => DataPath_RF_bus_reg_dataout_1430_port,
                           regs(1429) => DataPath_RF_bus_reg_dataout_1429_port,
                           regs(1428) => DataPath_RF_bus_reg_dataout_1428_port,
                           regs(1427) => DataPath_RF_bus_reg_dataout_1427_port,
                           regs(1426) => DataPath_RF_bus_reg_dataout_1426_port,
                           regs(1425) => DataPath_RF_bus_reg_dataout_1425_port,
                           regs(1424) => DataPath_RF_bus_reg_dataout_1424_port,
                           regs(1423) => DataPath_RF_bus_reg_dataout_1423_port,
                           regs(1422) => DataPath_RF_bus_reg_dataout_1422_port,
                           regs(1421) => DataPath_RF_bus_reg_dataout_1421_port,
                           regs(1420) => DataPath_RF_bus_reg_dataout_1420_port,
                           regs(1419) => DataPath_RF_bus_reg_dataout_1419_port,
                           regs(1418) => DataPath_RF_bus_reg_dataout_1418_port,
                           regs(1417) => DataPath_RF_bus_reg_dataout_1417_port,
                           regs(1416) => DataPath_RF_bus_reg_dataout_1416_port,
                           regs(1415) => DataPath_RF_bus_reg_dataout_1415_port,
                           regs(1414) => DataPath_RF_bus_reg_dataout_1414_port,
                           regs(1413) => DataPath_RF_bus_reg_dataout_1413_port,
                           regs(1412) => DataPath_RF_bus_reg_dataout_1412_port,
                           regs(1411) => DataPath_RF_bus_reg_dataout_1411_port,
                           regs(1410) => DataPath_RF_bus_reg_dataout_1410_port,
                           regs(1409) => DataPath_RF_bus_reg_dataout_1409_port,
                           regs(1408) => DataPath_RF_bus_reg_dataout_1408_port,
                           regs(1407) => DataPath_RF_bus_reg_dataout_1407_port,
                           regs(1406) => DataPath_RF_bus_reg_dataout_1406_port,
                           regs(1405) => DataPath_RF_bus_reg_dataout_1405_port,
                           regs(1404) => DataPath_RF_bus_reg_dataout_1404_port,
                           regs(1403) => DataPath_RF_bus_reg_dataout_1403_port,
                           regs(1402) => DataPath_RF_bus_reg_dataout_1402_port,
                           regs(1401) => DataPath_RF_bus_reg_dataout_1401_port,
                           regs(1400) => DataPath_RF_bus_reg_dataout_1400_port,
                           regs(1399) => DataPath_RF_bus_reg_dataout_1399_port,
                           regs(1398) => DataPath_RF_bus_reg_dataout_1398_port,
                           regs(1397) => DataPath_RF_bus_reg_dataout_1397_port,
                           regs(1396) => DataPath_RF_bus_reg_dataout_1396_port,
                           regs(1395) => DataPath_RF_bus_reg_dataout_1395_port,
                           regs(1394) => DataPath_RF_bus_reg_dataout_1394_port,
                           regs(1393) => DataPath_RF_bus_reg_dataout_1393_port,
                           regs(1392) => DataPath_RF_bus_reg_dataout_1392_port,
                           regs(1391) => DataPath_RF_bus_reg_dataout_1391_port,
                           regs(1390) => DataPath_RF_bus_reg_dataout_1390_port,
                           regs(1389) => DataPath_RF_bus_reg_dataout_1389_port,
                           regs(1388) => DataPath_RF_bus_reg_dataout_1388_port,
                           regs(1387) => DataPath_RF_bus_reg_dataout_1387_port,
                           regs(1386) => DataPath_RF_bus_reg_dataout_1386_port,
                           regs(1385) => DataPath_RF_bus_reg_dataout_1385_port,
                           regs(1384) => DataPath_RF_bus_reg_dataout_1384_port,
                           regs(1383) => DataPath_RF_bus_reg_dataout_1383_port,
                           regs(1382) => DataPath_RF_bus_reg_dataout_1382_port,
                           regs(1381) => DataPath_RF_bus_reg_dataout_1381_port,
                           regs(1380) => DataPath_RF_bus_reg_dataout_1380_port,
                           regs(1379) => DataPath_RF_bus_reg_dataout_1379_port,
                           regs(1378) => DataPath_RF_bus_reg_dataout_1378_port,
                           regs(1377) => DataPath_RF_bus_reg_dataout_1377_port,
                           regs(1376) => DataPath_RF_bus_reg_dataout_1376_port,
                           regs(1375) => DataPath_RF_bus_reg_dataout_1375_port,
                           regs(1374) => DataPath_RF_bus_reg_dataout_1374_port,
                           regs(1373) => DataPath_RF_bus_reg_dataout_1373_port,
                           regs(1372) => DataPath_RF_bus_reg_dataout_1372_port,
                           regs(1371) => DataPath_RF_bus_reg_dataout_1371_port,
                           regs(1370) => DataPath_RF_bus_reg_dataout_1370_port,
                           regs(1369) => DataPath_RF_bus_reg_dataout_1369_port,
                           regs(1368) => DataPath_RF_bus_reg_dataout_1368_port,
                           regs(1367) => DataPath_RF_bus_reg_dataout_1367_port,
                           regs(1366) => DataPath_RF_bus_reg_dataout_1366_port,
                           regs(1365) => DataPath_RF_bus_reg_dataout_1365_port,
                           regs(1364) => DataPath_RF_bus_reg_dataout_1364_port,
                           regs(1363) => DataPath_RF_bus_reg_dataout_1363_port,
                           regs(1362) => DataPath_RF_bus_reg_dataout_1362_port,
                           regs(1361) => DataPath_RF_bus_reg_dataout_1361_port,
                           regs(1360) => DataPath_RF_bus_reg_dataout_1360_port,
                           regs(1359) => DataPath_RF_bus_reg_dataout_1359_port,
                           regs(1358) => DataPath_RF_bus_reg_dataout_1358_port,
                           regs(1357) => DataPath_RF_bus_reg_dataout_1357_port,
                           regs(1356) => DataPath_RF_bus_reg_dataout_1356_port,
                           regs(1355) => DataPath_RF_bus_reg_dataout_1355_port,
                           regs(1354) => DataPath_RF_bus_reg_dataout_1354_port,
                           regs(1353) => DataPath_RF_bus_reg_dataout_1353_port,
                           regs(1352) => DataPath_RF_bus_reg_dataout_1352_port,
                           regs(1351) => DataPath_RF_bus_reg_dataout_1351_port,
                           regs(1350) => DataPath_RF_bus_reg_dataout_1350_port,
                           regs(1349) => DataPath_RF_bus_reg_dataout_1349_port,
                           regs(1348) => DataPath_RF_bus_reg_dataout_1348_port,
                           regs(1347) => DataPath_RF_bus_reg_dataout_1347_port,
                           regs(1346) => DataPath_RF_bus_reg_dataout_1346_port,
                           regs(1345) => DataPath_RF_bus_reg_dataout_1345_port,
                           regs(1344) => DataPath_RF_bus_reg_dataout_1344_port,
                           regs(1343) => DataPath_RF_bus_reg_dataout_1343_port,
                           regs(1342) => DataPath_RF_bus_reg_dataout_1342_port,
                           regs(1341) => DataPath_RF_bus_reg_dataout_1341_port,
                           regs(1340) => DataPath_RF_bus_reg_dataout_1340_port,
                           regs(1339) => DataPath_RF_bus_reg_dataout_1339_port,
                           regs(1338) => DataPath_RF_bus_reg_dataout_1338_port,
                           regs(1337) => DataPath_RF_bus_reg_dataout_1337_port,
                           regs(1336) => DataPath_RF_bus_reg_dataout_1336_port,
                           regs(1335) => DataPath_RF_bus_reg_dataout_1335_port,
                           regs(1334) => DataPath_RF_bus_reg_dataout_1334_port,
                           regs(1333) => DataPath_RF_bus_reg_dataout_1333_port,
                           regs(1332) => DataPath_RF_bus_reg_dataout_1332_port,
                           regs(1331) => DataPath_RF_bus_reg_dataout_1331_port,
                           regs(1330) => DataPath_RF_bus_reg_dataout_1330_port,
                           regs(1329) => DataPath_RF_bus_reg_dataout_1329_port,
                           regs(1328) => DataPath_RF_bus_reg_dataout_1328_port,
                           regs(1327) => DataPath_RF_bus_reg_dataout_1327_port,
                           regs(1326) => DataPath_RF_bus_reg_dataout_1326_port,
                           regs(1325) => DataPath_RF_bus_reg_dataout_1325_port,
                           regs(1324) => DataPath_RF_bus_reg_dataout_1324_port,
                           regs(1323) => DataPath_RF_bus_reg_dataout_1323_port,
                           regs(1322) => DataPath_RF_bus_reg_dataout_1322_port,
                           regs(1321) => DataPath_RF_bus_reg_dataout_1321_port,
                           regs(1320) => DataPath_RF_bus_reg_dataout_1320_port,
                           regs(1319) => DataPath_RF_bus_reg_dataout_1319_port,
                           regs(1318) => DataPath_RF_bus_reg_dataout_1318_port,
                           regs(1317) => DataPath_RF_bus_reg_dataout_1317_port,
                           regs(1316) => DataPath_RF_bus_reg_dataout_1316_port,
                           regs(1315) => DataPath_RF_bus_reg_dataout_1315_port,
                           regs(1314) => DataPath_RF_bus_reg_dataout_1314_port,
                           regs(1313) => DataPath_RF_bus_reg_dataout_1313_port,
                           regs(1312) => DataPath_RF_bus_reg_dataout_1312_port,
                           regs(1311) => DataPath_RF_bus_reg_dataout_1311_port,
                           regs(1310) => DataPath_RF_bus_reg_dataout_1310_port,
                           regs(1309) => DataPath_RF_bus_reg_dataout_1309_port,
                           regs(1308) => DataPath_RF_bus_reg_dataout_1308_port,
                           regs(1307) => DataPath_RF_bus_reg_dataout_1307_port,
                           regs(1306) => DataPath_RF_bus_reg_dataout_1306_port,
                           regs(1305) => DataPath_RF_bus_reg_dataout_1305_port,
                           regs(1304) => DataPath_RF_bus_reg_dataout_1304_port,
                           regs(1303) => DataPath_RF_bus_reg_dataout_1303_port,
                           regs(1302) => DataPath_RF_bus_reg_dataout_1302_port,
                           regs(1301) => DataPath_RF_bus_reg_dataout_1301_port,
                           regs(1300) => DataPath_RF_bus_reg_dataout_1300_port,
                           regs(1299) => DataPath_RF_bus_reg_dataout_1299_port,
                           regs(1298) => DataPath_RF_bus_reg_dataout_1298_port,
                           regs(1297) => DataPath_RF_bus_reg_dataout_1297_port,
                           regs(1296) => DataPath_RF_bus_reg_dataout_1296_port,
                           regs(1295) => DataPath_RF_bus_reg_dataout_1295_port,
                           regs(1294) => DataPath_RF_bus_reg_dataout_1294_port,
                           regs(1293) => DataPath_RF_bus_reg_dataout_1293_port,
                           regs(1292) => DataPath_RF_bus_reg_dataout_1292_port,
                           regs(1291) => DataPath_RF_bus_reg_dataout_1291_port,
                           regs(1290) => DataPath_RF_bus_reg_dataout_1290_port,
                           regs(1289) => DataPath_RF_bus_reg_dataout_1289_port,
                           regs(1288) => DataPath_RF_bus_reg_dataout_1288_port,
                           regs(1287) => DataPath_RF_bus_reg_dataout_1287_port,
                           regs(1286) => DataPath_RF_bus_reg_dataout_1286_port,
                           regs(1285) => DataPath_RF_bus_reg_dataout_1285_port,
                           regs(1284) => DataPath_RF_bus_reg_dataout_1284_port,
                           regs(1283) => DataPath_RF_bus_reg_dataout_1283_port,
                           regs(1282) => DataPath_RF_bus_reg_dataout_1282_port,
                           regs(1281) => DataPath_RF_bus_reg_dataout_1281_port,
                           regs(1280) => DataPath_RF_bus_reg_dataout_1280_port,
                           regs(1279) => DataPath_RF_bus_reg_dataout_1279_port,
                           regs(1278) => DataPath_RF_bus_reg_dataout_1278_port,
                           regs(1277) => DataPath_RF_bus_reg_dataout_1277_port,
                           regs(1276) => DataPath_RF_bus_reg_dataout_1276_port,
                           regs(1275) => DataPath_RF_bus_reg_dataout_1275_port,
                           regs(1274) => DataPath_RF_bus_reg_dataout_1274_port,
                           regs(1273) => DataPath_RF_bus_reg_dataout_1273_port,
                           regs(1272) => DataPath_RF_bus_reg_dataout_1272_port,
                           regs(1271) => DataPath_RF_bus_reg_dataout_1271_port,
                           regs(1270) => DataPath_RF_bus_reg_dataout_1270_port,
                           regs(1269) => DataPath_RF_bus_reg_dataout_1269_port,
                           regs(1268) => DataPath_RF_bus_reg_dataout_1268_port,
                           regs(1267) => DataPath_RF_bus_reg_dataout_1267_port,
                           regs(1266) => DataPath_RF_bus_reg_dataout_1266_port,
                           regs(1265) => DataPath_RF_bus_reg_dataout_1265_port,
                           regs(1264) => DataPath_RF_bus_reg_dataout_1264_port,
                           regs(1263) => DataPath_RF_bus_reg_dataout_1263_port,
                           regs(1262) => DataPath_RF_bus_reg_dataout_1262_port,
                           regs(1261) => DataPath_RF_bus_reg_dataout_1261_port,
                           regs(1260) => DataPath_RF_bus_reg_dataout_1260_port,
                           regs(1259) => DataPath_RF_bus_reg_dataout_1259_port,
                           regs(1258) => DataPath_RF_bus_reg_dataout_1258_port,
                           regs(1257) => DataPath_RF_bus_reg_dataout_1257_port,
                           regs(1256) => DataPath_RF_bus_reg_dataout_1256_port,
                           regs(1255) => DataPath_RF_bus_reg_dataout_1255_port,
                           regs(1254) => DataPath_RF_bus_reg_dataout_1254_port,
                           regs(1253) => DataPath_RF_bus_reg_dataout_1253_port,
                           regs(1252) => DataPath_RF_bus_reg_dataout_1252_port,
                           regs(1251) => DataPath_RF_bus_reg_dataout_1251_port,
                           regs(1250) => DataPath_RF_bus_reg_dataout_1250_port,
                           regs(1249) => DataPath_RF_bus_reg_dataout_1249_port,
                           regs(1248) => DataPath_RF_bus_reg_dataout_1248_port,
                           regs(1247) => DataPath_RF_bus_reg_dataout_1247_port,
                           regs(1246) => DataPath_RF_bus_reg_dataout_1246_port,
                           regs(1245) => DataPath_RF_bus_reg_dataout_1245_port,
                           regs(1244) => DataPath_RF_bus_reg_dataout_1244_port,
                           regs(1243) => DataPath_RF_bus_reg_dataout_1243_port,
                           regs(1242) => DataPath_RF_bus_reg_dataout_1242_port,
                           regs(1241) => DataPath_RF_bus_reg_dataout_1241_port,
                           regs(1240) => DataPath_RF_bus_reg_dataout_1240_port,
                           regs(1239) => DataPath_RF_bus_reg_dataout_1239_port,
                           regs(1238) => DataPath_RF_bus_reg_dataout_1238_port,
                           regs(1237) => DataPath_RF_bus_reg_dataout_1237_port,
                           regs(1236) => DataPath_RF_bus_reg_dataout_1236_port,
                           regs(1235) => DataPath_RF_bus_reg_dataout_1235_port,
                           regs(1234) => DataPath_RF_bus_reg_dataout_1234_port,
                           regs(1233) => DataPath_RF_bus_reg_dataout_1233_port,
                           regs(1232) => DataPath_RF_bus_reg_dataout_1232_port,
                           regs(1231) => DataPath_RF_bus_reg_dataout_1231_port,
                           regs(1230) => DataPath_RF_bus_reg_dataout_1230_port,
                           regs(1229) => DataPath_RF_bus_reg_dataout_1229_port,
                           regs(1228) => DataPath_RF_bus_reg_dataout_1228_port,
                           regs(1227) => DataPath_RF_bus_reg_dataout_1227_port,
                           regs(1226) => DataPath_RF_bus_reg_dataout_1226_port,
                           regs(1225) => DataPath_RF_bus_reg_dataout_1225_port,
                           regs(1224) => DataPath_RF_bus_reg_dataout_1224_port,
                           regs(1223) => DataPath_RF_bus_reg_dataout_1223_port,
                           regs(1222) => DataPath_RF_bus_reg_dataout_1222_port,
                           regs(1221) => DataPath_RF_bus_reg_dataout_1221_port,
                           regs(1220) => DataPath_RF_bus_reg_dataout_1220_port,
                           regs(1219) => DataPath_RF_bus_reg_dataout_1219_port,
                           regs(1218) => DataPath_RF_bus_reg_dataout_1218_port,
                           regs(1217) => DataPath_RF_bus_reg_dataout_1217_port,
                           regs(1216) => DataPath_RF_bus_reg_dataout_1216_port,
                           regs(1215) => DataPath_RF_bus_reg_dataout_1215_port,
                           regs(1214) => DataPath_RF_bus_reg_dataout_1214_port,
                           regs(1213) => DataPath_RF_bus_reg_dataout_1213_port,
                           regs(1212) => DataPath_RF_bus_reg_dataout_1212_port,
                           regs(1211) => DataPath_RF_bus_reg_dataout_1211_port,
                           regs(1210) => DataPath_RF_bus_reg_dataout_1210_port,
                           regs(1209) => DataPath_RF_bus_reg_dataout_1209_port,
                           regs(1208) => DataPath_RF_bus_reg_dataout_1208_port,
                           regs(1207) => DataPath_RF_bus_reg_dataout_1207_port,
                           regs(1206) => DataPath_RF_bus_reg_dataout_1206_port,
                           regs(1205) => DataPath_RF_bus_reg_dataout_1205_port,
                           regs(1204) => DataPath_RF_bus_reg_dataout_1204_port,
                           regs(1203) => DataPath_RF_bus_reg_dataout_1203_port,
                           regs(1202) => DataPath_RF_bus_reg_dataout_1202_port,
                           regs(1201) => DataPath_RF_bus_reg_dataout_1201_port,
                           regs(1200) => DataPath_RF_bus_reg_dataout_1200_port,
                           regs(1199) => DataPath_RF_bus_reg_dataout_1199_port,
                           regs(1198) => DataPath_RF_bus_reg_dataout_1198_port,
                           regs(1197) => DataPath_RF_bus_reg_dataout_1197_port,
                           regs(1196) => DataPath_RF_bus_reg_dataout_1196_port,
                           regs(1195) => DataPath_RF_bus_reg_dataout_1195_port,
                           regs(1194) => DataPath_RF_bus_reg_dataout_1194_port,
                           regs(1193) => DataPath_RF_bus_reg_dataout_1193_port,
                           regs(1192) => DataPath_RF_bus_reg_dataout_1192_port,
                           regs(1191) => DataPath_RF_bus_reg_dataout_1191_port,
                           regs(1190) => DataPath_RF_bus_reg_dataout_1190_port,
                           regs(1189) => DataPath_RF_bus_reg_dataout_1189_port,
                           regs(1188) => DataPath_RF_bus_reg_dataout_1188_port,
                           regs(1187) => DataPath_RF_bus_reg_dataout_1187_port,
                           regs(1186) => DataPath_RF_bus_reg_dataout_1186_port,
                           regs(1185) => DataPath_RF_bus_reg_dataout_1185_port,
                           regs(1184) => DataPath_RF_bus_reg_dataout_1184_port,
                           regs(1183) => DataPath_RF_bus_reg_dataout_1183_port,
                           regs(1182) => DataPath_RF_bus_reg_dataout_1182_port,
                           regs(1181) => DataPath_RF_bus_reg_dataout_1181_port,
                           regs(1180) => DataPath_RF_bus_reg_dataout_1180_port,
                           regs(1179) => DataPath_RF_bus_reg_dataout_1179_port,
                           regs(1178) => DataPath_RF_bus_reg_dataout_1178_port,
                           regs(1177) => DataPath_RF_bus_reg_dataout_1177_port,
                           regs(1176) => DataPath_RF_bus_reg_dataout_1176_port,
                           regs(1175) => DataPath_RF_bus_reg_dataout_1175_port,
                           regs(1174) => DataPath_RF_bus_reg_dataout_1174_port,
                           regs(1173) => DataPath_RF_bus_reg_dataout_1173_port,
                           regs(1172) => DataPath_RF_bus_reg_dataout_1172_port,
                           regs(1171) => DataPath_RF_bus_reg_dataout_1171_port,
                           regs(1170) => DataPath_RF_bus_reg_dataout_1170_port,
                           regs(1169) => DataPath_RF_bus_reg_dataout_1169_port,
                           regs(1168) => DataPath_RF_bus_reg_dataout_1168_port,
                           regs(1167) => DataPath_RF_bus_reg_dataout_1167_port,
                           regs(1166) => DataPath_RF_bus_reg_dataout_1166_port,
                           regs(1165) => DataPath_RF_bus_reg_dataout_1165_port,
                           regs(1164) => DataPath_RF_bus_reg_dataout_1164_port,
                           regs(1163) => DataPath_RF_bus_reg_dataout_1163_port,
                           regs(1162) => DataPath_RF_bus_reg_dataout_1162_port,
                           regs(1161) => DataPath_RF_bus_reg_dataout_1161_port,
                           regs(1160) => DataPath_RF_bus_reg_dataout_1160_port,
                           regs(1159) => DataPath_RF_bus_reg_dataout_1159_port,
                           regs(1158) => DataPath_RF_bus_reg_dataout_1158_port,
                           regs(1157) => DataPath_RF_bus_reg_dataout_1157_port,
                           regs(1156) => DataPath_RF_bus_reg_dataout_1156_port,
                           regs(1155) => DataPath_RF_bus_reg_dataout_1155_port,
                           regs(1154) => DataPath_RF_bus_reg_dataout_1154_port,
                           regs(1153) => DataPath_RF_bus_reg_dataout_1153_port,
                           regs(1152) => DataPath_RF_bus_reg_dataout_1152_port,
                           regs(1151) => DataPath_RF_bus_reg_dataout_1151_port,
                           regs(1150) => DataPath_RF_bus_reg_dataout_1150_port,
                           regs(1149) => DataPath_RF_bus_reg_dataout_1149_port,
                           regs(1148) => DataPath_RF_bus_reg_dataout_1148_port,
                           regs(1147) => DataPath_RF_bus_reg_dataout_1147_port,
                           regs(1146) => DataPath_RF_bus_reg_dataout_1146_port,
                           regs(1145) => DataPath_RF_bus_reg_dataout_1145_port,
                           regs(1144) => DataPath_RF_bus_reg_dataout_1144_port,
                           regs(1143) => DataPath_RF_bus_reg_dataout_1143_port,
                           regs(1142) => DataPath_RF_bus_reg_dataout_1142_port,
                           regs(1141) => DataPath_RF_bus_reg_dataout_1141_port,
                           regs(1140) => DataPath_RF_bus_reg_dataout_1140_port,
                           regs(1139) => DataPath_RF_bus_reg_dataout_1139_port,
                           regs(1138) => DataPath_RF_bus_reg_dataout_1138_port,
                           regs(1137) => DataPath_RF_bus_reg_dataout_1137_port,
                           regs(1136) => DataPath_RF_bus_reg_dataout_1136_port,
                           regs(1135) => DataPath_RF_bus_reg_dataout_1135_port,
                           regs(1134) => DataPath_RF_bus_reg_dataout_1134_port,
                           regs(1133) => DataPath_RF_bus_reg_dataout_1133_port,
                           regs(1132) => DataPath_RF_bus_reg_dataout_1132_port,
                           regs(1131) => DataPath_RF_bus_reg_dataout_1131_port,
                           regs(1130) => DataPath_RF_bus_reg_dataout_1130_port,
                           regs(1129) => DataPath_RF_bus_reg_dataout_1129_port,
                           regs(1128) => DataPath_RF_bus_reg_dataout_1128_port,
                           regs(1127) => DataPath_RF_bus_reg_dataout_1127_port,
                           regs(1126) => DataPath_RF_bus_reg_dataout_1126_port,
                           regs(1125) => DataPath_RF_bus_reg_dataout_1125_port,
                           regs(1124) => DataPath_RF_bus_reg_dataout_1124_port,
                           regs(1123) => DataPath_RF_bus_reg_dataout_1123_port,
                           regs(1122) => DataPath_RF_bus_reg_dataout_1122_port,
                           regs(1121) => DataPath_RF_bus_reg_dataout_1121_port,
                           regs(1120) => DataPath_RF_bus_reg_dataout_1120_port,
                           regs(1119) => DataPath_RF_bus_reg_dataout_1119_port,
                           regs(1118) => DataPath_RF_bus_reg_dataout_1118_port,
                           regs(1117) => DataPath_RF_bus_reg_dataout_1117_port,
                           regs(1116) => DataPath_RF_bus_reg_dataout_1116_port,
                           regs(1115) => DataPath_RF_bus_reg_dataout_1115_port,
                           regs(1114) => DataPath_RF_bus_reg_dataout_1114_port,
                           regs(1113) => DataPath_RF_bus_reg_dataout_1113_port,
                           regs(1112) => DataPath_RF_bus_reg_dataout_1112_port,
                           regs(1111) => DataPath_RF_bus_reg_dataout_1111_port,
                           regs(1110) => DataPath_RF_bus_reg_dataout_1110_port,
                           regs(1109) => DataPath_RF_bus_reg_dataout_1109_port,
                           regs(1108) => DataPath_RF_bus_reg_dataout_1108_port,
                           regs(1107) => DataPath_RF_bus_reg_dataout_1107_port,
                           regs(1106) => DataPath_RF_bus_reg_dataout_1106_port,
                           regs(1105) => DataPath_RF_bus_reg_dataout_1105_port,
                           regs(1104) => DataPath_RF_bus_reg_dataout_1104_port,
                           regs(1103) => DataPath_RF_bus_reg_dataout_1103_port,
                           regs(1102) => DataPath_RF_bus_reg_dataout_1102_port,
                           regs(1101) => DataPath_RF_bus_reg_dataout_1101_port,
                           regs(1100) => DataPath_RF_bus_reg_dataout_1100_port,
                           regs(1099) => DataPath_RF_bus_reg_dataout_1099_port,
                           regs(1098) => DataPath_RF_bus_reg_dataout_1098_port,
                           regs(1097) => DataPath_RF_bus_reg_dataout_1097_port,
                           regs(1096) => DataPath_RF_bus_reg_dataout_1096_port,
                           regs(1095) => DataPath_RF_bus_reg_dataout_1095_port,
                           regs(1094) => DataPath_RF_bus_reg_dataout_1094_port,
                           regs(1093) => DataPath_RF_bus_reg_dataout_1093_port,
                           regs(1092) => DataPath_RF_bus_reg_dataout_1092_port,
                           regs(1091) => DataPath_RF_bus_reg_dataout_1091_port,
                           regs(1090) => DataPath_RF_bus_reg_dataout_1090_port,
                           regs(1089) => DataPath_RF_bus_reg_dataout_1089_port,
                           regs(1088) => DataPath_RF_bus_reg_dataout_1088_port,
                           regs(1087) => DataPath_RF_bus_reg_dataout_1087_port,
                           regs(1086) => DataPath_RF_bus_reg_dataout_1086_port,
                           regs(1085) => DataPath_RF_bus_reg_dataout_1085_port,
                           regs(1084) => DataPath_RF_bus_reg_dataout_1084_port,
                           regs(1083) => DataPath_RF_bus_reg_dataout_1083_port,
                           regs(1082) => DataPath_RF_bus_reg_dataout_1082_port,
                           regs(1081) => DataPath_RF_bus_reg_dataout_1081_port,
                           regs(1080) => DataPath_RF_bus_reg_dataout_1080_port,
                           regs(1079) => DataPath_RF_bus_reg_dataout_1079_port,
                           regs(1078) => DataPath_RF_bus_reg_dataout_1078_port,
                           regs(1077) => DataPath_RF_bus_reg_dataout_1077_port,
                           regs(1076) => DataPath_RF_bus_reg_dataout_1076_port,
                           regs(1075) => DataPath_RF_bus_reg_dataout_1075_port,
                           regs(1074) => DataPath_RF_bus_reg_dataout_1074_port,
                           regs(1073) => DataPath_RF_bus_reg_dataout_1073_port,
                           regs(1072) => DataPath_RF_bus_reg_dataout_1072_port,
                           regs(1071) => DataPath_RF_bus_reg_dataout_1071_port,
                           regs(1070) => DataPath_RF_bus_reg_dataout_1070_port,
                           regs(1069) => DataPath_RF_bus_reg_dataout_1069_port,
                           regs(1068) => DataPath_RF_bus_reg_dataout_1068_port,
                           regs(1067) => DataPath_RF_bus_reg_dataout_1067_port,
                           regs(1066) => DataPath_RF_bus_reg_dataout_1066_port,
                           regs(1065) => DataPath_RF_bus_reg_dataout_1065_port,
                           regs(1064) => DataPath_RF_bus_reg_dataout_1064_port,
                           regs(1063) => DataPath_RF_bus_reg_dataout_1063_port,
                           regs(1062) => DataPath_RF_bus_reg_dataout_1062_port,
                           regs(1061) => DataPath_RF_bus_reg_dataout_1061_port,
                           regs(1060) => DataPath_RF_bus_reg_dataout_1060_port,
                           regs(1059) => DataPath_RF_bus_reg_dataout_1059_port,
                           regs(1058) => DataPath_RF_bus_reg_dataout_1058_port,
                           regs(1057) => DataPath_RF_bus_reg_dataout_1057_port,
                           regs(1056) => DataPath_RF_bus_reg_dataout_1056_port,
                           regs(1055) => DataPath_RF_bus_reg_dataout_1055_port,
                           regs(1054) => DataPath_RF_bus_reg_dataout_1054_port,
                           regs(1053) => DataPath_RF_bus_reg_dataout_1053_port,
                           regs(1052) => DataPath_RF_bus_reg_dataout_1052_port,
                           regs(1051) => DataPath_RF_bus_reg_dataout_1051_port,
                           regs(1050) => DataPath_RF_bus_reg_dataout_1050_port,
                           regs(1049) => DataPath_RF_bus_reg_dataout_1049_port,
                           regs(1048) => DataPath_RF_bus_reg_dataout_1048_port,
                           regs(1047) => DataPath_RF_bus_reg_dataout_1047_port,
                           regs(1046) => DataPath_RF_bus_reg_dataout_1046_port,
                           regs(1045) => DataPath_RF_bus_reg_dataout_1045_port,
                           regs(1044) => DataPath_RF_bus_reg_dataout_1044_port,
                           regs(1043) => DataPath_RF_bus_reg_dataout_1043_port,
                           regs(1042) => DataPath_RF_bus_reg_dataout_1042_port,
                           regs(1041) => DataPath_RF_bus_reg_dataout_1041_port,
                           regs(1040) => DataPath_RF_bus_reg_dataout_1040_port,
                           regs(1039) => DataPath_RF_bus_reg_dataout_1039_port,
                           regs(1038) => DataPath_RF_bus_reg_dataout_1038_port,
                           regs(1037) => DataPath_RF_bus_reg_dataout_1037_port,
                           regs(1036) => DataPath_RF_bus_reg_dataout_1036_port,
                           regs(1035) => DataPath_RF_bus_reg_dataout_1035_port,
                           regs(1034) => DataPath_RF_bus_reg_dataout_1034_port,
                           regs(1033) => DataPath_RF_bus_reg_dataout_1033_port,
                           regs(1032) => DataPath_RF_bus_reg_dataout_1032_port,
                           regs(1031) => DataPath_RF_bus_reg_dataout_1031_port,
                           regs(1030) => DataPath_RF_bus_reg_dataout_1030_port,
                           regs(1029) => DataPath_RF_bus_reg_dataout_1029_port,
                           regs(1028) => DataPath_RF_bus_reg_dataout_1028_port,
                           regs(1027) => DataPath_RF_bus_reg_dataout_1027_port,
                           regs(1026) => DataPath_RF_bus_reg_dataout_1026_port,
                           regs(1025) => DataPath_RF_bus_reg_dataout_1025_port,
                           regs(1024) => DataPath_RF_bus_reg_dataout_1024_port,
                           regs(1023) => DataPath_RF_bus_reg_dataout_1023_port,
                           regs(1022) => DataPath_RF_bus_reg_dataout_1022_port,
                           regs(1021) => DataPath_RF_bus_reg_dataout_1021_port,
                           regs(1020) => DataPath_RF_bus_reg_dataout_1020_port,
                           regs(1019) => DataPath_RF_bus_reg_dataout_1019_port,
                           regs(1018) => DataPath_RF_bus_reg_dataout_1018_port,
                           regs(1017) => DataPath_RF_bus_reg_dataout_1017_port,
                           regs(1016) => DataPath_RF_bus_reg_dataout_1016_port,
                           regs(1015) => DataPath_RF_bus_reg_dataout_1015_port,
                           regs(1014) => DataPath_RF_bus_reg_dataout_1014_port,
                           regs(1013) => DataPath_RF_bus_reg_dataout_1013_port,
                           regs(1012) => DataPath_RF_bus_reg_dataout_1012_port,
                           regs(1011) => DataPath_RF_bus_reg_dataout_1011_port,
                           regs(1010) => DataPath_RF_bus_reg_dataout_1010_port,
                           regs(1009) => DataPath_RF_bus_reg_dataout_1009_port,
                           regs(1008) => DataPath_RF_bus_reg_dataout_1008_port,
                           regs(1007) => DataPath_RF_bus_reg_dataout_1007_port,
                           regs(1006) => DataPath_RF_bus_reg_dataout_1006_port,
                           regs(1005) => DataPath_RF_bus_reg_dataout_1005_port,
                           regs(1004) => DataPath_RF_bus_reg_dataout_1004_port,
                           regs(1003) => DataPath_RF_bus_reg_dataout_1003_port,
                           regs(1002) => DataPath_RF_bus_reg_dataout_1002_port,
                           regs(1001) => DataPath_RF_bus_reg_dataout_1001_port,
                           regs(1000) => DataPath_RF_bus_reg_dataout_1000_port,
                           regs(999) => DataPath_RF_bus_reg_dataout_999_port, 
                           regs(998) => DataPath_RF_bus_reg_dataout_998_port, 
                           regs(997) => DataPath_RF_bus_reg_dataout_997_port, 
                           regs(996) => DataPath_RF_bus_reg_dataout_996_port, 
                           regs(995) => DataPath_RF_bus_reg_dataout_995_port, 
                           regs(994) => DataPath_RF_bus_reg_dataout_994_port, 
                           regs(993) => DataPath_RF_bus_reg_dataout_993_port, 
                           regs(992) => DataPath_RF_bus_reg_dataout_992_port, 
                           regs(991) => DataPath_RF_bus_reg_dataout_991_port, 
                           regs(990) => DataPath_RF_bus_reg_dataout_990_port, 
                           regs(989) => DataPath_RF_bus_reg_dataout_989_port, 
                           regs(988) => DataPath_RF_bus_reg_dataout_988_port, 
                           regs(987) => DataPath_RF_bus_reg_dataout_987_port, 
                           regs(986) => DataPath_RF_bus_reg_dataout_986_port, 
                           regs(985) => DataPath_RF_bus_reg_dataout_985_port, 
                           regs(984) => DataPath_RF_bus_reg_dataout_984_port, 
                           regs(983) => DataPath_RF_bus_reg_dataout_983_port, 
                           regs(982) => DataPath_RF_bus_reg_dataout_982_port, 
                           regs(981) => DataPath_RF_bus_reg_dataout_981_port, 
                           regs(980) => DataPath_RF_bus_reg_dataout_980_port, 
                           regs(979) => DataPath_RF_bus_reg_dataout_979_port, 
                           regs(978) => DataPath_RF_bus_reg_dataout_978_port, 
                           regs(977) => DataPath_RF_bus_reg_dataout_977_port, 
                           regs(976) => DataPath_RF_bus_reg_dataout_976_port, 
                           regs(975) => DataPath_RF_bus_reg_dataout_975_port, 
                           regs(974) => DataPath_RF_bus_reg_dataout_974_port, 
                           regs(973) => DataPath_RF_bus_reg_dataout_973_port, 
                           regs(972) => DataPath_RF_bus_reg_dataout_972_port, 
                           regs(971) => DataPath_RF_bus_reg_dataout_971_port, 
                           regs(970) => DataPath_RF_bus_reg_dataout_970_port, 
                           regs(969) => DataPath_RF_bus_reg_dataout_969_port, 
                           regs(968) => DataPath_RF_bus_reg_dataout_968_port, 
                           regs(967) => DataPath_RF_bus_reg_dataout_967_port, 
                           regs(966) => DataPath_RF_bus_reg_dataout_966_port, 
                           regs(965) => DataPath_RF_bus_reg_dataout_965_port, 
                           regs(964) => DataPath_RF_bus_reg_dataout_964_port, 
                           regs(963) => DataPath_RF_bus_reg_dataout_963_port, 
                           regs(962) => DataPath_RF_bus_reg_dataout_962_port, 
                           regs(961) => DataPath_RF_bus_reg_dataout_961_port, 
                           regs(960) => DataPath_RF_bus_reg_dataout_960_port, 
                           regs(959) => DataPath_RF_bus_reg_dataout_959_port, 
                           regs(958) => DataPath_RF_bus_reg_dataout_958_port, 
                           regs(957) => DataPath_RF_bus_reg_dataout_957_port, 
                           regs(956) => DataPath_RF_bus_reg_dataout_956_port, 
                           regs(955) => DataPath_RF_bus_reg_dataout_955_port, 
                           regs(954) => DataPath_RF_bus_reg_dataout_954_port, 
                           regs(953) => DataPath_RF_bus_reg_dataout_953_port, 
                           regs(952) => DataPath_RF_bus_reg_dataout_952_port, 
                           regs(951) => DataPath_RF_bus_reg_dataout_951_port, 
                           regs(950) => DataPath_RF_bus_reg_dataout_950_port, 
                           regs(949) => DataPath_RF_bus_reg_dataout_949_port, 
                           regs(948) => DataPath_RF_bus_reg_dataout_948_port, 
                           regs(947) => DataPath_RF_bus_reg_dataout_947_port, 
                           regs(946) => DataPath_RF_bus_reg_dataout_946_port, 
                           regs(945) => DataPath_RF_bus_reg_dataout_945_port, 
                           regs(944) => DataPath_RF_bus_reg_dataout_944_port, 
                           regs(943) => DataPath_RF_bus_reg_dataout_943_port, 
                           regs(942) => DataPath_RF_bus_reg_dataout_942_port, 
                           regs(941) => DataPath_RF_bus_reg_dataout_941_port, 
                           regs(940) => DataPath_RF_bus_reg_dataout_940_port, 
                           regs(939) => DataPath_RF_bus_reg_dataout_939_port, 
                           regs(938) => DataPath_RF_bus_reg_dataout_938_port, 
                           regs(937) => DataPath_RF_bus_reg_dataout_937_port, 
                           regs(936) => DataPath_RF_bus_reg_dataout_936_port, 
                           regs(935) => DataPath_RF_bus_reg_dataout_935_port, 
                           regs(934) => DataPath_RF_bus_reg_dataout_934_port, 
                           regs(933) => DataPath_RF_bus_reg_dataout_933_port, 
                           regs(932) => DataPath_RF_bus_reg_dataout_932_port, 
                           regs(931) => DataPath_RF_bus_reg_dataout_931_port, 
                           regs(930) => DataPath_RF_bus_reg_dataout_930_port, 
                           regs(929) => DataPath_RF_bus_reg_dataout_929_port, 
                           regs(928) => DataPath_RF_bus_reg_dataout_928_port, 
                           regs(927) => DataPath_RF_bus_reg_dataout_927_port, 
                           regs(926) => DataPath_RF_bus_reg_dataout_926_port, 
                           regs(925) => DataPath_RF_bus_reg_dataout_925_port, 
                           regs(924) => DataPath_RF_bus_reg_dataout_924_port, 
                           regs(923) => DataPath_RF_bus_reg_dataout_923_port, 
                           regs(922) => DataPath_RF_bus_reg_dataout_922_port, 
                           regs(921) => DataPath_RF_bus_reg_dataout_921_port, 
                           regs(920) => DataPath_RF_bus_reg_dataout_920_port, 
                           regs(919) => DataPath_RF_bus_reg_dataout_919_port, 
                           regs(918) => DataPath_RF_bus_reg_dataout_918_port, 
                           regs(917) => DataPath_RF_bus_reg_dataout_917_port, 
                           regs(916) => DataPath_RF_bus_reg_dataout_916_port, 
                           regs(915) => DataPath_RF_bus_reg_dataout_915_port, 
                           regs(914) => DataPath_RF_bus_reg_dataout_914_port, 
                           regs(913) => DataPath_RF_bus_reg_dataout_913_port, 
                           regs(912) => DataPath_RF_bus_reg_dataout_912_port, 
                           regs(911) => DataPath_RF_bus_reg_dataout_911_port, 
                           regs(910) => DataPath_RF_bus_reg_dataout_910_port, 
                           regs(909) => DataPath_RF_bus_reg_dataout_909_port, 
                           regs(908) => DataPath_RF_bus_reg_dataout_908_port, 
                           regs(907) => DataPath_RF_bus_reg_dataout_907_port, 
                           regs(906) => DataPath_RF_bus_reg_dataout_906_port, 
                           regs(905) => DataPath_RF_bus_reg_dataout_905_port, 
                           regs(904) => DataPath_RF_bus_reg_dataout_904_port, 
                           regs(903) => DataPath_RF_bus_reg_dataout_903_port, 
                           regs(902) => DataPath_RF_bus_reg_dataout_902_port, 
                           regs(901) => DataPath_RF_bus_reg_dataout_901_port, 
                           regs(900) => DataPath_RF_bus_reg_dataout_900_port, 
                           regs(899) => DataPath_RF_bus_reg_dataout_899_port, 
                           regs(898) => DataPath_RF_bus_reg_dataout_898_port, 
                           regs(897) => DataPath_RF_bus_reg_dataout_897_port, 
                           regs(896) => DataPath_RF_bus_reg_dataout_896_port, 
                           regs(895) => DataPath_RF_bus_reg_dataout_895_port, 
                           regs(894) => DataPath_RF_bus_reg_dataout_894_port, 
                           regs(893) => DataPath_RF_bus_reg_dataout_893_port, 
                           regs(892) => DataPath_RF_bus_reg_dataout_892_port, 
                           regs(891) => DataPath_RF_bus_reg_dataout_891_port, 
                           regs(890) => DataPath_RF_bus_reg_dataout_890_port, 
                           regs(889) => DataPath_RF_bus_reg_dataout_889_port, 
                           regs(888) => DataPath_RF_bus_reg_dataout_888_port, 
                           regs(887) => DataPath_RF_bus_reg_dataout_887_port, 
                           regs(886) => DataPath_RF_bus_reg_dataout_886_port, 
                           regs(885) => DataPath_RF_bus_reg_dataout_885_port, 
                           regs(884) => DataPath_RF_bus_reg_dataout_884_port, 
                           regs(883) => DataPath_RF_bus_reg_dataout_883_port, 
                           regs(882) => DataPath_RF_bus_reg_dataout_882_port, 
                           regs(881) => DataPath_RF_bus_reg_dataout_881_port, 
                           regs(880) => DataPath_RF_bus_reg_dataout_880_port, 
                           regs(879) => DataPath_RF_bus_reg_dataout_879_port, 
                           regs(878) => DataPath_RF_bus_reg_dataout_878_port, 
                           regs(877) => DataPath_RF_bus_reg_dataout_877_port, 
                           regs(876) => DataPath_RF_bus_reg_dataout_876_port, 
                           regs(875) => DataPath_RF_bus_reg_dataout_875_port, 
                           regs(874) => DataPath_RF_bus_reg_dataout_874_port, 
                           regs(873) => DataPath_RF_bus_reg_dataout_873_port, 
                           regs(872) => DataPath_RF_bus_reg_dataout_872_port, 
                           regs(871) => DataPath_RF_bus_reg_dataout_871_port, 
                           regs(870) => DataPath_RF_bus_reg_dataout_870_port, 
                           regs(869) => DataPath_RF_bus_reg_dataout_869_port, 
                           regs(868) => DataPath_RF_bus_reg_dataout_868_port, 
                           regs(867) => DataPath_RF_bus_reg_dataout_867_port, 
                           regs(866) => DataPath_RF_bus_reg_dataout_866_port, 
                           regs(865) => DataPath_RF_bus_reg_dataout_865_port, 
                           regs(864) => DataPath_RF_bus_reg_dataout_864_port, 
                           regs(863) => DataPath_RF_bus_reg_dataout_863_port, 
                           regs(862) => DataPath_RF_bus_reg_dataout_862_port, 
                           regs(861) => DataPath_RF_bus_reg_dataout_861_port, 
                           regs(860) => DataPath_RF_bus_reg_dataout_860_port, 
                           regs(859) => DataPath_RF_bus_reg_dataout_859_port, 
                           regs(858) => DataPath_RF_bus_reg_dataout_858_port, 
                           regs(857) => DataPath_RF_bus_reg_dataout_857_port, 
                           regs(856) => DataPath_RF_bus_reg_dataout_856_port, 
                           regs(855) => DataPath_RF_bus_reg_dataout_855_port, 
                           regs(854) => DataPath_RF_bus_reg_dataout_854_port, 
                           regs(853) => DataPath_RF_bus_reg_dataout_853_port, 
                           regs(852) => DataPath_RF_bus_reg_dataout_852_port, 
                           regs(851) => DataPath_RF_bus_reg_dataout_851_port, 
                           regs(850) => DataPath_RF_bus_reg_dataout_850_port, 
                           regs(849) => DataPath_RF_bus_reg_dataout_849_port, 
                           regs(848) => DataPath_RF_bus_reg_dataout_848_port, 
                           regs(847) => DataPath_RF_bus_reg_dataout_847_port, 
                           regs(846) => DataPath_RF_bus_reg_dataout_846_port, 
                           regs(845) => DataPath_RF_bus_reg_dataout_845_port, 
                           regs(844) => DataPath_RF_bus_reg_dataout_844_port, 
                           regs(843) => DataPath_RF_bus_reg_dataout_843_port, 
                           regs(842) => DataPath_RF_bus_reg_dataout_842_port, 
                           regs(841) => DataPath_RF_bus_reg_dataout_841_port, 
                           regs(840) => DataPath_RF_bus_reg_dataout_840_port, 
                           regs(839) => DataPath_RF_bus_reg_dataout_839_port, 
                           regs(838) => DataPath_RF_bus_reg_dataout_838_port, 
                           regs(837) => DataPath_RF_bus_reg_dataout_837_port, 
                           regs(836) => DataPath_RF_bus_reg_dataout_836_port, 
                           regs(835) => DataPath_RF_bus_reg_dataout_835_port, 
                           regs(834) => DataPath_RF_bus_reg_dataout_834_port, 
                           regs(833) => DataPath_RF_bus_reg_dataout_833_port, 
                           regs(832) => DataPath_RF_bus_reg_dataout_832_port, 
                           regs(831) => DataPath_RF_bus_reg_dataout_831_port, 
                           regs(830) => DataPath_RF_bus_reg_dataout_830_port, 
                           regs(829) => DataPath_RF_bus_reg_dataout_829_port, 
                           regs(828) => DataPath_RF_bus_reg_dataout_828_port, 
                           regs(827) => DataPath_RF_bus_reg_dataout_827_port, 
                           regs(826) => DataPath_RF_bus_reg_dataout_826_port, 
                           regs(825) => DataPath_RF_bus_reg_dataout_825_port, 
                           regs(824) => DataPath_RF_bus_reg_dataout_824_port, 
                           regs(823) => DataPath_RF_bus_reg_dataout_823_port, 
                           regs(822) => DataPath_RF_bus_reg_dataout_822_port, 
                           regs(821) => DataPath_RF_bus_reg_dataout_821_port, 
                           regs(820) => DataPath_RF_bus_reg_dataout_820_port, 
                           regs(819) => DataPath_RF_bus_reg_dataout_819_port, 
                           regs(818) => DataPath_RF_bus_reg_dataout_818_port, 
                           regs(817) => DataPath_RF_bus_reg_dataout_817_port, 
                           regs(816) => DataPath_RF_bus_reg_dataout_816_port, 
                           regs(815) => DataPath_RF_bus_reg_dataout_815_port, 
                           regs(814) => DataPath_RF_bus_reg_dataout_814_port, 
                           regs(813) => DataPath_RF_bus_reg_dataout_813_port, 
                           regs(812) => DataPath_RF_bus_reg_dataout_812_port, 
                           regs(811) => DataPath_RF_bus_reg_dataout_811_port, 
                           regs(810) => DataPath_RF_bus_reg_dataout_810_port, 
                           regs(809) => DataPath_RF_bus_reg_dataout_809_port, 
                           regs(808) => DataPath_RF_bus_reg_dataout_808_port, 
                           regs(807) => DataPath_RF_bus_reg_dataout_807_port, 
                           regs(806) => DataPath_RF_bus_reg_dataout_806_port, 
                           regs(805) => DataPath_RF_bus_reg_dataout_805_port, 
                           regs(804) => DataPath_RF_bus_reg_dataout_804_port, 
                           regs(803) => DataPath_RF_bus_reg_dataout_803_port, 
                           regs(802) => DataPath_RF_bus_reg_dataout_802_port, 
                           regs(801) => DataPath_RF_bus_reg_dataout_801_port, 
                           regs(800) => DataPath_RF_bus_reg_dataout_800_port, 
                           regs(799) => DataPath_RF_bus_reg_dataout_799_port, 
                           regs(798) => DataPath_RF_bus_reg_dataout_798_port, 
                           regs(797) => DataPath_RF_bus_reg_dataout_797_port, 
                           regs(796) => DataPath_RF_bus_reg_dataout_796_port, 
                           regs(795) => DataPath_RF_bus_reg_dataout_795_port, 
                           regs(794) => DataPath_RF_bus_reg_dataout_794_port, 
                           regs(793) => DataPath_RF_bus_reg_dataout_793_port, 
                           regs(792) => DataPath_RF_bus_reg_dataout_792_port, 
                           regs(791) => DataPath_RF_bus_reg_dataout_791_port, 
                           regs(790) => DataPath_RF_bus_reg_dataout_790_port, 
                           regs(789) => DataPath_RF_bus_reg_dataout_789_port, 
                           regs(788) => DataPath_RF_bus_reg_dataout_788_port, 
                           regs(787) => DataPath_RF_bus_reg_dataout_787_port, 
                           regs(786) => DataPath_RF_bus_reg_dataout_786_port, 
                           regs(785) => DataPath_RF_bus_reg_dataout_785_port, 
                           regs(784) => DataPath_RF_bus_reg_dataout_784_port, 
                           regs(783) => DataPath_RF_bus_reg_dataout_783_port, 
                           regs(782) => DataPath_RF_bus_reg_dataout_782_port, 
                           regs(781) => DataPath_RF_bus_reg_dataout_781_port, 
                           regs(780) => DataPath_RF_bus_reg_dataout_780_port, 
                           regs(779) => DataPath_RF_bus_reg_dataout_779_port, 
                           regs(778) => DataPath_RF_bus_reg_dataout_778_port, 
                           regs(777) => DataPath_RF_bus_reg_dataout_777_port, 
                           regs(776) => DataPath_RF_bus_reg_dataout_776_port, 
                           regs(775) => DataPath_RF_bus_reg_dataout_775_port, 
                           regs(774) => DataPath_RF_bus_reg_dataout_774_port, 
                           regs(773) => DataPath_RF_bus_reg_dataout_773_port, 
                           regs(772) => DataPath_RF_bus_reg_dataout_772_port, 
                           regs(771) => DataPath_RF_bus_reg_dataout_771_port, 
                           regs(770) => DataPath_RF_bus_reg_dataout_770_port, 
                           regs(769) => DataPath_RF_bus_reg_dataout_769_port, 
                           regs(768) => DataPath_RF_bus_reg_dataout_768_port, 
                           regs(767) => DataPath_RF_bus_reg_dataout_767_port, 
                           regs(766) => DataPath_RF_bus_reg_dataout_766_port, 
                           regs(765) => DataPath_RF_bus_reg_dataout_765_port, 
                           regs(764) => DataPath_RF_bus_reg_dataout_764_port, 
                           regs(763) => DataPath_RF_bus_reg_dataout_763_port, 
                           regs(762) => DataPath_RF_bus_reg_dataout_762_port, 
                           regs(761) => DataPath_RF_bus_reg_dataout_761_port, 
                           regs(760) => DataPath_RF_bus_reg_dataout_760_port, 
                           regs(759) => DataPath_RF_bus_reg_dataout_759_port, 
                           regs(758) => DataPath_RF_bus_reg_dataout_758_port, 
                           regs(757) => DataPath_RF_bus_reg_dataout_757_port, 
                           regs(756) => DataPath_RF_bus_reg_dataout_756_port, 
                           regs(755) => DataPath_RF_bus_reg_dataout_755_port, 
                           regs(754) => DataPath_RF_bus_reg_dataout_754_port, 
                           regs(753) => DataPath_RF_bus_reg_dataout_753_port, 
                           regs(752) => DataPath_RF_bus_reg_dataout_752_port, 
                           regs(751) => DataPath_RF_bus_reg_dataout_751_port, 
                           regs(750) => DataPath_RF_bus_reg_dataout_750_port, 
                           regs(749) => DataPath_RF_bus_reg_dataout_749_port, 
                           regs(748) => DataPath_RF_bus_reg_dataout_748_port, 
                           regs(747) => DataPath_RF_bus_reg_dataout_747_port, 
                           regs(746) => DataPath_RF_bus_reg_dataout_746_port, 
                           regs(745) => DataPath_RF_bus_reg_dataout_745_port, 
                           regs(744) => DataPath_RF_bus_reg_dataout_744_port, 
                           regs(743) => DataPath_RF_bus_reg_dataout_743_port, 
                           regs(742) => DataPath_RF_bus_reg_dataout_742_port, 
                           regs(741) => DataPath_RF_bus_reg_dataout_741_port, 
                           regs(740) => DataPath_RF_bus_reg_dataout_740_port, 
                           regs(739) => DataPath_RF_bus_reg_dataout_739_port, 
                           regs(738) => DataPath_RF_bus_reg_dataout_738_port, 
                           regs(737) => DataPath_RF_bus_reg_dataout_737_port, 
                           regs(736) => DataPath_RF_bus_reg_dataout_736_port, 
                           regs(735) => DataPath_RF_bus_reg_dataout_735_port, 
                           regs(734) => DataPath_RF_bus_reg_dataout_734_port, 
                           regs(733) => DataPath_RF_bus_reg_dataout_733_port, 
                           regs(732) => DataPath_RF_bus_reg_dataout_732_port, 
                           regs(731) => DataPath_RF_bus_reg_dataout_731_port, 
                           regs(730) => DataPath_RF_bus_reg_dataout_730_port, 
                           regs(729) => DataPath_RF_bus_reg_dataout_729_port, 
                           regs(728) => DataPath_RF_bus_reg_dataout_728_port, 
                           regs(727) => DataPath_RF_bus_reg_dataout_727_port, 
                           regs(726) => DataPath_RF_bus_reg_dataout_726_port, 
                           regs(725) => DataPath_RF_bus_reg_dataout_725_port, 
                           regs(724) => DataPath_RF_bus_reg_dataout_724_port, 
                           regs(723) => DataPath_RF_bus_reg_dataout_723_port, 
                           regs(722) => DataPath_RF_bus_reg_dataout_722_port, 
                           regs(721) => DataPath_RF_bus_reg_dataout_721_port, 
                           regs(720) => DataPath_RF_bus_reg_dataout_720_port, 
                           regs(719) => DataPath_RF_bus_reg_dataout_719_port, 
                           regs(718) => DataPath_RF_bus_reg_dataout_718_port, 
                           regs(717) => DataPath_RF_bus_reg_dataout_717_port, 
                           regs(716) => DataPath_RF_bus_reg_dataout_716_port, 
                           regs(715) => DataPath_RF_bus_reg_dataout_715_port, 
                           regs(714) => DataPath_RF_bus_reg_dataout_714_port, 
                           regs(713) => DataPath_RF_bus_reg_dataout_713_port, 
                           regs(712) => DataPath_RF_bus_reg_dataout_712_port, 
                           regs(711) => DataPath_RF_bus_reg_dataout_711_port, 
                           regs(710) => DataPath_RF_bus_reg_dataout_710_port, 
                           regs(709) => DataPath_RF_bus_reg_dataout_709_port, 
                           regs(708) => DataPath_RF_bus_reg_dataout_708_port, 
                           regs(707) => DataPath_RF_bus_reg_dataout_707_port, 
                           regs(706) => DataPath_RF_bus_reg_dataout_706_port, 
                           regs(705) => DataPath_RF_bus_reg_dataout_705_port, 
                           regs(704) => DataPath_RF_bus_reg_dataout_704_port, 
                           regs(703) => DataPath_RF_bus_reg_dataout_703_port, 
                           regs(702) => DataPath_RF_bus_reg_dataout_702_port, 
                           regs(701) => DataPath_RF_bus_reg_dataout_701_port, 
                           regs(700) => DataPath_RF_bus_reg_dataout_700_port, 
                           regs(699) => DataPath_RF_bus_reg_dataout_699_port, 
                           regs(698) => DataPath_RF_bus_reg_dataout_698_port, 
                           regs(697) => DataPath_RF_bus_reg_dataout_697_port, 
                           regs(696) => DataPath_RF_bus_reg_dataout_696_port, 
                           regs(695) => DataPath_RF_bus_reg_dataout_695_port, 
                           regs(694) => DataPath_RF_bus_reg_dataout_694_port, 
                           regs(693) => DataPath_RF_bus_reg_dataout_693_port, 
                           regs(692) => DataPath_RF_bus_reg_dataout_692_port, 
                           regs(691) => DataPath_RF_bus_reg_dataout_691_port, 
                           regs(690) => DataPath_RF_bus_reg_dataout_690_port, 
                           regs(689) => DataPath_RF_bus_reg_dataout_689_port, 
                           regs(688) => DataPath_RF_bus_reg_dataout_688_port, 
                           regs(687) => DataPath_RF_bus_reg_dataout_687_port, 
                           regs(686) => DataPath_RF_bus_reg_dataout_686_port, 
                           regs(685) => DataPath_RF_bus_reg_dataout_685_port, 
                           regs(684) => DataPath_RF_bus_reg_dataout_684_port, 
                           regs(683) => DataPath_RF_bus_reg_dataout_683_port, 
                           regs(682) => DataPath_RF_bus_reg_dataout_682_port, 
                           regs(681) => DataPath_RF_bus_reg_dataout_681_port, 
                           regs(680) => DataPath_RF_bus_reg_dataout_680_port, 
                           regs(679) => DataPath_RF_bus_reg_dataout_679_port, 
                           regs(678) => DataPath_RF_bus_reg_dataout_678_port, 
                           regs(677) => DataPath_RF_bus_reg_dataout_677_port, 
                           regs(676) => DataPath_RF_bus_reg_dataout_676_port, 
                           regs(675) => DataPath_RF_bus_reg_dataout_675_port, 
                           regs(674) => DataPath_RF_bus_reg_dataout_674_port, 
                           regs(673) => DataPath_RF_bus_reg_dataout_673_port, 
                           regs(672) => DataPath_RF_bus_reg_dataout_672_port, 
                           regs(671) => DataPath_RF_bus_reg_dataout_671_port, 
                           regs(670) => DataPath_RF_bus_reg_dataout_670_port, 
                           regs(669) => DataPath_RF_bus_reg_dataout_669_port, 
                           regs(668) => DataPath_RF_bus_reg_dataout_668_port, 
                           regs(667) => DataPath_RF_bus_reg_dataout_667_port, 
                           regs(666) => DataPath_RF_bus_reg_dataout_666_port, 
                           regs(665) => DataPath_RF_bus_reg_dataout_665_port, 
                           regs(664) => DataPath_RF_bus_reg_dataout_664_port, 
                           regs(663) => DataPath_RF_bus_reg_dataout_663_port, 
                           regs(662) => DataPath_RF_bus_reg_dataout_662_port, 
                           regs(661) => DataPath_RF_bus_reg_dataout_661_port, 
                           regs(660) => DataPath_RF_bus_reg_dataout_660_port, 
                           regs(659) => DataPath_RF_bus_reg_dataout_659_port, 
                           regs(658) => DataPath_RF_bus_reg_dataout_658_port, 
                           regs(657) => DataPath_RF_bus_reg_dataout_657_port, 
                           regs(656) => DataPath_RF_bus_reg_dataout_656_port, 
                           regs(655) => DataPath_RF_bus_reg_dataout_655_port, 
                           regs(654) => DataPath_RF_bus_reg_dataout_654_port, 
                           regs(653) => DataPath_RF_bus_reg_dataout_653_port, 
                           regs(652) => DataPath_RF_bus_reg_dataout_652_port, 
                           regs(651) => DataPath_RF_bus_reg_dataout_651_port, 
                           regs(650) => DataPath_RF_bus_reg_dataout_650_port, 
                           regs(649) => DataPath_RF_bus_reg_dataout_649_port, 
                           regs(648) => DataPath_RF_bus_reg_dataout_648_port, 
                           regs(647) => DataPath_RF_bus_reg_dataout_647_port, 
                           regs(646) => DataPath_RF_bus_reg_dataout_646_port, 
                           regs(645) => DataPath_RF_bus_reg_dataout_645_port, 
                           regs(644) => DataPath_RF_bus_reg_dataout_644_port, 
                           regs(643) => DataPath_RF_bus_reg_dataout_643_port, 
                           regs(642) => DataPath_RF_bus_reg_dataout_642_port, 
                           regs(641) => DataPath_RF_bus_reg_dataout_641_port, 
                           regs(640) => DataPath_RF_bus_reg_dataout_640_port, 
                           regs(639) => DataPath_RF_bus_reg_dataout_639_port, 
                           regs(638) => DataPath_RF_bus_reg_dataout_638_port, 
                           regs(637) => DataPath_RF_bus_reg_dataout_637_port, 
                           regs(636) => DataPath_RF_bus_reg_dataout_636_port, 
                           regs(635) => DataPath_RF_bus_reg_dataout_635_port, 
                           regs(634) => DataPath_RF_bus_reg_dataout_634_port, 
                           regs(633) => DataPath_RF_bus_reg_dataout_633_port, 
                           regs(632) => DataPath_RF_bus_reg_dataout_632_port, 
                           regs(631) => DataPath_RF_bus_reg_dataout_631_port, 
                           regs(630) => DataPath_RF_bus_reg_dataout_630_port, 
                           regs(629) => DataPath_RF_bus_reg_dataout_629_port, 
                           regs(628) => DataPath_RF_bus_reg_dataout_628_port, 
                           regs(627) => DataPath_RF_bus_reg_dataout_627_port, 
                           regs(626) => DataPath_RF_bus_reg_dataout_626_port, 
                           regs(625) => DataPath_RF_bus_reg_dataout_625_port, 
                           regs(624) => DataPath_RF_bus_reg_dataout_624_port, 
                           regs(623) => DataPath_RF_bus_reg_dataout_623_port, 
                           regs(622) => DataPath_RF_bus_reg_dataout_622_port, 
                           regs(621) => DataPath_RF_bus_reg_dataout_621_port, 
                           regs(620) => DataPath_RF_bus_reg_dataout_620_port, 
                           regs(619) => DataPath_RF_bus_reg_dataout_619_port, 
                           regs(618) => DataPath_RF_bus_reg_dataout_618_port, 
                           regs(617) => DataPath_RF_bus_reg_dataout_617_port, 
                           regs(616) => DataPath_RF_bus_reg_dataout_616_port, 
                           regs(615) => DataPath_RF_bus_reg_dataout_615_port, 
                           regs(614) => DataPath_RF_bus_reg_dataout_614_port, 
                           regs(613) => DataPath_RF_bus_reg_dataout_613_port, 
                           regs(612) => DataPath_RF_bus_reg_dataout_612_port, 
                           regs(611) => DataPath_RF_bus_reg_dataout_611_port, 
                           regs(610) => DataPath_RF_bus_reg_dataout_610_port, 
                           regs(609) => DataPath_RF_bus_reg_dataout_609_port, 
                           regs(608) => DataPath_RF_bus_reg_dataout_608_port, 
                           regs(607) => DataPath_RF_bus_reg_dataout_607_port, 
                           regs(606) => DataPath_RF_bus_reg_dataout_606_port, 
                           regs(605) => DataPath_RF_bus_reg_dataout_605_port, 
                           regs(604) => DataPath_RF_bus_reg_dataout_604_port, 
                           regs(603) => DataPath_RF_bus_reg_dataout_603_port, 
                           regs(602) => DataPath_RF_bus_reg_dataout_602_port, 
                           regs(601) => DataPath_RF_bus_reg_dataout_601_port, 
                           regs(600) => DataPath_RF_bus_reg_dataout_600_port, 
                           regs(599) => DataPath_RF_bus_reg_dataout_599_port, 
                           regs(598) => DataPath_RF_bus_reg_dataout_598_port, 
                           regs(597) => DataPath_RF_bus_reg_dataout_597_port, 
                           regs(596) => DataPath_RF_bus_reg_dataout_596_port, 
                           regs(595) => DataPath_RF_bus_reg_dataout_595_port, 
                           regs(594) => DataPath_RF_bus_reg_dataout_594_port, 
                           regs(593) => DataPath_RF_bus_reg_dataout_593_port, 
                           regs(592) => DataPath_RF_bus_reg_dataout_592_port, 
                           regs(591) => DataPath_RF_bus_reg_dataout_591_port, 
                           regs(590) => DataPath_RF_bus_reg_dataout_590_port, 
                           regs(589) => DataPath_RF_bus_reg_dataout_589_port, 
                           regs(588) => DataPath_RF_bus_reg_dataout_588_port, 
                           regs(587) => DataPath_RF_bus_reg_dataout_587_port, 
                           regs(586) => DataPath_RF_bus_reg_dataout_586_port, 
                           regs(585) => DataPath_RF_bus_reg_dataout_585_port, 
                           regs(584) => DataPath_RF_bus_reg_dataout_584_port, 
                           regs(583) => DataPath_RF_bus_reg_dataout_583_port, 
                           regs(582) => DataPath_RF_bus_reg_dataout_582_port, 
                           regs(581) => DataPath_RF_bus_reg_dataout_581_port, 
                           regs(580) => DataPath_RF_bus_reg_dataout_580_port, 
                           regs(579) => DataPath_RF_bus_reg_dataout_579_port, 
                           regs(578) => DataPath_RF_bus_reg_dataout_578_port, 
                           regs(577) => DataPath_RF_bus_reg_dataout_577_port, 
                           regs(576) => DataPath_RF_bus_reg_dataout_576_port, 
                           regs(575) => DataPath_RF_bus_reg_dataout_575_port, 
                           regs(574) => DataPath_RF_bus_reg_dataout_574_port, 
                           regs(573) => DataPath_RF_bus_reg_dataout_573_port, 
                           regs(572) => DataPath_RF_bus_reg_dataout_572_port, 
                           regs(571) => DataPath_RF_bus_reg_dataout_571_port, 
                           regs(570) => DataPath_RF_bus_reg_dataout_570_port, 
                           regs(569) => DataPath_RF_bus_reg_dataout_569_port, 
                           regs(568) => DataPath_RF_bus_reg_dataout_568_port, 
                           regs(567) => DataPath_RF_bus_reg_dataout_567_port, 
                           regs(566) => DataPath_RF_bus_reg_dataout_566_port, 
                           regs(565) => DataPath_RF_bus_reg_dataout_565_port, 
                           regs(564) => DataPath_RF_bus_reg_dataout_564_port, 
                           regs(563) => DataPath_RF_bus_reg_dataout_563_port, 
                           regs(562) => DataPath_RF_bus_reg_dataout_562_port, 
                           regs(561) => DataPath_RF_bus_reg_dataout_561_port, 
                           regs(560) => DataPath_RF_bus_reg_dataout_560_port, 
                           regs(559) => DataPath_RF_bus_reg_dataout_559_port, 
                           regs(558) => DataPath_RF_bus_reg_dataout_558_port, 
                           regs(557) => DataPath_RF_bus_reg_dataout_557_port, 
                           regs(556) => DataPath_RF_bus_reg_dataout_556_port, 
                           regs(555) => DataPath_RF_bus_reg_dataout_555_port, 
                           regs(554) => DataPath_RF_bus_reg_dataout_554_port, 
                           regs(553) => DataPath_RF_bus_reg_dataout_553_port, 
                           regs(552) => DataPath_RF_bus_reg_dataout_552_port, 
                           regs(551) => DataPath_RF_bus_reg_dataout_551_port, 
                           regs(550) => DataPath_RF_bus_reg_dataout_550_port, 
                           regs(549) => DataPath_RF_bus_reg_dataout_549_port, 
                           regs(548) => DataPath_RF_bus_reg_dataout_548_port, 
                           regs(547) => DataPath_RF_bus_reg_dataout_547_port, 
                           regs(546) => DataPath_RF_bus_reg_dataout_546_port, 
                           regs(545) => DataPath_RF_bus_reg_dataout_545_port, 
                           regs(544) => DataPath_RF_bus_reg_dataout_544_port, 
                           regs(543) => DataPath_RF_bus_reg_dataout_543_port, 
                           regs(542) => DataPath_RF_bus_reg_dataout_542_port, 
                           regs(541) => DataPath_RF_bus_reg_dataout_541_port, 
                           regs(540) => DataPath_RF_bus_reg_dataout_540_port, 
                           regs(539) => DataPath_RF_bus_reg_dataout_539_port, 
                           regs(538) => DataPath_RF_bus_reg_dataout_538_port, 
                           regs(537) => DataPath_RF_bus_reg_dataout_537_port, 
                           regs(536) => DataPath_RF_bus_reg_dataout_536_port, 
                           regs(535) => DataPath_RF_bus_reg_dataout_535_port, 
                           regs(534) => DataPath_RF_bus_reg_dataout_534_port, 
                           regs(533) => DataPath_RF_bus_reg_dataout_533_port, 
                           regs(532) => DataPath_RF_bus_reg_dataout_532_port, 
                           regs(531) => DataPath_RF_bus_reg_dataout_531_port, 
                           regs(530) => DataPath_RF_bus_reg_dataout_530_port, 
                           regs(529) => DataPath_RF_bus_reg_dataout_529_port, 
                           regs(528) => DataPath_RF_bus_reg_dataout_528_port, 
                           regs(527) => DataPath_RF_bus_reg_dataout_527_port, 
                           regs(526) => DataPath_RF_bus_reg_dataout_526_port, 
                           regs(525) => DataPath_RF_bus_reg_dataout_525_port, 
                           regs(524) => DataPath_RF_bus_reg_dataout_524_port, 
                           regs(523) => DataPath_RF_bus_reg_dataout_523_port, 
                           regs(522) => DataPath_RF_bus_reg_dataout_522_port, 
                           regs(521) => DataPath_RF_bus_reg_dataout_521_port, 
                           regs(520) => DataPath_RF_bus_reg_dataout_520_port, 
                           regs(519) => DataPath_RF_bus_reg_dataout_519_port, 
                           regs(518) => DataPath_RF_bus_reg_dataout_518_port, 
                           regs(517) => DataPath_RF_bus_reg_dataout_517_port, 
                           regs(516) => DataPath_RF_bus_reg_dataout_516_port, 
                           regs(515) => DataPath_RF_bus_reg_dataout_515_port, 
                           regs(514) => DataPath_RF_bus_reg_dataout_514_port, 
                           regs(513) => DataPath_RF_bus_reg_dataout_513_port, 
                           regs(512) => DataPath_RF_bus_reg_dataout_512_port, 
                           regs(511) => DataPath_RF_bus_reg_dataout_511_port, 
                           regs(510) => DataPath_RF_bus_reg_dataout_510_port, 
                           regs(509) => DataPath_RF_bus_reg_dataout_509_port, 
                           regs(508) => DataPath_RF_bus_reg_dataout_508_port, 
                           regs(507) => DataPath_RF_bus_reg_dataout_507_port, 
                           regs(506) => DataPath_RF_bus_reg_dataout_506_port, 
                           regs(505) => DataPath_RF_bus_reg_dataout_505_port, 
                           regs(504) => DataPath_RF_bus_reg_dataout_504_port, 
                           regs(503) => DataPath_RF_bus_reg_dataout_503_port, 
                           regs(502) => DataPath_RF_bus_reg_dataout_502_port, 
                           regs(501) => DataPath_RF_bus_reg_dataout_501_port, 
                           regs(500) => DataPath_RF_bus_reg_dataout_500_port, 
                           regs(499) => DataPath_RF_bus_reg_dataout_499_port, 
                           regs(498) => DataPath_RF_bus_reg_dataout_498_port, 
                           regs(497) => DataPath_RF_bus_reg_dataout_497_port, 
                           regs(496) => DataPath_RF_bus_reg_dataout_496_port, 
                           regs(495) => DataPath_RF_bus_reg_dataout_495_port, 
                           regs(494) => DataPath_RF_bus_reg_dataout_494_port, 
                           regs(493) => DataPath_RF_bus_reg_dataout_493_port, 
                           regs(492) => DataPath_RF_bus_reg_dataout_492_port, 
                           regs(491) => DataPath_RF_bus_reg_dataout_491_port, 
                           regs(490) => DataPath_RF_bus_reg_dataout_490_port, 
                           regs(489) => DataPath_RF_bus_reg_dataout_489_port, 
                           regs(488) => DataPath_RF_bus_reg_dataout_488_port, 
                           regs(487) => DataPath_RF_bus_reg_dataout_487_port, 
                           regs(486) => DataPath_RF_bus_reg_dataout_486_port, 
                           regs(485) => DataPath_RF_bus_reg_dataout_485_port, 
                           regs(484) => DataPath_RF_bus_reg_dataout_484_port, 
                           regs(483) => DataPath_RF_bus_reg_dataout_483_port, 
                           regs(482) => DataPath_RF_bus_reg_dataout_482_port, 
                           regs(481) => DataPath_RF_bus_reg_dataout_481_port, 
                           regs(480) => DataPath_RF_bus_reg_dataout_480_port, 
                           regs(479) => DataPath_RF_bus_reg_dataout_479_port, 
                           regs(478) => DataPath_RF_bus_reg_dataout_478_port, 
                           regs(477) => DataPath_RF_bus_reg_dataout_477_port, 
                           regs(476) => DataPath_RF_bus_reg_dataout_476_port, 
                           regs(475) => DataPath_RF_bus_reg_dataout_475_port, 
                           regs(474) => DataPath_RF_bus_reg_dataout_474_port, 
                           regs(473) => DataPath_RF_bus_reg_dataout_473_port, 
                           regs(472) => DataPath_RF_bus_reg_dataout_472_port, 
                           regs(471) => DataPath_RF_bus_reg_dataout_471_port, 
                           regs(470) => DataPath_RF_bus_reg_dataout_470_port, 
                           regs(469) => DataPath_RF_bus_reg_dataout_469_port, 
                           regs(468) => DataPath_RF_bus_reg_dataout_468_port, 
                           regs(467) => DataPath_RF_bus_reg_dataout_467_port, 
                           regs(466) => DataPath_RF_bus_reg_dataout_466_port, 
                           regs(465) => DataPath_RF_bus_reg_dataout_465_port, 
                           regs(464) => DataPath_RF_bus_reg_dataout_464_port, 
                           regs(463) => DataPath_RF_bus_reg_dataout_463_port, 
                           regs(462) => DataPath_RF_bus_reg_dataout_462_port, 
                           regs(461) => DataPath_RF_bus_reg_dataout_461_port, 
                           regs(460) => DataPath_RF_bus_reg_dataout_460_port, 
                           regs(459) => DataPath_RF_bus_reg_dataout_459_port, 
                           regs(458) => DataPath_RF_bus_reg_dataout_458_port, 
                           regs(457) => DataPath_RF_bus_reg_dataout_457_port, 
                           regs(456) => DataPath_RF_bus_reg_dataout_456_port, 
                           regs(455) => DataPath_RF_bus_reg_dataout_455_port, 
                           regs(454) => DataPath_RF_bus_reg_dataout_454_port, 
                           regs(453) => DataPath_RF_bus_reg_dataout_453_port, 
                           regs(452) => DataPath_RF_bus_reg_dataout_452_port, 
                           regs(451) => DataPath_RF_bus_reg_dataout_451_port, 
                           regs(450) => DataPath_RF_bus_reg_dataout_450_port, 
                           regs(449) => DataPath_RF_bus_reg_dataout_449_port, 
                           regs(448) => DataPath_RF_bus_reg_dataout_448_port, 
                           regs(447) => DataPath_RF_bus_reg_dataout_447_port, 
                           regs(446) => DataPath_RF_bus_reg_dataout_446_port, 
                           regs(445) => DataPath_RF_bus_reg_dataout_445_port, 
                           regs(444) => DataPath_RF_bus_reg_dataout_444_port, 
                           regs(443) => DataPath_RF_bus_reg_dataout_443_port, 
                           regs(442) => DataPath_RF_bus_reg_dataout_442_port, 
                           regs(441) => DataPath_RF_bus_reg_dataout_441_port, 
                           regs(440) => DataPath_RF_bus_reg_dataout_440_port, 
                           regs(439) => DataPath_RF_bus_reg_dataout_439_port, 
                           regs(438) => DataPath_RF_bus_reg_dataout_438_port, 
                           regs(437) => DataPath_RF_bus_reg_dataout_437_port, 
                           regs(436) => DataPath_RF_bus_reg_dataout_436_port, 
                           regs(435) => DataPath_RF_bus_reg_dataout_435_port, 
                           regs(434) => DataPath_RF_bus_reg_dataout_434_port, 
                           regs(433) => DataPath_RF_bus_reg_dataout_433_port, 
                           regs(432) => DataPath_RF_bus_reg_dataout_432_port, 
                           regs(431) => DataPath_RF_bus_reg_dataout_431_port, 
                           regs(430) => DataPath_RF_bus_reg_dataout_430_port, 
                           regs(429) => DataPath_RF_bus_reg_dataout_429_port, 
                           regs(428) => DataPath_RF_bus_reg_dataout_428_port, 
                           regs(427) => DataPath_RF_bus_reg_dataout_427_port, 
                           regs(426) => DataPath_RF_bus_reg_dataout_426_port, 
                           regs(425) => DataPath_RF_bus_reg_dataout_425_port, 
                           regs(424) => DataPath_RF_bus_reg_dataout_424_port, 
                           regs(423) => DataPath_RF_bus_reg_dataout_423_port, 
                           regs(422) => DataPath_RF_bus_reg_dataout_422_port, 
                           regs(421) => DataPath_RF_bus_reg_dataout_421_port, 
                           regs(420) => DataPath_RF_bus_reg_dataout_420_port, 
                           regs(419) => DataPath_RF_bus_reg_dataout_419_port, 
                           regs(418) => DataPath_RF_bus_reg_dataout_418_port, 
                           regs(417) => DataPath_RF_bus_reg_dataout_417_port, 
                           regs(416) => DataPath_RF_bus_reg_dataout_416_port, 
                           regs(415) => DataPath_RF_bus_reg_dataout_415_port, 
                           regs(414) => DataPath_RF_bus_reg_dataout_414_port, 
                           regs(413) => DataPath_RF_bus_reg_dataout_413_port, 
                           regs(412) => DataPath_RF_bus_reg_dataout_412_port, 
                           regs(411) => DataPath_RF_bus_reg_dataout_411_port, 
                           regs(410) => DataPath_RF_bus_reg_dataout_410_port, 
                           regs(409) => DataPath_RF_bus_reg_dataout_409_port, 
                           regs(408) => DataPath_RF_bus_reg_dataout_408_port, 
                           regs(407) => DataPath_RF_bus_reg_dataout_407_port, 
                           regs(406) => DataPath_RF_bus_reg_dataout_406_port, 
                           regs(405) => DataPath_RF_bus_reg_dataout_405_port, 
                           regs(404) => DataPath_RF_bus_reg_dataout_404_port, 
                           regs(403) => DataPath_RF_bus_reg_dataout_403_port, 
                           regs(402) => DataPath_RF_bus_reg_dataout_402_port, 
                           regs(401) => DataPath_RF_bus_reg_dataout_401_port, 
                           regs(400) => DataPath_RF_bus_reg_dataout_400_port, 
                           regs(399) => DataPath_RF_bus_reg_dataout_399_port, 
                           regs(398) => DataPath_RF_bus_reg_dataout_398_port, 
                           regs(397) => DataPath_RF_bus_reg_dataout_397_port, 
                           regs(396) => DataPath_RF_bus_reg_dataout_396_port, 
                           regs(395) => DataPath_RF_bus_reg_dataout_395_port, 
                           regs(394) => DataPath_RF_bus_reg_dataout_394_port, 
                           regs(393) => DataPath_RF_bus_reg_dataout_393_port, 
                           regs(392) => DataPath_RF_bus_reg_dataout_392_port, 
                           regs(391) => DataPath_RF_bus_reg_dataout_391_port, 
                           regs(390) => DataPath_RF_bus_reg_dataout_390_port, 
                           regs(389) => DataPath_RF_bus_reg_dataout_389_port, 
                           regs(388) => DataPath_RF_bus_reg_dataout_388_port, 
                           regs(387) => DataPath_RF_bus_reg_dataout_387_port, 
                           regs(386) => DataPath_RF_bus_reg_dataout_386_port, 
                           regs(385) => DataPath_RF_bus_reg_dataout_385_port, 
                           regs(384) => DataPath_RF_bus_reg_dataout_384_port, 
                           regs(383) => DataPath_RF_bus_reg_dataout_383_port, 
                           regs(382) => DataPath_RF_bus_reg_dataout_382_port, 
                           regs(381) => DataPath_RF_bus_reg_dataout_381_port, 
                           regs(380) => DataPath_RF_bus_reg_dataout_380_port, 
                           regs(379) => DataPath_RF_bus_reg_dataout_379_port, 
                           regs(378) => DataPath_RF_bus_reg_dataout_378_port, 
                           regs(377) => DataPath_RF_bus_reg_dataout_377_port, 
                           regs(376) => DataPath_RF_bus_reg_dataout_376_port, 
                           regs(375) => DataPath_RF_bus_reg_dataout_375_port, 
                           regs(374) => DataPath_RF_bus_reg_dataout_374_port, 
                           regs(373) => DataPath_RF_bus_reg_dataout_373_port, 
                           regs(372) => DataPath_RF_bus_reg_dataout_372_port, 
                           regs(371) => DataPath_RF_bus_reg_dataout_371_port, 
                           regs(370) => DataPath_RF_bus_reg_dataout_370_port, 
                           regs(369) => DataPath_RF_bus_reg_dataout_369_port, 
                           regs(368) => DataPath_RF_bus_reg_dataout_368_port, 
                           regs(367) => DataPath_RF_bus_reg_dataout_367_port, 
                           regs(366) => DataPath_RF_bus_reg_dataout_366_port, 
                           regs(365) => DataPath_RF_bus_reg_dataout_365_port, 
                           regs(364) => DataPath_RF_bus_reg_dataout_364_port, 
                           regs(363) => DataPath_RF_bus_reg_dataout_363_port, 
                           regs(362) => DataPath_RF_bus_reg_dataout_362_port, 
                           regs(361) => DataPath_RF_bus_reg_dataout_361_port, 
                           regs(360) => DataPath_RF_bus_reg_dataout_360_port, 
                           regs(359) => DataPath_RF_bus_reg_dataout_359_port, 
                           regs(358) => DataPath_RF_bus_reg_dataout_358_port, 
                           regs(357) => DataPath_RF_bus_reg_dataout_357_port, 
                           regs(356) => DataPath_RF_bus_reg_dataout_356_port, 
                           regs(355) => DataPath_RF_bus_reg_dataout_355_port, 
                           regs(354) => DataPath_RF_bus_reg_dataout_354_port, 
                           regs(353) => DataPath_RF_bus_reg_dataout_353_port, 
                           regs(352) => DataPath_RF_bus_reg_dataout_352_port, 
                           regs(351) => DataPath_RF_bus_reg_dataout_351_port, 
                           regs(350) => DataPath_RF_bus_reg_dataout_350_port, 
                           regs(349) => DataPath_RF_bus_reg_dataout_349_port, 
                           regs(348) => DataPath_RF_bus_reg_dataout_348_port, 
                           regs(347) => DataPath_RF_bus_reg_dataout_347_port, 
                           regs(346) => DataPath_RF_bus_reg_dataout_346_port, 
                           regs(345) => DataPath_RF_bus_reg_dataout_345_port, 
                           regs(344) => DataPath_RF_bus_reg_dataout_344_port, 
                           regs(343) => DataPath_RF_bus_reg_dataout_343_port, 
                           regs(342) => DataPath_RF_bus_reg_dataout_342_port, 
                           regs(341) => DataPath_RF_bus_reg_dataout_341_port, 
                           regs(340) => DataPath_RF_bus_reg_dataout_340_port, 
                           regs(339) => DataPath_RF_bus_reg_dataout_339_port, 
                           regs(338) => DataPath_RF_bus_reg_dataout_338_port, 
                           regs(337) => DataPath_RF_bus_reg_dataout_337_port, 
                           regs(336) => DataPath_RF_bus_reg_dataout_336_port, 
                           regs(335) => DataPath_RF_bus_reg_dataout_335_port, 
                           regs(334) => DataPath_RF_bus_reg_dataout_334_port, 
                           regs(333) => DataPath_RF_bus_reg_dataout_333_port, 
                           regs(332) => DataPath_RF_bus_reg_dataout_332_port, 
                           regs(331) => DataPath_RF_bus_reg_dataout_331_port, 
                           regs(330) => DataPath_RF_bus_reg_dataout_330_port, 
                           regs(329) => DataPath_RF_bus_reg_dataout_329_port, 
                           regs(328) => DataPath_RF_bus_reg_dataout_328_port, 
                           regs(327) => DataPath_RF_bus_reg_dataout_327_port, 
                           regs(326) => DataPath_RF_bus_reg_dataout_326_port, 
                           regs(325) => DataPath_RF_bus_reg_dataout_325_port, 
                           regs(324) => DataPath_RF_bus_reg_dataout_324_port, 
                           regs(323) => DataPath_RF_bus_reg_dataout_323_port, 
                           regs(322) => DataPath_RF_bus_reg_dataout_322_port, 
                           regs(321) => DataPath_RF_bus_reg_dataout_321_port, 
                           regs(320) => DataPath_RF_bus_reg_dataout_320_port, 
                           regs(319) => DataPath_RF_bus_reg_dataout_319_port, 
                           regs(318) => DataPath_RF_bus_reg_dataout_318_port, 
                           regs(317) => DataPath_RF_bus_reg_dataout_317_port, 
                           regs(316) => DataPath_RF_bus_reg_dataout_316_port, 
                           regs(315) => DataPath_RF_bus_reg_dataout_315_port, 
                           regs(314) => DataPath_RF_bus_reg_dataout_314_port, 
                           regs(313) => DataPath_RF_bus_reg_dataout_313_port, 
                           regs(312) => DataPath_RF_bus_reg_dataout_312_port, 
                           regs(311) => DataPath_RF_bus_reg_dataout_311_port, 
                           regs(310) => DataPath_RF_bus_reg_dataout_310_port, 
                           regs(309) => DataPath_RF_bus_reg_dataout_309_port, 
                           regs(308) => DataPath_RF_bus_reg_dataout_308_port, 
                           regs(307) => DataPath_RF_bus_reg_dataout_307_port, 
                           regs(306) => DataPath_RF_bus_reg_dataout_306_port, 
                           regs(305) => DataPath_RF_bus_reg_dataout_305_port, 
                           regs(304) => DataPath_RF_bus_reg_dataout_304_port, 
                           regs(303) => DataPath_RF_bus_reg_dataout_303_port, 
                           regs(302) => DataPath_RF_bus_reg_dataout_302_port, 
                           regs(301) => DataPath_RF_bus_reg_dataout_301_port, 
                           regs(300) => DataPath_RF_bus_reg_dataout_300_port, 
                           regs(299) => DataPath_RF_bus_reg_dataout_299_port, 
                           regs(298) => DataPath_RF_bus_reg_dataout_298_port, 
                           regs(297) => DataPath_RF_bus_reg_dataout_297_port, 
                           regs(296) => DataPath_RF_bus_reg_dataout_296_port, 
                           regs(295) => DataPath_RF_bus_reg_dataout_295_port, 
                           regs(294) => DataPath_RF_bus_reg_dataout_294_port, 
                           regs(293) => DataPath_RF_bus_reg_dataout_293_port, 
                           regs(292) => DataPath_RF_bus_reg_dataout_292_port, 
                           regs(291) => DataPath_RF_bus_reg_dataout_291_port, 
                           regs(290) => DataPath_RF_bus_reg_dataout_290_port, 
                           regs(289) => DataPath_RF_bus_reg_dataout_289_port, 
                           regs(288) => DataPath_RF_bus_reg_dataout_288_port, 
                           regs(287) => DataPath_RF_bus_reg_dataout_287_port, 
                           regs(286) => DataPath_RF_bus_reg_dataout_286_port, 
                           regs(285) => DataPath_RF_bus_reg_dataout_285_port, 
                           regs(284) => DataPath_RF_bus_reg_dataout_284_port, 
                           regs(283) => DataPath_RF_bus_reg_dataout_283_port, 
                           regs(282) => DataPath_RF_bus_reg_dataout_282_port, 
                           regs(281) => DataPath_RF_bus_reg_dataout_281_port, 
                           regs(280) => DataPath_RF_bus_reg_dataout_280_port, 
                           regs(279) => DataPath_RF_bus_reg_dataout_279_port, 
                           regs(278) => DataPath_RF_bus_reg_dataout_278_port, 
                           regs(277) => DataPath_RF_bus_reg_dataout_277_port, 
                           regs(276) => DataPath_RF_bus_reg_dataout_276_port, 
                           regs(275) => DataPath_RF_bus_reg_dataout_275_port, 
                           regs(274) => DataPath_RF_bus_reg_dataout_274_port, 
                           regs(273) => DataPath_RF_bus_reg_dataout_273_port, 
                           regs(272) => DataPath_RF_bus_reg_dataout_272_port, 
                           regs(271) => DataPath_RF_bus_reg_dataout_271_port, 
                           regs(270) => DataPath_RF_bus_reg_dataout_270_port, 
                           regs(269) => DataPath_RF_bus_reg_dataout_269_port, 
                           regs(268) => DataPath_RF_bus_reg_dataout_268_port, 
                           regs(267) => DataPath_RF_bus_reg_dataout_267_port, 
                           regs(266) => DataPath_RF_bus_reg_dataout_266_port, 
                           regs(265) => DataPath_RF_bus_reg_dataout_265_port, 
                           regs(264) => DataPath_RF_bus_reg_dataout_264_port, 
                           regs(263) => DataPath_RF_bus_reg_dataout_263_port, 
                           regs(262) => DataPath_RF_bus_reg_dataout_262_port, 
                           regs(261) => DataPath_RF_bus_reg_dataout_261_port, 
                           regs(260) => DataPath_RF_bus_reg_dataout_260_port, 
                           regs(259) => DataPath_RF_bus_reg_dataout_259_port, 
                           regs(258) => DataPath_RF_bus_reg_dataout_258_port, 
                           regs(257) => DataPath_RF_bus_reg_dataout_257_port, 
                           regs(256) => DataPath_RF_bus_reg_dataout_256_port, 
                           regs(255) => DataPath_RF_bus_reg_dataout_255_port, 
                           regs(254) => DataPath_RF_bus_reg_dataout_254_port, 
                           regs(253) => DataPath_RF_bus_reg_dataout_253_port, 
                           regs(252) => DataPath_RF_bus_reg_dataout_252_port, 
                           regs(251) => DataPath_RF_bus_reg_dataout_251_port, 
                           regs(250) => DataPath_RF_bus_reg_dataout_250_port, 
                           regs(249) => DataPath_RF_bus_reg_dataout_249_port, 
                           regs(248) => DataPath_RF_bus_reg_dataout_248_port, 
                           regs(247) => DataPath_RF_bus_reg_dataout_247_port, 
                           regs(246) => DataPath_RF_bus_reg_dataout_246_port, 
                           regs(245) => DataPath_RF_bus_reg_dataout_245_port, 
                           regs(244) => DataPath_RF_bus_reg_dataout_244_port, 
                           regs(243) => DataPath_RF_bus_reg_dataout_243_port, 
                           regs(242) => DataPath_RF_bus_reg_dataout_242_port, 
                           regs(241) => DataPath_RF_bus_reg_dataout_241_port, 
                           regs(240) => DataPath_RF_bus_reg_dataout_240_port, 
                           regs(239) => DataPath_RF_bus_reg_dataout_239_port, 
                           regs(238) => DataPath_RF_bus_reg_dataout_238_port, 
                           regs(237) => DataPath_RF_bus_reg_dataout_237_port, 
                           regs(236) => DataPath_RF_bus_reg_dataout_236_port, 
                           regs(235) => DataPath_RF_bus_reg_dataout_235_port, 
                           regs(234) => DataPath_RF_bus_reg_dataout_234_port, 
                           regs(233) => DataPath_RF_bus_reg_dataout_233_port, 
                           regs(232) => DataPath_RF_bus_reg_dataout_232_port, 
                           regs(231) => DataPath_RF_bus_reg_dataout_231_port, 
                           regs(230) => DataPath_RF_bus_reg_dataout_230_port, 
                           regs(229) => DataPath_RF_bus_reg_dataout_229_port, 
                           regs(228) => DataPath_RF_bus_reg_dataout_228_port, 
                           regs(227) => DataPath_RF_bus_reg_dataout_227_port, 
                           regs(226) => DataPath_RF_bus_reg_dataout_226_port, 
                           regs(225) => DataPath_RF_bus_reg_dataout_225_port, 
                           regs(224) => DataPath_RF_bus_reg_dataout_224_port, 
                           regs(223) => DataPath_RF_bus_reg_dataout_223_port, 
                           regs(222) => DataPath_RF_bus_reg_dataout_222_port, 
                           regs(221) => DataPath_RF_bus_reg_dataout_221_port, 
                           regs(220) => DataPath_RF_bus_reg_dataout_220_port, 
                           regs(219) => DataPath_RF_bus_reg_dataout_219_port, 
                           regs(218) => DataPath_RF_bus_reg_dataout_218_port, 
                           regs(217) => DataPath_RF_bus_reg_dataout_217_port, 
                           regs(216) => DataPath_RF_bus_reg_dataout_216_port, 
                           regs(215) => DataPath_RF_bus_reg_dataout_215_port, 
                           regs(214) => DataPath_RF_bus_reg_dataout_214_port, 
                           regs(213) => DataPath_RF_bus_reg_dataout_213_port, 
                           regs(212) => DataPath_RF_bus_reg_dataout_212_port, 
                           regs(211) => DataPath_RF_bus_reg_dataout_211_port, 
                           regs(210) => DataPath_RF_bus_reg_dataout_210_port, 
                           regs(209) => DataPath_RF_bus_reg_dataout_209_port, 
                           regs(208) => DataPath_RF_bus_reg_dataout_208_port, 
                           regs(207) => DataPath_RF_bus_reg_dataout_207_port, 
                           regs(206) => DataPath_RF_bus_reg_dataout_206_port, 
                           regs(205) => DataPath_RF_bus_reg_dataout_205_port, 
                           regs(204) => DataPath_RF_bus_reg_dataout_204_port, 
                           regs(203) => DataPath_RF_bus_reg_dataout_203_port, 
                           regs(202) => DataPath_RF_bus_reg_dataout_202_port, 
                           regs(201) => DataPath_RF_bus_reg_dataout_201_port, 
                           regs(200) => DataPath_RF_bus_reg_dataout_200_port, 
                           regs(199) => DataPath_RF_bus_reg_dataout_199_port, 
                           regs(198) => DataPath_RF_bus_reg_dataout_198_port, 
                           regs(197) => DataPath_RF_bus_reg_dataout_197_port, 
                           regs(196) => DataPath_RF_bus_reg_dataout_196_port, 
                           regs(195) => DataPath_RF_bus_reg_dataout_195_port, 
                           regs(194) => DataPath_RF_bus_reg_dataout_194_port, 
                           regs(193) => DataPath_RF_bus_reg_dataout_193_port, 
                           regs(192) => DataPath_RF_bus_reg_dataout_192_port, 
                           regs(191) => DataPath_RF_bus_reg_dataout_191_port, 
                           regs(190) => DataPath_RF_bus_reg_dataout_190_port, 
                           regs(189) => DataPath_RF_bus_reg_dataout_189_port, 
                           regs(188) => DataPath_RF_bus_reg_dataout_188_port, 
                           regs(187) => DataPath_RF_bus_reg_dataout_187_port, 
                           regs(186) => DataPath_RF_bus_reg_dataout_186_port, 
                           regs(185) => DataPath_RF_bus_reg_dataout_185_port, 
                           regs(184) => DataPath_RF_bus_reg_dataout_184_port, 
                           regs(183) => DataPath_RF_bus_reg_dataout_183_port, 
                           regs(182) => DataPath_RF_bus_reg_dataout_182_port, 
                           regs(181) => DataPath_RF_bus_reg_dataout_181_port, 
                           regs(180) => DataPath_RF_bus_reg_dataout_180_port, 
                           regs(179) => DataPath_RF_bus_reg_dataout_179_port, 
                           regs(178) => DataPath_RF_bus_reg_dataout_178_port, 
                           regs(177) => DataPath_RF_bus_reg_dataout_177_port, 
                           regs(176) => DataPath_RF_bus_reg_dataout_176_port, 
                           regs(175) => DataPath_RF_bus_reg_dataout_175_port, 
                           regs(174) => DataPath_RF_bus_reg_dataout_174_port, 
                           regs(173) => DataPath_RF_bus_reg_dataout_173_port, 
                           regs(172) => DataPath_RF_bus_reg_dataout_172_port, 
                           regs(171) => DataPath_RF_bus_reg_dataout_171_port, 
                           regs(170) => DataPath_RF_bus_reg_dataout_170_port, 
                           regs(169) => DataPath_RF_bus_reg_dataout_169_port, 
                           regs(168) => DataPath_RF_bus_reg_dataout_168_port, 
                           regs(167) => DataPath_RF_bus_reg_dataout_167_port, 
                           regs(166) => DataPath_RF_bus_reg_dataout_166_port, 
                           regs(165) => DataPath_RF_bus_reg_dataout_165_port, 
                           regs(164) => DataPath_RF_bus_reg_dataout_164_port, 
                           regs(163) => DataPath_RF_bus_reg_dataout_163_port, 
                           regs(162) => DataPath_RF_bus_reg_dataout_162_port, 
                           regs(161) => DataPath_RF_bus_reg_dataout_161_port, 
                           regs(160) => DataPath_RF_bus_reg_dataout_160_port, 
                           regs(159) => DataPath_RF_bus_reg_dataout_159_port, 
                           regs(158) => DataPath_RF_bus_reg_dataout_158_port, 
                           regs(157) => DataPath_RF_bus_reg_dataout_157_port, 
                           regs(156) => DataPath_RF_bus_reg_dataout_156_port, 
                           regs(155) => DataPath_RF_bus_reg_dataout_155_port, 
                           regs(154) => DataPath_RF_bus_reg_dataout_154_port, 
                           regs(153) => DataPath_RF_bus_reg_dataout_153_port, 
                           regs(152) => DataPath_RF_bus_reg_dataout_152_port, 
                           regs(151) => DataPath_RF_bus_reg_dataout_151_port, 
                           regs(150) => DataPath_RF_bus_reg_dataout_150_port, 
                           regs(149) => DataPath_RF_bus_reg_dataout_149_port, 
                           regs(148) => DataPath_RF_bus_reg_dataout_148_port, 
                           regs(147) => DataPath_RF_bus_reg_dataout_147_port, 
                           regs(146) => DataPath_RF_bus_reg_dataout_146_port, 
                           regs(145) => DataPath_RF_bus_reg_dataout_145_port, 
                           regs(144) => DataPath_RF_bus_reg_dataout_144_port, 
                           regs(143) => DataPath_RF_bus_reg_dataout_143_port, 
                           regs(142) => DataPath_RF_bus_reg_dataout_142_port, 
                           regs(141) => DataPath_RF_bus_reg_dataout_141_port, 
                           regs(140) => DataPath_RF_bus_reg_dataout_140_port, 
                           regs(139) => DataPath_RF_bus_reg_dataout_139_port, 
                           regs(138) => DataPath_RF_bus_reg_dataout_138_port, 
                           regs(137) => DataPath_RF_bus_reg_dataout_137_port, 
                           regs(136) => DataPath_RF_bus_reg_dataout_136_port, 
                           regs(135) => DataPath_RF_bus_reg_dataout_135_port, 
                           regs(134) => DataPath_RF_bus_reg_dataout_134_port, 
                           regs(133) => DataPath_RF_bus_reg_dataout_133_port, 
                           regs(132) => DataPath_RF_bus_reg_dataout_132_port, 
                           regs(131) => DataPath_RF_bus_reg_dataout_131_port, 
                           regs(130) => DataPath_RF_bus_reg_dataout_130_port, 
                           regs(129) => DataPath_RF_bus_reg_dataout_129_port, 
                           regs(128) => DataPath_RF_bus_reg_dataout_128_port, 
                           regs(127) => DataPath_RF_bus_reg_dataout_127_port, 
                           regs(126) => DataPath_RF_bus_reg_dataout_126_port, 
                           regs(125) => DataPath_RF_bus_reg_dataout_125_port, 
                           regs(124) => DataPath_RF_bus_reg_dataout_124_port, 
                           regs(123) => DataPath_RF_bus_reg_dataout_123_port, 
                           regs(122) => DataPath_RF_bus_reg_dataout_122_port, 
                           regs(121) => DataPath_RF_bus_reg_dataout_121_port, 
                           regs(120) => DataPath_RF_bus_reg_dataout_120_port, 
                           regs(119) => DataPath_RF_bus_reg_dataout_119_port, 
                           regs(118) => DataPath_RF_bus_reg_dataout_118_port, 
                           regs(117) => DataPath_RF_bus_reg_dataout_117_port, 
                           regs(116) => DataPath_RF_bus_reg_dataout_116_port, 
                           regs(115) => DataPath_RF_bus_reg_dataout_115_port, 
                           regs(114) => DataPath_RF_bus_reg_dataout_114_port, 
                           regs(113) => DataPath_RF_bus_reg_dataout_113_port, 
                           regs(112) => DataPath_RF_bus_reg_dataout_112_port, 
                           regs(111) => DataPath_RF_bus_reg_dataout_111_port, 
                           regs(110) => DataPath_RF_bus_reg_dataout_110_port, 
                           regs(109) => DataPath_RF_bus_reg_dataout_109_port, 
                           regs(108) => DataPath_RF_bus_reg_dataout_108_port, 
                           regs(107) => DataPath_RF_bus_reg_dataout_107_port, 
                           regs(106) => DataPath_RF_bus_reg_dataout_106_port, 
                           regs(105) => DataPath_RF_bus_reg_dataout_105_port, 
                           regs(104) => DataPath_RF_bus_reg_dataout_104_port, 
                           regs(103) => DataPath_RF_bus_reg_dataout_103_port, 
                           regs(102) => DataPath_RF_bus_reg_dataout_102_port, 
                           regs(101) => DataPath_RF_bus_reg_dataout_101_port, 
                           regs(100) => DataPath_RF_bus_reg_dataout_100_port, 
                           regs(99) => DataPath_RF_bus_reg_dataout_99_port, 
                           regs(98) => DataPath_RF_bus_reg_dataout_98_port, 
                           regs(97) => DataPath_RF_bus_reg_dataout_97_port, 
                           regs(96) => DataPath_RF_bus_reg_dataout_96_port, 
                           regs(95) => DataPath_RF_bus_reg_dataout_95_port, 
                           regs(94) => DataPath_RF_bus_reg_dataout_94_port, 
                           regs(93) => DataPath_RF_bus_reg_dataout_93_port, 
                           regs(92) => DataPath_RF_bus_reg_dataout_92_port, 
                           regs(91) => DataPath_RF_bus_reg_dataout_91_port, 
                           regs(90) => DataPath_RF_bus_reg_dataout_90_port, 
                           regs(89) => DataPath_RF_bus_reg_dataout_89_port, 
                           regs(88) => DataPath_RF_bus_reg_dataout_88_port, 
                           regs(87) => DataPath_RF_bus_reg_dataout_87_port, 
                           regs(86) => DataPath_RF_bus_reg_dataout_86_port, 
                           regs(85) => DataPath_RF_bus_reg_dataout_85_port, 
                           regs(84) => DataPath_RF_bus_reg_dataout_84_port, 
                           regs(83) => DataPath_RF_bus_reg_dataout_83_port, 
                           regs(82) => DataPath_RF_bus_reg_dataout_82_port, 
                           regs(81) => DataPath_RF_bus_reg_dataout_81_port, 
                           regs(80) => DataPath_RF_bus_reg_dataout_80_port, 
                           regs(79) => DataPath_RF_bus_reg_dataout_79_port, 
                           regs(78) => DataPath_RF_bus_reg_dataout_78_port, 
                           regs(77) => DataPath_RF_bus_reg_dataout_77_port, 
                           regs(76) => DataPath_RF_bus_reg_dataout_76_port, 
                           regs(75) => DataPath_RF_bus_reg_dataout_75_port, 
                           regs(74) => DataPath_RF_bus_reg_dataout_74_port, 
                           regs(73) => DataPath_RF_bus_reg_dataout_73_port, 
                           regs(72) => DataPath_RF_bus_reg_dataout_72_port, 
                           regs(71) => DataPath_RF_bus_reg_dataout_71_port, 
                           regs(70) => DataPath_RF_bus_reg_dataout_70_port, 
                           regs(69) => DataPath_RF_bus_reg_dataout_69_port, 
                           regs(68) => DataPath_RF_bus_reg_dataout_68_port, 
                           regs(67) => DataPath_RF_bus_reg_dataout_67_port, 
                           regs(66) => DataPath_RF_bus_reg_dataout_66_port, 
                           regs(65) => DataPath_RF_bus_reg_dataout_65_port, 
                           regs(64) => DataPath_RF_bus_reg_dataout_64_port, 
                           regs(63) => DataPath_RF_bus_reg_dataout_63_port, 
                           regs(62) => DataPath_RF_bus_reg_dataout_62_port, 
                           regs(61) => DataPath_RF_bus_reg_dataout_61_port, 
                           regs(60) => DataPath_RF_bus_reg_dataout_60_port, 
                           regs(59) => DataPath_RF_bus_reg_dataout_59_port, 
                           regs(58) => DataPath_RF_bus_reg_dataout_58_port, 
                           regs(57) => DataPath_RF_bus_reg_dataout_57_port, 
                           regs(56) => DataPath_RF_bus_reg_dataout_56_port, 
                           regs(55) => DataPath_RF_bus_reg_dataout_55_port, 
                           regs(54) => DataPath_RF_bus_reg_dataout_54_port, 
                           regs(53) => DataPath_RF_bus_reg_dataout_53_port, 
                           regs(52) => DataPath_RF_bus_reg_dataout_52_port, 
                           regs(51) => DataPath_RF_bus_reg_dataout_51_port, 
                           regs(50) => DataPath_RF_bus_reg_dataout_50_port, 
                           regs(49) => DataPath_RF_bus_reg_dataout_49_port, 
                           regs(48) => DataPath_RF_bus_reg_dataout_48_port, 
                           regs(47) => DataPath_RF_bus_reg_dataout_47_port, 
                           regs(46) => DataPath_RF_bus_reg_dataout_46_port, 
                           regs(45) => DataPath_RF_bus_reg_dataout_45_port, 
                           regs(44) => DataPath_RF_bus_reg_dataout_44_port, 
                           regs(43) => DataPath_RF_bus_reg_dataout_43_port, 
                           regs(42) => DataPath_RF_bus_reg_dataout_42_port, 
                           regs(41) => DataPath_RF_bus_reg_dataout_41_port, 
                           regs(40) => DataPath_RF_bus_reg_dataout_40_port, 
                           regs(39) => DataPath_RF_bus_reg_dataout_39_port, 
                           regs(38) => DataPath_RF_bus_reg_dataout_38_port, 
                           regs(37) => DataPath_RF_bus_reg_dataout_37_port, 
                           regs(36) => DataPath_RF_bus_reg_dataout_36_port, 
                           regs(35) => DataPath_RF_bus_reg_dataout_35_port, 
                           regs(34) => DataPath_RF_bus_reg_dataout_34_port, 
                           regs(33) => DataPath_RF_bus_reg_dataout_33_port, 
                           regs(32) => DataPath_RF_bus_reg_dataout_32_port, 
                           regs(31) => DataPath_RF_bus_reg_dataout_31_port, 
                           regs(30) => DataPath_RF_bus_reg_dataout_30_port, 
                           regs(29) => DataPath_RF_bus_reg_dataout_29_port, 
                           regs(28) => DataPath_RF_bus_reg_dataout_28_port, 
                           regs(27) => DataPath_RF_bus_reg_dataout_27_port, 
                           regs(26) => DataPath_RF_bus_reg_dataout_26_port, 
                           regs(25) => DataPath_RF_bus_reg_dataout_25_port, 
                           regs(24) => DataPath_RF_bus_reg_dataout_24_port, 
                           regs(23) => DataPath_RF_bus_reg_dataout_23_port, 
                           regs(22) => DataPath_RF_bus_reg_dataout_22_port, 
                           regs(21) => DataPath_RF_bus_reg_dataout_21_port, 
                           regs(20) => DataPath_RF_bus_reg_dataout_20_port, 
                           regs(19) => DataPath_RF_bus_reg_dataout_19_port, 
                           regs(18) => DataPath_RF_bus_reg_dataout_18_port, 
                           regs(17) => DataPath_RF_bus_reg_dataout_17_port, 
                           regs(16) => DataPath_RF_bus_reg_dataout_16_port, 
                           regs(15) => DataPath_RF_bus_reg_dataout_15_port, 
                           regs(14) => DataPath_RF_bus_reg_dataout_14_port, 
                           regs(13) => DataPath_RF_bus_reg_dataout_13_port, 
                           regs(12) => DataPath_RF_bus_reg_dataout_12_port, 
                           regs(11) => DataPath_RF_bus_reg_dataout_11_port, 
                           regs(10) => DataPath_RF_bus_reg_dataout_10_port, 
                           regs(9) => DataPath_RF_bus_reg_dataout_9_port, 
                           regs(8) => DataPath_RF_bus_reg_dataout_8_port, 
                           regs(7) => DataPath_RF_bus_reg_dataout_7_port, 
                           regs(6) => DataPath_RF_bus_reg_dataout_6_port, 
                           regs(5) => DataPath_RF_bus_reg_dataout_5_port, 
                           regs(4) => DataPath_RF_bus_reg_dataout_4_port, 
                           regs(3) => DataPath_RF_bus_reg_dataout_3_port, 
                           regs(2) => DataPath_RF_bus_reg_dataout_2_port, 
                           regs(1) => DataPath_RF_bus_reg_dataout_1_port, 
                           regs(0) => DataPath_RF_bus_reg_dataout_0_port, 
                           win(4) => DataPath_RF_c_swin_4_port, win(3) => 
                           DataPath_RF_c_swin_3_port, win(2) => 
                           DataPath_RF_c_swin_2_port, win(1) => 
                           DataPath_RF_c_swin_1_port, win(0) => 
                           DataPath_RF_c_swin_0_port, curr_proc_regs(511) => 
                           DataPath_RF_bus_sel_savedwin_data_511_port, 
                           curr_proc_regs(510) => 
                           DataPath_RF_bus_sel_savedwin_data_510_port, 
                           curr_proc_regs(509) => 
                           DataPath_RF_bus_sel_savedwin_data_509_port, 
                           curr_proc_regs(508) => 
                           DataPath_RF_bus_sel_savedwin_data_508_port, 
                           curr_proc_regs(507) => 
                           DataPath_RF_bus_sel_savedwin_data_507_port, 
                           curr_proc_regs(506) => 
                           DataPath_RF_bus_sel_savedwin_data_506_port, 
                           curr_proc_regs(505) => 
                           DataPath_RF_bus_sel_savedwin_data_505_port, 
                           curr_proc_regs(504) => 
                           DataPath_RF_bus_sel_savedwin_data_504_port, 
                           curr_proc_regs(503) => 
                           DataPath_RF_bus_sel_savedwin_data_503_port, 
                           curr_proc_regs(502) => 
                           DataPath_RF_bus_sel_savedwin_data_502_port, 
                           curr_proc_regs(501) => 
                           DataPath_RF_bus_sel_savedwin_data_501_port, 
                           curr_proc_regs(500) => 
                           DataPath_RF_bus_sel_savedwin_data_500_port, 
                           curr_proc_regs(499) => 
                           DataPath_RF_bus_sel_savedwin_data_499_port, 
                           curr_proc_regs(498) => 
                           DataPath_RF_bus_sel_savedwin_data_498_port, 
                           curr_proc_regs(497) => 
                           DataPath_RF_bus_sel_savedwin_data_497_port, 
                           curr_proc_regs(496) => 
                           DataPath_RF_bus_sel_savedwin_data_496_port, 
                           curr_proc_regs(495) => 
                           DataPath_RF_bus_sel_savedwin_data_495_port, 
                           curr_proc_regs(494) => 
                           DataPath_RF_bus_sel_savedwin_data_494_port, 
                           curr_proc_regs(493) => 
                           DataPath_RF_bus_sel_savedwin_data_493_port, 
                           curr_proc_regs(492) => 
                           DataPath_RF_bus_sel_savedwin_data_492_port, 
                           curr_proc_regs(491) => 
                           DataPath_RF_bus_sel_savedwin_data_491_port, 
                           curr_proc_regs(490) => 
                           DataPath_RF_bus_sel_savedwin_data_490_port, 
                           curr_proc_regs(489) => 
                           DataPath_RF_bus_sel_savedwin_data_489_port, 
                           curr_proc_regs(488) => 
                           DataPath_RF_bus_sel_savedwin_data_488_port, 
                           curr_proc_regs(487) => 
                           DataPath_RF_bus_sel_savedwin_data_487_port, 
                           curr_proc_regs(486) => 
                           DataPath_RF_bus_sel_savedwin_data_486_port, 
                           curr_proc_regs(485) => 
                           DataPath_RF_bus_sel_savedwin_data_485_port, 
                           curr_proc_regs(484) => 
                           DataPath_RF_bus_sel_savedwin_data_484_port, 
                           curr_proc_regs(483) => 
                           DataPath_RF_bus_sel_savedwin_data_483_port, 
                           curr_proc_regs(482) => 
                           DataPath_RF_bus_sel_savedwin_data_482_port, 
                           curr_proc_regs(481) => 
                           DataPath_RF_bus_sel_savedwin_data_481_port, 
                           curr_proc_regs(480) => 
                           DataPath_RF_bus_sel_savedwin_data_480_port, 
                           curr_proc_regs(479) => 
                           DataPath_RF_bus_sel_savedwin_data_479_port, 
                           curr_proc_regs(478) => 
                           DataPath_RF_bus_sel_savedwin_data_478_port, 
                           curr_proc_regs(477) => 
                           DataPath_RF_bus_sel_savedwin_data_477_port, 
                           curr_proc_regs(476) => 
                           DataPath_RF_bus_sel_savedwin_data_476_port, 
                           curr_proc_regs(475) => 
                           DataPath_RF_bus_sel_savedwin_data_475_port, 
                           curr_proc_regs(474) => 
                           DataPath_RF_bus_sel_savedwin_data_474_port, 
                           curr_proc_regs(473) => 
                           DataPath_RF_bus_sel_savedwin_data_473_port, 
                           curr_proc_regs(472) => 
                           DataPath_RF_bus_sel_savedwin_data_472_port, 
                           curr_proc_regs(471) => 
                           DataPath_RF_bus_sel_savedwin_data_471_port, 
                           curr_proc_regs(470) => 
                           DataPath_RF_bus_sel_savedwin_data_470_port, 
                           curr_proc_regs(469) => 
                           DataPath_RF_bus_sel_savedwin_data_469_port, 
                           curr_proc_regs(468) => 
                           DataPath_RF_bus_sel_savedwin_data_468_port, 
                           curr_proc_regs(467) => 
                           DataPath_RF_bus_sel_savedwin_data_467_port, 
                           curr_proc_regs(466) => 
                           DataPath_RF_bus_sel_savedwin_data_466_port, 
                           curr_proc_regs(465) => 
                           DataPath_RF_bus_sel_savedwin_data_465_port, 
                           curr_proc_regs(464) => 
                           DataPath_RF_bus_sel_savedwin_data_464_port, 
                           curr_proc_regs(463) => 
                           DataPath_RF_bus_sel_savedwin_data_463_port, 
                           curr_proc_regs(462) => 
                           DataPath_RF_bus_sel_savedwin_data_462_port, 
                           curr_proc_regs(461) => 
                           DataPath_RF_bus_sel_savedwin_data_461_port, 
                           curr_proc_regs(460) => 
                           DataPath_RF_bus_sel_savedwin_data_460_port, 
                           curr_proc_regs(459) => 
                           DataPath_RF_bus_sel_savedwin_data_459_port, 
                           curr_proc_regs(458) => 
                           DataPath_RF_bus_sel_savedwin_data_458_port, 
                           curr_proc_regs(457) => 
                           DataPath_RF_bus_sel_savedwin_data_457_port, 
                           curr_proc_regs(456) => 
                           DataPath_RF_bus_sel_savedwin_data_456_port, 
                           curr_proc_regs(455) => 
                           DataPath_RF_bus_sel_savedwin_data_455_port, 
                           curr_proc_regs(454) => 
                           DataPath_RF_bus_sel_savedwin_data_454_port, 
                           curr_proc_regs(453) => 
                           DataPath_RF_bus_sel_savedwin_data_453_port, 
                           curr_proc_regs(452) => 
                           DataPath_RF_bus_sel_savedwin_data_452_port, 
                           curr_proc_regs(451) => 
                           DataPath_RF_bus_sel_savedwin_data_451_port, 
                           curr_proc_regs(450) => 
                           DataPath_RF_bus_sel_savedwin_data_450_port, 
                           curr_proc_regs(449) => 
                           DataPath_RF_bus_sel_savedwin_data_449_port, 
                           curr_proc_regs(448) => 
                           DataPath_RF_bus_sel_savedwin_data_448_port, 
                           curr_proc_regs(447) => 
                           DataPath_RF_bus_sel_savedwin_data_447_port, 
                           curr_proc_regs(446) => 
                           DataPath_RF_bus_sel_savedwin_data_446_port, 
                           curr_proc_regs(445) => 
                           DataPath_RF_bus_sel_savedwin_data_445_port, 
                           curr_proc_regs(444) => 
                           DataPath_RF_bus_sel_savedwin_data_444_port, 
                           curr_proc_regs(443) => 
                           DataPath_RF_bus_sel_savedwin_data_443_port, 
                           curr_proc_regs(442) => 
                           DataPath_RF_bus_sel_savedwin_data_442_port, 
                           curr_proc_regs(441) => 
                           DataPath_RF_bus_sel_savedwin_data_441_port, 
                           curr_proc_regs(440) => 
                           DataPath_RF_bus_sel_savedwin_data_440_port, 
                           curr_proc_regs(439) => 
                           DataPath_RF_bus_sel_savedwin_data_439_port, 
                           curr_proc_regs(438) => 
                           DataPath_RF_bus_sel_savedwin_data_438_port, 
                           curr_proc_regs(437) => 
                           DataPath_RF_bus_sel_savedwin_data_437_port, 
                           curr_proc_regs(436) => 
                           DataPath_RF_bus_sel_savedwin_data_436_port, 
                           curr_proc_regs(435) => 
                           DataPath_RF_bus_sel_savedwin_data_435_port, 
                           curr_proc_regs(434) => 
                           DataPath_RF_bus_sel_savedwin_data_434_port, 
                           curr_proc_regs(433) => 
                           DataPath_RF_bus_sel_savedwin_data_433_port, 
                           curr_proc_regs(432) => 
                           DataPath_RF_bus_sel_savedwin_data_432_port, 
                           curr_proc_regs(431) => 
                           DataPath_RF_bus_sel_savedwin_data_431_port, 
                           curr_proc_regs(430) => 
                           DataPath_RF_bus_sel_savedwin_data_430_port, 
                           curr_proc_regs(429) => 
                           DataPath_RF_bus_sel_savedwin_data_429_port, 
                           curr_proc_regs(428) => 
                           DataPath_RF_bus_sel_savedwin_data_428_port, 
                           curr_proc_regs(427) => 
                           DataPath_RF_bus_sel_savedwin_data_427_port, 
                           curr_proc_regs(426) => 
                           DataPath_RF_bus_sel_savedwin_data_426_port, 
                           curr_proc_regs(425) => 
                           DataPath_RF_bus_sel_savedwin_data_425_port, 
                           curr_proc_regs(424) => 
                           DataPath_RF_bus_sel_savedwin_data_424_port, 
                           curr_proc_regs(423) => 
                           DataPath_RF_bus_sel_savedwin_data_423_port, 
                           curr_proc_regs(422) => 
                           DataPath_RF_bus_sel_savedwin_data_422_port, 
                           curr_proc_regs(421) => 
                           DataPath_RF_bus_sel_savedwin_data_421_port, 
                           curr_proc_regs(420) => 
                           DataPath_RF_bus_sel_savedwin_data_420_port, 
                           curr_proc_regs(419) => 
                           DataPath_RF_bus_sel_savedwin_data_419_port, 
                           curr_proc_regs(418) => 
                           DataPath_RF_bus_sel_savedwin_data_418_port, 
                           curr_proc_regs(417) => 
                           DataPath_RF_bus_sel_savedwin_data_417_port, 
                           curr_proc_regs(416) => 
                           DataPath_RF_bus_sel_savedwin_data_416_port, 
                           curr_proc_regs(415) => 
                           DataPath_RF_bus_sel_savedwin_data_415_port, 
                           curr_proc_regs(414) => 
                           DataPath_RF_bus_sel_savedwin_data_414_port, 
                           curr_proc_regs(413) => 
                           DataPath_RF_bus_sel_savedwin_data_413_port, 
                           curr_proc_regs(412) => 
                           DataPath_RF_bus_sel_savedwin_data_412_port, 
                           curr_proc_regs(411) => 
                           DataPath_RF_bus_sel_savedwin_data_411_port, 
                           curr_proc_regs(410) => 
                           DataPath_RF_bus_sel_savedwin_data_410_port, 
                           curr_proc_regs(409) => 
                           DataPath_RF_bus_sel_savedwin_data_409_port, 
                           curr_proc_regs(408) => 
                           DataPath_RF_bus_sel_savedwin_data_408_port, 
                           curr_proc_regs(407) => 
                           DataPath_RF_bus_sel_savedwin_data_407_port, 
                           curr_proc_regs(406) => 
                           DataPath_RF_bus_sel_savedwin_data_406_port, 
                           curr_proc_regs(405) => 
                           DataPath_RF_bus_sel_savedwin_data_405_port, 
                           curr_proc_regs(404) => 
                           DataPath_RF_bus_sel_savedwin_data_404_port, 
                           curr_proc_regs(403) => 
                           DataPath_RF_bus_sel_savedwin_data_403_port, 
                           curr_proc_regs(402) => 
                           DataPath_RF_bus_sel_savedwin_data_402_port, 
                           curr_proc_regs(401) => 
                           DataPath_RF_bus_sel_savedwin_data_401_port, 
                           curr_proc_regs(400) => 
                           DataPath_RF_bus_sel_savedwin_data_400_port, 
                           curr_proc_regs(399) => 
                           DataPath_RF_bus_sel_savedwin_data_399_port, 
                           curr_proc_regs(398) => 
                           DataPath_RF_bus_sel_savedwin_data_398_port, 
                           curr_proc_regs(397) => 
                           DataPath_RF_bus_sel_savedwin_data_397_port, 
                           curr_proc_regs(396) => 
                           DataPath_RF_bus_sel_savedwin_data_396_port, 
                           curr_proc_regs(395) => 
                           DataPath_RF_bus_sel_savedwin_data_395_port, 
                           curr_proc_regs(394) => 
                           DataPath_RF_bus_sel_savedwin_data_394_port, 
                           curr_proc_regs(393) => 
                           DataPath_RF_bus_sel_savedwin_data_393_port, 
                           curr_proc_regs(392) => 
                           DataPath_RF_bus_sel_savedwin_data_392_port, 
                           curr_proc_regs(391) => 
                           DataPath_RF_bus_sel_savedwin_data_391_port, 
                           curr_proc_regs(390) => 
                           DataPath_RF_bus_sel_savedwin_data_390_port, 
                           curr_proc_regs(389) => 
                           DataPath_RF_bus_sel_savedwin_data_389_port, 
                           curr_proc_regs(388) => 
                           DataPath_RF_bus_sel_savedwin_data_388_port, 
                           curr_proc_regs(387) => 
                           DataPath_RF_bus_sel_savedwin_data_387_port, 
                           curr_proc_regs(386) => 
                           DataPath_RF_bus_sel_savedwin_data_386_port, 
                           curr_proc_regs(385) => 
                           DataPath_RF_bus_sel_savedwin_data_385_port, 
                           curr_proc_regs(384) => 
                           DataPath_RF_bus_sel_savedwin_data_384_port, 
                           curr_proc_regs(383) => 
                           DataPath_RF_bus_sel_savedwin_data_383_port, 
                           curr_proc_regs(382) => 
                           DataPath_RF_bus_sel_savedwin_data_382_port, 
                           curr_proc_regs(381) => 
                           DataPath_RF_bus_sel_savedwin_data_381_port, 
                           curr_proc_regs(380) => 
                           DataPath_RF_bus_sel_savedwin_data_380_port, 
                           curr_proc_regs(379) => 
                           DataPath_RF_bus_sel_savedwin_data_379_port, 
                           curr_proc_regs(378) => 
                           DataPath_RF_bus_sel_savedwin_data_378_port, 
                           curr_proc_regs(377) => 
                           DataPath_RF_bus_sel_savedwin_data_377_port, 
                           curr_proc_regs(376) => 
                           DataPath_RF_bus_sel_savedwin_data_376_port, 
                           curr_proc_regs(375) => 
                           DataPath_RF_bus_sel_savedwin_data_375_port, 
                           curr_proc_regs(374) => 
                           DataPath_RF_bus_sel_savedwin_data_374_port, 
                           curr_proc_regs(373) => 
                           DataPath_RF_bus_sel_savedwin_data_373_port, 
                           curr_proc_regs(372) => 
                           DataPath_RF_bus_sel_savedwin_data_372_port, 
                           curr_proc_regs(371) => 
                           DataPath_RF_bus_sel_savedwin_data_371_port, 
                           curr_proc_regs(370) => 
                           DataPath_RF_bus_sel_savedwin_data_370_port, 
                           curr_proc_regs(369) => 
                           DataPath_RF_bus_sel_savedwin_data_369_port, 
                           curr_proc_regs(368) => 
                           DataPath_RF_bus_sel_savedwin_data_368_port, 
                           curr_proc_regs(367) => 
                           DataPath_RF_bus_sel_savedwin_data_367_port, 
                           curr_proc_regs(366) => 
                           DataPath_RF_bus_sel_savedwin_data_366_port, 
                           curr_proc_regs(365) => 
                           DataPath_RF_bus_sel_savedwin_data_365_port, 
                           curr_proc_regs(364) => 
                           DataPath_RF_bus_sel_savedwin_data_364_port, 
                           curr_proc_regs(363) => 
                           DataPath_RF_bus_sel_savedwin_data_363_port, 
                           curr_proc_regs(362) => 
                           DataPath_RF_bus_sel_savedwin_data_362_port, 
                           curr_proc_regs(361) => 
                           DataPath_RF_bus_sel_savedwin_data_361_port, 
                           curr_proc_regs(360) => 
                           DataPath_RF_bus_sel_savedwin_data_360_port, 
                           curr_proc_regs(359) => 
                           DataPath_RF_bus_sel_savedwin_data_359_port, 
                           curr_proc_regs(358) => 
                           DataPath_RF_bus_sel_savedwin_data_358_port, 
                           curr_proc_regs(357) => 
                           DataPath_RF_bus_sel_savedwin_data_357_port, 
                           curr_proc_regs(356) => 
                           DataPath_RF_bus_sel_savedwin_data_356_port, 
                           curr_proc_regs(355) => 
                           DataPath_RF_bus_sel_savedwin_data_355_port, 
                           curr_proc_regs(354) => 
                           DataPath_RF_bus_sel_savedwin_data_354_port, 
                           curr_proc_regs(353) => 
                           DataPath_RF_bus_sel_savedwin_data_353_port, 
                           curr_proc_regs(352) => 
                           DataPath_RF_bus_sel_savedwin_data_352_port, 
                           curr_proc_regs(351) => 
                           DataPath_RF_bus_sel_savedwin_data_351_port, 
                           curr_proc_regs(350) => 
                           DataPath_RF_bus_sel_savedwin_data_350_port, 
                           curr_proc_regs(349) => 
                           DataPath_RF_bus_sel_savedwin_data_349_port, 
                           curr_proc_regs(348) => 
                           DataPath_RF_bus_sel_savedwin_data_348_port, 
                           curr_proc_regs(347) => 
                           DataPath_RF_bus_sel_savedwin_data_347_port, 
                           curr_proc_regs(346) => 
                           DataPath_RF_bus_sel_savedwin_data_346_port, 
                           curr_proc_regs(345) => 
                           DataPath_RF_bus_sel_savedwin_data_345_port, 
                           curr_proc_regs(344) => 
                           DataPath_RF_bus_sel_savedwin_data_344_port, 
                           curr_proc_regs(343) => 
                           DataPath_RF_bus_sel_savedwin_data_343_port, 
                           curr_proc_regs(342) => 
                           DataPath_RF_bus_sel_savedwin_data_342_port, 
                           curr_proc_regs(341) => 
                           DataPath_RF_bus_sel_savedwin_data_341_port, 
                           curr_proc_regs(340) => 
                           DataPath_RF_bus_sel_savedwin_data_340_port, 
                           curr_proc_regs(339) => 
                           DataPath_RF_bus_sel_savedwin_data_339_port, 
                           curr_proc_regs(338) => 
                           DataPath_RF_bus_sel_savedwin_data_338_port, 
                           curr_proc_regs(337) => 
                           DataPath_RF_bus_sel_savedwin_data_337_port, 
                           curr_proc_regs(336) => 
                           DataPath_RF_bus_sel_savedwin_data_336_port, 
                           curr_proc_regs(335) => 
                           DataPath_RF_bus_sel_savedwin_data_335_port, 
                           curr_proc_regs(334) => 
                           DataPath_RF_bus_sel_savedwin_data_334_port, 
                           curr_proc_regs(333) => 
                           DataPath_RF_bus_sel_savedwin_data_333_port, 
                           curr_proc_regs(332) => 
                           DataPath_RF_bus_sel_savedwin_data_332_port, 
                           curr_proc_regs(331) => 
                           DataPath_RF_bus_sel_savedwin_data_331_port, 
                           curr_proc_regs(330) => 
                           DataPath_RF_bus_sel_savedwin_data_330_port, 
                           curr_proc_regs(329) => 
                           DataPath_RF_bus_sel_savedwin_data_329_port, 
                           curr_proc_regs(328) => 
                           DataPath_RF_bus_sel_savedwin_data_328_port, 
                           curr_proc_regs(327) => 
                           DataPath_RF_bus_sel_savedwin_data_327_port, 
                           curr_proc_regs(326) => 
                           DataPath_RF_bus_sel_savedwin_data_326_port, 
                           curr_proc_regs(325) => 
                           DataPath_RF_bus_sel_savedwin_data_325_port, 
                           curr_proc_regs(324) => 
                           DataPath_RF_bus_sel_savedwin_data_324_port, 
                           curr_proc_regs(323) => 
                           DataPath_RF_bus_sel_savedwin_data_323_port, 
                           curr_proc_regs(322) => 
                           DataPath_RF_bus_sel_savedwin_data_322_port, 
                           curr_proc_regs(321) => 
                           DataPath_RF_bus_sel_savedwin_data_321_port, 
                           curr_proc_regs(320) => 
                           DataPath_RF_bus_sel_savedwin_data_320_port, 
                           curr_proc_regs(319) => 
                           DataPath_RF_bus_sel_savedwin_data_319_port, 
                           curr_proc_regs(318) => 
                           DataPath_RF_bus_sel_savedwin_data_318_port, 
                           curr_proc_regs(317) => 
                           DataPath_RF_bus_sel_savedwin_data_317_port, 
                           curr_proc_regs(316) => 
                           DataPath_RF_bus_sel_savedwin_data_316_port, 
                           curr_proc_regs(315) => 
                           DataPath_RF_bus_sel_savedwin_data_315_port, 
                           curr_proc_regs(314) => 
                           DataPath_RF_bus_sel_savedwin_data_314_port, 
                           curr_proc_regs(313) => 
                           DataPath_RF_bus_sel_savedwin_data_313_port, 
                           curr_proc_regs(312) => 
                           DataPath_RF_bus_sel_savedwin_data_312_port, 
                           curr_proc_regs(311) => 
                           DataPath_RF_bus_sel_savedwin_data_311_port, 
                           curr_proc_regs(310) => 
                           DataPath_RF_bus_sel_savedwin_data_310_port, 
                           curr_proc_regs(309) => 
                           DataPath_RF_bus_sel_savedwin_data_309_port, 
                           curr_proc_regs(308) => 
                           DataPath_RF_bus_sel_savedwin_data_308_port, 
                           curr_proc_regs(307) => 
                           DataPath_RF_bus_sel_savedwin_data_307_port, 
                           curr_proc_regs(306) => 
                           DataPath_RF_bus_sel_savedwin_data_306_port, 
                           curr_proc_regs(305) => 
                           DataPath_RF_bus_sel_savedwin_data_305_port, 
                           curr_proc_regs(304) => 
                           DataPath_RF_bus_sel_savedwin_data_304_port, 
                           curr_proc_regs(303) => 
                           DataPath_RF_bus_sel_savedwin_data_303_port, 
                           curr_proc_regs(302) => 
                           DataPath_RF_bus_sel_savedwin_data_302_port, 
                           curr_proc_regs(301) => 
                           DataPath_RF_bus_sel_savedwin_data_301_port, 
                           curr_proc_regs(300) => 
                           DataPath_RF_bus_sel_savedwin_data_300_port, 
                           curr_proc_regs(299) => 
                           DataPath_RF_bus_sel_savedwin_data_299_port, 
                           curr_proc_regs(298) => 
                           DataPath_RF_bus_sel_savedwin_data_298_port, 
                           curr_proc_regs(297) => 
                           DataPath_RF_bus_sel_savedwin_data_297_port, 
                           curr_proc_regs(296) => 
                           DataPath_RF_bus_sel_savedwin_data_296_port, 
                           curr_proc_regs(295) => 
                           DataPath_RF_bus_sel_savedwin_data_295_port, 
                           curr_proc_regs(294) => 
                           DataPath_RF_bus_sel_savedwin_data_294_port, 
                           curr_proc_regs(293) => 
                           DataPath_RF_bus_sel_savedwin_data_293_port, 
                           curr_proc_regs(292) => 
                           DataPath_RF_bus_sel_savedwin_data_292_port, 
                           curr_proc_regs(291) => 
                           DataPath_RF_bus_sel_savedwin_data_291_port, 
                           curr_proc_regs(290) => 
                           DataPath_RF_bus_sel_savedwin_data_290_port, 
                           curr_proc_regs(289) => 
                           DataPath_RF_bus_sel_savedwin_data_289_port, 
                           curr_proc_regs(288) => 
                           DataPath_RF_bus_sel_savedwin_data_288_port, 
                           curr_proc_regs(287) => 
                           DataPath_RF_bus_sel_savedwin_data_287_port, 
                           curr_proc_regs(286) => 
                           DataPath_RF_bus_sel_savedwin_data_286_port, 
                           curr_proc_regs(285) => 
                           DataPath_RF_bus_sel_savedwin_data_285_port, 
                           curr_proc_regs(284) => 
                           DataPath_RF_bus_sel_savedwin_data_284_port, 
                           curr_proc_regs(283) => 
                           DataPath_RF_bus_sel_savedwin_data_283_port, 
                           curr_proc_regs(282) => 
                           DataPath_RF_bus_sel_savedwin_data_282_port, 
                           curr_proc_regs(281) => 
                           DataPath_RF_bus_sel_savedwin_data_281_port, 
                           curr_proc_regs(280) => 
                           DataPath_RF_bus_sel_savedwin_data_280_port, 
                           curr_proc_regs(279) => 
                           DataPath_RF_bus_sel_savedwin_data_279_port, 
                           curr_proc_regs(278) => 
                           DataPath_RF_bus_sel_savedwin_data_278_port, 
                           curr_proc_regs(277) => 
                           DataPath_RF_bus_sel_savedwin_data_277_port, 
                           curr_proc_regs(276) => 
                           DataPath_RF_bus_sel_savedwin_data_276_port, 
                           curr_proc_regs(275) => 
                           DataPath_RF_bus_sel_savedwin_data_275_port, 
                           curr_proc_regs(274) => 
                           DataPath_RF_bus_sel_savedwin_data_274_port, 
                           curr_proc_regs(273) => 
                           DataPath_RF_bus_sel_savedwin_data_273_port, 
                           curr_proc_regs(272) => 
                           DataPath_RF_bus_sel_savedwin_data_272_port, 
                           curr_proc_regs(271) => 
                           DataPath_RF_bus_sel_savedwin_data_271_port, 
                           curr_proc_regs(270) => 
                           DataPath_RF_bus_sel_savedwin_data_270_port, 
                           curr_proc_regs(269) => 
                           DataPath_RF_bus_sel_savedwin_data_269_port, 
                           curr_proc_regs(268) => 
                           DataPath_RF_bus_sel_savedwin_data_268_port, 
                           curr_proc_regs(267) => 
                           DataPath_RF_bus_sel_savedwin_data_267_port, 
                           curr_proc_regs(266) => 
                           DataPath_RF_bus_sel_savedwin_data_266_port, 
                           curr_proc_regs(265) => 
                           DataPath_RF_bus_sel_savedwin_data_265_port, 
                           curr_proc_regs(264) => 
                           DataPath_RF_bus_sel_savedwin_data_264_port, 
                           curr_proc_regs(263) => 
                           DataPath_RF_bus_sel_savedwin_data_263_port, 
                           curr_proc_regs(262) => 
                           DataPath_RF_bus_sel_savedwin_data_262_port, 
                           curr_proc_regs(261) => 
                           DataPath_RF_bus_sel_savedwin_data_261_port, 
                           curr_proc_regs(260) => 
                           DataPath_RF_bus_sel_savedwin_data_260_port, 
                           curr_proc_regs(259) => 
                           DataPath_RF_bus_sel_savedwin_data_259_port, 
                           curr_proc_regs(258) => 
                           DataPath_RF_bus_sel_savedwin_data_258_port, 
                           curr_proc_regs(257) => 
                           DataPath_RF_bus_sel_savedwin_data_257_port, 
                           curr_proc_regs(256) => 
                           DataPath_RF_bus_sel_savedwin_data_256_port, 
                           curr_proc_regs(255) => 
                           DataPath_RF_bus_sel_savedwin_data_255_port, 
                           curr_proc_regs(254) => 
                           DataPath_RF_bus_sel_savedwin_data_254_port, 
                           curr_proc_regs(253) => 
                           DataPath_RF_bus_sel_savedwin_data_253_port, 
                           curr_proc_regs(252) => 
                           DataPath_RF_bus_sel_savedwin_data_252_port, 
                           curr_proc_regs(251) => 
                           DataPath_RF_bus_sel_savedwin_data_251_port, 
                           curr_proc_regs(250) => 
                           DataPath_RF_bus_sel_savedwin_data_250_port, 
                           curr_proc_regs(249) => 
                           DataPath_RF_bus_sel_savedwin_data_249_port, 
                           curr_proc_regs(248) => 
                           DataPath_RF_bus_sel_savedwin_data_248_port, 
                           curr_proc_regs(247) => 
                           DataPath_RF_bus_sel_savedwin_data_247_port, 
                           curr_proc_regs(246) => 
                           DataPath_RF_bus_sel_savedwin_data_246_port, 
                           curr_proc_regs(245) => 
                           DataPath_RF_bus_sel_savedwin_data_245_port, 
                           curr_proc_regs(244) => 
                           DataPath_RF_bus_sel_savedwin_data_244_port, 
                           curr_proc_regs(243) => 
                           DataPath_RF_bus_sel_savedwin_data_243_port, 
                           curr_proc_regs(242) => 
                           DataPath_RF_bus_sel_savedwin_data_242_port, 
                           curr_proc_regs(241) => 
                           DataPath_RF_bus_sel_savedwin_data_241_port, 
                           curr_proc_regs(240) => 
                           DataPath_RF_bus_sel_savedwin_data_240_port, 
                           curr_proc_regs(239) => 
                           DataPath_RF_bus_sel_savedwin_data_239_port, 
                           curr_proc_regs(238) => 
                           DataPath_RF_bus_sel_savedwin_data_238_port, 
                           curr_proc_regs(237) => 
                           DataPath_RF_bus_sel_savedwin_data_237_port, 
                           curr_proc_regs(236) => 
                           DataPath_RF_bus_sel_savedwin_data_236_port, 
                           curr_proc_regs(235) => 
                           DataPath_RF_bus_sel_savedwin_data_235_port, 
                           curr_proc_regs(234) => 
                           DataPath_RF_bus_sel_savedwin_data_234_port, 
                           curr_proc_regs(233) => 
                           DataPath_RF_bus_sel_savedwin_data_233_port, 
                           curr_proc_regs(232) => 
                           DataPath_RF_bus_sel_savedwin_data_232_port, 
                           curr_proc_regs(231) => 
                           DataPath_RF_bus_sel_savedwin_data_231_port, 
                           curr_proc_regs(230) => 
                           DataPath_RF_bus_sel_savedwin_data_230_port, 
                           curr_proc_regs(229) => 
                           DataPath_RF_bus_sel_savedwin_data_229_port, 
                           curr_proc_regs(228) => 
                           DataPath_RF_bus_sel_savedwin_data_228_port, 
                           curr_proc_regs(227) => 
                           DataPath_RF_bus_sel_savedwin_data_227_port, 
                           curr_proc_regs(226) => 
                           DataPath_RF_bus_sel_savedwin_data_226_port, 
                           curr_proc_regs(225) => 
                           DataPath_RF_bus_sel_savedwin_data_225_port, 
                           curr_proc_regs(224) => 
                           DataPath_RF_bus_sel_savedwin_data_224_port, 
                           curr_proc_regs(223) => 
                           DataPath_RF_bus_sel_savedwin_data_223_port, 
                           curr_proc_regs(222) => 
                           DataPath_RF_bus_sel_savedwin_data_222_port, 
                           curr_proc_regs(221) => 
                           DataPath_RF_bus_sel_savedwin_data_221_port, 
                           curr_proc_regs(220) => 
                           DataPath_RF_bus_sel_savedwin_data_220_port, 
                           curr_proc_regs(219) => 
                           DataPath_RF_bus_sel_savedwin_data_219_port, 
                           curr_proc_regs(218) => 
                           DataPath_RF_bus_sel_savedwin_data_218_port, 
                           curr_proc_regs(217) => 
                           DataPath_RF_bus_sel_savedwin_data_217_port, 
                           curr_proc_regs(216) => 
                           DataPath_RF_bus_sel_savedwin_data_216_port, 
                           curr_proc_regs(215) => 
                           DataPath_RF_bus_sel_savedwin_data_215_port, 
                           curr_proc_regs(214) => 
                           DataPath_RF_bus_sel_savedwin_data_214_port, 
                           curr_proc_regs(213) => 
                           DataPath_RF_bus_sel_savedwin_data_213_port, 
                           curr_proc_regs(212) => 
                           DataPath_RF_bus_sel_savedwin_data_212_port, 
                           curr_proc_regs(211) => 
                           DataPath_RF_bus_sel_savedwin_data_211_port, 
                           curr_proc_regs(210) => 
                           DataPath_RF_bus_sel_savedwin_data_210_port, 
                           curr_proc_regs(209) => 
                           DataPath_RF_bus_sel_savedwin_data_209_port, 
                           curr_proc_regs(208) => 
                           DataPath_RF_bus_sel_savedwin_data_208_port, 
                           curr_proc_regs(207) => 
                           DataPath_RF_bus_sel_savedwin_data_207_port, 
                           curr_proc_regs(206) => 
                           DataPath_RF_bus_sel_savedwin_data_206_port, 
                           curr_proc_regs(205) => 
                           DataPath_RF_bus_sel_savedwin_data_205_port, 
                           curr_proc_regs(204) => 
                           DataPath_RF_bus_sel_savedwin_data_204_port, 
                           curr_proc_regs(203) => 
                           DataPath_RF_bus_sel_savedwin_data_203_port, 
                           curr_proc_regs(202) => 
                           DataPath_RF_bus_sel_savedwin_data_202_port, 
                           curr_proc_regs(201) => 
                           DataPath_RF_bus_sel_savedwin_data_201_port, 
                           curr_proc_regs(200) => 
                           DataPath_RF_bus_sel_savedwin_data_200_port, 
                           curr_proc_regs(199) => 
                           DataPath_RF_bus_sel_savedwin_data_199_port, 
                           curr_proc_regs(198) => 
                           DataPath_RF_bus_sel_savedwin_data_198_port, 
                           curr_proc_regs(197) => 
                           DataPath_RF_bus_sel_savedwin_data_197_port, 
                           curr_proc_regs(196) => 
                           DataPath_RF_bus_sel_savedwin_data_196_port, 
                           curr_proc_regs(195) => 
                           DataPath_RF_bus_sel_savedwin_data_195_port, 
                           curr_proc_regs(194) => 
                           DataPath_RF_bus_sel_savedwin_data_194_port, 
                           curr_proc_regs(193) => 
                           DataPath_RF_bus_sel_savedwin_data_193_port, 
                           curr_proc_regs(192) => 
                           DataPath_RF_bus_sel_savedwin_data_192_port, 
                           curr_proc_regs(191) => 
                           DataPath_RF_bus_sel_savedwin_data_191_port, 
                           curr_proc_regs(190) => 
                           DataPath_RF_bus_sel_savedwin_data_190_port, 
                           curr_proc_regs(189) => 
                           DataPath_RF_bus_sel_savedwin_data_189_port, 
                           curr_proc_regs(188) => 
                           DataPath_RF_bus_sel_savedwin_data_188_port, 
                           curr_proc_regs(187) => 
                           DataPath_RF_bus_sel_savedwin_data_187_port, 
                           curr_proc_regs(186) => 
                           DataPath_RF_bus_sel_savedwin_data_186_port, 
                           curr_proc_regs(185) => 
                           DataPath_RF_bus_sel_savedwin_data_185_port, 
                           curr_proc_regs(184) => 
                           DataPath_RF_bus_sel_savedwin_data_184_port, 
                           curr_proc_regs(183) => 
                           DataPath_RF_bus_sel_savedwin_data_183_port, 
                           curr_proc_regs(182) => 
                           DataPath_RF_bus_sel_savedwin_data_182_port, 
                           curr_proc_regs(181) => 
                           DataPath_RF_bus_sel_savedwin_data_181_port, 
                           curr_proc_regs(180) => 
                           DataPath_RF_bus_sel_savedwin_data_180_port, 
                           curr_proc_regs(179) => 
                           DataPath_RF_bus_sel_savedwin_data_179_port, 
                           curr_proc_regs(178) => 
                           DataPath_RF_bus_sel_savedwin_data_178_port, 
                           curr_proc_regs(177) => 
                           DataPath_RF_bus_sel_savedwin_data_177_port, 
                           curr_proc_regs(176) => 
                           DataPath_RF_bus_sel_savedwin_data_176_port, 
                           curr_proc_regs(175) => 
                           DataPath_RF_bus_sel_savedwin_data_175_port, 
                           curr_proc_regs(174) => 
                           DataPath_RF_bus_sel_savedwin_data_174_port, 
                           curr_proc_regs(173) => 
                           DataPath_RF_bus_sel_savedwin_data_173_port, 
                           curr_proc_regs(172) => 
                           DataPath_RF_bus_sel_savedwin_data_172_port, 
                           curr_proc_regs(171) => 
                           DataPath_RF_bus_sel_savedwin_data_171_port, 
                           curr_proc_regs(170) => 
                           DataPath_RF_bus_sel_savedwin_data_170_port, 
                           curr_proc_regs(169) => 
                           DataPath_RF_bus_sel_savedwin_data_169_port, 
                           curr_proc_regs(168) => 
                           DataPath_RF_bus_sel_savedwin_data_168_port, 
                           curr_proc_regs(167) => 
                           DataPath_RF_bus_sel_savedwin_data_167_port, 
                           curr_proc_regs(166) => 
                           DataPath_RF_bus_sel_savedwin_data_166_port, 
                           curr_proc_regs(165) => 
                           DataPath_RF_bus_sel_savedwin_data_165_port, 
                           curr_proc_regs(164) => 
                           DataPath_RF_bus_sel_savedwin_data_164_port, 
                           curr_proc_regs(163) => 
                           DataPath_RF_bus_sel_savedwin_data_163_port, 
                           curr_proc_regs(162) => 
                           DataPath_RF_bus_sel_savedwin_data_162_port, 
                           curr_proc_regs(161) => 
                           DataPath_RF_bus_sel_savedwin_data_161_port, 
                           curr_proc_regs(160) => 
                           DataPath_RF_bus_sel_savedwin_data_160_port, 
                           curr_proc_regs(159) => 
                           DataPath_RF_bus_sel_savedwin_data_159_port, 
                           curr_proc_regs(158) => 
                           DataPath_RF_bus_sel_savedwin_data_158_port, 
                           curr_proc_regs(157) => 
                           DataPath_RF_bus_sel_savedwin_data_157_port, 
                           curr_proc_regs(156) => 
                           DataPath_RF_bus_sel_savedwin_data_156_port, 
                           curr_proc_regs(155) => 
                           DataPath_RF_bus_sel_savedwin_data_155_port, 
                           curr_proc_regs(154) => 
                           DataPath_RF_bus_sel_savedwin_data_154_port, 
                           curr_proc_regs(153) => 
                           DataPath_RF_bus_sel_savedwin_data_153_port, 
                           curr_proc_regs(152) => 
                           DataPath_RF_bus_sel_savedwin_data_152_port, 
                           curr_proc_regs(151) => 
                           DataPath_RF_bus_sel_savedwin_data_151_port, 
                           curr_proc_regs(150) => 
                           DataPath_RF_bus_sel_savedwin_data_150_port, 
                           curr_proc_regs(149) => 
                           DataPath_RF_bus_sel_savedwin_data_149_port, 
                           curr_proc_regs(148) => 
                           DataPath_RF_bus_sel_savedwin_data_148_port, 
                           curr_proc_regs(147) => 
                           DataPath_RF_bus_sel_savedwin_data_147_port, 
                           curr_proc_regs(146) => 
                           DataPath_RF_bus_sel_savedwin_data_146_port, 
                           curr_proc_regs(145) => 
                           DataPath_RF_bus_sel_savedwin_data_145_port, 
                           curr_proc_regs(144) => 
                           DataPath_RF_bus_sel_savedwin_data_144_port, 
                           curr_proc_regs(143) => 
                           DataPath_RF_bus_sel_savedwin_data_143_port, 
                           curr_proc_regs(142) => 
                           DataPath_RF_bus_sel_savedwin_data_142_port, 
                           curr_proc_regs(141) => 
                           DataPath_RF_bus_sel_savedwin_data_141_port, 
                           curr_proc_regs(140) => 
                           DataPath_RF_bus_sel_savedwin_data_140_port, 
                           curr_proc_regs(139) => 
                           DataPath_RF_bus_sel_savedwin_data_139_port, 
                           curr_proc_regs(138) => 
                           DataPath_RF_bus_sel_savedwin_data_138_port, 
                           curr_proc_regs(137) => 
                           DataPath_RF_bus_sel_savedwin_data_137_port, 
                           curr_proc_regs(136) => 
                           DataPath_RF_bus_sel_savedwin_data_136_port, 
                           curr_proc_regs(135) => 
                           DataPath_RF_bus_sel_savedwin_data_135_port, 
                           curr_proc_regs(134) => 
                           DataPath_RF_bus_sel_savedwin_data_134_port, 
                           curr_proc_regs(133) => 
                           DataPath_RF_bus_sel_savedwin_data_133_port, 
                           curr_proc_regs(132) => 
                           DataPath_RF_bus_sel_savedwin_data_132_port, 
                           curr_proc_regs(131) => 
                           DataPath_RF_bus_sel_savedwin_data_131_port, 
                           curr_proc_regs(130) => 
                           DataPath_RF_bus_sel_savedwin_data_130_port, 
                           curr_proc_regs(129) => 
                           DataPath_RF_bus_sel_savedwin_data_129_port, 
                           curr_proc_regs(128) => 
                           DataPath_RF_bus_sel_savedwin_data_128_port, 
                           curr_proc_regs(127) => 
                           DataPath_RF_bus_sel_savedwin_data_127_port, 
                           curr_proc_regs(126) => 
                           DataPath_RF_bus_sel_savedwin_data_126_port, 
                           curr_proc_regs(125) => 
                           DataPath_RF_bus_sel_savedwin_data_125_port, 
                           curr_proc_regs(124) => 
                           DataPath_RF_bus_sel_savedwin_data_124_port, 
                           curr_proc_regs(123) => 
                           DataPath_RF_bus_sel_savedwin_data_123_port, 
                           curr_proc_regs(122) => 
                           DataPath_RF_bus_sel_savedwin_data_122_port, 
                           curr_proc_regs(121) => 
                           DataPath_RF_bus_sel_savedwin_data_121_port, 
                           curr_proc_regs(120) => 
                           DataPath_RF_bus_sel_savedwin_data_120_port, 
                           curr_proc_regs(119) => 
                           DataPath_RF_bus_sel_savedwin_data_119_port, 
                           curr_proc_regs(118) => 
                           DataPath_RF_bus_sel_savedwin_data_118_port, 
                           curr_proc_regs(117) => 
                           DataPath_RF_bus_sel_savedwin_data_117_port, 
                           curr_proc_regs(116) => 
                           DataPath_RF_bus_sel_savedwin_data_116_port, 
                           curr_proc_regs(115) => 
                           DataPath_RF_bus_sel_savedwin_data_115_port, 
                           curr_proc_regs(114) => 
                           DataPath_RF_bus_sel_savedwin_data_114_port, 
                           curr_proc_regs(113) => 
                           DataPath_RF_bus_sel_savedwin_data_113_port, 
                           curr_proc_regs(112) => 
                           DataPath_RF_bus_sel_savedwin_data_112_port, 
                           curr_proc_regs(111) => 
                           DataPath_RF_bus_sel_savedwin_data_111_port, 
                           curr_proc_regs(110) => 
                           DataPath_RF_bus_sel_savedwin_data_110_port, 
                           curr_proc_regs(109) => 
                           DataPath_RF_bus_sel_savedwin_data_109_port, 
                           curr_proc_regs(108) => 
                           DataPath_RF_bus_sel_savedwin_data_108_port, 
                           curr_proc_regs(107) => 
                           DataPath_RF_bus_sel_savedwin_data_107_port, 
                           curr_proc_regs(106) => 
                           DataPath_RF_bus_sel_savedwin_data_106_port, 
                           curr_proc_regs(105) => 
                           DataPath_RF_bus_sel_savedwin_data_105_port, 
                           curr_proc_regs(104) => 
                           DataPath_RF_bus_sel_savedwin_data_104_port, 
                           curr_proc_regs(103) => 
                           DataPath_RF_bus_sel_savedwin_data_103_port, 
                           curr_proc_regs(102) => 
                           DataPath_RF_bus_sel_savedwin_data_102_port, 
                           curr_proc_regs(101) => 
                           DataPath_RF_bus_sel_savedwin_data_101_port, 
                           curr_proc_regs(100) => 
                           DataPath_RF_bus_sel_savedwin_data_100_port, 
                           curr_proc_regs(99) => 
                           DataPath_RF_bus_sel_savedwin_data_99_port, 
                           curr_proc_regs(98) => 
                           DataPath_RF_bus_sel_savedwin_data_98_port, 
                           curr_proc_regs(97) => 
                           DataPath_RF_bus_sel_savedwin_data_97_port, 
                           curr_proc_regs(96) => 
                           DataPath_RF_bus_sel_savedwin_data_96_port, 
                           curr_proc_regs(95) => 
                           DataPath_RF_bus_sel_savedwin_data_95_port, 
                           curr_proc_regs(94) => 
                           DataPath_RF_bus_sel_savedwin_data_94_port, 
                           curr_proc_regs(93) => 
                           DataPath_RF_bus_sel_savedwin_data_93_port, 
                           curr_proc_regs(92) => 
                           DataPath_RF_bus_sel_savedwin_data_92_port, 
                           curr_proc_regs(91) => 
                           DataPath_RF_bus_sel_savedwin_data_91_port, 
                           curr_proc_regs(90) => 
                           DataPath_RF_bus_sel_savedwin_data_90_port, 
                           curr_proc_regs(89) => 
                           DataPath_RF_bus_sel_savedwin_data_89_port, 
                           curr_proc_regs(88) => 
                           DataPath_RF_bus_sel_savedwin_data_88_port, 
                           curr_proc_regs(87) => 
                           DataPath_RF_bus_sel_savedwin_data_87_port, 
                           curr_proc_regs(86) => 
                           DataPath_RF_bus_sel_savedwin_data_86_port, 
                           curr_proc_regs(85) => 
                           DataPath_RF_bus_sel_savedwin_data_85_port, 
                           curr_proc_regs(84) => 
                           DataPath_RF_bus_sel_savedwin_data_84_port, 
                           curr_proc_regs(83) => 
                           DataPath_RF_bus_sel_savedwin_data_83_port, 
                           curr_proc_regs(82) => 
                           DataPath_RF_bus_sel_savedwin_data_82_port, 
                           curr_proc_regs(81) => 
                           DataPath_RF_bus_sel_savedwin_data_81_port, 
                           curr_proc_regs(80) => 
                           DataPath_RF_bus_sel_savedwin_data_80_port, 
                           curr_proc_regs(79) => 
                           DataPath_RF_bus_sel_savedwin_data_79_port, 
                           curr_proc_regs(78) => 
                           DataPath_RF_bus_sel_savedwin_data_78_port, 
                           curr_proc_regs(77) => 
                           DataPath_RF_bus_sel_savedwin_data_77_port, 
                           curr_proc_regs(76) => 
                           DataPath_RF_bus_sel_savedwin_data_76_port, 
                           curr_proc_regs(75) => 
                           DataPath_RF_bus_sel_savedwin_data_75_port, 
                           curr_proc_regs(74) => 
                           DataPath_RF_bus_sel_savedwin_data_74_port, 
                           curr_proc_regs(73) => 
                           DataPath_RF_bus_sel_savedwin_data_73_port, 
                           curr_proc_regs(72) => 
                           DataPath_RF_bus_sel_savedwin_data_72_port, 
                           curr_proc_regs(71) => 
                           DataPath_RF_bus_sel_savedwin_data_71_port, 
                           curr_proc_regs(70) => 
                           DataPath_RF_bus_sel_savedwin_data_70_port, 
                           curr_proc_regs(69) => 
                           DataPath_RF_bus_sel_savedwin_data_69_port, 
                           curr_proc_regs(68) => 
                           DataPath_RF_bus_sel_savedwin_data_68_port, 
                           curr_proc_regs(67) => 
                           DataPath_RF_bus_sel_savedwin_data_67_port, 
                           curr_proc_regs(66) => 
                           DataPath_RF_bus_sel_savedwin_data_66_port, 
                           curr_proc_regs(65) => 
                           DataPath_RF_bus_sel_savedwin_data_65_port, 
                           curr_proc_regs(64) => 
                           DataPath_RF_bus_sel_savedwin_data_64_port, 
                           curr_proc_regs(63) => 
                           DataPath_RF_bus_sel_savedwin_data_63_port, 
                           curr_proc_regs(62) => 
                           DataPath_RF_bus_sel_savedwin_data_62_port, 
                           curr_proc_regs(61) => 
                           DataPath_RF_bus_sel_savedwin_data_61_port, 
                           curr_proc_regs(60) => 
                           DataPath_RF_bus_sel_savedwin_data_60_port, 
                           curr_proc_regs(59) => 
                           DataPath_RF_bus_sel_savedwin_data_59_port, 
                           curr_proc_regs(58) => 
                           DataPath_RF_bus_sel_savedwin_data_58_port, 
                           curr_proc_regs(57) => 
                           DataPath_RF_bus_sel_savedwin_data_57_port, 
                           curr_proc_regs(56) => 
                           DataPath_RF_bus_sel_savedwin_data_56_port, 
                           curr_proc_regs(55) => 
                           DataPath_RF_bus_sel_savedwin_data_55_port, 
                           curr_proc_regs(54) => 
                           DataPath_RF_bus_sel_savedwin_data_54_port, 
                           curr_proc_regs(53) => 
                           DataPath_RF_bus_sel_savedwin_data_53_port, 
                           curr_proc_regs(52) => 
                           DataPath_RF_bus_sel_savedwin_data_52_port, 
                           curr_proc_regs(51) => 
                           DataPath_RF_bus_sel_savedwin_data_51_port, 
                           curr_proc_regs(50) => 
                           DataPath_RF_bus_sel_savedwin_data_50_port, 
                           curr_proc_regs(49) => 
                           DataPath_RF_bus_sel_savedwin_data_49_port, 
                           curr_proc_regs(48) => 
                           DataPath_RF_bus_sel_savedwin_data_48_port, 
                           curr_proc_regs(47) => 
                           DataPath_RF_bus_sel_savedwin_data_47_port, 
                           curr_proc_regs(46) => 
                           DataPath_RF_bus_sel_savedwin_data_46_port, 
                           curr_proc_regs(45) => 
                           DataPath_RF_bus_sel_savedwin_data_45_port, 
                           curr_proc_regs(44) => 
                           DataPath_RF_bus_sel_savedwin_data_44_port, 
                           curr_proc_regs(43) => 
                           DataPath_RF_bus_sel_savedwin_data_43_port, 
                           curr_proc_regs(42) => 
                           DataPath_RF_bus_sel_savedwin_data_42_port, 
                           curr_proc_regs(41) => 
                           DataPath_RF_bus_sel_savedwin_data_41_port, 
                           curr_proc_regs(40) => 
                           DataPath_RF_bus_sel_savedwin_data_40_port, 
                           curr_proc_regs(39) => 
                           DataPath_RF_bus_sel_savedwin_data_39_port, 
                           curr_proc_regs(38) => 
                           DataPath_RF_bus_sel_savedwin_data_38_port, 
                           curr_proc_regs(37) => 
                           DataPath_RF_bus_sel_savedwin_data_37_port, 
                           curr_proc_regs(36) => 
                           DataPath_RF_bus_sel_savedwin_data_36_port, 
                           curr_proc_regs(35) => 
                           DataPath_RF_bus_sel_savedwin_data_35_port, 
                           curr_proc_regs(34) => 
                           DataPath_RF_bus_sel_savedwin_data_34_port, 
                           curr_proc_regs(33) => 
                           DataPath_RF_bus_sel_savedwin_data_33_port, 
                           curr_proc_regs(32) => 
                           DataPath_RF_bus_sel_savedwin_data_32_port, 
                           curr_proc_regs(31) => 
                           DataPath_RF_bus_sel_savedwin_data_31_port, 
                           curr_proc_regs(30) => 
                           DataPath_RF_bus_sel_savedwin_data_30_port, 
                           curr_proc_regs(29) => 
                           DataPath_RF_bus_sel_savedwin_data_29_port, 
                           curr_proc_regs(28) => 
                           DataPath_RF_bus_sel_savedwin_data_28_port, 
                           curr_proc_regs(27) => 
                           DataPath_RF_bus_sel_savedwin_data_27_port, 
                           curr_proc_regs(26) => 
                           DataPath_RF_bus_sel_savedwin_data_26_port, 
                           curr_proc_regs(25) => 
                           DataPath_RF_bus_sel_savedwin_data_25_port, 
                           curr_proc_regs(24) => 
                           DataPath_RF_bus_sel_savedwin_data_24_port, 
                           curr_proc_regs(23) => 
                           DataPath_RF_bus_sel_savedwin_data_23_port, 
                           curr_proc_regs(22) => 
                           DataPath_RF_bus_sel_savedwin_data_22_port, 
                           curr_proc_regs(21) => 
                           DataPath_RF_bus_sel_savedwin_data_21_port, 
                           curr_proc_regs(20) => 
                           DataPath_RF_bus_sel_savedwin_data_20_port, 
                           curr_proc_regs(19) => 
                           DataPath_RF_bus_sel_savedwin_data_19_port, 
                           curr_proc_regs(18) => 
                           DataPath_RF_bus_sel_savedwin_data_18_port, 
                           curr_proc_regs(17) => 
                           DataPath_RF_bus_sel_savedwin_data_17_port, 
                           curr_proc_regs(16) => 
                           DataPath_RF_bus_sel_savedwin_data_16_port, 
                           curr_proc_regs(15) => 
                           DataPath_RF_bus_sel_savedwin_data_15_port, 
                           curr_proc_regs(14) => 
                           DataPath_RF_bus_sel_savedwin_data_14_port, 
                           curr_proc_regs(13) => 
                           DataPath_RF_bus_sel_savedwin_data_13_port, 
                           curr_proc_regs(12) => 
                           DataPath_RF_bus_sel_savedwin_data_12_port, 
                           curr_proc_regs(11) => 
                           DataPath_RF_bus_sel_savedwin_data_11_port, 
                           curr_proc_regs(10) => 
                           DataPath_RF_bus_sel_savedwin_data_10_port, 
                           curr_proc_regs(9) => 
                           DataPath_RF_bus_sel_savedwin_data_9_port, 
                           curr_proc_regs(8) => 
                           DataPath_RF_bus_sel_savedwin_data_8_port, 
                           curr_proc_regs(7) => 
                           DataPath_RF_bus_sel_savedwin_data_7_port, 
                           curr_proc_regs(6) => 
                           DataPath_RF_bus_sel_savedwin_data_6_port, 
                           curr_proc_regs(5) => 
                           DataPath_RF_bus_sel_savedwin_data_5_port, 
                           curr_proc_regs(4) => 
                           DataPath_RF_bus_sel_savedwin_data_4_port, 
                           curr_proc_regs(3) => 
                           DataPath_RF_bus_sel_savedwin_data_3_port, 
                           curr_proc_regs(2) => 
                           DataPath_RF_bus_sel_savedwin_data_2_port, 
                           curr_proc_regs(1) => 
                           DataPath_RF_bus_sel_savedwin_data_1_port, 
                           curr_proc_regs(0) => 
                           DataPath_RF_bus_sel_savedwin_data_0_port);
   DataPath_RF_RDPORT1 : mux_N32_M5_1 port map( S(4) => i_ADD_RS2_4_port, S(3) 
                           => i_ADD_RS2_3_port, S(2) => i_ADD_RS2_2_port, S(1) 
                           => i_ADD_RS2_1_port, S(0) => i_ADD_RS2_0_port, 
                           Q(1023) => 
                           DataPath_RF_bus_selected_win_data_767_port, Q(1022) 
                           => DataPath_RF_bus_selected_win_data_766_port, 
                           Q(1021) => 
                           DataPath_RF_bus_selected_win_data_765_port, Q(1020) 
                           => DataPath_RF_bus_selected_win_data_764_port, 
                           Q(1019) => 
                           DataPath_RF_bus_selected_win_data_763_port, Q(1018) 
                           => DataPath_RF_bus_selected_win_data_762_port, 
                           Q(1017) => 
                           DataPath_RF_bus_selected_win_data_761_port, Q(1016) 
                           => DataPath_RF_bus_selected_win_data_760_port, 
                           Q(1015) => 
                           DataPath_RF_bus_selected_win_data_759_port, Q(1014) 
                           => DataPath_RF_bus_selected_win_data_758_port, 
                           Q(1013) => 
                           DataPath_RF_bus_selected_win_data_757_port, Q(1012) 
                           => DataPath_RF_bus_selected_win_data_756_port, 
                           Q(1011) => 
                           DataPath_RF_bus_selected_win_data_755_port, Q(1010) 
                           => DataPath_RF_bus_selected_win_data_754_port, 
                           Q(1009) => 
                           DataPath_RF_bus_selected_win_data_753_port, Q(1008) 
                           => DataPath_RF_bus_selected_win_data_752_port, 
                           Q(1007) => 
                           DataPath_RF_bus_selected_win_data_751_port, Q(1006) 
                           => DataPath_RF_bus_selected_win_data_750_port, 
                           Q(1005) => 
                           DataPath_RF_bus_selected_win_data_749_port, Q(1004) 
                           => DataPath_RF_bus_selected_win_data_748_port, 
                           Q(1003) => 
                           DataPath_RF_bus_selected_win_data_747_port, Q(1002) 
                           => DataPath_RF_bus_selected_win_data_746_port, 
                           Q(1001) => 
                           DataPath_RF_bus_selected_win_data_745_port, Q(1000) 
                           => DataPath_RF_bus_selected_win_data_744_port, 
                           Q(999) => DataPath_RF_bus_selected_win_data_743_port
                           , Q(998) => 
                           DataPath_RF_bus_selected_win_data_742_port, Q(997) 
                           => DataPath_RF_bus_selected_win_data_741_port, 
                           Q(996) => DataPath_RF_bus_selected_win_data_740_port
                           , Q(995) => 
                           DataPath_RF_bus_selected_win_data_739_port, Q(994) 
                           => DataPath_RF_bus_selected_win_data_738_port, 
                           Q(993) => DataPath_RF_bus_selected_win_data_737_port
                           , Q(992) => 
                           DataPath_RF_bus_selected_win_data_736_port, Q(991) 
                           => DataPath_RF_bus_selected_win_data_735_port, 
                           Q(990) => DataPath_RF_bus_selected_win_data_734_port
                           , Q(989) => 
                           DataPath_RF_bus_selected_win_data_733_port, Q(988) 
                           => DataPath_RF_bus_selected_win_data_732_port, 
                           Q(987) => DataPath_RF_bus_selected_win_data_731_port
                           , Q(986) => 
                           DataPath_RF_bus_selected_win_data_730_port, Q(985) 
                           => DataPath_RF_bus_selected_win_data_729_port, 
                           Q(984) => DataPath_RF_bus_selected_win_data_728_port
                           , Q(983) => 
                           DataPath_RF_bus_selected_win_data_727_port, Q(982) 
                           => DataPath_RF_bus_selected_win_data_726_port, 
                           Q(981) => DataPath_RF_bus_selected_win_data_725_port
                           , Q(980) => 
                           DataPath_RF_bus_selected_win_data_724_port, Q(979) 
                           => DataPath_RF_bus_selected_win_data_723_port, 
                           Q(978) => DataPath_RF_bus_selected_win_data_722_port
                           , Q(977) => 
                           DataPath_RF_bus_selected_win_data_721_port, Q(976) 
                           => DataPath_RF_bus_selected_win_data_720_port, 
                           Q(975) => DataPath_RF_bus_selected_win_data_719_port
                           , Q(974) => 
                           DataPath_RF_bus_selected_win_data_718_port, Q(973) 
                           => DataPath_RF_bus_selected_win_data_717_port, 
                           Q(972) => DataPath_RF_bus_selected_win_data_716_port
                           , Q(971) => 
                           DataPath_RF_bus_selected_win_data_715_port, Q(970) 
                           => DataPath_RF_bus_selected_win_data_714_port, 
                           Q(969) => DataPath_RF_bus_selected_win_data_713_port
                           , Q(968) => 
                           DataPath_RF_bus_selected_win_data_712_port, Q(967) 
                           => DataPath_RF_bus_selected_win_data_711_port, 
                           Q(966) => DataPath_RF_bus_selected_win_data_710_port
                           , Q(965) => 
                           DataPath_RF_bus_selected_win_data_709_port, Q(964) 
                           => DataPath_RF_bus_selected_win_data_708_port, 
                           Q(963) => DataPath_RF_bus_selected_win_data_707_port
                           , Q(962) => 
                           DataPath_RF_bus_selected_win_data_706_port, Q(961) 
                           => DataPath_RF_bus_selected_win_data_705_port, 
                           Q(960) => DataPath_RF_bus_selected_win_data_704_port
                           , Q(959) => 
                           DataPath_RF_bus_selected_win_data_703_port, Q(958) 
                           => DataPath_RF_bus_selected_win_data_702_port, 
                           Q(957) => DataPath_RF_bus_selected_win_data_701_port
                           , Q(956) => 
                           DataPath_RF_bus_selected_win_data_700_port, Q(955) 
                           => DataPath_RF_bus_selected_win_data_699_port, 
                           Q(954) => DataPath_RF_bus_selected_win_data_698_port
                           , Q(953) => 
                           DataPath_RF_bus_selected_win_data_697_port, Q(952) 
                           => DataPath_RF_bus_selected_win_data_696_port, 
                           Q(951) => DataPath_RF_bus_selected_win_data_695_port
                           , Q(950) => 
                           DataPath_RF_bus_selected_win_data_694_port, Q(949) 
                           => DataPath_RF_bus_selected_win_data_693_port, 
                           Q(948) => DataPath_RF_bus_selected_win_data_692_port
                           , Q(947) => 
                           DataPath_RF_bus_selected_win_data_691_port, Q(946) 
                           => DataPath_RF_bus_selected_win_data_690_port, 
                           Q(945) => DataPath_RF_bus_selected_win_data_689_port
                           , Q(944) => 
                           DataPath_RF_bus_selected_win_data_688_port, Q(943) 
                           => DataPath_RF_bus_selected_win_data_687_port, 
                           Q(942) => DataPath_RF_bus_selected_win_data_686_port
                           , Q(941) => 
                           DataPath_RF_bus_selected_win_data_685_port, Q(940) 
                           => DataPath_RF_bus_selected_win_data_684_port, 
                           Q(939) => DataPath_RF_bus_selected_win_data_683_port
                           , Q(938) => 
                           DataPath_RF_bus_selected_win_data_682_port, Q(937) 
                           => DataPath_RF_bus_selected_win_data_681_port, 
                           Q(936) => DataPath_RF_bus_selected_win_data_680_port
                           , Q(935) => 
                           DataPath_RF_bus_selected_win_data_679_port, Q(934) 
                           => DataPath_RF_bus_selected_win_data_678_port, 
                           Q(933) => DataPath_RF_bus_selected_win_data_677_port
                           , Q(932) => 
                           DataPath_RF_bus_selected_win_data_676_port, Q(931) 
                           => DataPath_RF_bus_selected_win_data_675_port, 
                           Q(930) => DataPath_RF_bus_selected_win_data_674_port
                           , Q(929) => 
                           DataPath_RF_bus_selected_win_data_673_port, Q(928) 
                           => DataPath_RF_bus_selected_win_data_672_port, 
                           Q(927) => DataPath_RF_bus_selected_win_data_671_port
                           , Q(926) => 
                           DataPath_RF_bus_selected_win_data_670_port, Q(925) 
                           => DataPath_RF_bus_selected_win_data_669_port, 
                           Q(924) => DataPath_RF_bus_selected_win_data_668_port
                           , Q(923) => 
                           DataPath_RF_bus_selected_win_data_667_port, Q(922) 
                           => DataPath_RF_bus_selected_win_data_666_port, 
                           Q(921) => DataPath_RF_bus_selected_win_data_665_port
                           , Q(920) => 
                           DataPath_RF_bus_selected_win_data_664_port, Q(919) 
                           => DataPath_RF_bus_selected_win_data_663_port, 
                           Q(918) => DataPath_RF_bus_selected_win_data_662_port
                           , Q(917) => 
                           DataPath_RF_bus_selected_win_data_661_port, Q(916) 
                           => DataPath_RF_bus_selected_win_data_660_port, 
                           Q(915) => DataPath_RF_bus_selected_win_data_659_port
                           , Q(914) => 
                           DataPath_RF_bus_selected_win_data_658_port, Q(913) 
                           => DataPath_RF_bus_selected_win_data_657_port, 
                           Q(912) => DataPath_RF_bus_selected_win_data_656_port
                           , Q(911) => 
                           DataPath_RF_bus_selected_win_data_655_port, Q(910) 
                           => DataPath_RF_bus_selected_win_data_654_port, 
                           Q(909) => DataPath_RF_bus_selected_win_data_653_port
                           , Q(908) => 
                           DataPath_RF_bus_selected_win_data_652_port, Q(907) 
                           => DataPath_RF_bus_selected_win_data_651_port, 
                           Q(906) => DataPath_RF_bus_selected_win_data_650_port
                           , Q(905) => 
                           DataPath_RF_bus_selected_win_data_649_port, Q(904) 
                           => DataPath_RF_bus_selected_win_data_648_port, 
                           Q(903) => DataPath_RF_bus_selected_win_data_647_port
                           , Q(902) => 
                           DataPath_RF_bus_selected_win_data_646_port, Q(901) 
                           => DataPath_RF_bus_selected_win_data_645_port, 
                           Q(900) => DataPath_RF_bus_selected_win_data_644_port
                           , Q(899) => 
                           DataPath_RF_bus_selected_win_data_643_port, Q(898) 
                           => DataPath_RF_bus_selected_win_data_642_port, 
                           Q(897) => DataPath_RF_bus_selected_win_data_641_port
                           , Q(896) => 
                           DataPath_RF_bus_selected_win_data_640_port, Q(895) 
                           => DataPath_RF_bus_selected_win_data_639_port, 
                           Q(894) => DataPath_RF_bus_selected_win_data_638_port
                           , Q(893) => 
                           DataPath_RF_bus_selected_win_data_637_port, Q(892) 
                           => DataPath_RF_bus_selected_win_data_636_port, 
                           Q(891) => DataPath_RF_bus_selected_win_data_635_port
                           , Q(890) => 
                           DataPath_RF_bus_selected_win_data_634_port, Q(889) 
                           => DataPath_RF_bus_selected_win_data_633_port, 
                           Q(888) => DataPath_RF_bus_selected_win_data_632_port
                           , Q(887) => 
                           DataPath_RF_bus_selected_win_data_631_port, Q(886) 
                           => DataPath_RF_bus_selected_win_data_630_port, 
                           Q(885) => DataPath_RF_bus_selected_win_data_629_port
                           , Q(884) => 
                           DataPath_RF_bus_selected_win_data_628_port, Q(883) 
                           => DataPath_RF_bus_selected_win_data_627_port, 
                           Q(882) => DataPath_RF_bus_selected_win_data_626_port
                           , Q(881) => 
                           DataPath_RF_bus_selected_win_data_625_port, Q(880) 
                           => DataPath_RF_bus_selected_win_data_624_port, 
                           Q(879) => DataPath_RF_bus_selected_win_data_623_port
                           , Q(878) => 
                           DataPath_RF_bus_selected_win_data_622_port, Q(877) 
                           => DataPath_RF_bus_selected_win_data_621_port, 
                           Q(876) => DataPath_RF_bus_selected_win_data_620_port
                           , Q(875) => 
                           DataPath_RF_bus_selected_win_data_619_port, Q(874) 
                           => DataPath_RF_bus_selected_win_data_618_port, 
                           Q(873) => DataPath_RF_bus_selected_win_data_617_port
                           , Q(872) => 
                           DataPath_RF_bus_selected_win_data_616_port, Q(871) 
                           => DataPath_RF_bus_selected_win_data_615_port, 
                           Q(870) => DataPath_RF_bus_selected_win_data_614_port
                           , Q(869) => 
                           DataPath_RF_bus_selected_win_data_613_port, Q(868) 
                           => DataPath_RF_bus_selected_win_data_612_port, 
                           Q(867) => DataPath_RF_bus_selected_win_data_611_port
                           , Q(866) => 
                           DataPath_RF_bus_selected_win_data_610_port, Q(865) 
                           => DataPath_RF_bus_selected_win_data_609_port, 
                           Q(864) => DataPath_RF_bus_selected_win_data_608_port
                           , Q(863) => 
                           DataPath_RF_bus_selected_win_data_607_port, Q(862) 
                           => DataPath_RF_bus_selected_win_data_606_port, 
                           Q(861) => DataPath_RF_bus_selected_win_data_605_port
                           , Q(860) => 
                           DataPath_RF_bus_selected_win_data_604_port, Q(859) 
                           => DataPath_RF_bus_selected_win_data_603_port, 
                           Q(858) => DataPath_RF_bus_selected_win_data_602_port
                           , Q(857) => 
                           DataPath_RF_bus_selected_win_data_601_port, Q(856) 
                           => DataPath_RF_bus_selected_win_data_600_port, 
                           Q(855) => DataPath_RF_bus_selected_win_data_599_port
                           , Q(854) => 
                           DataPath_RF_bus_selected_win_data_598_port, Q(853) 
                           => DataPath_RF_bus_selected_win_data_597_port, 
                           Q(852) => DataPath_RF_bus_selected_win_data_596_port
                           , Q(851) => 
                           DataPath_RF_bus_selected_win_data_595_port, Q(850) 
                           => DataPath_RF_bus_selected_win_data_594_port, 
                           Q(849) => DataPath_RF_bus_selected_win_data_593_port
                           , Q(848) => 
                           DataPath_RF_bus_selected_win_data_592_port, Q(847) 
                           => DataPath_RF_bus_selected_win_data_591_port, 
                           Q(846) => DataPath_RF_bus_selected_win_data_590_port
                           , Q(845) => 
                           DataPath_RF_bus_selected_win_data_589_port, Q(844) 
                           => DataPath_RF_bus_selected_win_data_588_port, 
                           Q(843) => DataPath_RF_bus_selected_win_data_587_port
                           , Q(842) => 
                           DataPath_RF_bus_selected_win_data_586_port, Q(841) 
                           => DataPath_RF_bus_selected_win_data_585_port, 
                           Q(840) => DataPath_RF_bus_selected_win_data_584_port
                           , Q(839) => 
                           DataPath_RF_bus_selected_win_data_583_port, Q(838) 
                           => DataPath_RF_bus_selected_win_data_582_port, 
                           Q(837) => DataPath_RF_bus_selected_win_data_581_port
                           , Q(836) => 
                           DataPath_RF_bus_selected_win_data_580_port, Q(835) 
                           => DataPath_RF_bus_selected_win_data_579_port, 
                           Q(834) => DataPath_RF_bus_selected_win_data_578_port
                           , Q(833) => 
                           DataPath_RF_bus_selected_win_data_577_port, Q(832) 
                           => DataPath_RF_bus_selected_win_data_576_port, 
                           Q(831) => DataPath_RF_bus_selected_win_data_575_port
                           , Q(830) => 
                           DataPath_RF_bus_selected_win_data_574_port, Q(829) 
                           => DataPath_RF_bus_selected_win_data_573_port, 
                           Q(828) => DataPath_RF_bus_selected_win_data_572_port
                           , Q(827) => 
                           DataPath_RF_bus_selected_win_data_571_port, Q(826) 
                           => DataPath_RF_bus_selected_win_data_570_port, 
                           Q(825) => DataPath_RF_bus_selected_win_data_569_port
                           , Q(824) => 
                           DataPath_RF_bus_selected_win_data_568_port, Q(823) 
                           => DataPath_RF_bus_selected_win_data_567_port, 
                           Q(822) => DataPath_RF_bus_selected_win_data_566_port
                           , Q(821) => 
                           DataPath_RF_bus_selected_win_data_565_port, Q(820) 
                           => DataPath_RF_bus_selected_win_data_564_port, 
                           Q(819) => DataPath_RF_bus_selected_win_data_563_port
                           , Q(818) => 
                           DataPath_RF_bus_selected_win_data_562_port, Q(817) 
                           => DataPath_RF_bus_selected_win_data_561_port, 
                           Q(816) => DataPath_RF_bus_selected_win_data_560_port
                           , Q(815) => 
                           DataPath_RF_bus_selected_win_data_559_port, Q(814) 
                           => DataPath_RF_bus_selected_win_data_558_port, 
                           Q(813) => DataPath_RF_bus_selected_win_data_557_port
                           , Q(812) => 
                           DataPath_RF_bus_selected_win_data_556_port, Q(811) 
                           => DataPath_RF_bus_selected_win_data_555_port, 
                           Q(810) => DataPath_RF_bus_selected_win_data_554_port
                           , Q(809) => 
                           DataPath_RF_bus_selected_win_data_553_port, Q(808) 
                           => DataPath_RF_bus_selected_win_data_552_port, 
                           Q(807) => DataPath_RF_bus_selected_win_data_551_port
                           , Q(806) => 
                           DataPath_RF_bus_selected_win_data_550_port, Q(805) 
                           => DataPath_RF_bus_selected_win_data_549_port, 
                           Q(804) => DataPath_RF_bus_selected_win_data_548_port
                           , Q(803) => 
                           DataPath_RF_bus_selected_win_data_547_port, Q(802) 
                           => DataPath_RF_bus_selected_win_data_546_port, 
                           Q(801) => DataPath_RF_bus_selected_win_data_545_port
                           , Q(800) => 
                           DataPath_RF_bus_selected_win_data_544_port, Q(799) 
                           => DataPath_RF_bus_selected_win_data_543_port, 
                           Q(798) => DataPath_RF_bus_selected_win_data_542_port
                           , Q(797) => 
                           DataPath_RF_bus_selected_win_data_541_port, Q(796) 
                           => DataPath_RF_bus_selected_win_data_540_port, 
                           Q(795) => DataPath_RF_bus_selected_win_data_539_port
                           , Q(794) => 
                           DataPath_RF_bus_selected_win_data_538_port, Q(793) 
                           => DataPath_RF_bus_selected_win_data_537_port, 
                           Q(792) => DataPath_RF_bus_selected_win_data_536_port
                           , Q(791) => 
                           DataPath_RF_bus_selected_win_data_535_port, Q(790) 
                           => DataPath_RF_bus_selected_win_data_534_port, 
                           Q(789) => DataPath_RF_bus_selected_win_data_533_port
                           , Q(788) => 
                           DataPath_RF_bus_selected_win_data_532_port, Q(787) 
                           => DataPath_RF_bus_selected_win_data_531_port, 
                           Q(786) => DataPath_RF_bus_selected_win_data_530_port
                           , Q(785) => 
                           DataPath_RF_bus_selected_win_data_529_port, Q(784) 
                           => DataPath_RF_bus_selected_win_data_528_port, 
                           Q(783) => DataPath_RF_bus_selected_win_data_527_port
                           , Q(782) => 
                           DataPath_RF_bus_selected_win_data_526_port, Q(781) 
                           => DataPath_RF_bus_selected_win_data_525_port, 
                           Q(780) => DataPath_RF_bus_selected_win_data_524_port
                           , Q(779) => 
                           DataPath_RF_bus_selected_win_data_523_port, Q(778) 
                           => DataPath_RF_bus_selected_win_data_522_port, 
                           Q(777) => DataPath_RF_bus_selected_win_data_521_port
                           , Q(776) => 
                           DataPath_RF_bus_selected_win_data_520_port, Q(775) 
                           => DataPath_RF_bus_selected_win_data_519_port, 
                           Q(774) => DataPath_RF_bus_selected_win_data_518_port
                           , Q(773) => 
                           DataPath_RF_bus_selected_win_data_517_port, Q(772) 
                           => DataPath_RF_bus_selected_win_data_516_port, 
                           Q(771) => DataPath_RF_bus_selected_win_data_515_port
                           , Q(770) => 
                           DataPath_RF_bus_selected_win_data_514_port, Q(769) 
                           => DataPath_RF_bus_selected_win_data_513_port, 
                           Q(768) => DataPath_RF_bus_selected_win_data_512_port
                           , Q(767) => 
                           DataPath_RF_bus_selected_win_data_511_port, Q(766) 
                           => DataPath_RF_bus_selected_win_data_510_port, 
                           Q(765) => DataPath_RF_bus_selected_win_data_509_port
                           , Q(764) => 
                           DataPath_RF_bus_selected_win_data_508_port, Q(763) 
                           => DataPath_RF_bus_selected_win_data_507_port, 
                           Q(762) => DataPath_RF_bus_selected_win_data_506_port
                           , Q(761) => 
                           DataPath_RF_bus_selected_win_data_505_port, Q(760) 
                           => DataPath_RF_bus_selected_win_data_504_port, 
                           Q(759) => DataPath_RF_bus_selected_win_data_503_port
                           , Q(758) => 
                           DataPath_RF_bus_selected_win_data_502_port, Q(757) 
                           => DataPath_RF_bus_selected_win_data_501_port, 
                           Q(756) => DataPath_RF_bus_selected_win_data_500_port
                           , Q(755) => 
                           DataPath_RF_bus_selected_win_data_499_port, Q(754) 
                           => DataPath_RF_bus_selected_win_data_498_port, 
                           Q(753) => DataPath_RF_bus_selected_win_data_497_port
                           , Q(752) => 
                           DataPath_RF_bus_selected_win_data_496_port, Q(751) 
                           => DataPath_RF_bus_selected_win_data_495_port, 
                           Q(750) => DataPath_RF_bus_selected_win_data_494_port
                           , Q(749) => 
                           DataPath_RF_bus_selected_win_data_493_port, Q(748) 
                           => DataPath_RF_bus_selected_win_data_492_port, 
                           Q(747) => DataPath_RF_bus_selected_win_data_491_port
                           , Q(746) => 
                           DataPath_RF_bus_selected_win_data_490_port, Q(745) 
                           => DataPath_RF_bus_selected_win_data_489_port, 
                           Q(744) => DataPath_RF_bus_selected_win_data_488_port
                           , Q(743) => 
                           DataPath_RF_bus_selected_win_data_487_port, Q(742) 
                           => DataPath_RF_bus_selected_win_data_486_port, 
                           Q(741) => DataPath_RF_bus_selected_win_data_485_port
                           , Q(740) => 
                           DataPath_RF_bus_selected_win_data_484_port, Q(739) 
                           => DataPath_RF_bus_selected_win_data_483_port, 
                           Q(738) => DataPath_RF_bus_selected_win_data_482_port
                           , Q(737) => 
                           DataPath_RF_bus_selected_win_data_481_port, Q(736) 
                           => DataPath_RF_bus_selected_win_data_480_port, 
                           Q(735) => DataPath_RF_bus_selected_win_data_479_port
                           , Q(734) => 
                           DataPath_RF_bus_selected_win_data_478_port, Q(733) 
                           => DataPath_RF_bus_selected_win_data_477_port, 
                           Q(732) => DataPath_RF_bus_selected_win_data_476_port
                           , Q(731) => 
                           DataPath_RF_bus_selected_win_data_475_port, Q(730) 
                           => DataPath_RF_bus_selected_win_data_474_port, 
                           Q(729) => DataPath_RF_bus_selected_win_data_473_port
                           , Q(728) => 
                           DataPath_RF_bus_selected_win_data_472_port, Q(727) 
                           => DataPath_RF_bus_selected_win_data_471_port, 
                           Q(726) => DataPath_RF_bus_selected_win_data_470_port
                           , Q(725) => 
                           DataPath_RF_bus_selected_win_data_469_port, Q(724) 
                           => DataPath_RF_bus_selected_win_data_468_port, 
                           Q(723) => DataPath_RF_bus_selected_win_data_467_port
                           , Q(722) => 
                           DataPath_RF_bus_selected_win_data_466_port, Q(721) 
                           => DataPath_RF_bus_selected_win_data_465_port, 
                           Q(720) => DataPath_RF_bus_selected_win_data_464_port
                           , Q(719) => 
                           DataPath_RF_bus_selected_win_data_463_port, Q(718) 
                           => DataPath_RF_bus_selected_win_data_462_port, 
                           Q(717) => DataPath_RF_bus_selected_win_data_461_port
                           , Q(716) => 
                           DataPath_RF_bus_selected_win_data_460_port, Q(715) 
                           => DataPath_RF_bus_selected_win_data_459_port, 
                           Q(714) => DataPath_RF_bus_selected_win_data_458_port
                           , Q(713) => 
                           DataPath_RF_bus_selected_win_data_457_port, Q(712) 
                           => DataPath_RF_bus_selected_win_data_456_port, 
                           Q(711) => DataPath_RF_bus_selected_win_data_455_port
                           , Q(710) => 
                           DataPath_RF_bus_selected_win_data_454_port, Q(709) 
                           => DataPath_RF_bus_selected_win_data_453_port, 
                           Q(708) => DataPath_RF_bus_selected_win_data_452_port
                           , Q(707) => 
                           DataPath_RF_bus_selected_win_data_451_port, Q(706) 
                           => DataPath_RF_bus_selected_win_data_450_port, 
                           Q(705) => DataPath_RF_bus_selected_win_data_449_port
                           , Q(704) => 
                           DataPath_RF_bus_selected_win_data_448_port, Q(703) 
                           => DataPath_RF_bus_selected_win_data_447_port, 
                           Q(702) => DataPath_RF_bus_selected_win_data_446_port
                           , Q(701) => 
                           DataPath_RF_bus_selected_win_data_445_port, Q(700) 
                           => DataPath_RF_bus_selected_win_data_444_port, 
                           Q(699) => DataPath_RF_bus_selected_win_data_443_port
                           , Q(698) => 
                           DataPath_RF_bus_selected_win_data_442_port, Q(697) 
                           => DataPath_RF_bus_selected_win_data_441_port, 
                           Q(696) => DataPath_RF_bus_selected_win_data_440_port
                           , Q(695) => 
                           DataPath_RF_bus_selected_win_data_439_port, Q(694) 
                           => DataPath_RF_bus_selected_win_data_438_port, 
                           Q(693) => DataPath_RF_bus_selected_win_data_437_port
                           , Q(692) => 
                           DataPath_RF_bus_selected_win_data_436_port, Q(691) 
                           => DataPath_RF_bus_selected_win_data_435_port, 
                           Q(690) => DataPath_RF_bus_selected_win_data_434_port
                           , Q(689) => 
                           DataPath_RF_bus_selected_win_data_433_port, Q(688) 
                           => DataPath_RF_bus_selected_win_data_432_port, 
                           Q(687) => DataPath_RF_bus_selected_win_data_431_port
                           , Q(686) => 
                           DataPath_RF_bus_selected_win_data_430_port, Q(685) 
                           => DataPath_RF_bus_selected_win_data_429_port, 
                           Q(684) => DataPath_RF_bus_selected_win_data_428_port
                           , Q(683) => 
                           DataPath_RF_bus_selected_win_data_427_port, Q(682) 
                           => DataPath_RF_bus_selected_win_data_426_port, 
                           Q(681) => DataPath_RF_bus_selected_win_data_425_port
                           , Q(680) => 
                           DataPath_RF_bus_selected_win_data_424_port, Q(679) 
                           => DataPath_RF_bus_selected_win_data_423_port, 
                           Q(678) => DataPath_RF_bus_selected_win_data_422_port
                           , Q(677) => 
                           DataPath_RF_bus_selected_win_data_421_port, Q(676) 
                           => DataPath_RF_bus_selected_win_data_420_port, 
                           Q(675) => DataPath_RF_bus_selected_win_data_419_port
                           , Q(674) => 
                           DataPath_RF_bus_selected_win_data_418_port, Q(673) 
                           => DataPath_RF_bus_selected_win_data_417_port, 
                           Q(672) => DataPath_RF_bus_selected_win_data_416_port
                           , Q(671) => 
                           DataPath_RF_bus_selected_win_data_415_port, Q(670) 
                           => DataPath_RF_bus_selected_win_data_414_port, 
                           Q(669) => DataPath_RF_bus_selected_win_data_413_port
                           , Q(668) => 
                           DataPath_RF_bus_selected_win_data_412_port, Q(667) 
                           => DataPath_RF_bus_selected_win_data_411_port, 
                           Q(666) => DataPath_RF_bus_selected_win_data_410_port
                           , Q(665) => 
                           DataPath_RF_bus_selected_win_data_409_port, Q(664) 
                           => DataPath_RF_bus_selected_win_data_408_port, 
                           Q(663) => DataPath_RF_bus_selected_win_data_407_port
                           , Q(662) => 
                           DataPath_RF_bus_selected_win_data_406_port, Q(661) 
                           => DataPath_RF_bus_selected_win_data_405_port, 
                           Q(660) => DataPath_RF_bus_selected_win_data_404_port
                           , Q(659) => 
                           DataPath_RF_bus_selected_win_data_403_port, Q(658) 
                           => DataPath_RF_bus_selected_win_data_402_port, 
                           Q(657) => DataPath_RF_bus_selected_win_data_401_port
                           , Q(656) => 
                           DataPath_RF_bus_selected_win_data_400_port, Q(655) 
                           => DataPath_RF_bus_selected_win_data_399_port, 
                           Q(654) => DataPath_RF_bus_selected_win_data_398_port
                           , Q(653) => 
                           DataPath_RF_bus_selected_win_data_397_port, Q(652) 
                           => DataPath_RF_bus_selected_win_data_396_port, 
                           Q(651) => DataPath_RF_bus_selected_win_data_395_port
                           , Q(650) => 
                           DataPath_RF_bus_selected_win_data_394_port, Q(649) 
                           => DataPath_RF_bus_selected_win_data_393_port, 
                           Q(648) => DataPath_RF_bus_selected_win_data_392_port
                           , Q(647) => 
                           DataPath_RF_bus_selected_win_data_391_port, Q(646) 
                           => DataPath_RF_bus_selected_win_data_390_port, 
                           Q(645) => DataPath_RF_bus_selected_win_data_389_port
                           , Q(644) => 
                           DataPath_RF_bus_selected_win_data_388_port, Q(643) 
                           => DataPath_RF_bus_selected_win_data_387_port, 
                           Q(642) => DataPath_RF_bus_selected_win_data_386_port
                           , Q(641) => 
                           DataPath_RF_bus_selected_win_data_385_port, Q(640) 
                           => DataPath_RF_bus_selected_win_data_384_port, 
                           Q(639) => DataPath_RF_bus_selected_win_data_383_port
                           , Q(638) => 
                           DataPath_RF_bus_selected_win_data_382_port, Q(637) 
                           => DataPath_RF_bus_selected_win_data_381_port, 
                           Q(636) => DataPath_RF_bus_selected_win_data_380_port
                           , Q(635) => 
                           DataPath_RF_bus_selected_win_data_379_port, Q(634) 
                           => DataPath_RF_bus_selected_win_data_378_port, 
                           Q(633) => DataPath_RF_bus_selected_win_data_377_port
                           , Q(632) => 
                           DataPath_RF_bus_selected_win_data_376_port, Q(631) 
                           => DataPath_RF_bus_selected_win_data_375_port, 
                           Q(630) => DataPath_RF_bus_selected_win_data_374_port
                           , Q(629) => 
                           DataPath_RF_bus_selected_win_data_373_port, Q(628) 
                           => DataPath_RF_bus_selected_win_data_372_port, 
                           Q(627) => DataPath_RF_bus_selected_win_data_371_port
                           , Q(626) => 
                           DataPath_RF_bus_selected_win_data_370_port, Q(625) 
                           => DataPath_RF_bus_selected_win_data_369_port, 
                           Q(624) => DataPath_RF_bus_selected_win_data_368_port
                           , Q(623) => 
                           DataPath_RF_bus_selected_win_data_367_port, Q(622) 
                           => DataPath_RF_bus_selected_win_data_366_port, 
                           Q(621) => DataPath_RF_bus_selected_win_data_365_port
                           , Q(620) => 
                           DataPath_RF_bus_selected_win_data_364_port, Q(619) 
                           => DataPath_RF_bus_selected_win_data_363_port, 
                           Q(618) => DataPath_RF_bus_selected_win_data_362_port
                           , Q(617) => 
                           DataPath_RF_bus_selected_win_data_361_port, Q(616) 
                           => DataPath_RF_bus_selected_win_data_360_port, 
                           Q(615) => DataPath_RF_bus_selected_win_data_359_port
                           , Q(614) => 
                           DataPath_RF_bus_selected_win_data_358_port, Q(613) 
                           => DataPath_RF_bus_selected_win_data_357_port, 
                           Q(612) => DataPath_RF_bus_selected_win_data_356_port
                           , Q(611) => 
                           DataPath_RF_bus_selected_win_data_355_port, Q(610) 
                           => DataPath_RF_bus_selected_win_data_354_port, 
                           Q(609) => DataPath_RF_bus_selected_win_data_353_port
                           , Q(608) => 
                           DataPath_RF_bus_selected_win_data_352_port, Q(607) 
                           => DataPath_RF_bus_selected_win_data_351_port, 
                           Q(606) => DataPath_RF_bus_selected_win_data_350_port
                           , Q(605) => 
                           DataPath_RF_bus_selected_win_data_349_port, Q(604) 
                           => DataPath_RF_bus_selected_win_data_348_port, 
                           Q(603) => DataPath_RF_bus_selected_win_data_347_port
                           , Q(602) => 
                           DataPath_RF_bus_selected_win_data_346_port, Q(601) 
                           => DataPath_RF_bus_selected_win_data_345_port, 
                           Q(600) => DataPath_RF_bus_selected_win_data_344_port
                           , Q(599) => 
                           DataPath_RF_bus_selected_win_data_343_port, Q(598) 
                           => DataPath_RF_bus_selected_win_data_342_port, 
                           Q(597) => DataPath_RF_bus_selected_win_data_341_port
                           , Q(596) => 
                           DataPath_RF_bus_selected_win_data_340_port, Q(595) 
                           => DataPath_RF_bus_selected_win_data_339_port, 
                           Q(594) => DataPath_RF_bus_selected_win_data_338_port
                           , Q(593) => 
                           DataPath_RF_bus_selected_win_data_337_port, Q(592) 
                           => DataPath_RF_bus_selected_win_data_336_port, 
                           Q(591) => DataPath_RF_bus_selected_win_data_335_port
                           , Q(590) => 
                           DataPath_RF_bus_selected_win_data_334_port, Q(589) 
                           => DataPath_RF_bus_selected_win_data_333_port, 
                           Q(588) => DataPath_RF_bus_selected_win_data_332_port
                           , Q(587) => 
                           DataPath_RF_bus_selected_win_data_331_port, Q(586) 
                           => DataPath_RF_bus_selected_win_data_330_port, 
                           Q(585) => DataPath_RF_bus_selected_win_data_329_port
                           , Q(584) => 
                           DataPath_RF_bus_selected_win_data_328_port, Q(583) 
                           => DataPath_RF_bus_selected_win_data_327_port, 
                           Q(582) => DataPath_RF_bus_selected_win_data_326_port
                           , Q(581) => 
                           DataPath_RF_bus_selected_win_data_325_port, Q(580) 
                           => DataPath_RF_bus_selected_win_data_324_port, 
                           Q(579) => DataPath_RF_bus_selected_win_data_323_port
                           , Q(578) => 
                           DataPath_RF_bus_selected_win_data_322_port, Q(577) 
                           => DataPath_RF_bus_selected_win_data_321_port, 
                           Q(576) => DataPath_RF_bus_selected_win_data_320_port
                           , Q(575) => 
                           DataPath_RF_bus_selected_win_data_319_port, Q(574) 
                           => DataPath_RF_bus_selected_win_data_318_port, 
                           Q(573) => DataPath_RF_bus_selected_win_data_317_port
                           , Q(572) => 
                           DataPath_RF_bus_selected_win_data_316_port, Q(571) 
                           => DataPath_RF_bus_selected_win_data_315_port, 
                           Q(570) => DataPath_RF_bus_selected_win_data_314_port
                           , Q(569) => 
                           DataPath_RF_bus_selected_win_data_313_port, Q(568) 
                           => DataPath_RF_bus_selected_win_data_312_port, 
                           Q(567) => DataPath_RF_bus_selected_win_data_311_port
                           , Q(566) => 
                           DataPath_RF_bus_selected_win_data_310_port, Q(565) 
                           => DataPath_RF_bus_selected_win_data_309_port, 
                           Q(564) => DataPath_RF_bus_selected_win_data_308_port
                           , Q(563) => 
                           DataPath_RF_bus_selected_win_data_307_port, Q(562) 
                           => DataPath_RF_bus_selected_win_data_306_port, 
                           Q(561) => DataPath_RF_bus_selected_win_data_305_port
                           , Q(560) => 
                           DataPath_RF_bus_selected_win_data_304_port, Q(559) 
                           => DataPath_RF_bus_selected_win_data_303_port, 
                           Q(558) => DataPath_RF_bus_selected_win_data_302_port
                           , Q(557) => 
                           DataPath_RF_bus_selected_win_data_301_port, Q(556) 
                           => DataPath_RF_bus_selected_win_data_300_port, 
                           Q(555) => DataPath_RF_bus_selected_win_data_299_port
                           , Q(554) => 
                           DataPath_RF_bus_selected_win_data_298_port, Q(553) 
                           => DataPath_RF_bus_selected_win_data_297_port, 
                           Q(552) => DataPath_RF_bus_selected_win_data_296_port
                           , Q(551) => 
                           DataPath_RF_bus_selected_win_data_295_port, Q(550) 
                           => DataPath_RF_bus_selected_win_data_294_port, 
                           Q(549) => DataPath_RF_bus_selected_win_data_293_port
                           , Q(548) => 
                           DataPath_RF_bus_selected_win_data_292_port, Q(547) 
                           => DataPath_RF_bus_selected_win_data_291_port, 
                           Q(546) => DataPath_RF_bus_selected_win_data_290_port
                           , Q(545) => 
                           DataPath_RF_bus_selected_win_data_289_port, Q(544) 
                           => DataPath_RF_bus_selected_win_data_288_port, 
                           Q(543) => DataPath_RF_bus_selected_win_data_287_port
                           , Q(542) => 
                           DataPath_RF_bus_selected_win_data_286_port, Q(541) 
                           => DataPath_RF_bus_selected_win_data_285_port, 
                           Q(540) => DataPath_RF_bus_selected_win_data_284_port
                           , Q(539) => 
                           DataPath_RF_bus_selected_win_data_283_port, Q(538) 
                           => DataPath_RF_bus_selected_win_data_282_port, 
                           Q(537) => DataPath_RF_bus_selected_win_data_281_port
                           , Q(536) => 
                           DataPath_RF_bus_selected_win_data_280_port, Q(535) 
                           => DataPath_RF_bus_selected_win_data_279_port, 
                           Q(534) => DataPath_RF_bus_selected_win_data_278_port
                           , Q(533) => 
                           DataPath_RF_bus_selected_win_data_277_port, Q(532) 
                           => DataPath_RF_bus_selected_win_data_276_port, 
                           Q(531) => DataPath_RF_bus_selected_win_data_275_port
                           , Q(530) => 
                           DataPath_RF_bus_selected_win_data_274_port, Q(529) 
                           => DataPath_RF_bus_selected_win_data_273_port, 
                           Q(528) => DataPath_RF_bus_selected_win_data_272_port
                           , Q(527) => 
                           DataPath_RF_bus_selected_win_data_271_port, Q(526) 
                           => DataPath_RF_bus_selected_win_data_270_port, 
                           Q(525) => DataPath_RF_bus_selected_win_data_269_port
                           , Q(524) => 
                           DataPath_RF_bus_selected_win_data_268_port, Q(523) 
                           => DataPath_RF_bus_selected_win_data_267_port, 
                           Q(522) => DataPath_RF_bus_selected_win_data_266_port
                           , Q(521) => 
                           DataPath_RF_bus_selected_win_data_265_port, Q(520) 
                           => DataPath_RF_bus_selected_win_data_264_port, 
                           Q(519) => DataPath_RF_bus_selected_win_data_263_port
                           , Q(518) => 
                           DataPath_RF_bus_selected_win_data_262_port, Q(517) 
                           => DataPath_RF_bus_selected_win_data_261_port, 
                           Q(516) => DataPath_RF_bus_selected_win_data_260_port
                           , Q(515) => 
                           DataPath_RF_bus_selected_win_data_259_port, Q(514) 
                           => DataPath_RF_bus_selected_win_data_258_port, 
                           Q(513) => DataPath_RF_bus_selected_win_data_257_port
                           , Q(512) => 
                           DataPath_RF_bus_selected_win_data_256_port, Q(511) 
                           => DataPath_RF_bus_selected_win_data_255_port, 
                           Q(510) => DataPath_RF_bus_selected_win_data_254_port
                           , Q(509) => 
                           DataPath_RF_bus_selected_win_data_253_port, Q(508) 
                           => DataPath_RF_bus_selected_win_data_252_port, 
                           Q(507) => DataPath_RF_bus_selected_win_data_251_port
                           , Q(506) => 
                           DataPath_RF_bus_selected_win_data_250_port, Q(505) 
                           => DataPath_RF_bus_selected_win_data_249_port, 
                           Q(504) => DataPath_RF_bus_selected_win_data_248_port
                           , Q(503) => 
                           DataPath_RF_bus_selected_win_data_247_port, Q(502) 
                           => DataPath_RF_bus_selected_win_data_246_port, 
                           Q(501) => DataPath_RF_bus_selected_win_data_245_port
                           , Q(500) => 
                           DataPath_RF_bus_selected_win_data_244_port, Q(499) 
                           => DataPath_RF_bus_selected_win_data_243_port, 
                           Q(498) => DataPath_RF_bus_selected_win_data_242_port
                           , Q(497) => 
                           DataPath_RF_bus_selected_win_data_241_port, Q(496) 
                           => DataPath_RF_bus_selected_win_data_240_port, 
                           Q(495) => DataPath_RF_bus_selected_win_data_239_port
                           , Q(494) => 
                           DataPath_RF_bus_selected_win_data_238_port, Q(493) 
                           => DataPath_RF_bus_selected_win_data_237_port, 
                           Q(492) => DataPath_RF_bus_selected_win_data_236_port
                           , Q(491) => 
                           DataPath_RF_bus_selected_win_data_235_port, Q(490) 
                           => DataPath_RF_bus_selected_win_data_234_port, 
                           Q(489) => DataPath_RF_bus_selected_win_data_233_port
                           , Q(488) => 
                           DataPath_RF_bus_selected_win_data_232_port, Q(487) 
                           => DataPath_RF_bus_selected_win_data_231_port, 
                           Q(486) => DataPath_RF_bus_selected_win_data_230_port
                           , Q(485) => 
                           DataPath_RF_bus_selected_win_data_229_port, Q(484) 
                           => DataPath_RF_bus_selected_win_data_228_port, 
                           Q(483) => DataPath_RF_bus_selected_win_data_227_port
                           , Q(482) => 
                           DataPath_RF_bus_selected_win_data_226_port, Q(481) 
                           => DataPath_RF_bus_selected_win_data_225_port, 
                           Q(480) => DataPath_RF_bus_selected_win_data_224_port
                           , Q(479) => 
                           DataPath_RF_bus_selected_win_data_223_port, Q(478) 
                           => DataPath_RF_bus_selected_win_data_222_port, 
                           Q(477) => DataPath_RF_bus_selected_win_data_221_port
                           , Q(476) => 
                           DataPath_RF_bus_selected_win_data_220_port, Q(475) 
                           => DataPath_RF_bus_selected_win_data_219_port, 
                           Q(474) => DataPath_RF_bus_selected_win_data_218_port
                           , Q(473) => 
                           DataPath_RF_bus_selected_win_data_217_port, Q(472) 
                           => DataPath_RF_bus_selected_win_data_216_port, 
                           Q(471) => DataPath_RF_bus_selected_win_data_215_port
                           , Q(470) => 
                           DataPath_RF_bus_selected_win_data_214_port, Q(469) 
                           => DataPath_RF_bus_selected_win_data_213_port, 
                           Q(468) => DataPath_RF_bus_selected_win_data_212_port
                           , Q(467) => 
                           DataPath_RF_bus_selected_win_data_211_port, Q(466) 
                           => DataPath_RF_bus_selected_win_data_210_port, 
                           Q(465) => DataPath_RF_bus_selected_win_data_209_port
                           , Q(464) => 
                           DataPath_RF_bus_selected_win_data_208_port, Q(463) 
                           => DataPath_RF_bus_selected_win_data_207_port, 
                           Q(462) => DataPath_RF_bus_selected_win_data_206_port
                           , Q(461) => 
                           DataPath_RF_bus_selected_win_data_205_port, Q(460) 
                           => DataPath_RF_bus_selected_win_data_204_port, 
                           Q(459) => DataPath_RF_bus_selected_win_data_203_port
                           , Q(458) => 
                           DataPath_RF_bus_selected_win_data_202_port, Q(457) 
                           => DataPath_RF_bus_selected_win_data_201_port, 
                           Q(456) => DataPath_RF_bus_selected_win_data_200_port
                           , Q(455) => 
                           DataPath_RF_bus_selected_win_data_199_port, Q(454) 
                           => DataPath_RF_bus_selected_win_data_198_port, 
                           Q(453) => DataPath_RF_bus_selected_win_data_197_port
                           , Q(452) => 
                           DataPath_RF_bus_selected_win_data_196_port, Q(451) 
                           => DataPath_RF_bus_selected_win_data_195_port, 
                           Q(450) => DataPath_RF_bus_selected_win_data_194_port
                           , Q(449) => 
                           DataPath_RF_bus_selected_win_data_193_port, Q(448) 
                           => DataPath_RF_bus_selected_win_data_192_port, 
                           Q(447) => DataPath_RF_bus_selected_win_data_191_port
                           , Q(446) => 
                           DataPath_RF_bus_selected_win_data_190_port, Q(445) 
                           => DataPath_RF_bus_selected_win_data_189_port, 
                           Q(444) => DataPath_RF_bus_selected_win_data_188_port
                           , Q(443) => 
                           DataPath_RF_bus_selected_win_data_187_port, Q(442) 
                           => DataPath_RF_bus_selected_win_data_186_port, 
                           Q(441) => DataPath_RF_bus_selected_win_data_185_port
                           , Q(440) => 
                           DataPath_RF_bus_selected_win_data_184_port, Q(439) 
                           => DataPath_RF_bus_selected_win_data_183_port, 
                           Q(438) => DataPath_RF_bus_selected_win_data_182_port
                           , Q(437) => 
                           DataPath_RF_bus_selected_win_data_181_port, Q(436) 
                           => DataPath_RF_bus_selected_win_data_180_port, 
                           Q(435) => DataPath_RF_bus_selected_win_data_179_port
                           , Q(434) => 
                           DataPath_RF_bus_selected_win_data_178_port, Q(433) 
                           => DataPath_RF_bus_selected_win_data_177_port, 
                           Q(432) => DataPath_RF_bus_selected_win_data_176_port
                           , Q(431) => 
                           DataPath_RF_bus_selected_win_data_175_port, Q(430) 
                           => DataPath_RF_bus_selected_win_data_174_port, 
                           Q(429) => DataPath_RF_bus_selected_win_data_173_port
                           , Q(428) => 
                           DataPath_RF_bus_selected_win_data_172_port, Q(427) 
                           => DataPath_RF_bus_selected_win_data_171_port, 
                           Q(426) => DataPath_RF_bus_selected_win_data_170_port
                           , Q(425) => 
                           DataPath_RF_bus_selected_win_data_169_port, Q(424) 
                           => DataPath_RF_bus_selected_win_data_168_port, 
                           Q(423) => DataPath_RF_bus_selected_win_data_167_port
                           , Q(422) => 
                           DataPath_RF_bus_selected_win_data_166_port, Q(421) 
                           => DataPath_RF_bus_selected_win_data_165_port, 
                           Q(420) => DataPath_RF_bus_selected_win_data_164_port
                           , Q(419) => 
                           DataPath_RF_bus_selected_win_data_163_port, Q(418) 
                           => DataPath_RF_bus_selected_win_data_162_port, 
                           Q(417) => DataPath_RF_bus_selected_win_data_161_port
                           , Q(416) => 
                           DataPath_RF_bus_selected_win_data_160_port, Q(415) 
                           => DataPath_RF_bus_selected_win_data_159_port, 
                           Q(414) => DataPath_RF_bus_selected_win_data_158_port
                           , Q(413) => 
                           DataPath_RF_bus_selected_win_data_157_port, Q(412) 
                           => DataPath_RF_bus_selected_win_data_156_port, 
                           Q(411) => DataPath_RF_bus_selected_win_data_155_port
                           , Q(410) => 
                           DataPath_RF_bus_selected_win_data_154_port, Q(409) 
                           => DataPath_RF_bus_selected_win_data_153_port, 
                           Q(408) => DataPath_RF_bus_selected_win_data_152_port
                           , Q(407) => 
                           DataPath_RF_bus_selected_win_data_151_port, Q(406) 
                           => DataPath_RF_bus_selected_win_data_150_port, 
                           Q(405) => DataPath_RF_bus_selected_win_data_149_port
                           , Q(404) => 
                           DataPath_RF_bus_selected_win_data_148_port, Q(403) 
                           => DataPath_RF_bus_selected_win_data_147_port, 
                           Q(402) => DataPath_RF_bus_selected_win_data_146_port
                           , Q(401) => 
                           DataPath_RF_bus_selected_win_data_145_port, Q(400) 
                           => DataPath_RF_bus_selected_win_data_144_port, 
                           Q(399) => DataPath_RF_bus_selected_win_data_143_port
                           , Q(398) => 
                           DataPath_RF_bus_selected_win_data_142_port, Q(397) 
                           => DataPath_RF_bus_selected_win_data_141_port, 
                           Q(396) => DataPath_RF_bus_selected_win_data_140_port
                           , Q(395) => 
                           DataPath_RF_bus_selected_win_data_139_port, Q(394) 
                           => DataPath_RF_bus_selected_win_data_138_port, 
                           Q(393) => DataPath_RF_bus_selected_win_data_137_port
                           , Q(392) => 
                           DataPath_RF_bus_selected_win_data_136_port, Q(391) 
                           => DataPath_RF_bus_selected_win_data_135_port, 
                           Q(390) => DataPath_RF_bus_selected_win_data_134_port
                           , Q(389) => 
                           DataPath_RF_bus_selected_win_data_133_port, Q(388) 
                           => DataPath_RF_bus_selected_win_data_132_port, 
                           Q(387) => DataPath_RF_bus_selected_win_data_131_port
                           , Q(386) => 
                           DataPath_RF_bus_selected_win_data_130_port, Q(385) 
                           => DataPath_RF_bus_selected_win_data_129_port, 
                           Q(384) => DataPath_RF_bus_selected_win_data_128_port
                           , Q(383) => 
                           DataPath_RF_bus_selected_win_data_127_port, Q(382) 
                           => DataPath_RF_bus_selected_win_data_126_port, 
                           Q(381) => DataPath_RF_bus_selected_win_data_125_port
                           , Q(380) => 
                           DataPath_RF_bus_selected_win_data_124_port, Q(379) 
                           => DataPath_RF_bus_selected_win_data_123_port, 
                           Q(378) => DataPath_RF_bus_selected_win_data_122_port
                           , Q(377) => 
                           DataPath_RF_bus_selected_win_data_121_port, Q(376) 
                           => DataPath_RF_bus_selected_win_data_120_port, 
                           Q(375) => DataPath_RF_bus_selected_win_data_119_port
                           , Q(374) => 
                           DataPath_RF_bus_selected_win_data_118_port, Q(373) 
                           => DataPath_RF_bus_selected_win_data_117_port, 
                           Q(372) => DataPath_RF_bus_selected_win_data_116_port
                           , Q(371) => 
                           DataPath_RF_bus_selected_win_data_115_port, Q(370) 
                           => DataPath_RF_bus_selected_win_data_114_port, 
                           Q(369) => DataPath_RF_bus_selected_win_data_113_port
                           , Q(368) => 
                           DataPath_RF_bus_selected_win_data_112_port, Q(367) 
                           => DataPath_RF_bus_selected_win_data_111_port, 
                           Q(366) => DataPath_RF_bus_selected_win_data_110_port
                           , Q(365) => 
                           DataPath_RF_bus_selected_win_data_109_port, Q(364) 
                           => DataPath_RF_bus_selected_win_data_108_port, 
                           Q(363) => DataPath_RF_bus_selected_win_data_107_port
                           , Q(362) => 
                           DataPath_RF_bus_selected_win_data_106_port, Q(361) 
                           => DataPath_RF_bus_selected_win_data_105_port, 
                           Q(360) => DataPath_RF_bus_selected_win_data_104_port
                           , Q(359) => 
                           DataPath_RF_bus_selected_win_data_103_port, Q(358) 
                           => DataPath_RF_bus_selected_win_data_102_port, 
                           Q(357) => DataPath_RF_bus_selected_win_data_101_port
                           , Q(356) => 
                           DataPath_RF_bus_selected_win_data_100_port, Q(355) 
                           => DataPath_RF_bus_selected_win_data_99_port, Q(354)
                           => DataPath_RF_bus_selected_win_data_98_port, Q(353)
                           => DataPath_RF_bus_selected_win_data_97_port, Q(352)
                           => DataPath_RF_bus_selected_win_data_96_port, Q(351)
                           => DataPath_RF_bus_selected_win_data_95_port, Q(350)
                           => DataPath_RF_bus_selected_win_data_94_port, Q(349)
                           => DataPath_RF_bus_selected_win_data_93_port, Q(348)
                           => DataPath_RF_bus_selected_win_data_92_port, Q(347)
                           => DataPath_RF_bus_selected_win_data_91_port, Q(346)
                           => DataPath_RF_bus_selected_win_data_90_port, Q(345)
                           => DataPath_RF_bus_selected_win_data_89_port, Q(344)
                           => DataPath_RF_bus_selected_win_data_88_port, Q(343)
                           => DataPath_RF_bus_selected_win_data_87_port, Q(342)
                           => DataPath_RF_bus_selected_win_data_86_port, Q(341)
                           => DataPath_RF_bus_selected_win_data_85_port, Q(340)
                           => DataPath_RF_bus_selected_win_data_84_port, Q(339)
                           => DataPath_RF_bus_selected_win_data_83_port, Q(338)
                           => DataPath_RF_bus_selected_win_data_82_port, Q(337)
                           => DataPath_RF_bus_selected_win_data_81_port, Q(336)
                           => DataPath_RF_bus_selected_win_data_80_port, Q(335)
                           => DataPath_RF_bus_selected_win_data_79_port, Q(334)
                           => DataPath_RF_bus_selected_win_data_78_port, Q(333)
                           => DataPath_RF_bus_selected_win_data_77_port, Q(332)
                           => DataPath_RF_bus_selected_win_data_76_port, Q(331)
                           => DataPath_RF_bus_selected_win_data_75_port, Q(330)
                           => DataPath_RF_bus_selected_win_data_74_port, Q(329)
                           => DataPath_RF_bus_selected_win_data_73_port, Q(328)
                           => DataPath_RF_bus_selected_win_data_72_port, Q(327)
                           => DataPath_RF_bus_selected_win_data_71_port, Q(326)
                           => DataPath_RF_bus_selected_win_data_70_port, Q(325)
                           => DataPath_RF_bus_selected_win_data_69_port, Q(324)
                           => DataPath_RF_bus_selected_win_data_68_port, Q(323)
                           => DataPath_RF_bus_selected_win_data_67_port, Q(322)
                           => DataPath_RF_bus_selected_win_data_66_port, Q(321)
                           => DataPath_RF_bus_selected_win_data_65_port, Q(320)
                           => DataPath_RF_bus_selected_win_data_64_port, Q(319)
                           => DataPath_RF_bus_selected_win_data_63_port, Q(318)
                           => DataPath_RF_bus_selected_win_data_62_port, Q(317)
                           => DataPath_RF_bus_selected_win_data_61_port, Q(316)
                           => DataPath_RF_bus_selected_win_data_60_port, Q(315)
                           => DataPath_RF_bus_selected_win_data_59_port, Q(314)
                           => DataPath_RF_bus_selected_win_data_58_port, Q(313)
                           => DataPath_RF_bus_selected_win_data_57_port, Q(312)
                           => DataPath_RF_bus_selected_win_data_56_port, Q(311)
                           => DataPath_RF_bus_selected_win_data_55_port, Q(310)
                           => DataPath_RF_bus_selected_win_data_54_port, Q(309)
                           => DataPath_RF_bus_selected_win_data_53_port, Q(308)
                           => DataPath_RF_bus_selected_win_data_52_port, Q(307)
                           => DataPath_RF_bus_selected_win_data_51_port, Q(306)
                           => DataPath_RF_bus_selected_win_data_50_port, Q(305)
                           => DataPath_RF_bus_selected_win_data_49_port, Q(304)
                           => DataPath_RF_bus_selected_win_data_48_port, Q(303)
                           => DataPath_RF_bus_selected_win_data_47_port, Q(302)
                           => DataPath_RF_bus_selected_win_data_46_port, Q(301)
                           => DataPath_RF_bus_selected_win_data_45_port, Q(300)
                           => DataPath_RF_bus_selected_win_data_44_port, Q(299)
                           => DataPath_RF_bus_selected_win_data_43_port, Q(298)
                           => DataPath_RF_bus_selected_win_data_42_port, Q(297)
                           => DataPath_RF_bus_selected_win_data_41_port, Q(296)
                           => DataPath_RF_bus_selected_win_data_40_port, Q(295)
                           => DataPath_RF_bus_selected_win_data_39_port, Q(294)
                           => DataPath_RF_bus_selected_win_data_38_port, Q(293)
                           => DataPath_RF_bus_selected_win_data_37_port, Q(292)
                           => DataPath_RF_bus_selected_win_data_36_port, Q(291)
                           => DataPath_RF_bus_selected_win_data_35_port, Q(290)
                           => DataPath_RF_bus_selected_win_data_34_port, Q(289)
                           => DataPath_RF_bus_selected_win_data_33_port, Q(288)
                           => DataPath_RF_bus_selected_win_data_32_port, Q(287)
                           => DataPath_RF_bus_selected_win_data_31_port, Q(286)
                           => DataPath_RF_bus_selected_win_data_30_port, Q(285)
                           => DataPath_RF_bus_selected_win_data_29_port, Q(284)
                           => DataPath_RF_bus_selected_win_data_28_port, Q(283)
                           => DataPath_RF_bus_selected_win_data_27_port, Q(282)
                           => DataPath_RF_bus_selected_win_data_26_port, Q(281)
                           => DataPath_RF_bus_selected_win_data_25_port, Q(280)
                           => DataPath_RF_bus_selected_win_data_24_port, Q(279)
                           => DataPath_RF_bus_selected_win_data_23_port, Q(278)
                           => DataPath_RF_bus_selected_win_data_22_port, Q(277)
                           => DataPath_RF_bus_selected_win_data_21_port, Q(276)
                           => DataPath_RF_bus_selected_win_data_20_port, Q(275)
                           => DataPath_RF_bus_selected_win_data_19_port, Q(274)
                           => DataPath_RF_bus_selected_win_data_18_port, Q(273)
                           => DataPath_RF_bus_selected_win_data_17_port, Q(272)
                           => DataPath_RF_bus_selected_win_data_16_port, Q(271)
                           => DataPath_RF_bus_selected_win_data_15_port, Q(270)
                           => DataPath_RF_bus_selected_win_data_14_port, Q(269)
                           => DataPath_RF_bus_selected_win_data_13_port, Q(268)
                           => DataPath_RF_bus_selected_win_data_12_port, Q(267)
                           => DataPath_RF_bus_selected_win_data_11_port, Q(266)
                           => DataPath_RF_bus_selected_win_data_10_port, Q(265)
                           => DataPath_RF_bus_selected_win_data_9_port, Q(264) 
                           => DataPath_RF_bus_selected_win_data_8_port, Q(263) 
                           => DataPath_RF_bus_selected_win_data_7_port, Q(262) 
                           => DataPath_RF_bus_selected_win_data_6_port, Q(261) 
                           => DataPath_RF_bus_selected_win_data_5_port, Q(260) 
                           => DataPath_RF_bus_selected_win_data_4_port, Q(259) 
                           => DataPath_RF_bus_selected_win_data_3_port, Q(258) 
                           => DataPath_RF_bus_selected_win_data_2_port, Q(257) 
                           => DataPath_RF_bus_selected_win_data_1_port, Q(256) 
                           => DataPath_RF_bus_selected_win_data_0_port, Q(255) 
                           => DataPath_RF_bus_complete_win_data_255_port, 
                           Q(254) => DataPath_RF_bus_complete_win_data_254_port
                           , Q(253) => 
                           DataPath_RF_bus_complete_win_data_253_port, Q(252) 
                           => DataPath_RF_bus_complete_win_data_252_port, 
                           Q(251) => DataPath_RF_bus_complete_win_data_251_port
                           , Q(250) => 
                           DataPath_RF_bus_complete_win_data_250_port, Q(249) 
                           => DataPath_RF_bus_complete_win_data_249_port, 
                           Q(248) => DataPath_RF_bus_complete_win_data_248_port
                           , Q(247) => 
                           DataPath_RF_bus_complete_win_data_247_port, Q(246) 
                           => DataPath_RF_bus_complete_win_data_246_port, 
                           Q(245) => DataPath_RF_bus_complete_win_data_245_port
                           , Q(244) => 
                           DataPath_RF_bus_complete_win_data_244_port, Q(243) 
                           => DataPath_RF_bus_complete_win_data_243_port, 
                           Q(242) => DataPath_RF_bus_complete_win_data_242_port
                           , Q(241) => 
                           DataPath_RF_bus_complete_win_data_241_port, Q(240) 
                           => DataPath_RF_bus_complete_win_data_240_port, 
                           Q(239) => DataPath_RF_bus_complete_win_data_239_port
                           , Q(238) => 
                           DataPath_RF_bus_complete_win_data_238_port, Q(237) 
                           => DataPath_RF_bus_complete_win_data_237_port, 
                           Q(236) => DataPath_RF_bus_complete_win_data_236_port
                           , Q(235) => 
                           DataPath_RF_bus_complete_win_data_235_port, Q(234) 
                           => DataPath_RF_bus_complete_win_data_234_port, 
                           Q(233) => DataPath_RF_bus_complete_win_data_233_port
                           , Q(232) => 
                           DataPath_RF_bus_complete_win_data_232_port, Q(231) 
                           => DataPath_RF_bus_complete_win_data_231_port, 
                           Q(230) => DataPath_RF_bus_complete_win_data_230_port
                           , Q(229) => 
                           DataPath_RF_bus_complete_win_data_229_port, Q(228) 
                           => DataPath_RF_bus_complete_win_data_228_port, 
                           Q(227) => DataPath_RF_bus_complete_win_data_227_port
                           , Q(226) => 
                           DataPath_RF_bus_complete_win_data_226_port, Q(225) 
                           => DataPath_RF_bus_complete_win_data_225_port, 
                           Q(224) => DataPath_RF_bus_complete_win_data_224_port
                           , Q(223) => 
                           DataPath_RF_bus_complete_win_data_223_port, Q(222) 
                           => DataPath_RF_bus_complete_win_data_222_port, 
                           Q(221) => DataPath_RF_bus_complete_win_data_221_port
                           , Q(220) => 
                           DataPath_RF_bus_complete_win_data_220_port, Q(219) 
                           => DataPath_RF_bus_complete_win_data_219_port, 
                           Q(218) => DataPath_RF_bus_complete_win_data_218_port
                           , Q(217) => 
                           DataPath_RF_bus_complete_win_data_217_port, Q(216) 
                           => DataPath_RF_bus_complete_win_data_216_port, 
                           Q(215) => DataPath_RF_bus_complete_win_data_215_port
                           , Q(214) => 
                           DataPath_RF_bus_complete_win_data_214_port, Q(213) 
                           => DataPath_RF_bus_complete_win_data_213_port, 
                           Q(212) => DataPath_RF_bus_complete_win_data_212_port
                           , Q(211) => 
                           DataPath_RF_bus_complete_win_data_211_port, Q(210) 
                           => DataPath_RF_bus_complete_win_data_210_port, 
                           Q(209) => DataPath_RF_bus_complete_win_data_209_port
                           , Q(208) => 
                           DataPath_RF_bus_complete_win_data_208_port, Q(207) 
                           => DataPath_RF_bus_complete_win_data_207_port, 
                           Q(206) => DataPath_RF_bus_complete_win_data_206_port
                           , Q(205) => 
                           DataPath_RF_bus_complete_win_data_205_port, Q(204) 
                           => DataPath_RF_bus_complete_win_data_204_port, 
                           Q(203) => DataPath_RF_bus_complete_win_data_203_port
                           , Q(202) => 
                           DataPath_RF_bus_complete_win_data_202_port, Q(201) 
                           => DataPath_RF_bus_complete_win_data_201_port, 
                           Q(200) => DataPath_RF_bus_complete_win_data_200_port
                           , Q(199) => 
                           DataPath_RF_bus_complete_win_data_199_port, Q(198) 
                           => DataPath_RF_bus_complete_win_data_198_port, 
                           Q(197) => DataPath_RF_bus_complete_win_data_197_port
                           , Q(196) => 
                           DataPath_RF_bus_complete_win_data_196_port, Q(195) 
                           => DataPath_RF_bus_complete_win_data_195_port, 
                           Q(194) => DataPath_RF_bus_complete_win_data_194_port
                           , Q(193) => 
                           DataPath_RF_bus_complete_win_data_193_port, Q(192) 
                           => DataPath_RF_bus_complete_win_data_192_port, 
                           Q(191) => DataPath_RF_bus_complete_win_data_191_port
                           , Q(190) => 
                           DataPath_RF_bus_complete_win_data_190_port, Q(189) 
                           => DataPath_RF_bus_complete_win_data_189_port, 
                           Q(188) => DataPath_RF_bus_complete_win_data_188_port
                           , Q(187) => 
                           DataPath_RF_bus_complete_win_data_187_port, Q(186) 
                           => DataPath_RF_bus_complete_win_data_186_port, 
                           Q(185) => DataPath_RF_bus_complete_win_data_185_port
                           , Q(184) => 
                           DataPath_RF_bus_complete_win_data_184_port, Q(183) 
                           => DataPath_RF_bus_complete_win_data_183_port, 
                           Q(182) => DataPath_RF_bus_complete_win_data_182_port
                           , Q(181) => 
                           DataPath_RF_bus_complete_win_data_181_port, Q(180) 
                           => DataPath_RF_bus_complete_win_data_180_port, 
                           Q(179) => DataPath_RF_bus_complete_win_data_179_port
                           , Q(178) => 
                           DataPath_RF_bus_complete_win_data_178_port, Q(177) 
                           => DataPath_RF_bus_complete_win_data_177_port, 
                           Q(176) => DataPath_RF_bus_complete_win_data_176_port
                           , Q(175) => 
                           DataPath_RF_bus_complete_win_data_175_port, Q(174) 
                           => DataPath_RF_bus_complete_win_data_174_port, 
                           Q(173) => DataPath_RF_bus_complete_win_data_173_port
                           , Q(172) => 
                           DataPath_RF_bus_complete_win_data_172_port, Q(171) 
                           => DataPath_RF_bus_complete_win_data_171_port, 
                           Q(170) => DataPath_RF_bus_complete_win_data_170_port
                           , Q(169) => 
                           DataPath_RF_bus_complete_win_data_169_port, Q(168) 
                           => DataPath_RF_bus_complete_win_data_168_port, 
                           Q(167) => DataPath_RF_bus_complete_win_data_167_port
                           , Q(166) => 
                           DataPath_RF_bus_complete_win_data_166_port, Q(165) 
                           => DataPath_RF_bus_complete_win_data_165_port, 
                           Q(164) => DataPath_RF_bus_complete_win_data_164_port
                           , Q(163) => 
                           DataPath_RF_bus_complete_win_data_163_port, Q(162) 
                           => DataPath_RF_bus_complete_win_data_162_port, 
                           Q(161) => DataPath_RF_bus_complete_win_data_161_port
                           , Q(160) => 
                           DataPath_RF_bus_complete_win_data_160_port, Q(159) 
                           => DataPath_RF_bus_complete_win_data_159_port, 
                           Q(158) => DataPath_RF_bus_complete_win_data_158_port
                           , Q(157) => 
                           DataPath_RF_bus_complete_win_data_157_port, Q(156) 
                           => DataPath_RF_bus_complete_win_data_156_port, 
                           Q(155) => DataPath_RF_bus_complete_win_data_155_port
                           , Q(154) => 
                           DataPath_RF_bus_complete_win_data_154_port, Q(153) 
                           => DataPath_RF_bus_complete_win_data_153_port, 
                           Q(152) => DataPath_RF_bus_complete_win_data_152_port
                           , Q(151) => 
                           DataPath_RF_bus_complete_win_data_151_port, Q(150) 
                           => DataPath_RF_bus_complete_win_data_150_port, 
                           Q(149) => DataPath_RF_bus_complete_win_data_149_port
                           , Q(148) => 
                           DataPath_RF_bus_complete_win_data_148_port, Q(147) 
                           => DataPath_RF_bus_complete_win_data_147_port, 
                           Q(146) => DataPath_RF_bus_complete_win_data_146_port
                           , Q(145) => 
                           DataPath_RF_bus_complete_win_data_145_port, Q(144) 
                           => DataPath_RF_bus_complete_win_data_144_port, 
                           Q(143) => DataPath_RF_bus_complete_win_data_143_port
                           , Q(142) => 
                           DataPath_RF_bus_complete_win_data_142_port, Q(141) 
                           => DataPath_RF_bus_complete_win_data_141_port, 
                           Q(140) => DataPath_RF_bus_complete_win_data_140_port
                           , Q(139) => 
                           DataPath_RF_bus_complete_win_data_139_port, Q(138) 
                           => DataPath_RF_bus_complete_win_data_138_port, 
                           Q(137) => DataPath_RF_bus_complete_win_data_137_port
                           , Q(136) => 
                           DataPath_RF_bus_complete_win_data_136_port, Q(135) 
                           => DataPath_RF_bus_complete_win_data_135_port, 
                           Q(134) => DataPath_RF_bus_complete_win_data_134_port
                           , Q(133) => 
                           DataPath_RF_bus_complete_win_data_133_port, Q(132) 
                           => DataPath_RF_bus_complete_win_data_132_port, 
                           Q(131) => DataPath_RF_bus_complete_win_data_131_port
                           , Q(130) => 
                           DataPath_RF_bus_complete_win_data_130_port, Q(129) 
                           => DataPath_RF_bus_complete_win_data_129_port, 
                           Q(128) => DataPath_RF_bus_complete_win_data_128_port
                           , Q(127) => 
                           DataPath_RF_bus_complete_win_data_127_port, Q(126) 
                           => DataPath_RF_bus_complete_win_data_126_port, 
                           Q(125) => DataPath_RF_bus_complete_win_data_125_port
                           , Q(124) => 
                           DataPath_RF_bus_complete_win_data_124_port, Q(123) 
                           => DataPath_RF_bus_complete_win_data_123_port, 
                           Q(122) => DataPath_RF_bus_complete_win_data_122_port
                           , Q(121) => 
                           DataPath_RF_bus_complete_win_data_121_port, Q(120) 
                           => DataPath_RF_bus_complete_win_data_120_port, 
                           Q(119) => DataPath_RF_bus_complete_win_data_119_port
                           , Q(118) => 
                           DataPath_RF_bus_complete_win_data_118_port, Q(117) 
                           => DataPath_RF_bus_complete_win_data_117_port, 
                           Q(116) => DataPath_RF_bus_complete_win_data_116_port
                           , Q(115) => 
                           DataPath_RF_bus_complete_win_data_115_port, Q(114) 
                           => DataPath_RF_bus_complete_win_data_114_port, 
                           Q(113) => DataPath_RF_bus_complete_win_data_113_port
                           , Q(112) => 
                           DataPath_RF_bus_complete_win_data_112_port, Q(111) 
                           => DataPath_RF_bus_complete_win_data_111_port, 
                           Q(110) => DataPath_RF_bus_complete_win_data_110_port
                           , Q(109) => 
                           DataPath_RF_bus_complete_win_data_109_port, Q(108) 
                           => DataPath_RF_bus_complete_win_data_108_port, 
                           Q(107) => DataPath_RF_bus_complete_win_data_107_port
                           , Q(106) => 
                           DataPath_RF_bus_complete_win_data_106_port, Q(105) 
                           => DataPath_RF_bus_complete_win_data_105_port, 
                           Q(104) => DataPath_RF_bus_complete_win_data_104_port
                           , Q(103) => 
                           DataPath_RF_bus_complete_win_data_103_port, Q(102) 
                           => DataPath_RF_bus_complete_win_data_102_port, 
                           Q(101) => DataPath_RF_bus_complete_win_data_101_port
                           , Q(100) => 
                           DataPath_RF_bus_complete_win_data_100_port, Q(99) =>
                           DataPath_RF_bus_complete_win_data_99_port, Q(98) => 
                           DataPath_RF_bus_complete_win_data_98_port, Q(97) => 
                           DataPath_RF_bus_complete_win_data_97_port, Q(96) => 
                           DataPath_RF_bus_complete_win_data_96_port, Q(95) => 
                           DataPath_RF_bus_complete_win_data_95_port, Q(94) => 
                           DataPath_RF_bus_complete_win_data_94_port, Q(93) => 
                           DataPath_RF_bus_complete_win_data_93_port, Q(92) => 
                           DataPath_RF_bus_complete_win_data_92_port, Q(91) => 
                           DataPath_RF_bus_complete_win_data_91_port, Q(90) => 
                           DataPath_RF_bus_complete_win_data_90_port, Q(89) => 
                           DataPath_RF_bus_complete_win_data_89_port, Q(88) => 
                           DataPath_RF_bus_complete_win_data_88_port, Q(87) => 
                           DataPath_RF_bus_complete_win_data_87_port, Q(86) => 
                           DataPath_RF_bus_complete_win_data_86_port, Q(85) => 
                           DataPath_RF_bus_complete_win_data_85_port, Q(84) => 
                           DataPath_RF_bus_complete_win_data_84_port, Q(83) => 
                           DataPath_RF_bus_complete_win_data_83_port, Q(82) => 
                           DataPath_RF_bus_complete_win_data_82_port, Q(81) => 
                           DataPath_RF_bus_complete_win_data_81_port, Q(80) => 
                           DataPath_RF_bus_complete_win_data_80_port, Q(79) => 
                           DataPath_RF_bus_complete_win_data_79_port, Q(78) => 
                           DataPath_RF_bus_complete_win_data_78_port, Q(77) => 
                           DataPath_RF_bus_complete_win_data_77_port, Q(76) => 
                           DataPath_RF_bus_complete_win_data_76_port, Q(75) => 
                           DataPath_RF_bus_complete_win_data_75_port, Q(74) => 
                           DataPath_RF_bus_complete_win_data_74_port, Q(73) => 
                           DataPath_RF_bus_complete_win_data_73_port, Q(72) => 
                           DataPath_RF_bus_complete_win_data_72_port, Q(71) => 
                           DataPath_RF_bus_complete_win_data_71_port, Q(70) => 
                           DataPath_RF_bus_complete_win_data_70_port, Q(69) => 
                           DataPath_RF_bus_complete_win_data_69_port, Q(68) => 
                           DataPath_RF_bus_complete_win_data_68_port, Q(67) => 
                           DataPath_RF_bus_complete_win_data_67_port, Q(66) => 
                           DataPath_RF_bus_complete_win_data_66_port, Q(65) => 
                           DataPath_RF_bus_complete_win_data_65_port, Q(64) => 
                           DataPath_RF_bus_complete_win_data_64_port, Q(63) => 
                           DataPath_RF_bus_complete_win_data_63_port, Q(62) => 
                           DataPath_RF_bus_complete_win_data_62_port, Q(61) => 
                           DataPath_RF_bus_complete_win_data_61_port, Q(60) => 
                           DataPath_RF_bus_complete_win_data_60_port, Q(59) => 
                           DataPath_RF_bus_complete_win_data_59_port, Q(58) => 
                           DataPath_RF_bus_complete_win_data_58_port, Q(57) => 
                           DataPath_RF_bus_complete_win_data_57_port, Q(56) => 
                           DataPath_RF_bus_complete_win_data_56_port, Q(55) => 
                           DataPath_RF_bus_complete_win_data_55_port, Q(54) => 
                           DataPath_RF_bus_complete_win_data_54_port, Q(53) => 
                           DataPath_RF_bus_complete_win_data_53_port, Q(52) => 
                           DataPath_RF_bus_complete_win_data_52_port, Q(51) => 
                           DataPath_RF_bus_complete_win_data_51_port, Q(50) => 
                           DataPath_RF_bus_complete_win_data_50_port, Q(49) => 
                           DataPath_RF_bus_complete_win_data_49_port, Q(48) => 
                           DataPath_RF_bus_complete_win_data_48_port, Q(47) => 
                           DataPath_RF_bus_complete_win_data_47_port, Q(46) => 
                           DataPath_RF_bus_complete_win_data_46_port, Q(45) => 
                           DataPath_RF_bus_complete_win_data_45_port, Q(44) => 
                           DataPath_RF_bus_complete_win_data_44_port, Q(43) => 
                           DataPath_RF_bus_complete_win_data_43_port, Q(42) => 
                           DataPath_RF_bus_complete_win_data_42_port, Q(41) => 
                           DataPath_RF_bus_complete_win_data_41_port, Q(40) => 
                           DataPath_RF_bus_complete_win_data_40_port, Q(39) => 
                           DataPath_RF_bus_complete_win_data_39_port, Q(38) => 
                           DataPath_RF_bus_complete_win_data_38_port, Q(37) => 
                           DataPath_RF_bus_complete_win_data_37_port, Q(36) => 
                           DataPath_RF_bus_complete_win_data_36_port, Q(35) => 
                           DataPath_RF_bus_complete_win_data_35_port, Q(34) => 
                           DataPath_RF_bus_complete_win_data_34_port, Q(33) => 
                           DataPath_RF_bus_complete_win_data_33_port, Q(32) => 
                           DataPath_RF_bus_complete_win_data_32_port, Q(31) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(30) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(29) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(28) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(27) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(26) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(25) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(24) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(23) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(22) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(21) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(20) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(19) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(18) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(17) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(16) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(15) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(14) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(13) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(12) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(11) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(10) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(9) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(8) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(7) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(6) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(5) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(4) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(3) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(2) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(1) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(0) => 
                           DataPath_RF_bus_complete_win_data_0_port, Y(31) => 
                           DataPath_RF_internal_out2_31_port, Y(30) => 
                           DataPath_RF_internal_out2_30_port, Y(29) => 
                           DataPath_RF_internal_out2_29_port, Y(28) => 
                           DataPath_RF_internal_out2_28_port, Y(27) => 
                           DataPath_RF_internal_out2_27_port, Y(26) => 
                           DataPath_RF_internal_out2_26_port, Y(25) => 
                           DataPath_RF_internal_out2_25_port, Y(24) => 
                           DataPath_RF_internal_out2_24_port, Y(23) => 
                           DataPath_RF_internal_out2_23_port, Y(22) => 
                           DataPath_RF_internal_out2_22_port, Y(21) => 
                           DataPath_RF_internal_out2_21_port, Y(20) => 
                           DataPath_RF_internal_out2_20_port, Y(19) => 
                           DataPath_RF_internal_out2_19_port, Y(18) => 
                           DataPath_RF_internal_out2_18_port, Y(17) => 
                           DataPath_RF_internal_out2_17_port, Y(16) => 
                           DataPath_RF_internal_out2_16_port, Y(15) => 
                           DataPath_RF_internal_out2_15_port, Y(14) => 
                           DataPath_RF_internal_out2_14_port, Y(13) => 
                           DataPath_RF_internal_out2_13_port, Y(12) => 
                           DataPath_RF_internal_out2_12_port, Y(11) => 
                           DataPath_RF_internal_out2_11_port, Y(10) => 
                           DataPath_RF_internal_out2_10_port, Y(9) => 
                           DataPath_RF_internal_out2_9_port, Y(8) => 
                           DataPath_RF_internal_out2_8_port, Y(7) => 
                           DataPath_RF_internal_out2_7_port, Y(6) => 
                           DataPath_RF_internal_out2_6_port, Y(5) => 
                           DataPath_RF_internal_out2_5_port, Y(4) => 
                           DataPath_RF_internal_out2_4_port, Y(3) => 
                           DataPath_RF_internal_out2_3_port, Y(2) => 
                           DataPath_RF_internal_out2_2_port, Y(1) => 
                           DataPath_RF_internal_out2_1_port, Y(0) => 
                           DataPath_RF_internal_out2_0_port);
   DataPath_RF_RDPORT0 : mux_N32_M5_0 port map( S(4) => i_ADD_RS1_4_port, S(3) 
                           => i_ADD_RS1_3_port, S(2) => i_ADD_RS1_2_port, S(1) 
                           => i_ADD_RS1_1_port, S(0) => i_ADD_RS1_0_port, 
                           Q(1023) => 
                           DataPath_RF_bus_selected_win_data_767_port, Q(1022) 
                           => DataPath_RF_bus_selected_win_data_766_port, 
                           Q(1021) => 
                           DataPath_RF_bus_selected_win_data_765_port, Q(1020) 
                           => DataPath_RF_bus_selected_win_data_764_port, 
                           Q(1019) => 
                           DataPath_RF_bus_selected_win_data_763_port, Q(1018) 
                           => DataPath_RF_bus_selected_win_data_762_port, 
                           Q(1017) => 
                           DataPath_RF_bus_selected_win_data_761_port, Q(1016) 
                           => DataPath_RF_bus_selected_win_data_760_port, 
                           Q(1015) => 
                           DataPath_RF_bus_selected_win_data_759_port, Q(1014) 
                           => DataPath_RF_bus_selected_win_data_758_port, 
                           Q(1013) => 
                           DataPath_RF_bus_selected_win_data_757_port, Q(1012) 
                           => DataPath_RF_bus_selected_win_data_756_port, 
                           Q(1011) => 
                           DataPath_RF_bus_selected_win_data_755_port, Q(1010) 
                           => DataPath_RF_bus_selected_win_data_754_port, 
                           Q(1009) => 
                           DataPath_RF_bus_selected_win_data_753_port, Q(1008) 
                           => DataPath_RF_bus_selected_win_data_752_port, 
                           Q(1007) => 
                           DataPath_RF_bus_selected_win_data_751_port, Q(1006) 
                           => DataPath_RF_bus_selected_win_data_750_port, 
                           Q(1005) => 
                           DataPath_RF_bus_selected_win_data_749_port, Q(1004) 
                           => DataPath_RF_bus_selected_win_data_748_port, 
                           Q(1003) => 
                           DataPath_RF_bus_selected_win_data_747_port, Q(1002) 
                           => DataPath_RF_bus_selected_win_data_746_port, 
                           Q(1001) => 
                           DataPath_RF_bus_selected_win_data_745_port, Q(1000) 
                           => DataPath_RF_bus_selected_win_data_744_port, 
                           Q(999) => DataPath_RF_bus_selected_win_data_743_port
                           , Q(998) => 
                           DataPath_RF_bus_selected_win_data_742_port, Q(997) 
                           => DataPath_RF_bus_selected_win_data_741_port, 
                           Q(996) => DataPath_RF_bus_selected_win_data_740_port
                           , Q(995) => 
                           DataPath_RF_bus_selected_win_data_739_port, Q(994) 
                           => DataPath_RF_bus_selected_win_data_738_port, 
                           Q(993) => DataPath_RF_bus_selected_win_data_737_port
                           , Q(992) => 
                           DataPath_RF_bus_selected_win_data_736_port, Q(991) 
                           => DataPath_RF_bus_selected_win_data_735_port, 
                           Q(990) => DataPath_RF_bus_selected_win_data_734_port
                           , Q(989) => 
                           DataPath_RF_bus_selected_win_data_733_port, Q(988) 
                           => DataPath_RF_bus_selected_win_data_732_port, 
                           Q(987) => DataPath_RF_bus_selected_win_data_731_port
                           , Q(986) => 
                           DataPath_RF_bus_selected_win_data_730_port, Q(985) 
                           => DataPath_RF_bus_selected_win_data_729_port, 
                           Q(984) => DataPath_RF_bus_selected_win_data_728_port
                           , Q(983) => 
                           DataPath_RF_bus_selected_win_data_727_port, Q(982) 
                           => DataPath_RF_bus_selected_win_data_726_port, 
                           Q(981) => DataPath_RF_bus_selected_win_data_725_port
                           , Q(980) => 
                           DataPath_RF_bus_selected_win_data_724_port, Q(979) 
                           => DataPath_RF_bus_selected_win_data_723_port, 
                           Q(978) => DataPath_RF_bus_selected_win_data_722_port
                           , Q(977) => 
                           DataPath_RF_bus_selected_win_data_721_port, Q(976) 
                           => DataPath_RF_bus_selected_win_data_720_port, 
                           Q(975) => DataPath_RF_bus_selected_win_data_719_port
                           , Q(974) => 
                           DataPath_RF_bus_selected_win_data_718_port, Q(973) 
                           => DataPath_RF_bus_selected_win_data_717_port, 
                           Q(972) => DataPath_RF_bus_selected_win_data_716_port
                           , Q(971) => 
                           DataPath_RF_bus_selected_win_data_715_port, Q(970) 
                           => DataPath_RF_bus_selected_win_data_714_port, 
                           Q(969) => DataPath_RF_bus_selected_win_data_713_port
                           , Q(968) => 
                           DataPath_RF_bus_selected_win_data_712_port, Q(967) 
                           => DataPath_RF_bus_selected_win_data_711_port, 
                           Q(966) => DataPath_RF_bus_selected_win_data_710_port
                           , Q(965) => 
                           DataPath_RF_bus_selected_win_data_709_port, Q(964) 
                           => DataPath_RF_bus_selected_win_data_708_port, 
                           Q(963) => DataPath_RF_bus_selected_win_data_707_port
                           , Q(962) => 
                           DataPath_RF_bus_selected_win_data_706_port, Q(961) 
                           => DataPath_RF_bus_selected_win_data_705_port, 
                           Q(960) => DataPath_RF_bus_selected_win_data_704_port
                           , Q(959) => 
                           DataPath_RF_bus_selected_win_data_703_port, Q(958) 
                           => DataPath_RF_bus_selected_win_data_702_port, 
                           Q(957) => DataPath_RF_bus_selected_win_data_701_port
                           , Q(956) => 
                           DataPath_RF_bus_selected_win_data_700_port, Q(955) 
                           => DataPath_RF_bus_selected_win_data_699_port, 
                           Q(954) => DataPath_RF_bus_selected_win_data_698_port
                           , Q(953) => 
                           DataPath_RF_bus_selected_win_data_697_port, Q(952) 
                           => DataPath_RF_bus_selected_win_data_696_port, 
                           Q(951) => DataPath_RF_bus_selected_win_data_695_port
                           , Q(950) => 
                           DataPath_RF_bus_selected_win_data_694_port, Q(949) 
                           => DataPath_RF_bus_selected_win_data_693_port, 
                           Q(948) => DataPath_RF_bus_selected_win_data_692_port
                           , Q(947) => 
                           DataPath_RF_bus_selected_win_data_691_port, Q(946) 
                           => DataPath_RF_bus_selected_win_data_690_port, 
                           Q(945) => DataPath_RF_bus_selected_win_data_689_port
                           , Q(944) => 
                           DataPath_RF_bus_selected_win_data_688_port, Q(943) 
                           => DataPath_RF_bus_selected_win_data_687_port, 
                           Q(942) => DataPath_RF_bus_selected_win_data_686_port
                           , Q(941) => 
                           DataPath_RF_bus_selected_win_data_685_port, Q(940) 
                           => DataPath_RF_bus_selected_win_data_684_port, 
                           Q(939) => DataPath_RF_bus_selected_win_data_683_port
                           , Q(938) => 
                           DataPath_RF_bus_selected_win_data_682_port, Q(937) 
                           => DataPath_RF_bus_selected_win_data_681_port, 
                           Q(936) => DataPath_RF_bus_selected_win_data_680_port
                           , Q(935) => 
                           DataPath_RF_bus_selected_win_data_679_port, Q(934) 
                           => DataPath_RF_bus_selected_win_data_678_port, 
                           Q(933) => DataPath_RF_bus_selected_win_data_677_port
                           , Q(932) => 
                           DataPath_RF_bus_selected_win_data_676_port, Q(931) 
                           => DataPath_RF_bus_selected_win_data_675_port, 
                           Q(930) => DataPath_RF_bus_selected_win_data_674_port
                           , Q(929) => 
                           DataPath_RF_bus_selected_win_data_673_port, Q(928) 
                           => DataPath_RF_bus_selected_win_data_672_port, 
                           Q(927) => DataPath_RF_bus_selected_win_data_671_port
                           , Q(926) => 
                           DataPath_RF_bus_selected_win_data_670_port, Q(925) 
                           => DataPath_RF_bus_selected_win_data_669_port, 
                           Q(924) => DataPath_RF_bus_selected_win_data_668_port
                           , Q(923) => 
                           DataPath_RF_bus_selected_win_data_667_port, Q(922) 
                           => DataPath_RF_bus_selected_win_data_666_port, 
                           Q(921) => DataPath_RF_bus_selected_win_data_665_port
                           , Q(920) => 
                           DataPath_RF_bus_selected_win_data_664_port, Q(919) 
                           => DataPath_RF_bus_selected_win_data_663_port, 
                           Q(918) => DataPath_RF_bus_selected_win_data_662_port
                           , Q(917) => 
                           DataPath_RF_bus_selected_win_data_661_port, Q(916) 
                           => DataPath_RF_bus_selected_win_data_660_port, 
                           Q(915) => DataPath_RF_bus_selected_win_data_659_port
                           , Q(914) => 
                           DataPath_RF_bus_selected_win_data_658_port, Q(913) 
                           => DataPath_RF_bus_selected_win_data_657_port, 
                           Q(912) => DataPath_RF_bus_selected_win_data_656_port
                           , Q(911) => 
                           DataPath_RF_bus_selected_win_data_655_port, Q(910) 
                           => DataPath_RF_bus_selected_win_data_654_port, 
                           Q(909) => DataPath_RF_bus_selected_win_data_653_port
                           , Q(908) => 
                           DataPath_RF_bus_selected_win_data_652_port, Q(907) 
                           => DataPath_RF_bus_selected_win_data_651_port, 
                           Q(906) => DataPath_RF_bus_selected_win_data_650_port
                           , Q(905) => 
                           DataPath_RF_bus_selected_win_data_649_port, Q(904) 
                           => DataPath_RF_bus_selected_win_data_648_port, 
                           Q(903) => DataPath_RF_bus_selected_win_data_647_port
                           , Q(902) => 
                           DataPath_RF_bus_selected_win_data_646_port, Q(901) 
                           => DataPath_RF_bus_selected_win_data_645_port, 
                           Q(900) => DataPath_RF_bus_selected_win_data_644_port
                           , Q(899) => 
                           DataPath_RF_bus_selected_win_data_643_port, Q(898) 
                           => DataPath_RF_bus_selected_win_data_642_port, 
                           Q(897) => DataPath_RF_bus_selected_win_data_641_port
                           , Q(896) => 
                           DataPath_RF_bus_selected_win_data_640_port, Q(895) 
                           => DataPath_RF_bus_selected_win_data_639_port, 
                           Q(894) => DataPath_RF_bus_selected_win_data_638_port
                           , Q(893) => 
                           DataPath_RF_bus_selected_win_data_637_port, Q(892) 
                           => DataPath_RF_bus_selected_win_data_636_port, 
                           Q(891) => DataPath_RF_bus_selected_win_data_635_port
                           , Q(890) => 
                           DataPath_RF_bus_selected_win_data_634_port, Q(889) 
                           => DataPath_RF_bus_selected_win_data_633_port, 
                           Q(888) => DataPath_RF_bus_selected_win_data_632_port
                           , Q(887) => 
                           DataPath_RF_bus_selected_win_data_631_port, Q(886) 
                           => DataPath_RF_bus_selected_win_data_630_port, 
                           Q(885) => DataPath_RF_bus_selected_win_data_629_port
                           , Q(884) => 
                           DataPath_RF_bus_selected_win_data_628_port, Q(883) 
                           => DataPath_RF_bus_selected_win_data_627_port, 
                           Q(882) => DataPath_RF_bus_selected_win_data_626_port
                           , Q(881) => 
                           DataPath_RF_bus_selected_win_data_625_port, Q(880) 
                           => DataPath_RF_bus_selected_win_data_624_port, 
                           Q(879) => DataPath_RF_bus_selected_win_data_623_port
                           , Q(878) => 
                           DataPath_RF_bus_selected_win_data_622_port, Q(877) 
                           => DataPath_RF_bus_selected_win_data_621_port, 
                           Q(876) => DataPath_RF_bus_selected_win_data_620_port
                           , Q(875) => 
                           DataPath_RF_bus_selected_win_data_619_port, Q(874) 
                           => DataPath_RF_bus_selected_win_data_618_port, 
                           Q(873) => DataPath_RF_bus_selected_win_data_617_port
                           , Q(872) => 
                           DataPath_RF_bus_selected_win_data_616_port, Q(871) 
                           => DataPath_RF_bus_selected_win_data_615_port, 
                           Q(870) => DataPath_RF_bus_selected_win_data_614_port
                           , Q(869) => 
                           DataPath_RF_bus_selected_win_data_613_port, Q(868) 
                           => DataPath_RF_bus_selected_win_data_612_port, 
                           Q(867) => DataPath_RF_bus_selected_win_data_611_port
                           , Q(866) => 
                           DataPath_RF_bus_selected_win_data_610_port, Q(865) 
                           => DataPath_RF_bus_selected_win_data_609_port, 
                           Q(864) => DataPath_RF_bus_selected_win_data_608_port
                           , Q(863) => 
                           DataPath_RF_bus_selected_win_data_607_port, Q(862) 
                           => DataPath_RF_bus_selected_win_data_606_port, 
                           Q(861) => DataPath_RF_bus_selected_win_data_605_port
                           , Q(860) => 
                           DataPath_RF_bus_selected_win_data_604_port, Q(859) 
                           => DataPath_RF_bus_selected_win_data_603_port, 
                           Q(858) => DataPath_RF_bus_selected_win_data_602_port
                           , Q(857) => 
                           DataPath_RF_bus_selected_win_data_601_port, Q(856) 
                           => DataPath_RF_bus_selected_win_data_600_port, 
                           Q(855) => DataPath_RF_bus_selected_win_data_599_port
                           , Q(854) => 
                           DataPath_RF_bus_selected_win_data_598_port, Q(853) 
                           => DataPath_RF_bus_selected_win_data_597_port, 
                           Q(852) => DataPath_RF_bus_selected_win_data_596_port
                           , Q(851) => 
                           DataPath_RF_bus_selected_win_data_595_port, Q(850) 
                           => DataPath_RF_bus_selected_win_data_594_port, 
                           Q(849) => DataPath_RF_bus_selected_win_data_593_port
                           , Q(848) => 
                           DataPath_RF_bus_selected_win_data_592_port, Q(847) 
                           => DataPath_RF_bus_selected_win_data_591_port, 
                           Q(846) => DataPath_RF_bus_selected_win_data_590_port
                           , Q(845) => 
                           DataPath_RF_bus_selected_win_data_589_port, Q(844) 
                           => DataPath_RF_bus_selected_win_data_588_port, 
                           Q(843) => DataPath_RF_bus_selected_win_data_587_port
                           , Q(842) => 
                           DataPath_RF_bus_selected_win_data_586_port, Q(841) 
                           => DataPath_RF_bus_selected_win_data_585_port, 
                           Q(840) => DataPath_RF_bus_selected_win_data_584_port
                           , Q(839) => 
                           DataPath_RF_bus_selected_win_data_583_port, Q(838) 
                           => DataPath_RF_bus_selected_win_data_582_port, 
                           Q(837) => DataPath_RF_bus_selected_win_data_581_port
                           , Q(836) => 
                           DataPath_RF_bus_selected_win_data_580_port, Q(835) 
                           => DataPath_RF_bus_selected_win_data_579_port, 
                           Q(834) => DataPath_RF_bus_selected_win_data_578_port
                           , Q(833) => 
                           DataPath_RF_bus_selected_win_data_577_port, Q(832) 
                           => DataPath_RF_bus_selected_win_data_576_port, 
                           Q(831) => DataPath_RF_bus_selected_win_data_575_port
                           , Q(830) => 
                           DataPath_RF_bus_selected_win_data_574_port, Q(829) 
                           => DataPath_RF_bus_selected_win_data_573_port, 
                           Q(828) => DataPath_RF_bus_selected_win_data_572_port
                           , Q(827) => 
                           DataPath_RF_bus_selected_win_data_571_port, Q(826) 
                           => DataPath_RF_bus_selected_win_data_570_port, 
                           Q(825) => DataPath_RF_bus_selected_win_data_569_port
                           , Q(824) => 
                           DataPath_RF_bus_selected_win_data_568_port, Q(823) 
                           => DataPath_RF_bus_selected_win_data_567_port, 
                           Q(822) => DataPath_RF_bus_selected_win_data_566_port
                           , Q(821) => 
                           DataPath_RF_bus_selected_win_data_565_port, Q(820) 
                           => DataPath_RF_bus_selected_win_data_564_port, 
                           Q(819) => DataPath_RF_bus_selected_win_data_563_port
                           , Q(818) => 
                           DataPath_RF_bus_selected_win_data_562_port, Q(817) 
                           => DataPath_RF_bus_selected_win_data_561_port, 
                           Q(816) => DataPath_RF_bus_selected_win_data_560_port
                           , Q(815) => 
                           DataPath_RF_bus_selected_win_data_559_port, Q(814) 
                           => DataPath_RF_bus_selected_win_data_558_port, 
                           Q(813) => DataPath_RF_bus_selected_win_data_557_port
                           , Q(812) => 
                           DataPath_RF_bus_selected_win_data_556_port, Q(811) 
                           => DataPath_RF_bus_selected_win_data_555_port, 
                           Q(810) => DataPath_RF_bus_selected_win_data_554_port
                           , Q(809) => 
                           DataPath_RF_bus_selected_win_data_553_port, Q(808) 
                           => DataPath_RF_bus_selected_win_data_552_port, 
                           Q(807) => DataPath_RF_bus_selected_win_data_551_port
                           , Q(806) => 
                           DataPath_RF_bus_selected_win_data_550_port, Q(805) 
                           => DataPath_RF_bus_selected_win_data_549_port, 
                           Q(804) => DataPath_RF_bus_selected_win_data_548_port
                           , Q(803) => 
                           DataPath_RF_bus_selected_win_data_547_port, Q(802) 
                           => DataPath_RF_bus_selected_win_data_546_port, 
                           Q(801) => DataPath_RF_bus_selected_win_data_545_port
                           , Q(800) => 
                           DataPath_RF_bus_selected_win_data_544_port, Q(799) 
                           => DataPath_RF_bus_selected_win_data_543_port, 
                           Q(798) => DataPath_RF_bus_selected_win_data_542_port
                           , Q(797) => 
                           DataPath_RF_bus_selected_win_data_541_port, Q(796) 
                           => DataPath_RF_bus_selected_win_data_540_port, 
                           Q(795) => DataPath_RF_bus_selected_win_data_539_port
                           , Q(794) => 
                           DataPath_RF_bus_selected_win_data_538_port, Q(793) 
                           => DataPath_RF_bus_selected_win_data_537_port, 
                           Q(792) => DataPath_RF_bus_selected_win_data_536_port
                           , Q(791) => 
                           DataPath_RF_bus_selected_win_data_535_port, Q(790) 
                           => DataPath_RF_bus_selected_win_data_534_port, 
                           Q(789) => DataPath_RF_bus_selected_win_data_533_port
                           , Q(788) => 
                           DataPath_RF_bus_selected_win_data_532_port, Q(787) 
                           => DataPath_RF_bus_selected_win_data_531_port, 
                           Q(786) => DataPath_RF_bus_selected_win_data_530_port
                           , Q(785) => 
                           DataPath_RF_bus_selected_win_data_529_port, Q(784) 
                           => DataPath_RF_bus_selected_win_data_528_port, 
                           Q(783) => DataPath_RF_bus_selected_win_data_527_port
                           , Q(782) => 
                           DataPath_RF_bus_selected_win_data_526_port, Q(781) 
                           => DataPath_RF_bus_selected_win_data_525_port, 
                           Q(780) => DataPath_RF_bus_selected_win_data_524_port
                           , Q(779) => 
                           DataPath_RF_bus_selected_win_data_523_port, Q(778) 
                           => DataPath_RF_bus_selected_win_data_522_port, 
                           Q(777) => DataPath_RF_bus_selected_win_data_521_port
                           , Q(776) => 
                           DataPath_RF_bus_selected_win_data_520_port, Q(775) 
                           => DataPath_RF_bus_selected_win_data_519_port, 
                           Q(774) => DataPath_RF_bus_selected_win_data_518_port
                           , Q(773) => 
                           DataPath_RF_bus_selected_win_data_517_port, Q(772) 
                           => DataPath_RF_bus_selected_win_data_516_port, 
                           Q(771) => DataPath_RF_bus_selected_win_data_515_port
                           , Q(770) => 
                           DataPath_RF_bus_selected_win_data_514_port, Q(769) 
                           => DataPath_RF_bus_selected_win_data_513_port, 
                           Q(768) => DataPath_RF_bus_selected_win_data_512_port
                           , Q(767) => 
                           DataPath_RF_bus_selected_win_data_511_port, Q(766) 
                           => DataPath_RF_bus_selected_win_data_510_port, 
                           Q(765) => DataPath_RF_bus_selected_win_data_509_port
                           , Q(764) => 
                           DataPath_RF_bus_selected_win_data_508_port, Q(763) 
                           => DataPath_RF_bus_selected_win_data_507_port, 
                           Q(762) => DataPath_RF_bus_selected_win_data_506_port
                           , Q(761) => 
                           DataPath_RF_bus_selected_win_data_505_port, Q(760) 
                           => DataPath_RF_bus_selected_win_data_504_port, 
                           Q(759) => DataPath_RF_bus_selected_win_data_503_port
                           , Q(758) => 
                           DataPath_RF_bus_selected_win_data_502_port, Q(757) 
                           => DataPath_RF_bus_selected_win_data_501_port, 
                           Q(756) => DataPath_RF_bus_selected_win_data_500_port
                           , Q(755) => 
                           DataPath_RF_bus_selected_win_data_499_port, Q(754) 
                           => DataPath_RF_bus_selected_win_data_498_port, 
                           Q(753) => DataPath_RF_bus_selected_win_data_497_port
                           , Q(752) => 
                           DataPath_RF_bus_selected_win_data_496_port, Q(751) 
                           => DataPath_RF_bus_selected_win_data_495_port, 
                           Q(750) => DataPath_RF_bus_selected_win_data_494_port
                           , Q(749) => 
                           DataPath_RF_bus_selected_win_data_493_port, Q(748) 
                           => DataPath_RF_bus_selected_win_data_492_port, 
                           Q(747) => DataPath_RF_bus_selected_win_data_491_port
                           , Q(746) => 
                           DataPath_RF_bus_selected_win_data_490_port, Q(745) 
                           => DataPath_RF_bus_selected_win_data_489_port, 
                           Q(744) => DataPath_RF_bus_selected_win_data_488_port
                           , Q(743) => 
                           DataPath_RF_bus_selected_win_data_487_port, Q(742) 
                           => DataPath_RF_bus_selected_win_data_486_port, 
                           Q(741) => DataPath_RF_bus_selected_win_data_485_port
                           , Q(740) => 
                           DataPath_RF_bus_selected_win_data_484_port, Q(739) 
                           => DataPath_RF_bus_selected_win_data_483_port, 
                           Q(738) => DataPath_RF_bus_selected_win_data_482_port
                           , Q(737) => 
                           DataPath_RF_bus_selected_win_data_481_port, Q(736) 
                           => DataPath_RF_bus_selected_win_data_480_port, 
                           Q(735) => DataPath_RF_bus_selected_win_data_479_port
                           , Q(734) => 
                           DataPath_RF_bus_selected_win_data_478_port, Q(733) 
                           => DataPath_RF_bus_selected_win_data_477_port, 
                           Q(732) => DataPath_RF_bus_selected_win_data_476_port
                           , Q(731) => 
                           DataPath_RF_bus_selected_win_data_475_port, Q(730) 
                           => DataPath_RF_bus_selected_win_data_474_port, 
                           Q(729) => DataPath_RF_bus_selected_win_data_473_port
                           , Q(728) => 
                           DataPath_RF_bus_selected_win_data_472_port, Q(727) 
                           => DataPath_RF_bus_selected_win_data_471_port, 
                           Q(726) => DataPath_RF_bus_selected_win_data_470_port
                           , Q(725) => 
                           DataPath_RF_bus_selected_win_data_469_port, Q(724) 
                           => DataPath_RF_bus_selected_win_data_468_port, 
                           Q(723) => DataPath_RF_bus_selected_win_data_467_port
                           , Q(722) => 
                           DataPath_RF_bus_selected_win_data_466_port, Q(721) 
                           => DataPath_RF_bus_selected_win_data_465_port, 
                           Q(720) => DataPath_RF_bus_selected_win_data_464_port
                           , Q(719) => 
                           DataPath_RF_bus_selected_win_data_463_port, Q(718) 
                           => DataPath_RF_bus_selected_win_data_462_port, 
                           Q(717) => DataPath_RF_bus_selected_win_data_461_port
                           , Q(716) => 
                           DataPath_RF_bus_selected_win_data_460_port, Q(715) 
                           => DataPath_RF_bus_selected_win_data_459_port, 
                           Q(714) => DataPath_RF_bus_selected_win_data_458_port
                           , Q(713) => 
                           DataPath_RF_bus_selected_win_data_457_port, Q(712) 
                           => DataPath_RF_bus_selected_win_data_456_port, 
                           Q(711) => DataPath_RF_bus_selected_win_data_455_port
                           , Q(710) => 
                           DataPath_RF_bus_selected_win_data_454_port, Q(709) 
                           => DataPath_RF_bus_selected_win_data_453_port, 
                           Q(708) => DataPath_RF_bus_selected_win_data_452_port
                           , Q(707) => 
                           DataPath_RF_bus_selected_win_data_451_port, Q(706) 
                           => DataPath_RF_bus_selected_win_data_450_port, 
                           Q(705) => DataPath_RF_bus_selected_win_data_449_port
                           , Q(704) => 
                           DataPath_RF_bus_selected_win_data_448_port, Q(703) 
                           => DataPath_RF_bus_selected_win_data_447_port, 
                           Q(702) => DataPath_RF_bus_selected_win_data_446_port
                           , Q(701) => 
                           DataPath_RF_bus_selected_win_data_445_port, Q(700) 
                           => DataPath_RF_bus_selected_win_data_444_port, 
                           Q(699) => DataPath_RF_bus_selected_win_data_443_port
                           , Q(698) => 
                           DataPath_RF_bus_selected_win_data_442_port, Q(697) 
                           => DataPath_RF_bus_selected_win_data_441_port, 
                           Q(696) => DataPath_RF_bus_selected_win_data_440_port
                           , Q(695) => 
                           DataPath_RF_bus_selected_win_data_439_port, Q(694) 
                           => DataPath_RF_bus_selected_win_data_438_port, 
                           Q(693) => DataPath_RF_bus_selected_win_data_437_port
                           , Q(692) => 
                           DataPath_RF_bus_selected_win_data_436_port, Q(691) 
                           => DataPath_RF_bus_selected_win_data_435_port, 
                           Q(690) => DataPath_RF_bus_selected_win_data_434_port
                           , Q(689) => 
                           DataPath_RF_bus_selected_win_data_433_port, Q(688) 
                           => DataPath_RF_bus_selected_win_data_432_port, 
                           Q(687) => DataPath_RF_bus_selected_win_data_431_port
                           , Q(686) => 
                           DataPath_RF_bus_selected_win_data_430_port, Q(685) 
                           => DataPath_RF_bus_selected_win_data_429_port, 
                           Q(684) => DataPath_RF_bus_selected_win_data_428_port
                           , Q(683) => 
                           DataPath_RF_bus_selected_win_data_427_port, Q(682) 
                           => DataPath_RF_bus_selected_win_data_426_port, 
                           Q(681) => DataPath_RF_bus_selected_win_data_425_port
                           , Q(680) => 
                           DataPath_RF_bus_selected_win_data_424_port, Q(679) 
                           => DataPath_RF_bus_selected_win_data_423_port, 
                           Q(678) => DataPath_RF_bus_selected_win_data_422_port
                           , Q(677) => 
                           DataPath_RF_bus_selected_win_data_421_port, Q(676) 
                           => DataPath_RF_bus_selected_win_data_420_port, 
                           Q(675) => DataPath_RF_bus_selected_win_data_419_port
                           , Q(674) => 
                           DataPath_RF_bus_selected_win_data_418_port, Q(673) 
                           => DataPath_RF_bus_selected_win_data_417_port, 
                           Q(672) => DataPath_RF_bus_selected_win_data_416_port
                           , Q(671) => 
                           DataPath_RF_bus_selected_win_data_415_port, Q(670) 
                           => DataPath_RF_bus_selected_win_data_414_port, 
                           Q(669) => DataPath_RF_bus_selected_win_data_413_port
                           , Q(668) => 
                           DataPath_RF_bus_selected_win_data_412_port, Q(667) 
                           => DataPath_RF_bus_selected_win_data_411_port, 
                           Q(666) => DataPath_RF_bus_selected_win_data_410_port
                           , Q(665) => 
                           DataPath_RF_bus_selected_win_data_409_port, Q(664) 
                           => DataPath_RF_bus_selected_win_data_408_port, 
                           Q(663) => DataPath_RF_bus_selected_win_data_407_port
                           , Q(662) => 
                           DataPath_RF_bus_selected_win_data_406_port, Q(661) 
                           => DataPath_RF_bus_selected_win_data_405_port, 
                           Q(660) => DataPath_RF_bus_selected_win_data_404_port
                           , Q(659) => 
                           DataPath_RF_bus_selected_win_data_403_port, Q(658) 
                           => DataPath_RF_bus_selected_win_data_402_port, 
                           Q(657) => DataPath_RF_bus_selected_win_data_401_port
                           , Q(656) => 
                           DataPath_RF_bus_selected_win_data_400_port, Q(655) 
                           => DataPath_RF_bus_selected_win_data_399_port, 
                           Q(654) => DataPath_RF_bus_selected_win_data_398_port
                           , Q(653) => 
                           DataPath_RF_bus_selected_win_data_397_port, Q(652) 
                           => DataPath_RF_bus_selected_win_data_396_port, 
                           Q(651) => DataPath_RF_bus_selected_win_data_395_port
                           , Q(650) => 
                           DataPath_RF_bus_selected_win_data_394_port, Q(649) 
                           => DataPath_RF_bus_selected_win_data_393_port, 
                           Q(648) => DataPath_RF_bus_selected_win_data_392_port
                           , Q(647) => 
                           DataPath_RF_bus_selected_win_data_391_port, Q(646) 
                           => DataPath_RF_bus_selected_win_data_390_port, 
                           Q(645) => DataPath_RF_bus_selected_win_data_389_port
                           , Q(644) => 
                           DataPath_RF_bus_selected_win_data_388_port, Q(643) 
                           => DataPath_RF_bus_selected_win_data_387_port, 
                           Q(642) => DataPath_RF_bus_selected_win_data_386_port
                           , Q(641) => 
                           DataPath_RF_bus_selected_win_data_385_port, Q(640) 
                           => DataPath_RF_bus_selected_win_data_384_port, 
                           Q(639) => DataPath_RF_bus_selected_win_data_383_port
                           , Q(638) => 
                           DataPath_RF_bus_selected_win_data_382_port, Q(637) 
                           => DataPath_RF_bus_selected_win_data_381_port, 
                           Q(636) => DataPath_RF_bus_selected_win_data_380_port
                           , Q(635) => 
                           DataPath_RF_bus_selected_win_data_379_port, Q(634) 
                           => DataPath_RF_bus_selected_win_data_378_port, 
                           Q(633) => DataPath_RF_bus_selected_win_data_377_port
                           , Q(632) => 
                           DataPath_RF_bus_selected_win_data_376_port, Q(631) 
                           => DataPath_RF_bus_selected_win_data_375_port, 
                           Q(630) => DataPath_RF_bus_selected_win_data_374_port
                           , Q(629) => 
                           DataPath_RF_bus_selected_win_data_373_port, Q(628) 
                           => DataPath_RF_bus_selected_win_data_372_port, 
                           Q(627) => DataPath_RF_bus_selected_win_data_371_port
                           , Q(626) => 
                           DataPath_RF_bus_selected_win_data_370_port, Q(625) 
                           => DataPath_RF_bus_selected_win_data_369_port, 
                           Q(624) => DataPath_RF_bus_selected_win_data_368_port
                           , Q(623) => 
                           DataPath_RF_bus_selected_win_data_367_port, Q(622) 
                           => DataPath_RF_bus_selected_win_data_366_port, 
                           Q(621) => DataPath_RF_bus_selected_win_data_365_port
                           , Q(620) => 
                           DataPath_RF_bus_selected_win_data_364_port, Q(619) 
                           => DataPath_RF_bus_selected_win_data_363_port, 
                           Q(618) => DataPath_RF_bus_selected_win_data_362_port
                           , Q(617) => 
                           DataPath_RF_bus_selected_win_data_361_port, Q(616) 
                           => DataPath_RF_bus_selected_win_data_360_port, 
                           Q(615) => DataPath_RF_bus_selected_win_data_359_port
                           , Q(614) => 
                           DataPath_RF_bus_selected_win_data_358_port, Q(613) 
                           => DataPath_RF_bus_selected_win_data_357_port, 
                           Q(612) => DataPath_RF_bus_selected_win_data_356_port
                           , Q(611) => 
                           DataPath_RF_bus_selected_win_data_355_port, Q(610) 
                           => DataPath_RF_bus_selected_win_data_354_port, 
                           Q(609) => DataPath_RF_bus_selected_win_data_353_port
                           , Q(608) => 
                           DataPath_RF_bus_selected_win_data_352_port, Q(607) 
                           => DataPath_RF_bus_selected_win_data_351_port, 
                           Q(606) => DataPath_RF_bus_selected_win_data_350_port
                           , Q(605) => 
                           DataPath_RF_bus_selected_win_data_349_port, Q(604) 
                           => DataPath_RF_bus_selected_win_data_348_port, 
                           Q(603) => DataPath_RF_bus_selected_win_data_347_port
                           , Q(602) => 
                           DataPath_RF_bus_selected_win_data_346_port, Q(601) 
                           => DataPath_RF_bus_selected_win_data_345_port, 
                           Q(600) => DataPath_RF_bus_selected_win_data_344_port
                           , Q(599) => 
                           DataPath_RF_bus_selected_win_data_343_port, Q(598) 
                           => DataPath_RF_bus_selected_win_data_342_port, 
                           Q(597) => DataPath_RF_bus_selected_win_data_341_port
                           , Q(596) => 
                           DataPath_RF_bus_selected_win_data_340_port, Q(595) 
                           => DataPath_RF_bus_selected_win_data_339_port, 
                           Q(594) => DataPath_RF_bus_selected_win_data_338_port
                           , Q(593) => 
                           DataPath_RF_bus_selected_win_data_337_port, Q(592) 
                           => DataPath_RF_bus_selected_win_data_336_port, 
                           Q(591) => DataPath_RF_bus_selected_win_data_335_port
                           , Q(590) => 
                           DataPath_RF_bus_selected_win_data_334_port, Q(589) 
                           => DataPath_RF_bus_selected_win_data_333_port, 
                           Q(588) => DataPath_RF_bus_selected_win_data_332_port
                           , Q(587) => 
                           DataPath_RF_bus_selected_win_data_331_port, Q(586) 
                           => DataPath_RF_bus_selected_win_data_330_port, 
                           Q(585) => DataPath_RF_bus_selected_win_data_329_port
                           , Q(584) => 
                           DataPath_RF_bus_selected_win_data_328_port, Q(583) 
                           => DataPath_RF_bus_selected_win_data_327_port, 
                           Q(582) => DataPath_RF_bus_selected_win_data_326_port
                           , Q(581) => 
                           DataPath_RF_bus_selected_win_data_325_port, Q(580) 
                           => DataPath_RF_bus_selected_win_data_324_port, 
                           Q(579) => DataPath_RF_bus_selected_win_data_323_port
                           , Q(578) => 
                           DataPath_RF_bus_selected_win_data_322_port, Q(577) 
                           => DataPath_RF_bus_selected_win_data_321_port, 
                           Q(576) => DataPath_RF_bus_selected_win_data_320_port
                           , Q(575) => 
                           DataPath_RF_bus_selected_win_data_319_port, Q(574) 
                           => DataPath_RF_bus_selected_win_data_318_port, 
                           Q(573) => DataPath_RF_bus_selected_win_data_317_port
                           , Q(572) => 
                           DataPath_RF_bus_selected_win_data_316_port, Q(571) 
                           => DataPath_RF_bus_selected_win_data_315_port, 
                           Q(570) => DataPath_RF_bus_selected_win_data_314_port
                           , Q(569) => 
                           DataPath_RF_bus_selected_win_data_313_port, Q(568) 
                           => DataPath_RF_bus_selected_win_data_312_port, 
                           Q(567) => DataPath_RF_bus_selected_win_data_311_port
                           , Q(566) => 
                           DataPath_RF_bus_selected_win_data_310_port, Q(565) 
                           => DataPath_RF_bus_selected_win_data_309_port, 
                           Q(564) => DataPath_RF_bus_selected_win_data_308_port
                           , Q(563) => 
                           DataPath_RF_bus_selected_win_data_307_port, Q(562) 
                           => DataPath_RF_bus_selected_win_data_306_port, 
                           Q(561) => DataPath_RF_bus_selected_win_data_305_port
                           , Q(560) => 
                           DataPath_RF_bus_selected_win_data_304_port, Q(559) 
                           => DataPath_RF_bus_selected_win_data_303_port, 
                           Q(558) => DataPath_RF_bus_selected_win_data_302_port
                           , Q(557) => 
                           DataPath_RF_bus_selected_win_data_301_port, Q(556) 
                           => DataPath_RF_bus_selected_win_data_300_port, 
                           Q(555) => DataPath_RF_bus_selected_win_data_299_port
                           , Q(554) => 
                           DataPath_RF_bus_selected_win_data_298_port, Q(553) 
                           => DataPath_RF_bus_selected_win_data_297_port, 
                           Q(552) => DataPath_RF_bus_selected_win_data_296_port
                           , Q(551) => 
                           DataPath_RF_bus_selected_win_data_295_port, Q(550) 
                           => DataPath_RF_bus_selected_win_data_294_port, 
                           Q(549) => DataPath_RF_bus_selected_win_data_293_port
                           , Q(548) => 
                           DataPath_RF_bus_selected_win_data_292_port, Q(547) 
                           => DataPath_RF_bus_selected_win_data_291_port, 
                           Q(546) => DataPath_RF_bus_selected_win_data_290_port
                           , Q(545) => 
                           DataPath_RF_bus_selected_win_data_289_port, Q(544) 
                           => DataPath_RF_bus_selected_win_data_288_port, 
                           Q(543) => DataPath_RF_bus_selected_win_data_287_port
                           , Q(542) => 
                           DataPath_RF_bus_selected_win_data_286_port, Q(541) 
                           => DataPath_RF_bus_selected_win_data_285_port, 
                           Q(540) => DataPath_RF_bus_selected_win_data_284_port
                           , Q(539) => 
                           DataPath_RF_bus_selected_win_data_283_port, Q(538) 
                           => DataPath_RF_bus_selected_win_data_282_port, 
                           Q(537) => DataPath_RF_bus_selected_win_data_281_port
                           , Q(536) => 
                           DataPath_RF_bus_selected_win_data_280_port, Q(535) 
                           => DataPath_RF_bus_selected_win_data_279_port, 
                           Q(534) => DataPath_RF_bus_selected_win_data_278_port
                           , Q(533) => 
                           DataPath_RF_bus_selected_win_data_277_port, Q(532) 
                           => DataPath_RF_bus_selected_win_data_276_port, 
                           Q(531) => DataPath_RF_bus_selected_win_data_275_port
                           , Q(530) => 
                           DataPath_RF_bus_selected_win_data_274_port, Q(529) 
                           => DataPath_RF_bus_selected_win_data_273_port, 
                           Q(528) => DataPath_RF_bus_selected_win_data_272_port
                           , Q(527) => 
                           DataPath_RF_bus_selected_win_data_271_port, Q(526) 
                           => DataPath_RF_bus_selected_win_data_270_port, 
                           Q(525) => DataPath_RF_bus_selected_win_data_269_port
                           , Q(524) => 
                           DataPath_RF_bus_selected_win_data_268_port, Q(523) 
                           => DataPath_RF_bus_selected_win_data_267_port, 
                           Q(522) => DataPath_RF_bus_selected_win_data_266_port
                           , Q(521) => 
                           DataPath_RF_bus_selected_win_data_265_port, Q(520) 
                           => DataPath_RF_bus_selected_win_data_264_port, 
                           Q(519) => DataPath_RF_bus_selected_win_data_263_port
                           , Q(518) => 
                           DataPath_RF_bus_selected_win_data_262_port, Q(517) 
                           => DataPath_RF_bus_selected_win_data_261_port, 
                           Q(516) => DataPath_RF_bus_selected_win_data_260_port
                           , Q(515) => 
                           DataPath_RF_bus_selected_win_data_259_port, Q(514) 
                           => DataPath_RF_bus_selected_win_data_258_port, 
                           Q(513) => DataPath_RF_bus_selected_win_data_257_port
                           , Q(512) => 
                           DataPath_RF_bus_selected_win_data_256_port, Q(511) 
                           => DataPath_RF_bus_selected_win_data_255_port, 
                           Q(510) => DataPath_RF_bus_selected_win_data_254_port
                           , Q(509) => 
                           DataPath_RF_bus_selected_win_data_253_port, Q(508) 
                           => DataPath_RF_bus_selected_win_data_252_port, 
                           Q(507) => DataPath_RF_bus_selected_win_data_251_port
                           , Q(506) => 
                           DataPath_RF_bus_selected_win_data_250_port, Q(505) 
                           => DataPath_RF_bus_selected_win_data_249_port, 
                           Q(504) => DataPath_RF_bus_selected_win_data_248_port
                           , Q(503) => 
                           DataPath_RF_bus_selected_win_data_247_port, Q(502) 
                           => DataPath_RF_bus_selected_win_data_246_port, 
                           Q(501) => DataPath_RF_bus_selected_win_data_245_port
                           , Q(500) => 
                           DataPath_RF_bus_selected_win_data_244_port, Q(499) 
                           => DataPath_RF_bus_selected_win_data_243_port, 
                           Q(498) => DataPath_RF_bus_selected_win_data_242_port
                           , Q(497) => 
                           DataPath_RF_bus_selected_win_data_241_port, Q(496) 
                           => DataPath_RF_bus_selected_win_data_240_port, 
                           Q(495) => DataPath_RF_bus_selected_win_data_239_port
                           , Q(494) => 
                           DataPath_RF_bus_selected_win_data_238_port, Q(493) 
                           => DataPath_RF_bus_selected_win_data_237_port, 
                           Q(492) => DataPath_RF_bus_selected_win_data_236_port
                           , Q(491) => 
                           DataPath_RF_bus_selected_win_data_235_port, Q(490) 
                           => DataPath_RF_bus_selected_win_data_234_port, 
                           Q(489) => DataPath_RF_bus_selected_win_data_233_port
                           , Q(488) => 
                           DataPath_RF_bus_selected_win_data_232_port, Q(487) 
                           => DataPath_RF_bus_selected_win_data_231_port, 
                           Q(486) => DataPath_RF_bus_selected_win_data_230_port
                           , Q(485) => 
                           DataPath_RF_bus_selected_win_data_229_port, Q(484) 
                           => DataPath_RF_bus_selected_win_data_228_port, 
                           Q(483) => DataPath_RF_bus_selected_win_data_227_port
                           , Q(482) => 
                           DataPath_RF_bus_selected_win_data_226_port, Q(481) 
                           => DataPath_RF_bus_selected_win_data_225_port, 
                           Q(480) => DataPath_RF_bus_selected_win_data_224_port
                           , Q(479) => 
                           DataPath_RF_bus_selected_win_data_223_port, Q(478) 
                           => DataPath_RF_bus_selected_win_data_222_port, 
                           Q(477) => DataPath_RF_bus_selected_win_data_221_port
                           , Q(476) => 
                           DataPath_RF_bus_selected_win_data_220_port, Q(475) 
                           => DataPath_RF_bus_selected_win_data_219_port, 
                           Q(474) => DataPath_RF_bus_selected_win_data_218_port
                           , Q(473) => 
                           DataPath_RF_bus_selected_win_data_217_port, Q(472) 
                           => DataPath_RF_bus_selected_win_data_216_port, 
                           Q(471) => DataPath_RF_bus_selected_win_data_215_port
                           , Q(470) => 
                           DataPath_RF_bus_selected_win_data_214_port, Q(469) 
                           => DataPath_RF_bus_selected_win_data_213_port, 
                           Q(468) => DataPath_RF_bus_selected_win_data_212_port
                           , Q(467) => 
                           DataPath_RF_bus_selected_win_data_211_port, Q(466) 
                           => DataPath_RF_bus_selected_win_data_210_port, 
                           Q(465) => DataPath_RF_bus_selected_win_data_209_port
                           , Q(464) => 
                           DataPath_RF_bus_selected_win_data_208_port, Q(463) 
                           => DataPath_RF_bus_selected_win_data_207_port, 
                           Q(462) => DataPath_RF_bus_selected_win_data_206_port
                           , Q(461) => 
                           DataPath_RF_bus_selected_win_data_205_port, Q(460) 
                           => DataPath_RF_bus_selected_win_data_204_port, 
                           Q(459) => DataPath_RF_bus_selected_win_data_203_port
                           , Q(458) => 
                           DataPath_RF_bus_selected_win_data_202_port, Q(457) 
                           => DataPath_RF_bus_selected_win_data_201_port, 
                           Q(456) => DataPath_RF_bus_selected_win_data_200_port
                           , Q(455) => 
                           DataPath_RF_bus_selected_win_data_199_port, Q(454) 
                           => DataPath_RF_bus_selected_win_data_198_port, 
                           Q(453) => DataPath_RF_bus_selected_win_data_197_port
                           , Q(452) => 
                           DataPath_RF_bus_selected_win_data_196_port, Q(451) 
                           => DataPath_RF_bus_selected_win_data_195_port, 
                           Q(450) => DataPath_RF_bus_selected_win_data_194_port
                           , Q(449) => 
                           DataPath_RF_bus_selected_win_data_193_port, Q(448) 
                           => DataPath_RF_bus_selected_win_data_192_port, 
                           Q(447) => DataPath_RF_bus_selected_win_data_191_port
                           , Q(446) => 
                           DataPath_RF_bus_selected_win_data_190_port, Q(445) 
                           => DataPath_RF_bus_selected_win_data_189_port, 
                           Q(444) => DataPath_RF_bus_selected_win_data_188_port
                           , Q(443) => 
                           DataPath_RF_bus_selected_win_data_187_port, Q(442) 
                           => DataPath_RF_bus_selected_win_data_186_port, 
                           Q(441) => DataPath_RF_bus_selected_win_data_185_port
                           , Q(440) => 
                           DataPath_RF_bus_selected_win_data_184_port, Q(439) 
                           => DataPath_RF_bus_selected_win_data_183_port, 
                           Q(438) => DataPath_RF_bus_selected_win_data_182_port
                           , Q(437) => 
                           DataPath_RF_bus_selected_win_data_181_port, Q(436) 
                           => DataPath_RF_bus_selected_win_data_180_port, 
                           Q(435) => DataPath_RF_bus_selected_win_data_179_port
                           , Q(434) => 
                           DataPath_RF_bus_selected_win_data_178_port, Q(433) 
                           => DataPath_RF_bus_selected_win_data_177_port, 
                           Q(432) => DataPath_RF_bus_selected_win_data_176_port
                           , Q(431) => 
                           DataPath_RF_bus_selected_win_data_175_port, Q(430) 
                           => DataPath_RF_bus_selected_win_data_174_port, 
                           Q(429) => DataPath_RF_bus_selected_win_data_173_port
                           , Q(428) => 
                           DataPath_RF_bus_selected_win_data_172_port, Q(427) 
                           => DataPath_RF_bus_selected_win_data_171_port, 
                           Q(426) => DataPath_RF_bus_selected_win_data_170_port
                           , Q(425) => 
                           DataPath_RF_bus_selected_win_data_169_port, Q(424) 
                           => DataPath_RF_bus_selected_win_data_168_port, 
                           Q(423) => DataPath_RF_bus_selected_win_data_167_port
                           , Q(422) => 
                           DataPath_RF_bus_selected_win_data_166_port, Q(421) 
                           => DataPath_RF_bus_selected_win_data_165_port, 
                           Q(420) => DataPath_RF_bus_selected_win_data_164_port
                           , Q(419) => 
                           DataPath_RF_bus_selected_win_data_163_port, Q(418) 
                           => DataPath_RF_bus_selected_win_data_162_port, 
                           Q(417) => DataPath_RF_bus_selected_win_data_161_port
                           , Q(416) => 
                           DataPath_RF_bus_selected_win_data_160_port, Q(415) 
                           => DataPath_RF_bus_selected_win_data_159_port, 
                           Q(414) => DataPath_RF_bus_selected_win_data_158_port
                           , Q(413) => 
                           DataPath_RF_bus_selected_win_data_157_port, Q(412) 
                           => DataPath_RF_bus_selected_win_data_156_port, 
                           Q(411) => DataPath_RF_bus_selected_win_data_155_port
                           , Q(410) => 
                           DataPath_RF_bus_selected_win_data_154_port, Q(409) 
                           => DataPath_RF_bus_selected_win_data_153_port, 
                           Q(408) => DataPath_RF_bus_selected_win_data_152_port
                           , Q(407) => 
                           DataPath_RF_bus_selected_win_data_151_port, Q(406) 
                           => DataPath_RF_bus_selected_win_data_150_port, 
                           Q(405) => DataPath_RF_bus_selected_win_data_149_port
                           , Q(404) => 
                           DataPath_RF_bus_selected_win_data_148_port, Q(403) 
                           => DataPath_RF_bus_selected_win_data_147_port, 
                           Q(402) => DataPath_RF_bus_selected_win_data_146_port
                           , Q(401) => 
                           DataPath_RF_bus_selected_win_data_145_port, Q(400) 
                           => DataPath_RF_bus_selected_win_data_144_port, 
                           Q(399) => DataPath_RF_bus_selected_win_data_143_port
                           , Q(398) => 
                           DataPath_RF_bus_selected_win_data_142_port, Q(397) 
                           => DataPath_RF_bus_selected_win_data_141_port, 
                           Q(396) => DataPath_RF_bus_selected_win_data_140_port
                           , Q(395) => 
                           DataPath_RF_bus_selected_win_data_139_port, Q(394) 
                           => DataPath_RF_bus_selected_win_data_138_port, 
                           Q(393) => DataPath_RF_bus_selected_win_data_137_port
                           , Q(392) => 
                           DataPath_RF_bus_selected_win_data_136_port, Q(391) 
                           => DataPath_RF_bus_selected_win_data_135_port, 
                           Q(390) => DataPath_RF_bus_selected_win_data_134_port
                           , Q(389) => 
                           DataPath_RF_bus_selected_win_data_133_port, Q(388) 
                           => DataPath_RF_bus_selected_win_data_132_port, 
                           Q(387) => DataPath_RF_bus_selected_win_data_131_port
                           , Q(386) => 
                           DataPath_RF_bus_selected_win_data_130_port, Q(385) 
                           => DataPath_RF_bus_selected_win_data_129_port, 
                           Q(384) => DataPath_RF_bus_selected_win_data_128_port
                           , Q(383) => 
                           DataPath_RF_bus_selected_win_data_127_port, Q(382) 
                           => DataPath_RF_bus_selected_win_data_126_port, 
                           Q(381) => DataPath_RF_bus_selected_win_data_125_port
                           , Q(380) => 
                           DataPath_RF_bus_selected_win_data_124_port, Q(379) 
                           => DataPath_RF_bus_selected_win_data_123_port, 
                           Q(378) => DataPath_RF_bus_selected_win_data_122_port
                           , Q(377) => 
                           DataPath_RF_bus_selected_win_data_121_port, Q(376) 
                           => DataPath_RF_bus_selected_win_data_120_port, 
                           Q(375) => DataPath_RF_bus_selected_win_data_119_port
                           , Q(374) => 
                           DataPath_RF_bus_selected_win_data_118_port, Q(373) 
                           => DataPath_RF_bus_selected_win_data_117_port, 
                           Q(372) => DataPath_RF_bus_selected_win_data_116_port
                           , Q(371) => 
                           DataPath_RF_bus_selected_win_data_115_port, Q(370) 
                           => DataPath_RF_bus_selected_win_data_114_port, 
                           Q(369) => DataPath_RF_bus_selected_win_data_113_port
                           , Q(368) => 
                           DataPath_RF_bus_selected_win_data_112_port, Q(367) 
                           => DataPath_RF_bus_selected_win_data_111_port, 
                           Q(366) => DataPath_RF_bus_selected_win_data_110_port
                           , Q(365) => 
                           DataPath_RF_bus_selected_win_data_109_port, Q(364) 
                           => DataPath_RF_bus_selected_win_data_108_port, 
                           Q(363) => DataPath_RF_bus_selected_win_data_107_port
                           , Q(362) => 
                           DataPath_RF_bus_selected_win_data_106_port, Q(361) 
                           => DataPath_RF_bus_selected_win_data_105_port, 
                           Q(360) => DataPath_RF_bus_selected_win_data_104_port
                           , Q(359) => 
                           DataPath_RF_bus_selected_win_data_103_port, Q(358) 
                           => DataPath_RF_bus_selected_win_data_102_port, 
                           Q(357) => DataPath_RF_bus_selected_win_data_101_port
                           , Q(356) => 
                           DataPath_RF_bus_selected_win_data_100_port, Q(355) 
                           => DataPath_RF_bus_selected_win_data_99_port, Q(354)
                           => DataPath_RF_bus_selected_win_data_98_port, Q(353)
                           => DataPath_RF_bus_selected_win_data_97_port, Q(352)
                           => DataPath_RF_bus_selected_win_data_96_port, Q(351)
                           => DataPath_RF_bus_selected_win_data_95_port, Q(350)
                           => DataPath_RF_bus_selected_win_data_94_port, Q(349)
                           => DataPath_RF_bus_selected_win_data_93_port, Q(348)
                           => DataPath_RF_bus_selected_win_data_92_port, Q(347)
                           => DataPath_RF_bus_selected_win_data_91_port, Q(346)
                           => DataPath_RF_bus_selected_win_data_90_port, Q(345)
                           => DataPath_RF_bus_selected_win_data_89_port, Q(344)
                           => DataPath_RF_bus_selected_win_data_88_port, Q(343)
                           => DataPath_RF_bus_selected_win_data_87_port, Q(342)
                           => DataPath_RF_bus_selected_win_data_86_port, Q(341)
                           => DataPath_RF_bus_selected_win_data_85_port, Q(340)
                           => DataPath_RF_bus_selected_win_data_84_port, Q(339)
                           => DataPath_RF_bus_selected_win_data_83_port, Q(338)
                           => DataPath_RF_bus_selected_win_data_82_port, Q(337)
                           => DataPath_RF_bus_selected_win_data_81_port, Q(336)
                           => DataPath_RF_bus_selected_win_data_80_port, Q(335)
                           => DataPath_RF_bus_selected_win_data_79_port, Q(334)
                           => DataPath_RF_bus_selected_win_data_78_port, Q(333)
                           => DataPath_RF_bus_selected_win_data_77_port, Q(332)
                           => DataPath_RF_bus_selected_win_data_76_port, Q(331)
                           => DataPath_RF_bus_selected_win_data_75_port, Q(330)
                           => DataPath_RF_bus_selected_win_data_74_port, Q(329)
                           => DataPath_RF_bus_selected_win_data_73_port, Q(328)
                           => DataPath_RF_bus_selected_win_data_72_port, Q(327)
                           => DataPath_RF_bus_selected_win_data_71_port, Q(326)
                           => DataPath_RF_bus_selected_win_data_70_port, Q(325)
                           => DataPath_RF_bus_selected_win_data_69_port, Q(324)
                           => DataPath_RF_bus_selected_win_data_68_port, Q(323)
                           => DataPath_RF_bus_selected_win_data_67_port, Q(322)
                           => DataPath_RF_bus_selected_win_data_66_port, Q(321)
                           => DataPath_RF_bus_selected_win_data_65_port, Q(320)
                           => DataPath_RF_bus_selected_win_data_64_port, Q(319)
                           => DataPath_RF_bus_selected_win_data_63_port, Q(318)
                           => DataPath_RF_bus_selected_win_data_62_port, Q(317)
                           => DataPath_RF_bus_selected_win_data_61_port, Q(316)
                           => DataPath_RF_bus_selected_win_data_60_port, Q(315)
                           => DataPath_RF_bus_selected_win_data_59_port, Q(314)
                           => DataPath_RF_bus_selected_win_data_58_port, Q(313)
                           => DataPath_RF_bus_selected_win_data_57_port, Q(312)
                           => DataPath_RF_bus_selected_win_data_56_port, Q(311)
                           => DataPath_RF_bus_selected_win_data_55_port, Q(310)
                           => DataPath_RF_bus_selected_win_data_54_port, Q(309)
                           => DataPath_RF_bus_selected_win_data_53_port, Q(308)
                           => DataPath_RF_bus_selected_win_data_52_port, Q(307)
                           => DataPath_RF_bus_selected_win_data_51_port, Q(306)
                           => DataPath_RF_bus_selected_win_data_50_port, Q(305)
                           => DataPath_RF_bus_selected_win_data_49_port, Q(304)
                           => DataPath_RF_bus_selected_win_data_48_port, Q(303)
                           => DataPath_RF_bus_selected_win_data_47_port, Q(302)
                           => DataPath_RF_bus_selected_win_data_46_port, Q(301)
                           => DataPath_RF_bus_selected_win_data_45_port, Q(300)
                           => DataPath_RF_bus_selected_win_data_44_port, Q(299)
                           => DataPath_RF_bus_selected_win_data_43_port, Q(298)
                           => DataPath_RF_bus_selected_win_data_42_port, Q(297)
                           => DataPath_RF_bus_selected_win_data_41_port, Q(296)
                           => DataPath_RF_bus_selected_win_data_40_port, Q(295)
                           => DataPath_RF_bus_selected_win_data_39_port, Q(294)
                           => DataPath_RF_bus_selected_win_data_38_port, Q(293)
                           => DataPath_RF_bus_selected_win_data_37_port, Q(292)
                           => DataPath_RF_bus_selected_win_data_36_port, Q(291)
                           => DataPath_RF_bus_selected_win_data_35_port, Q(290)
                           => DataPath_RF_bus_selected_win_data_34_port, Q(289)
                           => DataPath_RF_bus_selected_win_data_33_port, Q(288)
                           => DataPath_RF_bus_selected_win_data_32_port, Q(287)
                           => DataPath_RF_bus_selected_win_data_31_port, Q(286)
                           => DataPath_RF_bus_selected_win_data_30_port, Q(285)
                           => DataPath_RF_bus_selected_win_data_29_port, Q(284)
                           => DataPath_RF_bus_selected_win_data_28_port, Q(283)
                           => DataPath_RF_bus_selected_win_data_27_port, Q(282)
                           => DataPath_RF_bus_selected_win_data_26_port, Q(281)
                           => DataPath_RF_bus_selected_win_data_25_port, Q(280)
                           => DataPath_RF_bus_selected_win_data_24_port, Q(279)
                           => DataPath_RF_bus_selected_win_data_23_port, Q(278)
                           => DataPath_RF_bus_selected_win_data_22_port, Q(277)
                           => DataPath_RF_bus_selected_win_data_21_port, Q(276)
                           => DataPath_RF_bus_selected_win_data_20_port, Q(275)
                           => DataPath_RF_bus_selected_win_data_19_port, Q(274)
                           => DataPath_RF_bus_selected_win_data_18_port, Q(273)
                           => DataPath_RF_bus_selected_win_data_17_port, Q(272)
                           => DataPath_RF_bus_selected_win_data_16_port, Q(271)
                           => DataPath_RF_bus_selected_win_data_15_port, Q(270)
                           => DataPath_RF_bus_selected_win_data_14_port, Q(269)
                           => DataPath_RF_bus_selected_win_data_13_port, Q(268)
                           => DataPath_RF_bus_selected_win_data_12_port, Q(267)
                           => DataPath_RF_bus_selected_win_data_11_port, Q(266)
                           => DataPath_RF_bus_selected_win_data_10_port, Q(265)
                           => DataPath_RF_bus_selected_win_data_9_port, Q(264) 
                           => DataPath_RF_bus_selected_win_data_8_port, Q(263) 
                           => DataPath_RF_bus_selected_win_data_7_port, Q(262) 
                           => DataPath_RF_bus_selected_win_data_6_port, Q(261) 
                           => DataPath_RF_bus_selected_win_data_5_port, Q(260) 
                           => DataPath_RF_bus_selected_win_data_4_port, Q(259) 
                           => DataPath_RF_bus_selected_win_data_3_port, Q(258) 
                           => DataPath_RF_bus_selected_win_data_2_port, Q(257) 
                           => DataPath_RF_bus_selected_win_data_1_port, Q(256) 
                           => DataPath_RF_bus_selected_win_data_0_port, Q(255) 
                           => DataPath_RF_bus_complete_win_data_255_port, 
                           Q(254) => DataPath_RF_bus_complete_win_data_254_port
                           , Q(253) => 
                           DataPath_RF_bus_complete_win_data_253_port, Q(252) 
                           => DataPath_RF_bus_complete_win_data_252_port, 
                           Q(251) => DataPath_RF_bus_complete_win_data_251_port
                           , Q(250) => 
                           DataPath_RF_bus_complete_win_data_250_port, Q(249) 
                           => DataPath_RF_bus_complete_win_data_249_port, 
                           Q(248) => DataPath_RF_bus_complete_win_data_248_port
                           , Q(247) => 
                           DataPath_RF_bus_complete_win_data_247_port, Q(246) 
                           => DataPath_RF_bus_complete_win_data_246_port, 
                           Q(245) => DataPath_RF_bus_complete_win_data_245_port
                           , Q(244) => 
                           DataPath_RF_bus_complete_win_data_244_port, Q(243) 
                           => DataPath_RF_bus_complete_win_data_243_port, 
                           Q(242) => DataPath_RF_bus_complete_win_data_242_port
                           , Q(241) => 
                           DataPath_RF_bus_complete_win_data_241_port, Q(240) 
                           => DataPath_RF_bus_complete_win_data_240_port, 
                           Q(239) => DataPath_RF_bus_complete_win_data_239_port
                           , Q(238) => 
                           DataPath_RF_bus_complete_win_data_238_port, Q(237) 
                           => DataPath_RF_bus_complete_win_data_237_port, 
                           Q(236) => DataPath_RF_bus_complete_win_data_236_port
                           , Q(235) => 
                           DataPath_RF_bus_complete_win_data_235_port, Q(234) 
                           => DataPath_RF_bus_complete_win_data_234_port, 
                           Q(233) => DataPath_RF_bus_complete_win_data_233_port
                           , Q(232) => 
                           DataPath_RF_bus_complete_win_data_232_port, Q(231) 
                           => DataPath_RF_bus_complete_win_data_231_port, 
                           Q(230) => DataPath_RF_bus_complete_win_data_230_port
                           , Q(229) => 
                           DataPath_RF_bus_complete_win_data_229_port, Q(228) 
                           => DataPath_RF_bus_complete_win_data_228_port, 
                           Q(227) => DataPath_RF_bus_complete_win_data_227_port
                           , Q(226) => 
                           DataPath_RF_bus_complete_win_data_226_port, Q(225) 
                           => DataPath_RF_bus_complete_win_data_225_port, 
                           Q(224) => DataPath_RF_bus_complete_win_data_224_port
                           , Q(223) => 
                           DataPath_RF_bus_complete_win_data_223_port, Q(222) 
                           => DataPath_RF_bus_complete_win_data_222_port, 
                           Q(221) => DataPath_RF_bus_complete_win_data_221_port
                           , Q(220) => 
                           DataPath_RF_bus_complete_win_data_220_port, Q(219) 
                           => DataPath_RF_bus_complete_win_data_219_port, 
                           Q(218) => DataPath_RF_bus_complete_win_data_218_port
                           , Q(217) => 
                           DataPath_RF_bus_complete_win_data_217_port, Q(216) 
                           => DataPath_RF_bus_complete_win_data_216_port, 
                           Q(215) => DataPath_RF_bus_complete_win_data_215_port
                           , Q(214) => 
                           DataPath_RF_bus_complete_win_data_214_port, Q(213) 
                           => DataPath_RF_bus_complete_win_data_213_port, 
                           Q(212) => DataPath_RF_bus_complete_win_data_212_port
                           , Q(211) => 
                           DataPath_RF_bus_complete_win_data_211_port, Q(210) 
                           => DataPath_RF_bus_complete_win_data_210_port, 
                           Q(209) => DataPath_RF_bus_complete_win_data_209_port
                           , Q(208) => 
                           DataPath_RF_bus_complete_win_data_208_port, Q(207) 
                           => DataPath_RF_bus_complete_win_data_207_port, 
                           Q(206) => DataPath_RF_bus_complete_win_data_206_port
                           , Q(205) => 
                           DataPath_RF_bus_complete_win_data_205_port, Q(204) 
                           => DataPath_RF_bus_complete_win_data_204_port, 
                           Q(203) => DataPath_RF_bus_complete_win_data_203_port
                           , Q(202) => 
                           DataPath_RF_bus_complete_win_data_202_port, Q(201) 
                           => DataPath_RF_bus_complete_win_data_201_port, 
                           Q(200) => DataPath_RF_bus_complete_win_data_200_port
                           , Q(199) => 
                           DataPath_RF_bus_complete_win_data_199_port, Q(198) 
                           => DataPath_RF_bus_complete_win_data_198_port, 
                           Q(197) => DataPath_RF_bus_complete_win_data_197_port
                           , Q(196) => 
                           DataPath_RF_bus_complete_win_data_196_port, Q(195) 
                           => DataPath_RF_bus_complete_win_data_195_port, 
                           Q(194) => DataPath_RF_bus_complete_win_data_194_port
                           , Q(193) => 
                           DataPath_RF_bus_complete_win_data_193_port, Q(192) 
                           => DataPath_RF_bus_complete_win_data_192_port, 
                           Q(191) => DataPath_RF_bus_complete_win_data_191_port
                           , Q(190) => 
                           DataPath_RF_bus_complete_win_data_190_port, Q(189) 
                           => DataPath_RF_bus_complete_win_data_189_port, 
                           Q(188) => DataPath_RF_bus_complete_win_data_188_port
                           , Q(187) => 
                           DataPath_RF_bus_complete_win_data_187_port, Q(186) 
                           => DataPath_RF_bus_complete_win_data_186_port, 
                           Q(185) => DataPath_RF_bus_complete_win_data_185_port
                           , Q(184) => 
                           DataPath_RF_bus_complete_win_data_184_port, Q(183) 
                           => DataPath_RF_bus_complete_win_data_183_port, 
                           Q(182) => DataPath_RF_bus_complete_win_data_182_port
                           , Q(181) => 
                           DataPath_RF_bus_complete_win_data_181_port, Q(180) 
                           => DataPath_RF_bus_complete_win_data_180_port, 
                           Q(179) => DataPath_RF_bus_complete_win_data_179_port
                           , Q(178) => 
                           DataPath_RF_bus_complete_win_data_178_port, Q(177) 
                           => DataPath_RF_bus_complete_win_data_177_port, 
                           Q(176) => DataPath_RF_bus_complete_win_data_176_port
                           , Q(175) => 
                           DataPath_RF_bus_complete_win_data_175_port, Q(174) 
                           => DataPath_RF_bus_complete_win_data_174_port, 
                           Q(173) => DataPath_RF_bus_complete_win_data_173_port
                           , Q(172) => 
                           DataPath_RF_bus_complete_win_data_172_port, Q(171) 
                           => DataPath_RF_bus_complete_win_data_171_port, 
                           Q(170) => DataPath_RF_bus_complete_win_data_170_port
                           , Q(169) => 
                           DataPath_RF_bus_complete_win_data_169_port, Q(168) 
                           => DataPath_RF_bus_complete_win_data_168_port, 
                           Q(167) => DataPath_RF_bus_complete_win_data_167_port
                           , Q(166) => 
                           DataPath_RF_bus_complete_win_data_166_port, Q(165) 
                           => DataPath_RF_bus_complete_win_data_165_port, 
                           Q(164) => DataPath_RF_bus_complete_win_data_164_port
                           , Q(163) => 
                           DataPath_RF_bus_complete_win_data_163_port, Q(162) 
                           => DataPath_RF_bus_complete_win_data_162_port, 
                           Q(161) => DataPath_RF_bus_complete_win_data_161_port
                           , Q(160) => 
                           DataPath_RF_bus_complete_win_data_160_port, Q(159) 
                           => DataPath_RF_bus_complete_win_data_159_port, 
                           Q(158) => DataPath_RF_bus_complete_win_data_158_port
                           , Q(157) => 
                           DataPath_RF_bus_complete_win_data_157_port, Q(156) 
                           => DataPath_RF_bus_complete_win_data_156_port, 
                           Q(155) => DataPath_RF_bus_complete_win_data_155_port
                           , Q(154) => 
                           DataPath_RF_bus_complete_win_data_154_port, Q(153) 
                           => DataPath_RF_bus_complete_win_data_153_port, 
                           Q(152) => DataPath_RF_bus_complete_win_data_152_port
                           , Q(151) => 
                           DataPath_RF_bus_complete_win_data_151_port, Q(150) 
                           => DataPath_RF_bus_complete_win_data_150_port, 
                           Q(149) => DataPath_RF_bus_complete_win_data_149_port
                           , Q(148) => 
                           DataPath_RF_bus_complete_win_data_148_port, Q(147) 
                           => DataPath_RF_bus_complete_win_data_147_port, 
                           Q(146) => DataPath_RF_bus_complete_win_data_146_port
                           , Q(145) => 
                           DataPath_RF_bus_complete_win_data_145_port, Q(144) 
                           => DataPath_RF_bus_complete_win_data_144_port, 
                           Q(143) => DataPath_RF_bus_complete_win_data_143_port
                           , Q(142) => 
                           DataPath_RF_bus_complete_win_data_142_port, Q(141) 
                           => DataPath_RF_bus_complete_win_data_141_port, 
                           Q(140) => DataPath_RF_bus_complete_win_data_140_port
                           , Q(139) => 
                           DataPath_RF_bus_complete_win_data_139_port, Q(138) 
                           => DataPath_RF_bus_complete_win_data_138_port, 
                           Q(137) => DataPath_RF_bus_complete_win_data_137_port
                           , Q(136) => 
                           DataPath_RF_bus_complete_win_data_136_port, Q(135) 
                           => DataPath_RF_bus_complete_win_data_135_port, 
                           Q(134) => DataPath_RF_bus_complete_win_data_134_port
                           , Q(133) => 
                           DataPath_RF_bus_complete_win_data_133_port, Q(132) 
                           => DataPath_RF_bus_complete_win_data_132_port, 
                           Q(131) => DataPath_RF_bus_complete_win_data_131_port
                           , Q(130) => 
                           DataPath_RF_bus_complete_win_data_130_port, Q(129) 
                           => DataPath_RF_bus_complete_win_data_129_port, 
                           Q(128) => DataPath_RF_bus_complete_win_data_128_port
                           , Q(127) => 
                           DataPath_RF_bus_complete_win_data_127_port, Q(126) 
                           => DataPath_RF_bus_complete_win_data_126_port, 
                           Q(125) => DataPath_RF_bus_complete_win_data_125_port
                           , Q(124) => 
                           DataPath_RF_bus_complete_win_data_124_port, Q(123) 
                           => DataPath_RF_bus_complete_win_data_123_port, 
                           Q(122) => DataPath_RF_bus_complete_win_data_122_port
                           , Q(121) => 
                           DataPath_RF_bus_complete_win_data_121_port, Q(120) 
                           => DataPath_RF_bus_complete_win_data_120_port, 
                           Q(119) => DataPath_RF_bus_complete_win_data_119_port
                           , Q(118) => 
                           DataPath_RF_bus_complete_win_data_118_port, Q(117) 
                           => DataPath_RF_bus_complete_win_data_117_port, 
                           Q(116) => DataPath_RF_bus_complete_win_data_116_port
                           , Q(115) => 
                           DataPath_RF_bus_complete_win_data_115_port, Q(114) 
                           => DataPath_RF_bus_complete_win_data_114_port, 
                           Q(113) => DataPath_RF_bus_complete_win_data_113_port
                           , Q(112) => 
                           DataPath_RF_bus_complete_win_data_112_port, Q(111) 
                           => DataPath_RF_bus_complete_win_data_111_port, 
                           Q(110) => DataPath_RF_bus_complete_win_data_110_port
                           , Q(109) => 
                           DataPath_RF_bus_complete_win_data_109_port, Q(108) 
                           => DataPath_RF_bus_complete_win_data_108_port, 
                           Q(107) => DataPath_RF_bus_complete_win_data_107_port
                           , Q(106) => 
                           DataPath_RF_bus_complete_win_data_106_port, Q(105) 
                           => DataPath_RF_bus_complete_win_data_105_port, 
                           Q(104) => DataPath_RF_bus_complete_win_data_104_port
                           , Q(103) => 
                           DataPath_RF_bus_complete_win_data_103_port, Q(102) 
                           => DataPath_RF_bus_complete_win_data_102_port, 
                           Q(101) => DataPath_RF_bus_complete_win_data_101_port
                           , Q(100) => 
                           DataPath_RF_bus_complete_win_data_100_port, Q(99) =>
                           DataPath_RF_bus_complete_win_data_99_port, Q(98) => 
                           DataPath_RF_bus_complete_win_data_98_port, Q(97) => 
                           DataPath_RF_bus_complete_win_data_97_port, Q(96) => 
                           DataPath_RF_bus_complete_win_data_96_port, Q(95) => 
                           DataPath_RF_bus_complete_win_data_95_port, Q(94) => 
                           DataPath_RF_bus_complete_win_data_94_port, Q(93) => 
                           DataPath_RF_bus_complete_win_data_93_port, Q(92) => 
                           DataPath_RF_bus_complete_win_data_92_port, Q(91) => 
                           DataPath_RF_bus_complete_win_data_91_port, Q(90) => 
                           DataPath_RF_bus_complete_win_data_90_port, Q(89) => 
                           DataPath_RF_bus_complete_win_data_89_port, Q(88) => 
                           DataPath_RF_bus_complete_win_data_88_port, Q(87) => 
                           DataPath_RF_bus_complete_win_data_87_port, Q(86) => 
                           DataPath_RF_bus_complete_win_data_86_port, Q(85) => 
                           DataPath_RF_bus_complete_win_data_85_port, Q(84) => 
                           DataPath_RF_bus_complete_win_data_84_port, Q(83) => 
                           DataPath_RF_bus_complete_win_data_83_port, Q(82) => 
                           DataPath_RF_bus_complete_win_data_82_port, Q(81) => 
                           DataPath_RF_bus_complete_win_data_81_port, Q(80) => 
                           DataPath_RF_bus_complete_win_data_80_port, Q(79) => 
                           DataPath_RF_bus_complete_win_data_79_port, Q(78) => 
                           DataPath_RF_bus_complete_win_data_78_port, Q(77) => 
                           DataPath_RF_bus_complete_win_data_77_port, Q(76) => 
                           DataPath_RF_bus_complete_win_data_76_port, Q(75) => 
                           DataPath_RF_bus_complete_win_data_75_port, Q(74) => 
                           DataPath_RF_bus_complete_win_data_74_port, Q(73) => 
                           DataPath_RF_bus_complete_win_data_73_port, Q(72) => 
                           DataPath_RF_bus_complete_win_data_72_port, Q(71) => 
                           DataPath_RF_bus_complete_win_data_71_port, Q(70) => 
                           DataPath_RF_bus_complete_win_data_70_port, Q(69) => 
                           DataPath_RF_bus_complete_win_data_69_port, Q(68) => 
                           DataPath_RF_bus_complete_win_data_68_port, Q(67) => 
                           DataPath_RF_bus_complete_win_data_67_port, Q(66) => 
                           DataPath_RF_bus_complete_win_data_66_port, Q(65) => 
                           DataPath_RF_bus_complete_win_data_65_port, Q(64) => 
                           DataPath_RF_bus_complete_win_data_64_port, Q(63) => 
                           DataPath_RF_bus_complete_win_data_63_port, Q(62) => 
                           DataPath_RF_bus_complete_win_data_62_port, Q(61) => 
                           DataPath_RF_bus_complete_win_data_61_port, Q(60) => 
                           DataPath_RF_bus_complete_win_data_60_port, Q(59) => 
                           DataPath_RF_bus_complete_win_data_59_port, Q(58) => 
                           DataPath_RF_bus_complete_win_data_58_port, Q(57) => 
                           DataPath_RF_bus_complete_win_data_57_port, Q(56) => 
                           DataPath_RF_bus_complete_win_data_56_port, Q(55) => 
                           DataPath_RF_bus_complete_win_data_55_port, Q(54) => 
                           DataPath_RF_bus_complete_win_data_54_port, Q(53) => 
                           DataPath_RF_bus_complete_win_data_53_port, Q(52) => 
                           DataPath_RF_bus_complete_win_data_52_port, Q(51) => 
                           DataPath_RF_bus_complete_win_data_51_port, Q(50) => 
                           DataPath_RF_bus_complete_win_data_50_port, Q(49) => 
                           DataPath_RF_bus_complete_win_data_49_port, Q(48) => 
                           DataPath_RF_bus_complete_win_data_48_port, Q(47) => 
                           DataPath_RF_bus_complete_win_data_47_port, Q(46) => 
                           DataPath_RF_bus_complete_win_data_46_port, Q(45) => 
                           DataPath_RF_bus_complete_win_data_45_port, Q(44) => 
                           DataPath_RF_bus_complete_win_data_44_port, Q(43) => 
                           DataPath_RF_bus_complete_win_data_43_port, Q(42) => 
                           DataPath_RF_bus_complete_win_data_42_port, Q(41) => 
                           DataPath_RF_bus_complete_win_data_41_port, Q(40) => 
                           DataPath_RF_bus_complete_win_data_40_port, Q(39) => 
                           DataPath_RF_bus_complete_win_data_39_port, Q(38) => 
                           DataPath_RF_bus_complete_win_data_38_port, Q(37) => 
                           DataPath_RF_bus_complete_win_data_37_port, Q(36) => 
                           DataPath_RF_bus_complete_win_data_36_port, Q(35) => 
                           DataPath_RF_bus_complete_win_data_35_port, Q(34) => 
                           DataPath_RF_bus_complete_win_data_34_port, Q(33) => 
                           DataPath_RF_bus_complete_win_data_33_port, Q(32) => 
                           DataPath_RF_bus_complete_win_data_32_port, Q(31) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(30) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(29) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(28) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(27) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(26) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(25) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(24) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(23) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(22) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(21) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(20) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(19) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(18) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(17) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(16) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(15) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(14) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(13) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(12) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(11) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(10) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(9) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(8) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(7) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(6) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(5) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(4) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(3) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(2) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(1) => 
                           DataPath_RF_bus_complete_win_data_0_port, Q(0) => 
                           DataPath_RF_bus_complete_win_data_0_port, Y(31) => 
                           DataPath_RF_internal_out1_31_port, Y(30) => 
                           DataPath_RF_internal_out1_30_port, Y(29) => 
                           DataPath_RF_internal_out1_29_port, Y(28) => 
                           DataPath_RF_internal_out1_28_port, Y(27) => 
                           DataPath_RF_internal_out1_27_port, Y(26) => 
                           DataPath_RF_internal_out1_26_port, Y(25) => 
                           DataPath_RF_internal_out1_25_port, Y(24) => 
                           DataPath_RF_internal_out1_24_port, Y(23) => 
                           DataPath_RF_internal_out1_23_port, Y(22) => 
                           DataPath_RF_internal_out1_22_port, Y(21) => 
                           DataPath_RF_internal_out1_21_port, Y(20) => 
                           DataPath_RF_internal_out1_20_port, Y(19) => 
                           DataPath_RF_internal_out1_19_port, Y(18) => 
                           DataPath_RF_internal_out1_18_port, Y(17) => 
                           DataPath_RF_internal_out1_17_port, Y(16) => 
                           DataPath_RF_internal_out1_16_port, Y(15) => 
                           DataPath_RF_internal_out1_15_port, Y(14) => 
                           DataPath_RF_internal_out1_14_port, Y(13) => 
                           DataPath_RF_internal_out1_13_port, Y(12) => 
                           DataPath_RF_internal_out1_12_port, Y(11) => 
                           DataPath_RF_internal_out1_11_port, Y(10) => 
                           DataPath_RF_internal_out1_10_port, Y(9) => 
                           DataPath_RF_internal_out1_9_port, Y(8) => 
                           DataPath_RF_internal_out1_8_port, Y(7) => 
                           DataPath_RF_internal_out1_7_port, Y(6) => 
                           DataPath_RF_internal_out1_6_port, Y(5) => 
                           DataPath_RF_internal_out1_5_port, Y(4) => 
                           DataPath_RF_internal_out1_4_port, Y(3) => 
                           DataPath_RF_internal_out1_3_port, Y(2) => 
                           DataPath_RF_internal_out1_2_port, Y(1) => 
                           DataPath_RF_internal_out1_1_port, Y(0) => 
                           DataPath_RF_internal_out1_0_port);
   DataPath_RF_SEL_BLK : select_block_NBIT_DATA32_N8_F5 port map( regs(2559) =>
                           DataPath_RF_bus_reg_dataout_2559_port, regs(2558) =>
                           DataPath_RF_bus_reg_dataout_2558_port, regs(2557) =>
                           DataPath_RF_bus_reg_dataout_2557_port, regs(2556) =>
                           DataPath_RF_bus_reg_dataout_2556_port, regs(2555) =>
                           DataPath_RF_bus_reg_dataout_2555_port, regs(2554) =>
                           DataPath_RF_bus_reg_dataout_2554_port, regs(2553) =>
                           DataPath_RF_bus_reg_dataout_2553_port, regs(2552) =>
                           DataPath_RF_bus_reg_dataout_2552_port, regs(2551) =>
                           DataPath_RF_bus_reg_dataout_2551_port, regs(2550) =>
                           DataPath_RF_bus_reg_dataout_2550_port, regs(2549) =>
                           DataPath_RF_bus_reg_dataout_2549_port, regs(2548) =>
                           DataPath_RF_bus_reg_dataout_2548_port, regs(2547) =>
                           DataPath_RF_bus_reg_dataout_2547_port, regs(2546) =>
                           DataPath_RF_bus_reg_dataout_2546_port, regs(2545) =>
                           DataPath_RF_bus_reg_dataout_2545_port, regs(2544) =>
                           DataPath_RF_bus_reg_dataout_2544_port, regs(2543) =>
                           DataPath_RF_bus_reg_dataout_2543_port, regs(2542) =>
                           DataPath_RF_bus_reg_dataout_2542_port, regs(2541) =>
                           DataPath_RF_bus_reg_dataout_2541_port, regs(2540) =>
                           DataPath_RF_bus_reg_dataout_2540_port, regs(2539) =>
                           DataPath_RF_bus_reg_dataout_2539_port, regs(2538) =>
                           DataPath_RF_bus_reg_dataout_2538_port, regs(2537) =>
                           DataPath_RF_bus_reg_dataout_2537_port, regs(2536) =>
                           DataPath_RF_bus_reg_dataout_2536_port, regs(2535) =>
                           DataPath_RF_bus_reg_dataout_2535_port, regs(2534) =>
                           DataPath_RF_bus_reg_dataout_2534_port, regs(2533) =>
                           DataPath_RF_bus_reg_dataout_2533_port, regs(2532) =>
                           DataPath_RF_bus_reg_dataout_2532_port, regs(2531) =>
                           DataPath_RF_bus_reg_dataout_2531_port, regs(2530) =>
                           DataPath_RF_bus_reg_dataout_2530_port, regs(2529) =>
                           DataPath_RF_bus_reg_dataout_2529_port, regs(2528) =>
                           DataPath_RF_bus_reg_dataout_2528_port, regs(2527) =>
                           DataPath_RF_bus_reg_dataout_2527_port, regs(2526) =>
                           DataPath_RF_bus_reg_dataout_2526_port, regs(2525) =>
                           DataPath_RF_bus_reg_dataout_2525_port, regs(2524) =>
                           DataPath_RF_bus_reg_dataout_2524_port, regs(2523) =>
                           DataPath_RF_bus_reg_dataout_2523_port, regs(2522) =>
                           DataPath_RF_bus_reg_dataout_2522_port, regs(2521) =>
                           DataPath_RF_bus_reg_dataout_2521_port, regs(2520) =>
                           DataPath_RF_bus_reg_dataout_2520_port, regs(2519) =>
                           DataPath_RF_bus_reg_dataout_2519_port, regs(2518) =>
                           DataPath_RF_bus_reg_dataout_2518_port, regs(2517) =>
                           DataPath_RF_bus_reg_dataout_2517_port, regs(2516) =>
                           DataPath_RF_bus_reg_dataout_2516_port, regs(2515) =>
                           DataPath_RF_bus_reg_dataout_2515_port, regs(2514) =>
                           DataPath_RF_bus_reg_dataout_2514_port, regs(2513) =>
                           DataPath_RF_bus_reg_dataout_2513_port, regs(2512) =>
                           DataPath_RF_bus_reg_dataout_2512_port, regs(2511) =>
                           DataPath_RF_bus_reg_dataout_2511_port, regs(2510) =>
                           DataPath_RF_bus_reg_dataout_2510_port, regs(2509) =>
                           DataPath_RF_bus_reg_dataout_2509_port, regs(2508) =>
                           DataPath_RF_bus_reg_dataout_2508_port, regs(2507) =>
                           DataPath_RF_bus_reg_dataout_2507_port, regs(2506) =>
                           DataPath_RF_bus_reg_dataout_2506_port, regs(2505) =>
                           DataPath_RF_bus_reg_dataout_2505_port, regs(2504) =>
                           DataPath_RF_bus_reg_dataout_2504_port, regs(2503) =>
                           DataPath_RF_bus_reg_dataout_2503_port, regs(2502) =>
                           DataPath_RF_bus_reg_dataout_2502_port, regs(2501) =>
                           DataPath_RF_bus_reg_dataout_2501_port, regs(2500) =>
                           DataPath_RF_bus_reg_dataout_2500_port, regs(2499) =>
                           DataPath_RF_bus_reg_dataout_2499_port, regs(2498) =>
                           DataPath_RF_bus_reg_dataout_2498_port, regs(2497) =>
                           DataPath_RF_bus_reg_dataout_2497_port, regs(2496) =>
                           DataPath_RF_bus_reg_dataout_2496_port, regs(2495) =>
                           DataPath_RF_bus_reg_dataout_2495_port, regs(2494) =>
                           DataPath_RF_bus_reg_dataout_2494_port, regs(2493) =>
                           DataPath_RF_bus_reg_dataout_2493_port, regs(2492) =>
                           DataPath_RF_bus_reg_dataout_2492_port, regs(2491) =>
                           DataPath_RF_bus_reg_dataout_2491_port, regs(2490) =>
                           DataPath_RF_bus_reg_dataout_2490_port, regs(2489) =>
                           DataPath_RF_bus_reg_dataout_2489_port, regs(2488) =>
                           DataPath_RF_bus_reg_dataout_2488_port, regs(2487) =>
                           DataPath_RF_bus_reg_dataout_2487_port, regs(2486) =>
                           DataPath_RF_bus_reg_dataout_2486_port, regs(2485) =>
                           DataPath_RF_bus_reg_dataout_2485_port, regs(2484) =>
                           DataPath_RF_bus_reg_dataout_2484_port, regs(2483) =>
                           DataPath_RF_bus_reg_dataout_2483_port, regs(2482) =>
                           DataPath_RF_bus_reg_dataout_2482_port, regs(2481) =>
                           DataPath_RF_bus_reg_dataout_2481_port, regs(2480) =>
                           DataPath_RF_bus_reg_dataout_2480_port, regs(2479) =>
                           DataPath_RF_bus_reg_dataout_2479_port, regs(2478) =>
                           DataPath_RF_bus_reg_dataout_2478_port, regs(2477) =>
                           DataPath_RF_bus_reg_dataout_2477_port, regs(2476) =>
                           DataPath_RF_bus_reg_dataout_2476_port, regs(2475) =>
                           DataPath_RF_bus_reg_dataout_2475_port, regs(2474) =>
                           DataPath_RF_bus_reg_dataout_2474_port, regs(2473) =>
                           DataPath_RF_bus_reg_dataout_2473_port, regs(2472) =>
                           DataPath_RF_bus_reg_dataout_2472_port, regs(2471) =>
                           DataPath_RF_bus_reg_dataout_2471_port, regs(2470) =>
                           DataPath_RF_bus_reg_dataout_2470_port, regs(2469) =>
                           DataPath_RF_bus_reg_dataout_2469_port, regs(2468) =>
                           DataPath_RF_bus_reg_dataout_2468_port, regs(2467) =>
                           DataPath_RF_bus_reg_dataout_2467_port, regs(2466) =>
                           DataPath_RF_bus_reg_dataout_2466_port, regs(2465) =>
                           DataPath_RF_bus_reg_dataout_2465_port, regs(2464) =>
                           DataPath_RF_bus_reg_dataout_2464_port, regs(2463) =>
                           DataPath_RF_bus_reg_dataout_2463_port, regs(2462) =>
                           DataPath_RF_bus_reg_dataout_2462_port, regs(2461) =>
                           DataPath_RF_bus_reg_dataout_2461_port, regs(2460) =>
                           DataPath_RF_bus_reg_dataout_2460_port, regs(2459) =>
                           DataPath_RF_bus_reg_dataout_2459_port, regs(2458) =>
                           DataPath_RF_bus_reg_dataout_2458_port, regs(2457) =>
                           DataPath_RF_bus_reg_dataout_2457_port, regs(2456) =>
                           DataPath_RF_bus_reg_dataout_2456_port, regs(2455) =>
                           DataPath_RF_bus_reg_dataout_2455_port, regs(2454) =>
                           DataPath_RF_bus_reg_dataout_2454_port, regs(2453) =>
                           DataPath_RF_bus_reg_dataout_2453_port, regs(2452) =>
                           DataPath_RF_bus_reg_dataout_2452_port, regs(2451) =>
                           DataPath_RF_bus_reg_dataout_2451_port, regs(2450) =>
                           DataPath_RF_bus_reg_dataout_2450_port, regs(2449) =>
                           DataPath_RF_bus_reg_dataout_2449_port, regs(2448) =>
                           DataPath_RF_bus_reg_dataout_2448_port, regs(2447) =>
                           DataPath_RF_bus_reg_dataout_2447_port, regs(2446) =>
                           DataPath_RF_bus_reg_dataout_2446_port, regs(2445) =>
                           DataPath_RF_bus_reg_dataout_2445_port, regs(2444) =>
                           DataPath_RF_bus_reg_dataout_2444_port, regs(2443) =>
                           DataPath_RF_bus_reg_dataout_2443_port, regs(2442) =>
                           DataPath_RF_bus_reg_dataout_2442_port, regs(2441) =>
                           DataPath_RF_bus_reg_dataout_2441_port, regs(2440) =>
                           DataPath_RF_bus_reg_dataout_2440_port, regs(2439) =>
                           DataPath_RF_bus_reg_dataout_2439_port, regs(2438) =>
                           DataPath_RF_bus_reg_dataout_2438_port, regs(2437) =>
                           DataPath_RF_bus_reg_dataout_2437_port, regs(2436) =>
                           DataPath_RF_bus_reg_dataout_2436_port, regs(2435) =>
                           DataPath_RF_bus_reg_dataout_2435_port, regs(2434) =>
                           DataPath_RF_bus_reg_dataout_2434_port, regs(2433) =>
                           DataPath_RF_bus_reg_dataout_2433_port, regs(2432) =>
                           DataPath_RF_bus_reg_dataout_2432_port, regs(2431) =>
                           DataPath_RF_bus_reg_dataout_2431_port, regs(2430) =>
                           DataPath_RF_bus_reg_dataout_2430_port, regs(2429) =>
                           DataPath_RF_bus_reg_dataout_2429_port, regs(2428) =>
                           DataPath_RF_bus_reg_dataout_2428_port, regs(2427) =>
                           DataPath_RF_bus_reg_dataout_2427_port, regs(2426) =>
                           DataPath_RF_bus_reg_dataout_2426_port, regs(2425) =>
                           DataPath_RF_bus_reg_dataout_2425_port, regs(2424) =>
                           DataPath_RF_bus_reg_dataout_2424_port, regs(2423) =>
                           DataPath_RF_bus_reg_dataout_2423_port, regs(2422) =>
                           DataPath_RF_bus_reg_dataout_2422_port, regs(2421) =>
                           DataPath_RF_bus_reg_dataout_2421_port, regs(2420) =>
                           DataPath_RF_bus_reg_dataout_2420_port, regs(2419) =>
                           DataPath_RF_bus_reg_dataout_2419_port, regs(2418) =>
                           DataPath_RF_bus_reg_dataout_2418_port, regs(2417) =>
                           DataPath_RF_bus_reg_dataout_2417_port, regs(2416) =>
                           DataPath_RF_bus_reg_dataout_2416_port, regs(2415) =>
                           DataPath_RF_bus_reg_dataout_2415_port, regs(2414) =>
                           DataPath_RF_bus_reg_dataout_2414_port, regs(2413) =>
                           DataPath_RF_bus_reg_dataout_2413_port, regs(2412) =>
                           DataPath_RF_bus_reg_dataout_2412_port, regs(2411) =>
                           DataPath_RF_bus_reg_dataout_2411_port, regs(2410) =>
                           DataPath_RF_bus_reg_dataout_2410_port, regs(2409) =>
                           DataPath_RF_bus_reg_dataout_2409_port, regs(2408) =>
                           DataPath_RF_bus_reg_dataout_2408_port, regs(2407) =>
                           DataPath_RF_bus_reg_dataout_2407_port, regs(2406) =>
                           DataPath_RF_bus_reg_dataout_2406_port, regs(2405) =>
                           DataPath_RF_bus_reg_dataout_2405_port, regs(2404) =>
                           DataPath_RF_bus_reg_dataout_2404_port, regs(2403) =>
                           DataPath_RF_bus_reg_dataout_2403_port, regs(2402) =>
                           DataPath_RF_bus_reg_dataout_2402_port, regs(2401) =>
                           DataPath_RF_bus_reg_dataout_2401_port, regs(2400) =>
                           DataPath_RF_bus_reg_dataout_2400_port, regs(2399) =>
                           DataPath_RF_bus_reg_dataout_2399_port, regs(2398) =>
                           DataPath_RF_bus_reg_dataout_2398_port, regs(2397) =>
                           DataPath_RF_bus_reg_dataout_2397_port, regs(2396) =>
                           DataPath_RF_bus_reg_dataout_2396_port, regs(2395) =>
                           DataPath_RF_bus_reg_dataout_2395_port, regs(2394) =>
                           DataPath_RF_bus_reg_dataout_2394_port, regs(2393) =>
                           DataPath_RF_bus_reg_dataout_2393_port, regs(2392) =>
                           DataPath_RF_bus_reg_dataout_2392_port, regs(2391) =>
                           DataPath_RF_bus_reg_dataout_2391_port, regs(2390) =>
                           DataPath_RF_bus_reg_dataout_2390_port, regs(2389) =>
                           DataPath_RF_bus_reg_dataout_2389_port, regs(2388) =>
                           DataPath_RF_bus_reg_dataout_2388_port, regs(2387) =>
                           DataPath_RF_bus_reg_dataout_2387_port, regs(2386) =>
                           DataPath_RF_bus_reg_dataout_2386_port, regs(2385) =>
                           DataPath_RF_bus_reg_dataout_2385_port, regs(2384) =>
                           DataPath_RF_bus_reg_dataout_2384_port, regs(2383) =>
                           DataPath_RF_bus_reg_dataout_2383_port, regs(2382) =>
                           DataPath_RF_bus_reg_dataout_2382_port, regs(2381) =>
                           DataPath_RF_bus_reg_dataout_2381_port, regs(2380) =>
                           DataPath_RF_bus_reg_dataout_2380_port, regs(2379) =>
                           DataPath_RF_bus_reg_dataout_2379_port, regs(2378) =>
                           DataPath_RF_bus_reg_dataout_2378_port, regs(2377) =>
                           DataPath_RF_bus_reg_dataout_2377_port, regs(2376) =>
                           DataPath_RF_bus_reg_dataout_2376_port, regs(2375) =>
                           DataPath_RF_bus_reg_dataout_2375_port, regs(2374) =>
                           DataPath_RF_bus_reg_dataout_2374_port, regs(2373) =>
                           DataPath_RF_bus_reg_dataout_2373_port, regs(2372) =>
                           DataPath_RF_bus_reg_dataout_2372_port, regs(2371) =>
                           DataPath_RF_bus_reg_dataout_2371_port, regs(2370) =>
                           DataPath_RF_bus_reg_dataout_2370_port, regs(2369) =>
                           DataPath_RF_bus_reg_dataout_2369_port, regs(2368) =>
                           DataPath_RF_bus_reg_dataout_2368_port, regs(2367) =>
                           DataPath_RF_bus_reg_dataout_2367_port, regs(2366) =>
                           DataPath_RF_bus_reg_dataout_2366_port, regs(2365) =>
                           DataPath_RF_bus_reg_dataout_2365_port, regs(2364) =>
                           DataPath_RF_bus_reg_dataout_2364_port, regs(2363) =>
                           DataPath_RF_bus_reg_dataout_2363_port, regs(2362) =>
                           DataPath_RF_bus_reg_dataout_2362_port, regs(2361) =>
                           DataPath_RF_bus_reg_dataout_2361_port, regs(2360) =>
                           DataPath_RF_bus_reg_dataout_2360_port, regs(2359) =>
                           DataPath_RF_bus_reg_dataout_2359_port, regs(2358) =>
                           DataPath_RF_bus_reg_dataout_2358_port, regs(2357) =>
                           DataPath_RF_bus_reg_dataout_2357_port, regs(2356) =>
                           DataPath_RF_bus_reg_dataout_2356_port, regs(2355) =>
                           DataPath_RF_bus_reg_dataout_2355_port, regs(2354) =>
                           DataPath_RF_bus_reg_dataout_2354_port, regs(2353) =>
                           DataPath_RF_bus_reg_dataout_2353_port, regs(2352) =>
                           DataPath_RF_bus_reg_dataout_2352_port, regs(2351) =>
                           DataPath_RF_bus_reg_dataout_2351_port, regs(2350) =>
                           DataPath_RF_bus_reg_dataout_2350_port, regs(2349) =>
                           DataPath_RF_bus_reg_dataout_2349_port, regs(2348) =>
                           DataPath_RF_bus_reg_dataout_2348_port, regs(2347) =>
                           DataPath_RF_bus_reg_dataout_2347_port, regs(2346) =>
                           DataPath_RF_bus_reg_dataout_2346_port, regs(2345) =>
                           DataPath_RF_bus_reg_dataout_2345_port, regs(2344) =>
                           DataPath_RF_bus_reg_dataout_2344_port, regs(2343) =>
                           DataPath_RF_bus_reg_dataout_2343_port, regs(2342) =>
                           DataPath_RF_bus_reg_dataout_2342_port, regs(2341) =>
                           DataPath_RF_bus_reg_dataout_2341_port, regs(2340) =>
                           DataPath_RF_bus_reg_dataout_2340_port, regs(2339) =>
                           DataPath_RF_bus_reg_dataout_2339_port, regs(2338) =>
                           DataPath_RF_bus_reg_dataout_2338_port, regs(2337) =>
                           DataPath_RF_bus_reg_dataout_2337_port, regs(2336) =>
                           DataPath_RF_bus_reg_dataout_2336_port, regs(2335) =>
                           DataPath_RF_bus_reg_dataout_2335_port, regs(2334) =>
                           DataPath_RF_bus_reg_dataout_2334_port, regs(2333) =>
                           DataPath_RF_bus_reg_dataout_2333_port, regs(2332) =>
                           DataPath_RF_bus_reg_dataout_2332_port, regs(2331) =>
                           DataPath_RF_bus_reg_dataout_2331_port, regs(2330) =>
                           DataPath_RF_bus_reg_dataout_2330_port, regs(2329) =>
                           DataPath_RF_bus_reg_dataout_2329_port, regs(2328) =>
                           DataPath_RF_bus_reg_dataout_2328_port, regs(2327) =>
                           DataPath_RF_bus_reg_dataout_2327_port, regs(2326) =>
                           DataPath_RF_bus_reg_dataout_2326_port, regs(2325) =>
                           DataPath_RF_bus_reg_dataout_2325_port, regs(2324) =>
                           DataPath_RF_bus_reg_dataout_2324_port, regs(2323) =>
                           DataPath_RF_bus_reg_dataout_2323_port, regs(2322) =>
                           DataPath_RF_bus_reg_dataout_2322_port, regs(2321) =>
                           DataPath_RF_bus_reg_dataout_2321_port, regs(2320) =>
                           DataPath_RF_bus_reg_dataout_2320_port, regs(2319) =>
                           DataPath_RF_bus_reg_dataout_2319_port, regs(2318) =>
                           DataPath_RF_bus_reg_dataout_2318_port, regs(2317) =>
                           DataPath_RF_bus_reg_dataout_2317_port, regs(2316) =>
                           DataPath_RF_bus_reg_dataout_2316_port, regs(2315) =>
                           DataPath_RF_bus_reg_dataout_2315_port, regs(2314) =>
                           DataPath_RF_bus_reg_dataout_2314_port, regs(2313) =>
                           DataPath_RF_bus_reg_dataout_2313_port, regs(2312) =>
                           DataPath_RF_bus_reg_dataout_2312_port, regs(2311) =>
                           DataPath_RF_bus_reg_dataout_2311_port, regs(2310) =>
                           DataPath_RF_bus_reg_dataout_2310_port, regs(2309) =>
                           DataPath_RF_bus_reg_dataout_2309_port, regs(2308) =>
                           DataPath_RF_bus_reg_dataout_2308_port, regs(2307) =>
                           DataPath_RF_bus_reg_dataout_2307_port, regs(2306) =>
                           DataPath_RF_bus_reg_dataout_2306_port, regs(2305) =>
                           DataPath_RF_bus_reg_dataout_2305_port, regs(2304) =>
                           DataPath_RF_bus_reg_dataout_2304_port, regs(2303) =>
                           DataPath_RF_bus_reg_dataout_2303_port, regs(2302) =>
                           DataPath_RF_bus_reg_dataout_2302_port, regs(2301) =>
                           DataPath_RF_bus_reg_dataout_2301_port, regs(2300) =>
                           DataPath_RF_bus_reg_dataout_2300_port, regs(2299) =>
                           DataPath_RF_bus_reg_dataout_2299_port, regs(2298) =>
                           DataPath_RF_bus_reg_dataout_2298_port, regs(2297) =>
                           DataPath_RF_bus_reg_dataout_2297_port, regs(2296) =>
                           DataPath_RF_bus_reg_dataout_2296_port, regs(2295) =>
                           DataPath_RF_bus_reg_dataout_2295_port, regs(2294) =>
                           DataPath_RF_bus_reg_dataout_2294_port, regs(2293) =>
                           DataPath_RF_bus_reg_dataout_2293_port, regs(2292) =>
                           DataPath_RF_bus_reg_dataout_2292_port, regs(2291) =>
                           DataPath_RF_bus_reg_dataout_2291_port, regs(2290) =>
                           DataPath_RF_bus_reg_dataout_2290_port, regs(2289) =>
                           DataPath_RF_bus_reg_dataout_2289_port, regs(2288) =>
                           DataPath_RF_bus_reg_dataout_2288_port, regs(2287) =>
                           DataPath_RF_bus_reg_dataout_2287_port, regs(2286) =>
                           DataPath_RF_bus_reg_dataout_2286_port, regs(2285) =>
                           DataPath_RF_bus_reg_dataout_2285_port, regs(2284) =>
                           DataPath_RF_bus_reg_dataout_2284_port, regs(2283) =>
                           DataPath_RF_bus_reg_dataout_2283_port, regs(2282) =>
                           DataPath_RF_bus_reg_dataout_2282_port, regs(2281) =>
                           DataPath_RF_bus_reg_dataout_2281_port, regs(2280) =>
                           DataPath_RF_bus_reg_dataout_2280_port, regs(2279) =>
                           DataPath_RF_bus_reg_dataout_2279_port, regs(2278) =>
                           DataPath_RF_bus_reg_dataout_2278_port, regs(2277) =>
                           DataPath_RF_bus_reg_dataout_2277_port, regs(2276) =>
                           DataPath_RF_bus_reg_dataout_2276_port, regs(2275) =>
                           DataPath_RF_bus_reg_dataout_2275_port, regs(2274) =>
                           DataPath_RF_bus_reg_dataout_2274_port, regs(2273) =>
                           DataPath_RF_bus_reg_dataout_2273_port, regs(2272) =>
                           DataPath_RF_bus_reg_dataout_2272_port, regs(2271) =>
                           DataPath_RF_bus_reg_dataout_2271_port, regs(2270) =>
                           DataPath_RF_bus_reg_dataout_2270_port, regs(2269) =>
                           DataPath_RF_bus_reg_dataout_2269_port, regs(2268) =>
                           DataPath_RF_bus_reg_dataout_2268_port, regs(2267) =>
                           DataPath_RF_bus_reg_dataout_2267_port, regs(2266) =>
                           DataPath_RF_bus_reg_dataout_2266_port, regs(2265) =>
                           DataPath_RF_bus_reg_dataout_2265_port, regs(2264) =>
                           DataPath_RF_bus_reg_dataout_2264_port, regs(2263) =>
                           DataPath_RF_bus_reg_dataout_2263_port, regs(2262) =>
                           DataPath_RF_bus_reg_dataout_2262_port, regs(2261) =>
                           DataPath_RF_bus_reg_dataout_2261_port, regs(2260) =>
                           DataPath_RF_bus_reg_dataout_2260_port, regs(2259) =>
                           DataPath_RF_bus_reg_dataout_2259_port, regs(2258) =>
                           DataPath_RF_bus_reg_dataout_2258_port, regs(2257) =>
                           DataPath_RF_bus_reg_dataout_2257_port, regs(2256) =>
                           DataPath_RF_bus_reg_dataout_2256_port, regs(2255) =>
                           DataPath_RF_bus_reg_dataout_2255_port, regs(2254) =>
                           DataPath_RF_bus_reg_dataout_2254_port, regs(2253) =>
                           DataPath_RF_bus_reg_dataout_2253_port, regs(2252) =>
                           DataPath_RF_bus_reg_dataout_2252_port, regs(2251) =>
                           DataPath_RF_bus_reg_dataout_2251_port, regs(2250) =>
                           DataPath_RF_bus_reg_dataout_2250_port, regs(2249) =>
                           DataPath_RF_bus_reg_dataout_2249_port, regs(2248) =>
                           DataPath_RF_bus_reg_dataout_2248_port, regs(2247) =>
                           DataPath_RF_bus_reg_dataout_2247_port, regs(2246) =>
                           DataPath_RF_bus_reg_dataout_2246_port, regs(2245) =>
                           DataPath_RF_bus_reg_dataout_2245_port, regs(2244) =>
                           DataPath_RF_bus_reg_dataout_2244_port, regs(2243) =>
                           DataPath_RF_bus_reg_dataout_2243_port, regs(2242) =>
                           DataPath_RF_bus_reg_dataout_2242_port, regs(2241) =>
                           DataPath_RF_bus_reg_dataout_2241_port, regs(2240) =>
                           DataPath_RF_bus_reg_dataout_2240_port, regs(2239) =>
                           DataPath_RF_bus_reg_dataout_2239_port, regs(2238) =>
                           DataPath_RF_bus_reg_dataout_2238_port, regs(2237) =>
                           DataPath_RF_bus_reg_dataout_2237_port, regs(2236) =>
                           DataPath_RF_bus_reg_dataout_2236_port, regs(2235) =>
                           DataPath_RF_bus_reg_dataout_2235_port, regs(2234) =>
                           DataPath_RF_bus_reg_dataout_2234_port, regs(2233) =>
                           DataPath_RF_bus_reg_dataout_2233_port, regs(2232) =>
                           DataPath_RF_bus_reg_dataout_2232_port, regs(2231) =>
                           DataPath_RF_bus_reg_dataout_2231_port, regs(2230) =>
                           DataPath_RF_bus_reg_dataout_2230_port, regs(2229) =>
                           DataPath_RF_bus_reg_dataout_2229_port, regs(2228) =>
                           DataPath_RF_bus_reg_dataout_2228_port, regs(2227) =>
                           DataPath_RF_bus_reg_dataout_2227_port, regs(2226) =>
                           DataPath_RF_bus_reg_dataout_2226_port, regs(2225) =>
                           DataPath_RF_bus_reg_dataout_2225_port, regs(2224) =>
                           DataPath_RF_bus_reg_dataout_2224_port, regs(2223) =>
                           DataPath_RF_bus_reg_dataout_2223_port, regs(2222) =>
                           DataPath_RF_bus_reg_dataout_2222_port, regs(2221) =>
                           DataPath_RF_bus_reg_dataout_2221_port, regs(2220) =>
                           DataPath_RF_bus_reg_dataout_2220_port, regs(2219) =>
                           DataPath_RF_bus_reg_dataout_2219_port, regs(2218) =>
                           DataPath_RF_bus_reg_dataout_2218_port, regs(2217) =>
                           DataPath_RF_bus_reg_dataout_2217_port, regs(2216) =>
                           DataPath_RF_bus_reg_dataout_2216_port, regs(2215) =>
                           DataPath_RF_bus_reg_dataout_2215_port, regs(2214) =>
                           DataPath_RF_bus_reg_dataout_2214_port, regs(2213) =>
                           DataPath_RF_bus_reg_dataout_2213_port, regs(2212) =>
                           DataPath_RF_bus_reg_dataout_2212_port, regs(2211) =>
                           DataPath_RF_bus_reg_dataout_2211_port, regs(2210) =>
                           DataPath_RF_bus_reg_dataout_2210_port, regs(2209) =>
                           DataPath_RF_bus_reg_dataout_2209_port, regs(2208) =>
                           DataPath_RF_bus_reg_dataout_2208_port, regs(2207) =>
                           DataPath_RF_bus_reg_dataout_2207_port, regs(2206) =>
                           DataPath_RF_bus_reg_dataout_2206_port, regs(2205) =>
                           DataPath_RF_bus_reg_dataout_2205_port, regs(2204) =>
                           DataPath_RF_bus_reg_dataout_2204_port, regs(2203) =>
                           DataPath_RF_bus_reg_dataout_2203_port, regs(2202) =>
                           DataPath_RF_bus_reg_dataout_2202_port, regs(2201) =>
                           DataPath_RF_bus_reg_dataout_2201_port, regs(2200) =>
                           DataPath_RF_bus_reg_dataout_2200_port, regs(2199) =>
                           DataPath_RF_bus_reg_dataout_2199_port, regs(2198) =>
                           DataPath_RF_bus_reg_dataout_2198_port, regs(2197) =>
                           DataPath_RF_bus_reg_dataout_2197_port, regs(2196) =>
                           DataPath_RF_bus_reg_dataout_2196_port, regs(2195) =>
                           DataPath_RF_bus_reg_dataout_2195_port, regs(2194) =>
                           DataPath_RF_bus_reg_dataout_2194_port, regs(2193) =>
                           DataPath_RF_bus_reg_dataout_2193_port, regs(2192) =>
                           DataPath_RF_bus_reg_dataout_2192_port, regs(2191) =>
                           DataPath_RF_bus_reg_dataout_2191_port, regs(2190) =>
                           DataPath_RF_bus_reg_dataout_2190_port, regs(2189) =>
                           DataPath_RF_bus_reg_dataout_2189_port, regs(2188) =>
                           DataPath_RF_bus_reg_dataout_2188_port, regs(2187) =>
                           DataPath_RF_bus_reg_dataout_2187_port, regs(2186) =>
                           DataPath_RF_bus_reg_dataout_2186_port, regs(2185) =>
                           DataPath_RF_bus_reg_dataout_2185_port, regs(2184) =>
                           DataPath_RF_bus_reg_dataout_2184_port, regs(2183) =>
                           DataPath_RF_bus_reg_dataout_2183_port, regs(2182) =>
                           DataPath_RF_bus_reg_dataout_2182_port, regs(2181) =>
                           DataPath_RF_bus_reg_dataout_2181_port, regs(2180) =>
                           DataPath_RF_bus_reg_dataout_2180_port, regs(2179) =>
                           DataPath_RF_bus_reg_dataout_2179_port, regs(2178) =>
                           DataPath_RF_bus_reg_dataout_2178_port, regs(2177) =>
                           DataPath_RF_bus_reg_dataout_2177_port, regs(2176) =>
                           DataPath_RF_bus_reg_dataout_2176_port, regs(2175) =>
                           DataPath_RF_bus_reg_dataout_2175_port, regs(2174) =>
                           DataPath_RF_bus_reg_dataout_2174_port, regs(2173) =>
                           DataPath_RF_bus_reg_dataout_2173_port, regs(2172) =>
                           DataPath_RF_bus_reg_dataout_2172_port, regs(2171) =>
                           DataPath_RF_bus_reg_dataout_2171_port, regs(2170) =>
                           DataPath_RF_bus_reg_dataout_2170_port, regs(2169) =>
                           DataPath_RF_bus_reg_dataout_2169_port, regs(2168) =>
                           DataPath_RF_bus_reg_dataout_2168_port, regs(2167) =>
                           DataPath_RF_bus_reg_dataout_2167_port, regs(2166) =>
                           DataPath_RF_bus_reg_dataout_2166_port, regs(2165) =>
                           DataPath_RF_bus_reg_dataout_2165_port, regs(2164) =>
                           DataPath_RF_bus_reg_dataout_2164_port, regs(2163) =>
                           DataPath_RF_bus_reg_dataout_2163_port, regs(2162) =>
                           DataPath_RF_bus_reg_dataout_2162_port, regs(2161) =>
                           DataPath_RF_bus_reg_dataout_2161_port, regs(2160) =>
                           DataPath_RF_bus_reg_dataout_2160_port, regs(2159) =>
                           DataPath_RF_bus_reg_dataout_2159_port, regs(2158) =>
                           DataPath_RF_bus_reg_dataout_2158_port, regs(2157) =>
                           DataPath_RF_bus_reg_dataout_2157_port, regs(2156) =>
                           DataPath_RF_bus_reg_dataout_2156_port, regs(2155) =>
                           DataPath_RF_bus_reg_dataout_2155_port, regs(2154) =>
                           DataPath_RF_bus_reg_dataout_2154_port, regs(2153) =>
                           DataPath_RF_bus_reg_dataout_2153_port, regs(2152) =>
                           DataPath_RF_bus_reg_dataout_2152_port, regs(2151) =>
                           DataPath_RF_bus_reg_dataout_2151_port, regs(2150) =>
                           DataPath_RF_bus_reg_dataout_2150_port, regs(2149) =>
                           DataPath_RF_bus_reg_dataout_2149_port, regs(2148) =>
                           DataPath_RF_bus_reg_dataout_2148_port, regs(2147) =>
                           DataPath_RF_bus_reg_dataout_2147_port, regs(2146) =>
                           DataPath_RF_bus_reg_dataout_2146_port, regs(2145) =>
                           DataPath_RF_bus_reg_dataout_2145_port, regs(2144) =>
                           DataPath_RF_bus_reg_dataout_2144_port, regs(2143) =>
                           DataPath_RF_bus_reg_dataout_2143_port, regs(2142) =>
                           DataPath_RF_bus_reg_dataout_2142_port, regs(2141) =>
                           DataPath_RF_bus_reg_dataout_2141_port, regs(2140) =>
                           DataPath_RF_bus_reg_dataout_2140_port, regs(2139) =>
                           DataPath_RF_bus_reg_dataout_2139_port, regs(2138) =>
                           DataPath_RF_bus_reg_dataout_2138_port, regs(2137) =>
                           DataPath_RF_bus_reg_dataout_2137_port, regs(2136) =>
                           DataPath_RF_bus_reg_dataout_2136_port, regs(2135) =>
                           DataPath_RF_bus_reg_dataout_2135_port, regs(2134) =>
                           DataPath_RF_bus_reg_dataout_2134_port, regs(2133) =>
                           DataPath_RF_bus_reg_dataout_2133_port, regs(2132) =>
                           DataPath_RF_bus_reg_dataout_2132_port, regs(2131) =>
                           DataPath_RF_bus_reg_dataout_2131_port, regs(2130) =>
                           DataPath_RF_bus_reg_dataout_2130_port, regs(2129) =>
                           DataPath_RF_bus_reg_dataout_2129_port, regs(2128) =>
                           DataPath_RF_bus_reg_dataout_2128_port, regs(2127) =>
                           DataPath_RF_bus_reg_dataout_2127_port, regs(2126) =>
                           DataPath_RF_bus_reg_dataout_2126_port, regs(2125) =>
                           DataPath_RF_bus_reg_dataout_2125_port, regs(2124) =>
                           DataPath_RF_bus_reg_dataout_2124_port, regs(2123) =>
                           DataPath_RF_bus_reg_dataout_2123_port, regs(2122) =>
                           DataPath_RF_bus_reg_dataout_2122_port, regs(2121) =>
                           DataPath_RF_bus_reg_dataout_2121_port, regs(2120) =>
                           DataPath_RF_bus_reg_dataout_2120_port, regs(2119) =>
                           DataPath_RF_bus_reg_dataout_2119_port, regs(2118) =>
                           DataPath_RF_bus_reg_dataout_2118_port, regs(2117) =>
                           DataPath_RF_bus_reg_dataout_2117_port, regs(2116) =>
                           DataPath_RF_bus_reg_dataout_2116_port, regs(2115) =>
                           DataPath_RF_bus_reg_dataout_2115_port, regs(2114) =>
                           DataPath_RF_bus_reg_dataout_2114_port, regs(2113) =>
                           DataPath_RF_bus_reg_dataout_2113_port, regs(2112) =>
                           DataPath_RF_bus_reg_dataout_2112_port, regs(2111) =>
                           DataPath_RF_bus_reg_dataout_2111_port, regs(2110) =>
                           DataPath_RF_bus_reg_dataout_2110_port, regs(2109) =>
                           DataPath_RF_bus_reg_dataout_2109_port, regs(2108) =>
                           DataPath_RF_bus_reg_dataout_2108_port, regs(2107) =>
                           DataPath_RF_bus_reg_dataout_2107_port, regs(2106) =>
                           DataPath_RF_bus_reg_dataout_2106_port, regs(2105) =>
                           DataPath_RF_bus_reg_dataout_2105_port, regs(2104) =>
                           DataPath_RF_bus_reg_dataout_2104_port, regs(2103) =>
                           DataPath_RF_bus_reg_dataout_2103_port, regs(2102) =>
                           DataPath_RF_bus_reg_dataout_2102_port, regs(2101) =>
                           DataPath_RF_bus_reg_dataout_2101_port, regs(2100) =>
                           DataPath_RF_bus_reg_dataout_2100_port, regs(2099) =>
                           DataPath_RF_bus_reg_dataout_2099_port, regs(2098) =>
                           DataPath_RF_bus_reg_dataout_2098_port, regs(2097) =>
                           DataPath_RF_bus_reg_dataout_2097_port, regs(2096) =>
                           DataPath_RF_bus_reg_dataout_2096_port, regs(2095) =>
                           DataPath_RF_bus_reg_dataout_2095_port, regs(2094) =>
                           DataPath_RF_bus_reg_dataout_2094_port, regs(2093) =>
                           DataPath_RF_bus_reg_dataout_2093_port, regs(2092) =>
                           DataPath_RF_bus_reg_dataout_2092_port, regs(2091) =>
                           DataPath_RF_bus_reg_dataout_2091_port, regs(2090) =>
                           DataPath_RF_bus_reg_dataout_2090_port, regs(2089) =>
                           DataPath_RF_bus_reg_dataout_2089_port, regs(2088) =>
                           DataPath_RF_bus_reg_dataout_2088_port, regs(2087) =>
                           DataPath_RF_bus_reg_dataout_2087_port, regs(2086) =>
                           DataPath_RF_bus_reg_dataout_2086_port, regs(2085) =>
                           DataPath_RF_bus_reg_dataout_2085_port, regs(2084) =>
                           DataPath_RF_bus_reg_dataout_2084_port, regs(2083) =>
                           DataPath_RF_bus_reg_dataout_2083_port, regs(2082) =>
                           DataPath_RF_bus_reg_dataout_2082_port, regs(2081) =>
                           DataPath_RF_bus_reg_dataout_2081_port, regs(2080) =>
                           DataPath_RF_bus_reg_dataout_2080_port, regs(2079) =>
                           DataPath_RF_bus_reg_dataout_2079_port, regs(2078) =>
                           DataPath_RF_bus_reg_dataout_2078_port, regs(2077) =>
                           DataPath_RF_bus_reg_dataout_2077_port, regs(2076) =>
                           DataPath_RF_bus_reg_dataout_2076_port, regs(2075) =>
                           DataPath_RF_bus_reg_dataout_2075_port, regs(2074) =>
                           DataPath_RF_bus_reg_dataout_2074_port, regs(2073) =>
                           DataPath_RF_bus_reg_dataout_2073_port, regs(2072) =>
                           DataPath_RF_bus_reg_dataout_2072_port, regs(2071) =>
                           DataPath_RF_bus_reg_dataout_2071_port, regs(2070) =>
                           DataPath_RF_bus_reg_dataout_2070_port, regs(2069) =>
                           DataPath_RF_bus_reg_dataout_2069_port, regs(2068) =>
                           DataPath_RF_bus_reg_dataout_2068_port, regs(2067) =>
                           DataPath_RF_bus_reg_dataout_2067_port, regs(2066) =>
                           DataPath_RF_bus_reg_dataout_2066_port, regs(2065) =>
                           DataPath_RF_bus_reg_dataout_2065_port, regs(2064) =>
                           DataPath_RF_bus_reg_dataout_2064_port, regs(2063) =>
                           DataPath_RF_bus_reg_dataout_2063_port, regs(2062) =>
                           DataPath_RF_bus_reg_dataout_2062_port, regs(2061) =>
                           DataPath_RF_bus_reg_dataout_2061_port, regs(2060) =>
                           DataPath_RF_bus_reg_dataout_2060_port, regs(2059) =>
                           DataPath_RF_bus_reg_dataout_2059_port, regs(2058) =>
                           DataPath_RF_bus_reg_dataout_2058_port, regs(2057) =>
                           DataPath_RF_bus_reg_dataout_2057_port, regs(2056) =>
                           DataPath_RF_bus_reg_dataout_2056_port, regs(2055) =>
                           DataPath_RF_bus_reg_dataout_2055_port, regs(2054) =>
                           DataPath_RF_bus_reg_dataout_2054_port, regs(2053) =>
                           DataPath_RF_bus_reg_dataout_2053_port, regs(2052) =>
                           DataPath_RF_bus_reg_dataout_2052_port, regs(2051) =>
                           DataPath_RF_bus_reg_dataout_2051_port, regs(2050) =>
                           DataPath_RF_bus_reg_dataout_2050_port, regs(2049) =>
                           DataPath_RF_bus_reg_dataout_2049_port, regs(2048) =>
                           DataPath_RF_bus_reg_dataout_2048_port, regs(2047) =>
                           DataPath_RF_bus_reg_dataout_2047_port, regs(2046) =>
                           DataPath_RF_bus_reg_dataout_2046_port, regs(2045) =>
                           DataPath_RF_bus_reg_dataout_2045_port, regs(2044) =>
                           DataPath_RF_bus_reg_dataout_2044_port, regs(2043) =>
                           DataPath_RF_bus_reg_dataout_2043_port, regs(2042) =>
                           DataPath_RF_bus_reg_dataout_2042_port, regs(2041) =>
                           DataPath_RF_bus_reg_dataout_2041_port, regs(2040) =>
                           DataPath_RF_bus_reg_dataout_2040_port, regs(2039) =>
                           DataPath_RF_bus_reg_dataout_2039_port, regs(2038) =>
                           DataPath_RF_bus_reg_dataout_2038_port, regs(2037) =>
                           DataPath_RF_bus_reg_dataout_2037_port, regs(2036) =>
                           DataPath_RF_bus_reg_dataout_2036_port, regs(2035) =>
                           DataPath_RF_bus_reg_dataout_2035_port, regs(2034) =>
                           DataPath_RF_bus_reg_dataout_2034_port, regs(2033) =>
                           DataPath_RF_bus_reg_dataout_2033_port, regs(2032) =>
                           DataPath_RF_bus_reg_dataout_2032_port, regs(2031) =>
                           DataPath_RF_bus_reg_dataout_2031_port, regs(2030) =>
                           DataPath_RF_bus_reg_dataout_2030_port, regs(2029) =>
                           DataPath_RF_bus_reg_dataout_2029_port, regs(2028) =>
                           DataPath_RF_bus_reg_dataout_2028_port, regs(2027) =>
                           DataPath_RF_bus_reg_dataout_2027_port, regs(2026) =>
                           DataPath_RF_bus_reg_dataout_2026_port, regs(2025) =>
                           DataPath_RF_bus_reg_dataout_2025_port, regs(2024) =>
                           DataPath_RF_bus_reg_dataout_2024_port, regs(2023) =>
                           DataPath_RF_bus_reg_dataout_2023_port, regs(2022) =>
                           DataPath_RF_bus_reg_dataout_2022_port, regs(2021) =>
                           DataPath_RF_bus_reg_dataout_2021_port, regs(2020) =>
                           DataPath_RF_bus_reg_dataout_2020_port, regs(2019) =>
                           DataPath_RF_bus_reg_dataout_2019_port, regs(2018) =>
                           DataPath_RF_bus_reg_dataout_2018_port, regs(2017) =>
                           DataPath_RF_bus_reg_dataout_2017_port, regs(2016) =>
                           DataPath_RF_bus_reg_dataout_2016_port, regs(2015) =>
                           DataPath_RF_bus_reg_dataout_2015_port, regs(2014) =>
                           DataPath_RF_bus_reg_dataout_2014_port, regs(2013) =>
                           DataPath_RF_bus_reg_dataout_2013_port, regs(2012) =>
                           DataPath_RF_bus_reg_dataout_2012_port, regs(2011) =>
                           DataPath_RF_bus_reg_dataout_2011_port, regs(2010) =>
                           DataPath_RF_bus_reg_dataout_2010_port, regs(2009) =>
                           DataPath_RF_bus_reg_dataout_2009_port, regs(2008) =>
                           DataPath_RF_bus_reg_dataout_2008_port, regs(2007) =>
                           DataPath_RF_bus_reg_dataout_2007_port, regs(2006) =>
                           DataPath_RF_bus_reg_dataout_2006_port, regs(2005) =>
                           DataPath_RF_bus_reg_dataout_2005_port, regs(2004) =>
                           DataPath_RF_bus_reg_dataout_2004_port, regs(2003) =>
                           DataPath_RF_bus_reg_dataout_2003_port, regs(2002) =>
                           DataPath_RF_bus_reg_dataout_2002_port, regs(2001) =>
                           DataPath_RF_bus_reg_dataout_2001_port, regs(2000) =>
                           DataPath_RF_bus_reg_dataout_2000_port, regs(1999) =>
                           DataPath_RF_bus_reg_dataout_1999_port, regs(1998) =>
                           DataPath_RF_bus_reg_dataout_1998_port, regs(1997) =>
                           DataPath_RF_bus_reg_dataout_1997_port, regs(1996) =>
                           DataPath_RF_bus_reg_dataout_1996_port, regs(1995) =>
                           DataPath_RF_bus_reg_dataout_1995_port, regs(1994) =>
                           DataPath_RF_bus_reg_dataout_1994_port, regs(1993) =>
                           DataPath_RF_bus_reg_dataout_1993_port, regs(1992) =>
                           DataPath_RF_bus_reg_dataout_1992_port, regs(1991) =>
                           DataPath_RF_bus_reg_dataout_1991_port, regs(1990) =>
                           DataPath_RF_bus_reg_dataout_1990_port, regs(1989) =>
                           DataPath_RF_bus_reg_dataout_1989_port, regs(1988) =>
                           DataPath_RF_bus_reg_dataout_1988_port, regs(1987) =>
                           DataPath_RF_bus_reg_dataout_1987_port, regs(1986) =>
                           DataPath_RF_bus_reg_dataout_1986_port, regs(1985) =>
                           DataPath_RF_bus_reg_dataout_1985_port, regs(1984) =>
                           DataPath_RF_bus_reg_dataout_1984_port, regs(1983) =>
                           DataPath_RF_bus_reg_dataout_1983_port, regs(1982) =>
                           DataPath_RF_bus_reg_dataout_1982_port, regs(1981) =>
                           DataPath_RF_bus_reg_dataout_1981_port, regs(1980) =>
                           DataPath_RF_bus_reg_dataout_1980_port, regs(1979) =>
                           DataPath_RF_bus_reg_dataout_1979_port, regs(1978) =>
                           DataPath_RF_bus_reg_dataout_1978_port, regs(1977) =>
                           DataPath_RF_bus_reg_dataout_1977_port, regs(1976) =>
                           DataPath_RF_bus_reg_dataout_1976_port, regs(1975) =>
                           DataPath_RF_bus_reg_dataout_1975_port, regs(1974) =>
                           DataPath_RF_bus_reg_dataout_1974_port, regs(1973) =>
                           DataPath_RF_bus_reg_dataout_1973_port, regs(1972) =>
                           DataPath_RF_bus_reg_dataout_1972_port, regs(1971) =>
                           DataPath_RF_bus_reg_dataout_1971_port, regs(1970) =>
                           DataPath_RF_bus_reg_dataout_1970_port, regs(1969) =>
                           DataPath_RF_bus_reg_dataout_1969_port, regs(1968) =>
                           DataPath_RF_bus_reg_dataout_1968_port, regs(1967) =>
                           DataPath_RF_bus_reg_dataout_1967_port, regs(1966) =>
                           DataPath_RF_bus_reg_dataout_1966_port, regs(1965) =>
                           DataPath_RF_bus_reg_dataout_1965_port, regs(1964) =>
                           DataPath_RF_bus_reg_dataout_1964_port, regs(1963) =>
                           DataPath_RF_bus_reg_dataout_1963_port, regs(1962) =>
                           DataPath_RF_bus_reg_dataout_1962_port, regs(1961) =>
                           DataPath_RF_bus_reg_dataout_1961_port, regs(1960) =>
                           DataPath_RF_bus_reg_dataout_1960_port, regs(1959) =>
                           DataPath_RF_bus_reg_dataout_1959_port, regs(1958) =>
                           DataPath_RF_bus_reg_dataout_1958_port, regs(1957) =>
                           DataPath_RF_bus_reg_dataout_1957_port, regs(1956) =>
                           DataPath_RF_bus_reg_dataout_1956_port, regs(1955) =>
                           DataPath_RF_bus_reg_dataout_1955_port, regs(1954) =>
                           DataPath_RF_bus_reg_dataout_1954_port, regs(1953) =>
                           DataPath_RF_bus_reg_dataout_1953_port, regs(1952) =>
                           DataPath_RF_bus_reg_dataout_1952_port, regs(1951) =>
                           DataPath_RF_bus_reg_dataout_1951_port, regs(1950) =>
                           DataPath_RF_bus_reg_dataout_1950_port, regs(1949) =>
                           DataPath_RF_bus_reg_dataout_1949_port, regs(1948) =>
                           DataPath_RF_bus_reg_dataout_1948_port, regs(1947) =>
                           DataPath_RF_bus_reg_dataout_1947_port, regs(1946) =>
                           DataPath_RF_bus_reg_dataout_1946_port, regs(1945) =>
                           DataPath_RF_bus_reg_dataout_1945_port, regs(1944) =>
                           DataPath_RF_bus_reg_dataout_1944_port, regs(1943) =>
                           DataPath_RF_bus_reg_dataout_1943_port, regs(1942) =>
                           DataPath_RF_bus_reg_dataout_1942_port, regs(1941) =>
                           DataPath_RF_bus_reg_dataout_1941_port, regs(1940) =>
                           DataPath_RF_bus_reg_dataout_1940_port, regs(1939) =>
                           DataPath_RF_bus_reg_dataout_1939_port, regs(1938) =>
                           DataPath_RF_bus_reg_dataout_1938_port, regs(1937) =>
                           DataPath_RF_bus_reg_dataout_1937_port, regs(1936) =>
                           DataPath_RF_bus_reg_dataout_1936_port, regs(1935) =>
                           DataPath_RF_bus_reg_dataout_1935_port, regs(1934) =>
                           DataPath_RF_bus_reg_dataout_1934_port, regs(1933) =>
                           DataPath_RF_bus_reg_dataout_1933_port, regs(1932) =>
                           DataPath_RF_bus_reg_dataout_1932_port, regs(1931) =>
                           DataPath_RF_bus_reg_dataout_1931_port, regs(1930) =>
                           DataPath_RF_bus_reg_dataout_1930_port, regs(1929) =>
                           DataPath_RF_bus_reg_dataout_1929_port, regs(1928) =>
                           DataPath_RF_bus_reg_dataout_1928_port, regs(1927) =>
                           DataPath_RF_bus_reg_dataout_1927_port, regs(1926) =>
                           DataPath_RF_bus_reg_dataout_1926_port, regs(1925) =>
                           DataPath_RF_bus_reg_dataout_1925_port, regs(1924) =>
                           DataPath_RF_bus_reg_dataout_1924_port, regs(1923) =>
                           DataPath_RF_bus_reg_dataout_1923_port, regs(1922) =>
                           DataPath_RF_bus_reg_dataout_1922_port, regs(1921) =>
                           DataPath_RF_bus_reg_dataout_1921_port, regs(1920) =>
                           DataPath_RF_bus_reg_dataout_1920_port, regs(1919) =>
                           DataPath_RF_bus_reg_dataout_1919_port, regs(1918) =>
                           DataPath_RF_bus_reg_dataout_1918_port, regs(1917) =>
                           DataPath_RF_bus_reg_dataout_1917_port, regs(1916) =>
                           DataPath_RF_bus_reg_dataout_1916_port, regs(1915) =>
                           DataPath_RF_bus_reg_dataout_1915_port, regs(1914) =>
                           DataPath_RF_bus_reg_dataout_1914_port, regs(1913) =>
                           DataPath_RF_bus_reg_dataout_1913_port, regs(1912) =>
                           DataPath_RF_bus_reg_dataout_1912_port, regs(1911) =>
                           DataPath_RF_bus_reg_dataout_1911_port, regs(1910) =>
                           DataPath_RF_bus_reg_dataout_1910_port, regs(1909) =>
                           DataPath_RF_bus_reg_dataout_1909_port, regs(1908) =>
                           DataPath_RF_bus_reg_dataout_1908_port, regs(1907) =>
                           DataPath_RF_bus_reg_dataout_1907_port, regs(1906) =>
                           DataPath_RF_bus_reg_dataout_1906_port, regs(1905) =>
                           DataPath_RF_bus_reg_dataout_1905_port, regs(1904) =>
                           DataPath_RF_bus_reg_dataout_1904_port, regs(1903) =>
                           DataPath_RF_bus_reg_dataout_1903_port, regs(1902) =>
                           DataPath_RF_bus_reg_dataout_1902_port, regs(1901) =>
                           DataPath_RF_bus_reg_dataout_1901_port, regs(1900) =>
                           DataPath_RF_bus_reg_dataout_1900_port, regs(1899) =>
                           DataPath_RF_bus_reg_dataout_1899_port, regs(1898) =>
                           DataPath_RF_bus_reg_dataout_1898_port, regs(1897) =>
                           DataPath_RF_bus_reg_dataout_1897_port, regs(1896) =>
                           DataPath_RF_bus_reg_dataout_1896_port, regs(1895) =>
                           DataPath_RF_bus_reg_dataout_1895_port, regs(1894) =>
                           DataPath_RF_bus_reg_dataout_1894_port, regs(1893) =>
                           DataPath_RF_bus_reg_dataout_1893_port, regs(1892) =>
                           DataPath_RF_bus_reg_dataout_1892_port, regs(1891) =>
                           DataPath_RF_bus_reg_dataout_1891_port, regs(1890) =>
                           DataPath_RF_bus_reg_dataout_1890_port, regs(1889) =>
                           DataPath_RF_bus_reg_dataout_1889_port, regs(1888) =>
                           DataPath_RF_bus_reg_dataout_1888_port, regs(1887) =>
                           DataPath_RF_bus_reg_dataout_1887_port, regs(1886) =>
                           DataPath_RF_bus_reg_dataout_1886_port, regs(1885) =>
                           DataPath_RF_bus_reg_dataout_1885_port, regs(1884) =>
                           DataPath_RF_bus_reg_dataout_1884_port, regs(1883) =>
                           DataPath_RF_bus_reg_dataout_1883_port, regs(1882) =>
                           DataPath_RF_bus_reg_dataout_1882_port, regs(1881) =>
                           DataPath_RF_bus_reg_dataout_1881_port, regs(1880) =>
                           DataPath_RF_bus_reg_dataout_1880_port, regs(1879) =>
                           DataPath_RF_bus_reg_dataout_1879_port, regs(1878) =>
                           DataPath_RF_bus_reg_dataout_1878_port, regs(1877) =>
                           DataPath_RF_bus_reg_dataout_1877_port, regs(1876) =>
                           DataPath_RF_bus_reg_dataout_1876_port, regs(1875) =>
                           DataPath_RF_bus_reg_dataout_1875_port, regs(1874) =>
                           DataPath_RF_bus_reg_dataout_1874_port, regs(1873) =>
                           DataPath_RF_bus_reg_dataout_1873_port, regs(1872) =>
                           DataPath_RF_bus_reg_dataout_1872_port, regs(1871) =>
                           DataPath_RF_bus_reg_dataout_1871_port, regs(1870) =>
                           DataPath_RF_bus_reg_dataout_1870_port, regs(1869) =>
                           DataPath_RF_bus_reg_dataout_1869_port, regs(1868) =>
                           DataPath_RF_bus_reg_dataout_1868_port, regs(1867) =>
                           DataPath_RF_bus_reg_dataout_1867_port, regs(1866) =>
                           DataPath_RF_bus_reg_dataout_1866_port, regs(1865) =>
                           DataPath_RF_bus_reg_dataout_1865_port, regs(1864) =>
                           DataPath_RF_bus_reg_dataout_1864_port, regs(1863) =>
                           DataPath_RF_bus_reg_dataout_1863_port, regs(1862) =>
                           DataPath_RF_bus_reg_dataout_1862_port, regs(1861) =>
                           DataPath_RF_bus_reg_dataout_1861_port, regs(1860) =>
                           DataPath_RF_bus_reg_dataout_1860_port, regs(1859) =>
                           DataPath_RF_bus_reg_dataout_1859_port, regs(1858) =>
                           DataPath_RF_bus_reg_dataout_1858_port, regs(1857) =>
                           DataPath_RF_bus_reg_dataout_1857_port, regs(1856) =>
                           DataPath_RF_bus_reg_dataout_1856_port, regs(1855) =>
                           DataPath_RF_bus_reg_dataout_1855_port, regs(1854) =>
                           DataPath_RF_bus_reg_dataout_1854_port, regs(1853) =>
                           DataPath_RF_bus_reg_dataout_1853_port, regs(1852) =>
                           DataPath_RF_bus_reg_dataout_1852_port, regs(1851) =>
                           DataPath_RF_bus_reg_dataout_1851_port, regs(1850) =>
                           DataPath_RF_bus_reg_dataout_1850_port, regs(1849) =>
                           DataPath_RF_bus_reg_dataout_1849_port, regs(1848) =>
                           DataPath_RF_bus_reg_dataout_1848_port, regs(1847) =>
                           DataPath_RF_bus_reg_dataout_1847_port, regs(1846) =>
                           DataPath_RF_bus_reg_dataout_1846_port, regs(1845) =>
                           DataPath_RF_bus_reg_dataout_1845_port, regs(1844) =>
                           DataPath_RF_bus_reg_dataout_1844_port, regs(1843) =>
                           DataPath_RF_bus_reg_dataout_1843_port, regs(1842) =>
                           DataPath_RF_bus_reg_dataout_1842_port, regs(1841) =>
                           DataPath_RF_bus_reg_dataout_1841_port, regs(1840) =>
                           DataPath_RF_bus_reg_dataout_1840_port, regs(1839) =>
                           DataPath_RF_bus_reg_dataout_1839_port, regs(1838) =>
                           DataPath_RF_bus_reg_dataout_1838_port, regs(1837) =>
                           DataPath_RF_bus_reg_dataout_1837_port, regs(1836) =>
                           DataPath_RF_bus_reg_dataout_1836_port, regs(1835) =>
                           DataPath_RF_bus_reg_dataout_1835_port, regs(1834) =>
                           DataPath_RF_bus_reg_dataout_1834_port, regs(1833) =>
                           DataPath_RF_bus_reg_dataout_1833_port, regs(1832) =>
                           DataPath_RF_bus_reg_dataout_1832_port, regs(1831) =>
                           DataPath_RF_bus_reg_dataout_1831_port, regs(1830) =>
                           DataPath_RF_bus_reg_dataout_1830_port, regs(1829) =>
                           DataPath_RF_bus_reg_dataout_1829_port, regs(1828) =>
                           DataPath_RF_bus_reg_dataout_1828_port, regs(1827) =>
                           DataPath_RF_bus_reg_dataout_1827_port, regs(1826) =>
                           DataPath_RF_bus_reg_dataout_1826_port, regs(1825) =>
                           DataPath_RF_bus_reg_dataout_1825_port, regs(1824) =>
                           DataPath_RF_bus_reg_dataout_1824_port, regs(1823) =>
                           DataPath_RF_bus_reg_dataout_1823_port, regs(1822) =>
                           DataPath_RF_bus_reg_dataout_1822_port, regs(1821) =>
                           DataPath_RF_bus_reg_dataout_1821_port, regs(1820) =>
                           DataPath_RF_bus_reg_dataout_1820_port, regs(1819) =>
                           DataPath_RF_bus_reg_dataout_1819_port, regs(1818) =>
                           DataPath_RF_bus_reg_dataout_1818_port, regs(1817) =>
                           DataPath_RF_bus_reg_dataout_1817_port, regs(1816) =>
                           DataPath_RF_bus_reg_dataout_1816_port, regs(1815) =>
                           DataPath_RF_bus_reg_dataout_1815_port, regs(1814) =>
                           DataPath_RF_bus_reg_dataout_1814_port, regs(1813) =>
                           DataPath_RF_bus_reg_dataout_1813_port, regs(1812) =>
                           DataPath_RF_bus_reg_dataout_1812_port, regs(1811) =>
                           DataPath_RF_bus_reg_dataout_1811_port, regs(1810) =>
                           DataPath_RF_bus_reg_dataout_1810_port, regs(1809) =>
                           DataPath_RF_bus_reg_dataout_1809_port, regs(1808) =>
                           DataPath_RF_bus_reg_dataout_1808_port, regs(1807) =>
                           DataPath_RF_bus_reg_dataout_1807_port, regs(1806) =>
                           DataPath_RF_bus_reg_dataout_1806_port, regs(1805) =>
                           DataPath_RF_bus_reg_dataout_1805_port, regs(1804) =>
                           DataPath_RF_bus_reg_dataout_1804_port, regs(1803) =>
                           DataPath_RF_bus_reg_dataout_1803_port, regs(1802) =>
                           DataPath_RF_bus_reg_dataout_1802_port, regs(1801) =>
                           DataPath_RF_bus_reg_dataout_1801_port, regs(1800) =>
                           DataPath_RF_bus_reg_dataout_1800_port, regs(1799) =>
                           DataPath_RF_bus_reg_dataout_1799_port, regs(1798) =>
                           DataPath_RF_bus_reg_dataout_1798_port, regs(1797) =>
                           DataPath_RF_bus_reg_dataout_1797_port, regs(1796) =>
                           DataPath_RF_bus_reg_dataout_1796_port, regs(1795) =>
                           DataPath_RF_bus_reg_dataout_1795_port, regs(1794) =>
                           DataPath_RF_bus_reg_dataout_1794_port, regs(1793) =>
                           DataPath_RF_bus_reg_dataout_1793_port, regs(1792) =>
                           DataPath_RF_bus_reg_dataout_1792_port, regs(1791) =>
                           DataPath_RF_bus_reg_dataout_1791_port, regs(1790) =>
                           DataPath_RF_bus_reg_dataout_1790_port, regs(1789) =>
                           DataPath_RF_bus_reg_dataout_1789_port, regs(1788) =>
                           DataPath_RF_bus_reg_dataout_1788_port, regs(1787) =>
                           DataPath_RF_bus_reg_dataout_1787_port, regs(1786) =>
                           DataPath_RF_bus_reg_dataout_1786_port, regs(1785) =>
                           DataPath_RF_bus_reg_dataout_1785_port, regs(1784) =>
                           DataPath_RF_bus_reg_dataout_1784_port, regs(1783) =>
                           DataPath_RF_bus_reg_dataout_1783_port, regs(1782) =>
                           DataPath_RF_bus_reg_dataout_1782_port, regs(1781) =>
                           DataPath_RF_bus_reg_dataout_1781_port, regs(1780) =>
                           DataPath_RF_bus_reg_dataout_1780_port, regs(1779) =>
                           DataPath_RF_bus_reg_dataout_1779_port, regs(1778) =>
                           DataPath_RF_bus_reg_dataout_1778_port, regs(1777) =>
                           DataPath_RF_bus_reg_dataout_1777_port, regs(1776) =>
                           DataPath_RF_bus_reg_dataout_1776_port, regs(1775) =>
                           DataPath_RF_bus_reg_dataout_1775_port, regs(1774) =>
                           DataPath_RF_bus_reg_dataout_1774_port, regs(1773) =>
                           DataPath_RF_bus_reg_dataout_1773_port, regs(1772) =>
                           DataPath_RF_bus_reg_dataout_1772_port, regs(1771) =>
                           DataPath_RF_bus_reg_dataout_1771_port, regs(1770) =>
                           DataPath_RF_bus_reg_dataout_1770_port, regs(1769) =>
                           DataPath_RF_bus_reg_dataout_1769_port, regs(1768) =>
                           DataPath_RF_bus_reg_dataout_1768_port, regs(1767) =>
                           DataPath_RF_bus_reg_dataout_1767_port, regs(1766) =>
                           DataPath_RF_bus_reg_dataout_1766_port, regs(1765) =>
                           DataPath_RF_bus_reg_dataout_1765_port, regs(1764) =>
                           DataPath_RF_bus_reg_dataout_1764_port, regs(1763) =>
                           DataPath_RF_bus_reg_dataout_1763_port, regs(1762) =>
                           DataPath_RF_bus_reg_dataout_1762_port, regs(1761) =>
                           DataPath_RF_bus_reg_dataout_1761_port, regs(1760) =>
                           DataPath_RF_bus_reg_dataout_1760_port, regs(1759) =>
                           DataPath_RF_bus_reg_dataout_1759_port, regs(1758) =>
                           DataPath_RF_bus_reg_dataout_1758_port, regs(1757) =>
                           DataPath_RF_bus_reg_dataout_1757_port, regs(1756) =>
                           DataPath_RF_bus_reg_dataout_1756_port, regs(1755) =>
                           DataPath_RF_bus_reg_dataout_1755_port, regs(1754) =>
                           DataPath_RF_bus_reg_dataout_1754_port, regs(1753) =>
                           DataPath_RF_bus_reg_dataout_1753_port, regs(1752) =>
                           DataPath_RF_bus_reg_dataout_1752_port, regs(1751) =>
                           DataPath_RF_bus_reg_dataout_1751_port, regs(1750) =>
                           DataPath_RF_bus_reg_dataout_1750_port, regs(1749) =>
                           DataPath_RF_bus_reg_dataout_1749_port, regs(1748) =>
                           DataPath_RF_bus_reg_dataout_1748_port, regs(1747) =>
                           DataPath_RF_bus_reg_dataout_1747_port, regs(1746) =>
                           DataPath_RF_bus_reg_dataout_1746_port, regs(1745) =>
                           DataPath_RF_bus_reg_dataout_1745_port, regs(1744) =>
                           DataPath_RF_bus_reg_dataout_1744_port, regs(1743) =>
                           DataPath_RF_bus_reg_dataout_1743_port, regs(1742) =>
                           DataPath_RF_bus_reg_dataout_1742_port, regs(1741) =>
                           DataPath_RF_bus_reg_dataout_1741_port, regs(1740) =>
                           DataPath_RF_bus_reg_dataout_1740_port, regs(1739) =>
                           DataPath_RF_bus_reg_dataout_1739_port, regs(1738) =>
                           DataPath_RF_bus_reg_dataout_1738_port, regs(1737) =>
                           DataPath_RF_bus_reg_dataout_1737_port, regs(1736) =>
                           DataPath_RF_bus_reg_dataout_1736_port, regs(1735) =>
                           DataPath_RF_bus_reg_dataout_1735_port, regs(1734) =>
                           DataPath_RF_bus_reg_dataout_1734_port, regs(1733) =>
                           DataPath_RF_bus_reg_dataout_1733_port, regs(1732) =>
                           DataPath_RF_bus_reg_dataout_1732_port, regs(1731) =>
                           DataPath_RF_bus_reg_dataout_1731_port, regs(1730) =>
                           DataPath_RF_bus_reg_dataout_1730_port, regs(1729) =>
                           DataPath_RF_bus_reg_dataout_1729_port, regs(1728) =>
                           DataPath_RF_bus_reg_dataout_1728_port, regs(1727) =>
                           DataPath_RF_bus_reg_dataout_1727_port, regs(1726) =>
                           DataPath_RF_bus_reg_dataout_1726_port, regs(1725) =>
                           DataPath_RF_bus_reg_dataout_1725_port, regs(1724) =>
                           DataPath_RF_bus_reg_dataout_1724_port, regs(1723) =>
                           DataPath_RF_bus_reg_dataout_1723_port, regs(1722) =>
                           DataPath_RF_bus_reg_dataout_1722_port, regs(1721) =>
                           DataPath_RF_bus_reg_dataout_1721_port, regs(1720) =>
                           DataPath_RF_bus_reg_dataout_1720_port, regs(1719) =>
                           DataPath_RF_bus_reg_dataout_1719_port, regs(1718) =>
                           DataPath_RF_bus_reg_dataout_1718_port, regs(1717) =>
                           DataPath_RF_bus_reg_dataout_1717_port, regs(1716) =>
                           DataPath_RF_bus_reg_dataout_1716_port, regs(1715) =>
                           DataPath_RF_bus_reg_dataout_1715_port, regs(1714) =>
                           DataPath_RF_bus_reg_dataout_1714_port, regs(1713) =>
                           DataPath_RF_bus_reg_dataout_1713_port, regs(1712) =>
                           DataPath_RF_bus_reg_dataout_1712_port, regs(1711) =>
                           DataPath_RF_bus_reg_dataout_1711_port, regs(1710) =>
                           DataPath_RF_bus_reg_dataout_1710_port, regs(1709) =>
                           DataPath_RF_bus_reg_dataout_1709_port, regs(1708) =>
                           DataPath_RF_bus_reg_dataout_1708_port, regs(1707) =>
                           DataPath_RF_bus_reg_dataout_1707_port, regs(1706) =>
                           DataPath_RF_bus_reg_dataout_1706_port, regs(1705) =>
                           DataPath_RF_bus_reg_dataout_1705_port, regs(1704) =>
                           DataPath_RF_bus_reg_dataout_1704_port, regs(1703) =>
                           DataPath_RF_bus_reg_dataout_1703_port, regs(1702) =>
                           DataPath_RF_bus_reg_dataout_1702_port, regs(1701) =>
                           DataPath_RF_bus_reg_dataout_1701_port, regs(1700) =>
                           DataPath_RF_bus_reg_dataout_1700_port, regs(1699) =>
                           DataPath_RF_bus_reg_dataout_1699_port, regs(1698) =>
                           DataPath_RF_bus_reg_dataout_1698_port, regs(1697) =>
                           DataPath_RF_bus_reg_dataout_1697_port, regs(1696) =>
                           DataPath_RF_bus_reg_dataout_1696_port, regs(1695) =>
                           DataPath_RF_bus_reg_dataout_1695_port, regs(1694) =>
                           DataPath_RF_bus_reg_dataout_1694_port, regs(1693) =>
                           DataPath_RF_bus_reg_dataout_1693_port, regs(1692) =>
                           DataPath_RF_bus_reg_dataout_1692_port, regs(1691) =>
                           DataPath_RF_bus_reg_dataout_1691_port, regs(1690) =>
                           DataPath_RF_bus_reg_dataout_1690_port, regs(1689) =>
                           DataPath_RF_bus_reg_dataout_1689_port, regs(1688) =>
                           DataPath_RF_bus_reg_dataout_1688_port, regs(1687) =>
                           DataPath_RF_bus_reg_dataout_1687_port, regs(1686) =>
                           DataPath_RF_bus_reg_dataout_1686_port, regs(1685) =>
                           DataPath_RF_bus_reg_dataout_1685_port, regs(1684) =>
                           DataPath_RF_bus_reg_dataout_1684_port, regs(1683) =>
                           DataPath_RF_bus_reg_dataout_1683_port, regs(1682) =>
                           DataPath_RF_bus_reg_dataout_1682_port, regs(1681) =>
                           DataPath_RF_bus_reg_dataout_1681_port, regs(1680) =>
                           DataPath_RF_bus_reg_dataout_1680_port, regs(1679) =>
                           DataPath_RF_bus_reg_dataout_1679_port, regs(1678) =>
                           DataPath_RF_bus_reg_dataout_1678_port, regs(1677) =>
                           DataPath_RF_bus_reg_dataout_1677_port, regs(1676) =>
                           DataPath_RF_bus_reg_dataout_1676_port, regs(1675) =>
                           DataPath_RF_bus_reg_dataout_1675_port, regs(1674) =>
                           DataPath_RF_bus_reg_dataout_1674_port, regs(1673) =>
                           DataPath_RF_bus_reg_dataout_1673_port, regs(1672) =>
                           DataPath_RF_bus_reg_dataout_1672_port, regs(1671) =>
                           DataPath_RF_bus_reg_dataout_1671_port, regs(1670) =>
                           DataPath_RF_bus_reg_dataout_1670_port, regs(1669) =>
                           DataPath_RF_bus_reg_dataout_1669_port, regs(1668) =>
                           DataPath_RF_bus_reg_dataout_1668_port, regs(1667) =>
                           DataPath_RF_bus_reg_dataout_1667_port, regs(1666) =>
                           DataPath_RF_bus_reg_dataout_1666_port, regs(1665) =>
                           DataPath_RF_bus_reg_dataout_1665_port, regs(1664) =>
                           DataPath_RF_bus_reg_dataout_1664_port, regs(1663) =>
                           DataPath_RF_bus_reg_dataout_1663_port, regs(1662) =>
                           DataPath_RF_bus_reg_dataout_1662_port, regs(1661) =>
                           DataPath_RF_bus_reg_dataout_1661_port, regs(1660) =>
                           DataPath_RF_bus_reg_dataout_1660_port, regs(1659) =>
                           DataPath_RF_bus_reg_dataout_1659_port, regs(1658) =>
                           DataPath_RF_bus_reg_dataout_1658_port, regs(1657) =>
                           DataPath_RF_bus_reg_dataout_1657_port, regs(1656) =>
                           DataPath_RF_bus_reg_dataout_1656_port, regs(1655) =>
                           DataPath_RF_bus_reg_dataout_1655_port, regs(1654) =>
                           DataPath_RF_bus_reg_dataout_1654_port, regs(1653) =>
                           DataPath_RF_bus_reg_dataout_1653_port, regs(1652) =>
                           DataPath_RF_bus_reg_dataout_1652_port, regs(1651) =>
                           DataPath_RF_bus_reg_dataout_1651_port, regs(1650) =>
                           DataPath_RF_bus_reg_dataout_1650_port, regs(1649) =>
                           DataPath_RF_bus_reg_dataout_1649_port, regs(1648) =>
                           DataPath_RF_bus_reg_dataout_1648_port, regs(1647) =>
                           DataPath_RF_bus_reg_dataout_1647_port, regs(1646) =>
                           DataPath_RF_bus_reg_dataout_1646_port, regs(1645) =>
                           DataPath_RF_bus_reg_dataout_1645_port, regs(1644) =>
                           DataPath_RF_bus_reg_dataout_1644_port, regs(1643) =>
                           DataPath_RF_bus_reg_dataout_1643_port, regs(1642) =>
                           DataPath_RF_bus_reg_dataout_1642_port, regs(1641) =>
                           DataPath_RF_bus_reg_dataout_1641_port, regs(1640) =>
                           DataPath_RF_bus_reg_dataout_1640_port, regs(1639) =>
                           DataPath_RF_bus_reg_dataout_1639_port, regs(1638) =>
                           DataPath_RF_bus_reg_dataout_1638_port, regs(1637) =>
                           DataPath_RF_bus_reg_dataout_1637_port, regs(1636) =>
                           DataPath_RF_bus_reg_dataout_1636_port, regs(1635) =>
                           DataPath_RF_bus_reg_dataout_1635_port, regs(1634) =>
                           DataPath_RF_bus_reg_dataout_1634_port, regs(1633) =>
                           DataPath_RF_bus_reg_dataout_1633_port, regs(1632) =>
                           DataPath_RF_bus_reg_dataout_1632_port, regs(1631) =>
                           DataPath_RF_bus_reg_dataout_1631_port, regs(1630) =>
                           DataPath_RF_bus_reg_dataout_1630_port, regs(1629) =>
                           DataPath_RF_bus_reg_dataout_1629_port, regs(1628) =>
                           DataPath_RF_bus_reg_dataout_1628_port, regs(1627) =>
                           DataPath_RF_bus_reg_dataout_1627_port, regs(1626) =>
                           DataPath_RF_bus_reg_dataout_1626_port, regs(1625) =>
                           DataPath_RF_bus_reg_dataout_1625_port, regs(1624) =>
                           DataPath_RF_bus_reg_dataout_1624_port, regs(1623) =>
                           DataPath_RF_bus_reg_dataout_1623_port, regs(1622) =>
                           DataPath_RF_bus_reg_dataout_1622_port, regs(1621) =>
                           DataPath_RF_bus_reg_dataout_1621_port, regs(1620) =>
                           DataPath_RF_bus_reg_dataout_1620_port, regs(1619) =>
                           DataPath_RF_bus_reg_dataout_1619_port, regs(1618) =>
                           DataPath_RF_bus_reg_dataout_1618_port, regs(1617) =>
                           DataPath_RF_bus_reg_dataout_1617_port, regs(1616) =>
                           DataPath_RF_bus_reg_dataout_1616_port, regs(1615) =>
                           DataPath_RF_bus_reg_dataout_1615_port, regs(1614) =>
                           DataPath_RF_bus_reg_dataout_1614_port, regs(1613) =>
                           DataPath_RF_bus_reg_dataout_1613_port, regs(1612) =>
                           DataPath_RF_bus_reg_dataout_1612_port, regs(1611) =>
                           DataPath_RF_bus_reg_dataout_1611_port, regs(1610) =>
                           DataPath_RF_bus_reg_dataout_1610_port, regs(1609) =>
                           DataPath_RF_bus_reg_dataout_1609_port, regs(1608) =>
                           DataPath_RF_bus_reg_dataout_1608_port, regs(1607) =>
                           DataPath_RF_bus_reg_dataout_1607_port, regs(1606) =>
                           DataPath_RF_bus_reg_dataout_1606_port, regs(1605) =>
                           DataPath_RF_bus_reg_dataout_1605_port, regs(1604) =>
                           DataPath_RF_bus_reg_dataout_1604_port, regs(1603) =>
                           DataPath_RF_bus_reg_dataout_1603_port, regs(1602) =>
                           DataPath_RF_bus_reg_dataout_1602_port, regs(1601) =>
                           DataPath_RF_bus_reg_dataout_1601_port, regs(1600) =>
                           DataPath_RF_bus_reg_dataout_1600_port, regs(1599) =>
                           DataPath_RF_bus_reg_dataout_1599_port, regs(1598) =>
                           DataPath_RF_bus_reg_dataout_1598_port, regs(1597) =>
                           DataPath_RF_bus_reg_dataout_1597_port, regs(1596) =>
                           DataPath_RF_bus_reg_dataout_1596_port, regs(1595) =>
                           DataPath_RF_bus_reg_dataout_1595_port, regs(1594) =>
                           DataPath_RF_bus_reg_dataout_1594_port, regs(1593) =>
                           DataPath_RF_bus_reg_dataout_1593_port, regs(1592) =>
                           DataPath_RF_bus_reg_dataout_1592_port, regs(1591) =>
                           DataPath_RF_bus_reg_dataout_1591_port, regs(1590) =>
                           DataPath_RF_bus_reg_dataout_1590_port, regs(1589) =>
                           DataPath_RF_bus_reg_dataout_1589_port, regs(1588) =>
                           DataPath_RF_bus_reg_dataout_1588_port, regs(1587) =>
                           DataPath_RF_bus_reg_dataout_1587_port, regs(1586) =>
                           DataPath_RF_bus_reg_dataout_1586_port, regs(1585) =>
                           DataPath_RF_bus_reg_dataout_1585_port, regs(1584) =>
                           DataPath_RF_bus_reg_dataout_1584_port, regs(1583) =>
                           DataPath_RF_bus_reg_dataout_1583_port, regs(1582) =>
                           DataPath_RF_bus_reg_dataout_1582_port, regs(1581) =>
                           DataPath_RF_bus_reg_dataout_1581_port, regs(1580) =>
                           DataPath_RF_bus_reg_dataout_1580_port, regs(1579) =>
                           DataPath_RF_bus_reg_dataout_1579_port, regs(1578) =>
                           DataPath_RF_bus_reg_dataout_1578_port, regs(1577) =>
                           DataPath_RF_bus_reg_dataout_1577_port, regs(1576) =>
                           DataPath_RF_bus_reg_dataout_1576_port, regs(1575) =>
                           DataPath_RF_bus_reg_dataout_1575_port, regs(1574) =>
                           DataPath_RF_bus_reg_dataout_1574_port, regs(1573) =>
                           DataPath_RF_bus_reg_dataout_1573_port, regs(1572) =>
                           DataPath_RF_bus_reg_dataout_1572_port, regs(1571) =>
                           DataPath_RF_bus_reg_dataout_1571_port, regs(1570) =>
                           DataPath_RF_bus_reg_dataout_1570_port, regs(1569) =>
                           DataPath_RF_bus_reg_dataout_1569_port, regs(1568) =>
                           DataPath_RF_bus_reg_dataout_1568_port, regs(1567) =>
                           DataPath_RF_bus_reg_dataout_1567_port, regs(1566) =>
                           DataPath_RF_bus_reg_dataout_1566_port, regs(1565) =>
                           DataPath_RF_bus_reg_dataout_1565_port, regs(1564) =>
                           DataPath_RF_bus_reg_dataout_1564_port, regs(1563) =>
                           DataPath_RF_bus_reg_dataout_1563_port, regs(1562) =>
                           DataPath_RF_bus_reg_dataout_1562_port, regs(1561) =>
                           DataPath_RF_bus_reg_dataout_1561_port, regs(1560) =>
                           DataPath_RF_bus_reg_dataout_1560_port, regs(1559) =>
                           DataPath_RF_bus_reg_dataout_1559_port, regs(1558) =>
                           DataPath_RF_bus_reg_dataout_1558_port, regs(1557) =>
                           DataPath_RF_bus_reg_dataout_1557_port, regs(1556) =>
                           DataPath_RF_bus_reg_dataout_1556_port, regs(1555) =>
                           DataPath_RF_bus_reg_dataout_1555_port, regs(1554) =>
                           DataPath_RF_bus_reg_dataout_1554_port, regs(1553) =>
                           DataPath_RF_bus_reg_dataout_1553_port, regs(1552) =>
                           DataPath_RF_bus_reg_dataout_1552_port, regs(1551) =>
                           DataPath_RF_bus_reg_dataout_1551_port, regs(1550) =>
                           DataPath_RF_bus_reg_dataout_1550_port, regs(1549) =>
                           DataPath_RF_bus_reg_dataout_1549_port, regs(1548) =>
                           DataPath_RF_bus_reg_dataout_1548_port, regs(1547) =>
                           DataPath_RF_bus_reg_dataout_1547_port, regs(1546) =>
                           DataPath_RF_bus_reg_dataout_1546_port, regs(1545) =>
                           DataPath_RF_bus_reg_dataout_1545_port, regs(1544) =>
                           DataPath_RF_bus_reg_dataout_1544_port, regs(1543) =>
                           DataPath_RF_bus_reg_dataout_1543_port, regs(1542) =>
                           DataPath_RF_bus_reg_dataout_1542_port, regs(1541) =>
                           DataPath_RF_bus_reg_dataout_1541_port, regs(1540) =>
                           DataPath_RF_bus_reg_dataout_1540_port, regs(1539) =>
                           DataPath_RF_bus_reg_dataout_1539_port, regs(1538) =>
                           DataPath_RF_bus_reg_dataout_1538_port, regs(1537) =>
                           DataPath_RF_bus_reg_dataout_1537_port, regs(1536) =>
                           DataPath_RF_bus_reg_dataout_1536_port, regs(1535) =>
                           DataPath_RF_bus_reg_dataout_1535_port, regs(1534) =>
                           DataPath_RF_bus_reg_dataout_1534_port, regs(1533) =>
                           DataPath_RF_bus_reg_dataout_1533_port, regs(1532) =>
                           DataPath_RF_bus_reg_dataout_1532_port, regs(1531) =>
                           DataPath_RF_bus_reg_dataout_1531_port, regs(1530) =>
                           DataPath_RF_bus_reg_dataout_1530_port, regs(1529) =>
                           DataPath_RF_bus_reg_dataout_1529_port, regs(1528) =>
                           DataPath_RF_bus_reg_dataout_1528_port, regs(1527) =>
                           DataPath_RF_bus_reg_dataout_1527_port, regs(1526) =>
                           DataPath_RF_bus_reg_dataout_1526_port, regs(1525) =>
                           DataPath_RF_bus_reg_dataout_1525_port, regs(1524) =>
                           DataPath_RF_bus_reg_dataout_1524_port, regs(1523) =>
                           DataPath_RF_bus_reg_dataout_1523_port, regs(1522) =>
                           DataPath_RF_bus_reg_dataout_1522_port, regs(1521) =>
                           DataPath_RF_bus_reg_dataout_1521_port, regs(1520) =>
                           DataPath_RF_bus_reg_dataout_1520_port, regs(1519) =>
                           DataPath_RF_bus_reg_dataout_1519_port, regs(1518) =>
                           DataPath_RF_bus_reg_dataout_1518_port, regs(1517) =>
                           DataPath_RF_bus_reg_dataout_1517_port, regs(1516) =>
                           DataPath_RF_bus_reg_dataout_1516_port, regs(1515) =>
                           DataPath_RF_bus_reg_dataout_1515_port, regs(1514) =>
                           DataPath_RF_bus_reg_dataout_1514_port, regs(1513) =>
                           DataPath_RF_bus_reg_dataout_1513_port, regs(1512) =>
                           DataPath_RF_bus_reg_dataout_1512_port, regs(1511) =>
                           DataPath_RF_bus_reg_dataout_1511_port, regs(1510) =>
                           DataPath_RF_bus_reg_dataout_1510_port, regs(1509) =>
                           DataPath_RF_bus_reg_dataout_1509_port, regs(1508) =>
                           DataPath_RF_bus_reg_dataout_1508_port, regs(1507) =>
                           DataPath_RF_bus_reg_dataout_1507_port, regs(1506) =>
                           DataPath_RF_bus_reg_dataout_1506_port, regs(1505) =>
                           DataPath_RF_bus_reg_dataout_1505_port, regs(1504) =>
                           DataPath_RF_bus_reg_dataout_1504_port, regs(1503) =>
                           DataPath_RF_bus_reg_dataout_1503_port, regs(1502) =>
                           DataPath_RF_bus_reg_dataout_1502_port, regs(1501) =>
                           DataPath_RF_bus_reg_dataout_1501_port, regs(1500) =>
                           DataPath_RF_bus_reg_dataout_1500_port, regs(1499) =>
                           DataPath_RF_bus_reg_dataout_1499_port, regs(1498) =>
                           DataPath_RF_bus_reg_dataout_1498_port, regs(1497) =>
                           DataPath_RF_bus_reg_dataout_1497_port, regs(1496) =>
                           DataPath_RF_bus_reg_dataout_1496_port, regs(1495) =>
                           DataPath_RF_bus_reg_dataout_1495_port, regs(1494) =>
                           DataPath_RF_bus_reg_dataout_1494_port, regs(1493) =>
                           DataPath_RF_bus_reg_dataout_1493_port, regs(1492) =>
                           DataPath_RF_bus_reg_dataout_1492_port, regs(1491) =>
                           DataPath_RF_bus_reg_dataout_1491_port, regs(1490) =>
                           DataPath_RF_bus_reg_dataout_1490_port, regs(1489) =>
                           DataPath_RF_bus_reg_dataout_1489_port, regs(1488) =>
                           DataPath_RF_bus_reg_dataout_1488_port, regs(1487) =>
                           DataPath_RF_bus_reg_dataout_1487_port, regs(1486) =>
                           DataPath_RF_bus_reg_dataout_1486_port, regs(1485) =>
                           DataPath_RF_bus_reg_dataout_1485_port, regs(1484) =>
                           DataPath_RF_bus_reg_dataout_1484_port, regs(1483) =>
                           DataPath_RF_bus_reg_dataout_1483_port, regs(1482) =>
                           DataPath_RF_bus_reg_dataout_1482_port, regs(1481) =>
                           DataPath_RF_bus_reg_dataout_1481_port, regs(1480) =>
                           DataPath_RF_bus_reg_dataout_1480_port, regs(1479) =>
                           DataPath_RF_bus_reg_dataout_1479_port, regs(1478) =>
                           DataPath_RF_bus_reg_dataout_1478_port, regs(1477) =>
                           DataPath_RF_bus_reg_dataout_1477_port, regs(1476) =>
                           DataPath_RF_bus_reg_dataout_1476_port, regs(1475) =>
                           DataPath_RF_bus_reg_dataout_1475_port, regs(1474) =>
                           DataPath_RF_bus_reg_dataout_1474_port, regs(1473) =>
                           DataPath_RF_bus_reg_dataout_1473_port, regs(1472) =>
                           DataPath_RF_bus_reg_dataout_1472_port, regs(1471) =>
                           DataPath_RF_bus_reg_dataout_1471_port, regs(1470) =>
                           DataPath_RF_bus_reg_dataout_1470_port, regs(1469) =>
                           DataPath_RF_bus_reg_dataout_1469_port, regs(1468) =>
                           DataPath_RF_bus_reg_dataout_1468_port, regs(1467) =>
                           DataPath_RF_bus_reg_dataout_1467_port, regs(1466) =>
                           DataPath_RF_bus_reg_dataout_1466_port, regs(1465) =>
                           DataPath_RF_bus_reg_dataout_1465_port, regs(1464) =>
                           DataPath_RF_bus_reg_dataout_1464_port, regs(1463) =>
                           DataPath_RF_bus_reg_dataout_1463_port, regs(1462) =>
                           DataPath_RF_bus_reg_dataout_1462_port, regs(1461) =>
                           DataPath_RF_bus_reg_dataout_1461_port, regs(1460) =>
                           DataPath_RF_bus_reg_dataout_1460_port, regs(1459) =>
                           DataPath_RF_bus_reg_dataout_1459_port, regs(1458) =>
                           DataPath_RF_bus_reg_dataout_1458_port, regs(1457) =>
                           DataPath_RF_bus_reg_dataout_1457_port, regs(1456) =>
                           DataPath_RF_bus_reg_dataout_1456_port, regs(1455) =>
                           DataPath_RF_bus_reg_dataout_1455_port, regs(1454) =>
                           DataPath_RF_bus_reg_dataout_1454_port, regs(1453) =>
                           DataPath_RF_bus_reg_dataout_1453_port, regs(1452) =>
                           DataPath_RF_bus_reg_dataout_1452_port, regs(1451) =>
                           DataPath_RF_bus_reg_dataout_1451_port, regs(1450) =>
                           DataPath_RF_bus_reg_dataout_1450_port, regs(1449) =>
                           DataPath_RF_bus_reg_dataout_1449_port, regs(1448) =>
                           DataPath_RF_bus_reg_dataout_1448_port, regs(1447) =>
                           DataPath_RF_bus_reg_dataout_1447_port, regs(1446) =>
                           DataPath_RF_bus_reg_dataout_1446_port, regs(1445) =>
                           DataPath_RF_bus_reg_dataout_1445_port, regs(1444) =>
                           DataPath_RF_bus_reg_dataout_1444_port, regs(1443) =>
                           DataPath_RF_bus_reg_dataout_1443_port, regs(1442) =>
                           DataPath_RF_bus_reg_dataout_1442_port, regs(1441) =>
                           DataPath_RF_bus_reg_dataout_1441_port, regs(1440) =>
                           DataPath_RF_bus_reg_dataout_1440_port, regs(1439) =>
                           DataPath_RF_bus_reg_dataout_1439_port, regs(1438) =>
                           DataPath_RF_bus_reg_dataout_1438_port, regs(1437) =>
                           DataPath_RF_bus_reg_dataout_1437_port, regs(1436) =>
                           DataPath_RF_bus_reg_dataout_1436_port, regs(1435) =>
                           DataPath_RF_bus_reg_dataout_1435_port, regs(1434) =>
                           DataPath_RF_bus_reg_dataout_1434_port, regs(1433) =>
                           DataPath_RF_bus_reg_dataout_1433_port, regs(1432) =>
                           DataPath_RF_bus_reg_dataout_1432_port, regs(1431) =>
                           DataPath_RF_bus_reg_dataout_1431_port, regs(1430) =>
                           DataPath_RF_bus_reg_dataout_1430_port, regs(1429) =>
                           DataPath_RF_bus_reg_dataout_1429_port, regs(1428) =>
                           DataPath_RF_bus_reg_dataout_1428_port, regs(1427) =>
                           DataPath_RF_bus_reg_dataout_1427_port, regs(1426) =>
                           DataPath_RF_bus_reg_dataout_1426_port, regs(1425) =>
                           DataPath_RF_bus_reg_dataout_1425_port, regs(1424) =>
                           DataPath_RF_bus_reg_dataout_1424_port, regs(1423) =>
                           DataPath_RF_bus_reg_dataout_1423_port, regs(1422) =>
                           DataPath_RF_bus_reg_dataout_1422_port, regs(1421) =>
                           DataPath_RF_bus_reg_dataout_1421_port, regs(1420) =>
                           DataPath_RF_bus_reg_dataout_1420_port, regs(1419) =>
                           DataPath_RF_bus_reg_dataout_1419_port, regs(1418) =>
                           DataPath_RF_bus_reg_dataout_1418_port, regs(1417) =>
                           DataPath_RF_bus_reg_dataout_1417_port, regs(1416) =>
                           DataPath_RF_bus_reg_dataout_1416_port, regs(1415) =>
                           DataPath_RF_bus_reg_dataout_1415_port, regs(1414) =>
                           DataPath_RF_bus_reg_dataout_1414_port, regs(1413) =>
                           DataPath_RF_bus_reg_dataout_1413_port, regs(1412) =>
                           DataPath_RF_bus_reg_dataout_1412_port, regs(1411) =>
                           DataPath_RF_bus_reg_dataout_1411_port, regs(1410) =>
                           DataPath_RF_bus_reg_dataout_1410_port, regs(1409) =>
                           DataPath_RF_bus_reg_dataout_1409_port, regs(1408) =>
                           DataPath_RF_bus_reg_dataout_1408_port, regs(1407) =>
                           DataPath_RF_bus_reg_dataout_1407_port, regs(1406) =>
                           DataPath_RF_bus_reg_dataout_1406_port, regs(1405) =>
                           DataPath_RF_bus_reg_dataout_1405_port, regs(1404) =>
                           DataPath_RF_bus_reg_dataout_1404_port, regs(1403) =>
                           DataPath_RF_bus_reg_dataout_1403_port, regs(1402) =>
                           DataPath_RF_bus_reg_dataout_1402_port, regs(1401) =>
                           DataPath_RF_bus_reg_dataout_1401_port, regs(1400) =>
                           DataPath_RF_bus_reg_dataout_1400_port, regs(1399) =>
                           DataPath_RF_bus_reg_dataout_1399_port, regs(1398) =>
                           DataPath_RF_bus_reg_dataout_1398_port, regs(1397) =>
                           DataPath_RF_bus_reg_dataout_1397_port, regs(1396) =>
                           DataPath_RF_bus_reg_dataout_1396_port, regs(1395) =>
                           DataPath_RF_bus_reg_dataout_1395_port, regs(1394) =>
                           DataPath_RF_bus_reg_dataout_1394_port, regs(1393) =>
                           DataPath_RF_bus_reg_dataout_1393_port, regs(1392) =>
                           DataPath_RF_bus_reg_dataout_1392_port, regs(1391) =>
                           DataPath_RF_bus_reg_dataout_1391_port, regs(1390) =>
                           DataPath_RF_bus_reg_dataout_1390_port, regs(1389) =>
                           DataPath_RF_bus_reg_dataout_1389_port, regs(1388) =>
                           DataPath_RF_bus_reg_dataout_1388_port, regs(1387) =>
                           DataPath_RF_bus_reg_dataout_1387_port, regs(1386) =>
                           DataPath_RF_bus_reg_dataout_1386_port, regs(1385) =>
                           DataPath_RF_bus_reg_dataout_1385_port, regs(1384) =>
                           DataPath_RF_bus_reg_dataout_1384_port, regs(1383) =>
                           DataPath_RF_bus_reg_dataout_1383_port, regs(1382) =>
                           DataPath_RF_bus_reg_dataout_1382_port, regs(1381) =>
                           DataPath_RF_bus_reg_dataout_1381_port, regs(1380) =>
                           DataPath_RF_bus_reg_dataout_1380_port, regs(1379) =>
                           DataPath_RF_bus_reg_dataout_1379_port, regs(1378) =>
                           DataPath_RF_bus_reg_dataout_1378_port, regs(1377) =>
                           DataPath_RF_bus_reg_dataout_1377_port, regs(1376) =>
                           DataPath_RF_bus_reg_dataout_1376_port, regs(1375) =>
                           DataPath_RF_bus_reg_dataout_1375_port, regs(1374) =>
                           DataPath_RF_bus_reg_dataout_1374_port, regs(1373) =>
                           DataPath_RF_bus_reg_dataout_1373_port, regs(1372) =>
                           DataPath_RF_bus_reg_dataout_1372_port, regs(1371) =>
                           DataPath_RF_bus_reg_dataout_1371_port, regs(1370) =>
                           DataPath_RF_bus_reg_dataout_1370_port, regs(1369) =>
                           DataPath_RF_bus_reg_dataout_1369_port, regs(1368) =>
                           DataPath_RF_bus_reg_dataout_1368_port, regs(1367) =>
                           DataPath_RF_bus_reg_dataout_1367_port, regs(1366) =>
                           DataPath_RF_bus_reg_dataout_1366_port, regs(1365) =>
                           DataPath_RF_bus_reg_dataout_1365_port, regs(1364) =>
                           DataPath_RF_bus_reg_dataout_1364_port, regs(1363) =>
                           DataPath_RF_bus_reg_dataout_1363_port, regs(1362) =>
                           DataPath_RF_bus_reg_dataout_1362_port, regs(1361) =>
                           DataPath_RF_bus_reg_dataout_1361_port, regs(1360) =>
                           DataPath_RF_bus_reg_dataout_1360_port, regs(1359) =>
                           DataPath_RF_bus_reg_dataout_1359_port, regs(1358) =>
                           DataPath_RF_bus_reg_dataout_1358_port, regs(1357) =>
                           DataPath_RF_bus_reg_dataout_1357_port, regs(1356) =>
                           DataPath_RF_bus_reg_dataout_1356_port, regs(1355) =>
                           DataPath_RF_bus_reg_dataout_1355_port, regs(1354) =>
                           DataPath_RF_bus_reg_dataout_1354_port, regs(1353) =>
                           DataPath_RF_bus_reg_dataout_1353_port, regs(1352) =>
                           DataPath_RF_bus_reg_dataout_1352_port, regs(1351) =>
                           DataPath_RF_bus_reg_dataout_1351_port, regs(1350) =>
                           DataPath_RF_bus_reg_dataout_1350_port, regs(1349) =>
                           DataPath_RF_bus_reg_dataout_1349_port, regs(1348) =>
                           DataPath_RF_bus_reg_dataout_1348_port, regs(1347) =>
                           DataPath_RF_bus_reg_dataout_1347_port, regs(1346) =>
                           DataPath_RF_bus_reg_dataout_1346_port, regs(1345) =>
                           DataPath_RF_bus_reg_dataout_1345_port, regs(1344) =>
                           DataPath_RF_bus_reg_dataout_1344_port, regs(1343) =>
                           DataPath_RF_bus_reg_dataout_1343_port, regs(1342) =>
                           DataPath_RF_bus_reg_dataout_1342_port, regs(1341) =>
                           DataPath_RF_bus_reg_dataout_1341_port, regs(1340) =>
                           DataPath_RF_bus_reg_dataout_1340_port, regs(1339) =>
                           DataPath_RF_bus_reg_dataout_1339_port, regs(1338) =>
                           DataPath_RF_bus_reg_dataout_1338_port, regs(1337) =>
                           DataPath_RF_bus_reg_dataout_1337_port, regs(1336) =>
                           DataPath_RF_bus_reg_dataout_1336_port, regs(1335) =>
                           DataPath_RF_bus_reg_dataout_1335_port, regs(1334) =>
                           DataPath_RF_bus_reg_dataout_1334_port, regs(1333) =>
                           DataPath_RF_bus_reg_dataout_1333_port, regs(1332) =>
                           DataPath_RF_bus_reg_dataout_1332_port, regs(1331) =>
                           DataPath_RF_bus_reg_dataout_1331_port, regs(1330) =>
                           DataPath_RF_bus_reg_dataout_1330_port, regs(1329) =>
                           DataPath_RF_bus_reg_dataout_1329_port, regs(1328) =>
                           DataPath_RF_bus_reg_dataout_1328_port, regs(1327) =>
                           DataPath_RF_bus_reg_dataout_1327_port, regs(1326) =>
                           DataPath_RF_bus_reg_dataout_1326_port, regs(1325) =>
                           DataPath_RF_bus_reg_dataout_1325_port, regs(1324) =>
                           DataPath_RF_bus_reg_dataout_1324_port, regs(1323) =>
                           DataPath_RF_bus_reg_dataout_1323_port, regs(1322) =>
                           DataPath_RF_bus_reg_dataout_1322_port, regs(1321) =>
                           DataPath_RF_bus_reg_dataout_1321_port, regs(1320) =>
                           DataPath_RF_bus_reg_dataout_1320_port, regs(1319) =>
                           DataPath_RF_bus_reg_dataout_1319_port, regs(1318) =>
                           DataPath_RF_bus_reg_dataout_1318_port, regs(1317) =>
                           DataPath_RF_bus_reg_dataout_1317_port, regs(1316) =>
                           DataPath_RF_bus_reg_dataout_1316_port, regs(1315) =>
                           DataPath_RF_bus_reg_dataout_1315_port, regs(1314) =>
                           DataPath_RF_bus_reg_dataout_1314_port, regs(1313) =>
                           DataPath_RF_bus_reg_dataout_1313_port, regs(1312) =>
                           DataPath_RF_bus_reg_dataout_1312_port, regs(1311) =>
                           DataPath_RF_bus_reg_dataout_1311_port, regs(1310) =>
                           DataPath_RF_bus_reg_dataout_1310_port, regs(1309) =>
                           DataPath_RF_bus_reg_dataout_1309_port, regs(1308) =>
                           DataPath_RF_bus_reg_dataout_1308_port, regs(1307) =>
                           DataPath_RF_bus_reg_dataout_1307_port, regs(1306) =>
                           DataPath_RF_bus_reg_dataout_1306_port, regs(1305) =>
                           DataPath_RF_bus_reg_dataout_1305_port, regs(1304) =>
                           DataPath_RF_bus_reg_dataout_1304_port, regs(1303) =>
                           DataPath_RF_bus_reg_dataout_1303_port, regs(1302) =>
                           DataPath_RF_bus_reg_dataout_1302_port, regs(1301) =>
                           DataPath_RF_bus_reg_dataout_1301_port, regs(1300) =>
                           DataPath_RF_bus_reg_dataout_1300_port, regs(1299) =>
                           DataPath_RF_bus_reg_dataout_1299_port, regs(1298) =>
                           DataPath_RF_bus_reg_dataout_1298_port, regs(1297) =>
                           DataPath_RF_bus_reg_dataout_1297_port, regs(1296) =>
                           DataPath_RF_bus_reg_dataout_1296_port, regs(1295) =>
                           DataPath_RF_bus_reg_dataout_1295_port, regs(1294) =>
                           DataPath_RF_bus_reg_dataout_1294_port, regs(1293) =>
                           DataPath_RF_bus_reg_dataout_1293_port, regs(1292) =>
                           DataPath_RF_bus_reg_dataout_1292_port, regs(1291) =>
                           DataPath_RF_bus_reg_dataout_1291_port, regs(1290) =>
                           DataPath_RF_bus_reg_dataout_1290_port, regs(1289) =>
                           DataPath_RF_bus_reg_dataout_1289_port, regs(1288) =>
                           DataPath_RF_bus_reg_dataout_1288_port, regs(1287) =>
                           DataPath_RF_bus_reg_dataout_1287_port, regs(1286) =>
                           DataPath_RF_bus_reg_dataout_1286_port, regs(1285) =>
                           DataPath_RF_bus_reg_dataout_1285_port, regs(1284) =>
                           DataPath_RF_bus_reg_dataout_1284_port, regs(1283) =>
                           DataPath_RF_bus_reg_dataout_1283_port, regs(1282) =>
                           DataPath_RF_bus_reg_dataout_1282_port, regs(1281) =>
                           DataPath_RF_bus_reg_dataout_1281_port, regs(1280) =>
                           DataPath_RF_bus_reg_dataout_1280_port, regs(1279) =>
                           DataPath_RF_bus_reg_dataout_1279_port, regs(1278) =>
                           DataPath_RF_bus_reg_dataout_1278_port, regs(1277) =>
                           DataPath_RF_bus_reg_dataout_1277_port, regs(1276) =>
                           DataPath_RF_bus_reg_dataout_1276_port, regs(1275) =>
                           DataPath_RF_bus_reg_dataout_1275_port, regs(1274) =>
                           DataPath_RF_bus_reg_dataout_1274_port, regs(1273) =>
                           DataPath_RF_bus_reg_dataout_1273_port, regs(1272) =>
                           DataPath_RF_bus_reg_dataout_1272_port, regs(1271) =>
                           DataPath_RF_bus_reg_dataout_1271_port, regs(1270) =>
                           DataPath_RF_bus_reg_dataout_1270_port, regs(1269) =>
                           DataPath_RF_bus_reg_dataout_1269_port, regs(1268) =>
                           DataPath_RF_bus_reg_dataout_1268_port, regs(1267) =>
                           DataPath_RF_bus_reg_dataout_1267_port, regs(1266) =>
                           DataPath_RF_bus_reg_dataout_1266_port, regs(1265) =>
                           DataPath_RF_bus_reg_dataout_1265_port, regs(1264) =>
                           DataPath_RF_bus_reg_dataout_1264_port, regs(1263) =>
                           DataPath_RF_bus_reg_dataout_1263_port, regs(1262) =>
                           DataPath_RF_bus_reg_dataout_1262_port, regs(1261) =>
                           DataPath_RF_bus_reg_dataout_1261_port, regs(1260) =>
                           DataPath_RF_bus_reg_dataout_1260_port, regs(1259) =>
                           DataPath_RF_bus_reg_dataout_1259_port, regs(1258) =>
                           DataPath_RF_bus_reg_dataout_1258_port, regs(1257) =>
                           DataPath_RF_bus_reg_dataout_1257_port, regs(1256) =>
                           DataPath_RF_bus_reg_dataout_1256_port, regs(1255) =>
                           DataPath_RF_bus_reg_dataout_1255_port, regs(1254) =>
                           DataPath_RF_bus_reg_dataout_1254_port, regs(1253) =>
                           DataPath_RF_bus_reg_dataout_1253_port, regs(1252) =>
                           DataPath_RF_bus_reg_dataout_1252_port, regs(1251) =>
                           DataPath_RF_bus_reg_dataout_1251_port, regs(1250) =>
                           DataPath_RF_bus_reg_dataout_1250_port, regs(1249) =>
                           DataPath_RF_bus_reg_dataout_1249_port, regs(1248) =>
                           DataPath_RF_bus_reg_dataout_1248_port, regs(1247) =>
                           DataPath_RF_bus_reg_dataout_1247_port, regs(1246) =>
                           DataPath_RF_bus_reg_dataout_1246_port, regs(1245) =>
                           DataPath_RF_bus_reg_dataout_1245_port, regs(1244) =>
                           DataPath_RF_bus_reg_dataout_1244_port, regs(1243) =>
                           DataPath_RF_bus_reg_dataout_1243_port, regs(1242) =>
                           DataPath_RF_bus_reg_dataout_1242_port, regs(1241) =>
                           DataPath_RF_bus_reg_dataout_1241_port, regs(1240) =>
                           DataPath_RF_bus_reg_dataout_1240_port, regs(1239) =>
                           DataPath_RF_bus_reg_dataout_1239_port, regs(1238) =>
                           DataPath_RF_bus_reg_dataout_1238_port, regs(1237) =>
                           DataPath_RF_bus_reg_dataout_1237_port, regs(1236) =>
                           DataPath_RF_bus_reg_dataout_1236_port, regs(1235) =>
                           DataPath_RF_bus_reg_dataout_1235_port, regs(1234) =>
                           DataPath_RF_bus_reg_dataout_1234_port, regs(1233) =>
                           DataPath_RF_bus_reg_dataout_1233_port, regs(1232) =>
                           DataPath_RF_bus_reg_dataout_1232_port, regs(1231) =>
                           DataPath_RF_bus_reg_dataout_1231_port, regs(1230) =>
                           DataPath_RF_bus_reg_dataout_1230_port, regs(1229) =>
                           DataPath_RF_bus_reg_dataout_1229_port, regs(1228) =>
                           DataPath_RF_bus_reg_dataout_1228_port, regs(1227) =>
                           DataPath_RF_bus_reg_dataout_1227_port, regs(1226) =>
                           DataPath_RF_bus_reg_dataout_1226_port, regs(1225) =>
                           DataPath_RF_bus_reg_dataout_1225_port, regs(1224) =>
                           DataPath_RF_bus_reg_dataout_1224_port, regs(1223) =>
                           DataPath_RF_bus_reg_dataout_1223_port, regs(1222) =>
                           DataPath_RF_bus_reg_dataout_1222_port, regs(1221) =>
                           DataPath_RF_bus_reg_dataout_1221_port, regs(1220) =>
                           DataPath_RF_bus_reg_dataout_1220_port, regs(1219) =>
                           DataPath_RF_bus_reg_dataout_1219_port, regs(1218) =>
                           DataPath_RF_bus_reg_dataout_1218_port, regs(1217) =>
                           DataPath_RF_bus_reg_dataout_1217_port, regs(1216) =>
                           DataPath_RF_bus_reg_dataout_1216_port, regs(1215) =>
                           DataPath_RF_bus_reg_dataout_1215_port, regs(1214) =>
                           DataPath_RF_bus_reg_dataout_1214_port, regs(1213) =>
                           DataPath_RF_bus_reg_dataout_1213_port, regs(1212) =>
                           DataPath_RF_bus_reg_dataout_1212_port, regs(1211) =>
                           DataPath_RF_bus_reg_dataout_1211_port, regs(1210) =>
                           DataPath_RF_bus_reg_dataout_1210_port, regs(1209) =>
                           DataPath_RF_bus_reg_dataout_1209_port, regs(1208) =>
                           DataPath_RF_bus_reg_dataout_1208_port, regs(1207) =>
                           DataPath_RF_bus_reg_dataout_1207_port, regs(1206) =>
                           DataPath_RF_bus_reg_dataout_1206_port, regs(1205) =>
                           DataPath_RF_bus_reg_dataout_1205_port, regs(1204) =>
                           DataPath_RF_bus_reg_dataout_1204_port, regs(1203) =>
                           DataPath_RF_bus_reg_dataout_1203_port, regs(1202) =>
                           DataPath_RF_bus_reg_dataout_1202_port, regs(1201) =>
                           DataPath_RF_bus_reg_dataout_1201_port, regs(1200) =>
                           DataPath_RF_bus_reg_dataout_1200_port, regs(1199) =>
                           DataPath_RF_bus_reg_dataout_1199_port, regs(1198) =>
                           DataPath_RF_bus_reg_dataout_1198_port, regs(1197) =>
                           DataPath_RF_bus_reg_dataout_1197_port, regs(1196) =>
                           DataPath_RF_bus_reg_dataout_1196_port, regs(1195) =>
                           DataPath_RF_bus_reg_dataout_1195_port, regs(1194) =>
                           DataPath_RF_bus_reg_dataout_1194_port, regs(1193) =>
                           DataPath_RF_bus_reg_dataout_1193_port, regs(1192) =>
                           DataPath_RF_bus_reg_dataout_1192_port, regs(1191) =>
                           DataPath_RF_bus_reg_dataout_1191_port, regs(1190) =>
                           DataPath_RF_bus_reg_dataout_1190_port, regs(1189) =>
                           DataPath_RF_bus_reg_dataout_1189_port, regs(1188) =>
                           DataPath_RF_bus_reg_dataout_1188_port, regs(1187) =>
                           DataPath_RF_bus_reg_dataout_1187_port, regs(1186) =>
                           DataPath_RF_bus_reg_dataout_1186_port, regs(1185) =>
                           DataPath_RF_bus_reg_dataout_1185_port, regs(1184) =>
                           DataPath_RF_bus_reg_dataout_1184_port, regs(1183) =>
                           DataPath_RF_bus_reg_dataout_1183_port, regs(1182) =>
                           DataPath_RF_bus_reg_dataout_1182_port, regs(1181) =>
                           DataPath_RF_bus_reg_dataout_1181_port, regs(1180) =>
                           DataPath_RF_bus_reg_dataout_1180_port, regs(1179) =>
                           DataPath_RF_bus_reg_dataout_1179_port, regs(1178) =>
                           DataPath_RF_bus_reg_dataout_1178_port, regs(1177) =>
                           DataPath_RF_bus_reg_dataout_1177_port, regs(1176) =>
                           DataPath_RF_bus_reg_dataout_1176_port, regs(1175) =>
                           DataPath_RF_bus_reg_dataout_1175_port, regs(1174) =>
                           DataPath_RF_bus_reg_dataout_1174_port, regs(1173) =>
                           DataPath_RF_bus_reg_dataout_1173_port, regs(1172) =>
                           DataPath_RF_bus_reg_dataout_1172_port, regs(1171) =>
                           DataPath_RF_bus_reg_dataout_1171_port, regs(1170) =>
                           DataPath_RF_bus_reg_dataout_1170_port, regs(1169) =>
                           DataPath_RF_bus_reg_dataout_1169_port, regs(1168) =>
                           DataPath_RF_bus_reg_dataout_1168_port, regs(1167) =>
                           DataPath_RF_bus_reg_dataout_1167_port, regs(1166) =>
                           DataPath_RF_bus_reg_dataout_1166_port, regs(1165) =>
                           DataPath_RF_bus_reg_dataout_1165_port, regs(1164) =>
                           DataPath_RF_bus_reg_dataout_1164_port, regs(1163) =>
                           DataPath_RF_bus_reg_dataout_1163_port, regs(1162) =>
                           DataPath_RF_bus_reg_dataout_1162_port, regs(1161) =>
                           DataPath_RF_bus_reg_dataout_1161_port, regs(1160) =>
                           DataPath_RF_bus_reg_dataout_1160_port, regs(1159) =>
                           DataPath_RF_bus_reg_dataout_1159_port, regs(1158) =>
                           DataPath_RF_bus_reg_dataout_1158_port, regs(1157) =>
                           DataPath_RF_bus_reg_dataout_1157_port, regs(1156) =>
                           DataPath_RF_bus_reg_dataout_1156_port, regs(1155) =>
                           DataPath_RF_bus_reg_dataout_1155_port, regs(1154) =>
                           DataPath_RF_bus_reg_dataout_1154_port, regs(1153) =>
                           DataPath_RF_bus_reg_dataout_1153_port, regs(1152) =>
                           DataPath_RF_bus_reg_dataout_1152_port, regs(1151) =>
                           DataPath_RF_bus_reg_dataout_1151_port, regs(1150) =>
                           DataPath_RF_bus_reg_dataout_1150_port, regs(1149) =>
                           DataPath_RF_bus_reg_dataout_1149_port, regs(1148) =>
                           DataPath_RF_bus_reg_dataout_1148_port, regs(1147) =>
                           DataPath_RF_bus_reg_dataout_1147_port, regs(1146) =>
                           DataPath_RF_bus_reg_dataout_1146_port, regs(1145) =>
                           DataPath_RF_bus_reg_dataout_1145_port, regs(1144) =>
                           DataPath_RF_bus_reg_dataout_1144_port, regs(1143) =>
                           DataPath_RF_bus_reg_dataout_1143_port, regs(1142) =>
                           DataPath_RF_bus_reg_dataout_1142_port, regs(1141) =>
                           DataPath_RF_bus_reg_dataout_1141_port, regs(1140) =>
                           DataPath_RF_bus_reg_dataout_1140_port, regs(1139) =>
                           DataPath_RF_bus_reg_dataout_1139_port, regs(1138) =>
                           DataPath_RF_bus_reg_dataout_1138_port, regs(1137) =>
                           DataPath_RF_bus_reg_dataout_1137_port, regs(1136) =>
                           DataPath_RF_bus_reg_dataout_1136_port, regs(1135) =>
                           DataPath_RF_bus_reg_dataout_1135_port, regs(1134) =>
                           DataPath_RF_bus_reg_dataout_1134_port, regs(1133) =>
                           DataPath_RF_bus_reg_dataout_1133_port, regs(1132) =>
                           DataPath_RF_bus_reg_dataout_1132_port, regs(1131) =>
                           DataPath_RF_bus_reg_dataout_1131_port, regs(1130) =>
                           DataPath_RF_bus_reg_dataout_1130_port, regs(1129) =>
                           DataPath_RF_bus_reg_dataout_1129_port, regs(1128) =>
                           DataPath_RF_bus_reg_dataout_1128_port, regs(1127) =>
                           DataPath_RF_bus_reg_dataout_1127_port, regs(1126) =>
                           DataPath_RF_bus_reg_dataout_1126_port, regs(1125) =>
                           DataPath_RF_bus_reg_dataout_1125_port, regs(1124) =>
                           DataPath_RF_bus_reg_dataout_1124_port, regs(1123) =>
                           DataPath_RF_bus_reg_dataout_1123_port, regs(1122) =>
                           DataPath_RF_bus_reg_dataout_1122_port, regs(1121) =>
                           DataPath_RF_bus_reg_dataout_1121_port, regs(1120) =>
                           DataPath_RF_bus_reg_dataout_1120_port, regs(1119) =>
                           DataPath_RF_bus_reg_dataout_1119_port, regs(1118) =>
                           DataPath_RF_bus_reg_dataout_1118_port, regs(1117) =>
                           DataPath_RF_bus_reg_dataout_1117_port, regs(1116) =>
                           DataPath_RF_bus_reg_dataout_1116_port, regs(1115) =>
                           DataPath_RF_bus_reg_dataout_1115_port, regs(1114) =>
                           DataPath_RF_bus_reg_dataout_1114_port, regs(1113) =>
                           DataPath_RF_bus_reg_dataout_1113_port, regs(1112) =>
                           DataPath_RF_bus_reg_dataout_1112_port, regs(1111) =>
                           DataPath_RF_bus_reg_dataout_1111_port, regs(1110) =>
                           DataPath_RF_bus_reg_dataout_1110_port, regs(1109) =>
                           DataPath_RF_bus_reg_dataout_1109_port, regs(1108) =>
                           DataPath_RF_bus_reg_dataout_1108_port, regs(1107) =>
                           DataPath_RF_bus_reg_dataout_1107_port, regs(1106) =>
                           DataPath_RF_bus_reg_dataout_1106_port, regs(1105) =>
                           DataPath_RF_bus_reg_dataout_1105_port, regs(1104) =>
                           DataPath_RF_bus_reg_dataout_1104_port, regs(1103) =>
                           DataPath_RF_bus_reg_dataout_1103_port, regs(1102) =>
                           DataPath_RF_bus_reg_dataout_1102_port, regs(1101) =>
                           DataPath_RF_bus_reg_dataout_1101_port, regs(1100) =>
                           DataPath_RF_bus_reg_dataout_1100_port, regs(1099) =>
                           DataPath_RF_bus_reg_dataout_1099_port, regs(1098) =>
                           DataPath_RF_bus_reg_dataout_1098_port, regs(1097) =>
                           DataPath_RF_bus_reg_dataout_1097_port, regs(1096) =>
                           DataPath_RF_bus_reg_dataout_1096_port, regs(1095) =>
                           DataPath_RF_bus_reg_dataout_1095_port, regs(1094) =>
                           DataPath_RF_bus_reg_dataout_1094_port, regs(1093) =>
                           DataPath_RF_bus_reg_dataout_1093_port, regs(1092) =>
                           DataPath_RF_bus_reg_dataout_1092_port, regs(1091) =>
                           DataPath_RF_bus_reg_dataout_1091_port, regs(1090) =>
                           DataPath_RF_bus_reg_dataout_1090_port, regs(1089) =>
                           DataPath_RF_bus_reg_dataout_1089_port, regs(1088) =>
                           DataPath_RF_bus_reg_dataout_1088_port, regs(1087) =>
                           DataPath_RF_bus_reg_dataout_1087_port, regs(1086) =>
                           DataPath_RF_bus_reg_dataout_1086_port, regs(1085) =>
                           DataPath_RF_bus_reg_dataout_1085_port, regs(1084) =>
                           DataPath_RF_bus_reg_dataout_1084_port, regs(1083) =>
                           DataPath_RF_bus_reg_dataout_1083_port, regs(1082) =>
                           DataPath_RF_bus_reg_dataout_1082_port, regs(1081) =>
                           DataPath_RF_bus_reg_dataout_1081_port, regs(1080) =>
                           DataPath_RF_bus_reg_dataout_1080_port, regs(1079) =>
                           DataPath_RF_bus_reg_dataout_1079_port, regs(1078) =>
                           DataPath_RF_bus_reg_dataout_1078_port, regs(1077) =>
                           DataPath_RF_bus_reg_dataout_1077_port, regs(1076) =>
                           DataPath_RF_bus_reg_dataout_1076_port, regs(1075) =>
                           DataPath_RF_bus_reg_dataout_1075_port, regs(1074) =>
                           DataPath_RF_bus_reg_dataout_1074_port, regs(1073) =>
                           DataPath_RF_bus_reg_dataout_1073_port, regs(1072) =>
                           DataPath_RF_bus_reg_dataout_1072_port, regs(1071) =>
                           DataPath_RF_bus_reg_dataout_1071_port, regs(1070) =>
                           DataPath_RF_bus_reg_dataout_1070_port, regs(1069) =>
                           DataPath_RF_bus_reg_dataout_1069_port, regs(1068) =>
                           DataPath_RF_bus_reg_dataout_1068_port, regs(1067) =>
                           DataPath_RF_bus_reg_dataout_1067_port, regs(1066) =>
                           DataPath_RF_bus_reg_dataout_1066_port, regs(1065) =>
                           DataPath_RF_bus_reg_dataout_1065_port, regs(1064) =>
                           DataPath_RF_bus_reg_dataout_1064_port, regs(1063) =>
                           DataPath_RF_bus_reg_dataout_1063_port, regs(1062) =>
                           DataPath_RF_bus_reg_dataout_1062_port, regs(1061) =>
                           DataPath_RF_bus_reg_dataout_1061_port, regs(1060) =>
                           DataPath_RF_bus_reg_dataout_1060_port, regs(1059) =>
                           DataPath_RF_bus_reg_dataout_1059_port, regs(1058) =>
                           DataPath_RF_bus_reg_dataout_1058_port, regs(1057) =>
                           DataPath_RF_bus_reg_dataout_1057_port, regs(1056) =>
                           DataPath_RF_bus_reg_dataout_1056_port, regs(1055) =>
                           DataPath_RF_bus_reg_dataout_1055_port, regs(1054) =>
                           DataPath_RF_bus_reg_dataout_1054_port, regs(1053) =>
                           DataPath_RF_bus_reg_dataout_1053_port, regs(1052) =>
                           DataPath_RF_bus_reg_dataout_1052_port, regs(1051) =>
                           DataPath_RF_bus_reg_dataout_1051_port, regs(1050) =>
                           DataPath_RF_bus_reg_dataout_1050_port, regs(1049) =>
                           DataPath_RF_bus_reg_dataout_1049_port, regs(1048) =>
                           DataPath_RF_bus_reg_dataout_1048_port, regs(1047) =>
                           DataPath_RF_bus_reg_dataout_1047_port, regs(1046) =>
                           DataPath_RF_bus_reg_dataout_1046_port, regs(1045) =>
                           DataPath_RF_bus_reg_dataout_1045_port, regs(1044) =>
                           DataPath_RF_bus_reg_dataout_1044_port, regs(1043) =>
                           DataPath_RF_bus_reg_dataout_1043_port, regs(1042) =>
                           DataPath_RF_bus_reg_dataout_1042_port, regs(1041) =>
                           DataPath_RF_bus_reg_dataout_1041_port, regs(1040) =>
                           DataPath_RF_bus_reg_dataout_1040_port, regs(1039) =>
                           DataPath_RF_bus_reg_dataout_1039_port, regs(1038) =>
                           DataPath_RF_bus_reg_dataout_1038_port, regs(1037) =>
                           DataPath_RF_bus_reg_dataout_1037_port, regs(1036) =>
                           DataPath_RF_bus_reg_dataout_1036_port, regs(1035) =>
                           DataPath_RF_bus_reg_dataout_1035_port, regs(1034) =>
                           DataPath_RF_bus_reg_dataout_1034_port, regs(1033) =>
                           DataPath_RF_bus_reg_dataout_1033_port, regs(1032) =>
                           DataPath_RF_bus_reg_dataout_1032_port, regs(1031) =>
                           DataPath_RF_bus_reg_dataout_1031_port, regs(1030) =>
                           DataPath_RF_bus_reg_dataout_1030_port, regs(1029) =>
                           DataPath_RF_bus_reg_dataout_1029_port, regs(1028) =>
                           DataPath_RF_bus_reg_dataout_1028_port, regs(1027) =>
                           DataPath_RF_bus_reg_dataout_1027_port, regs(1026) =>
                           DataPath_RF_bus_reg_dataout_1026_port, regs(1025) =>
                           DataPath_RF_bus_reg_dataout_1025_port, regs(1024) =>
                           DataPath_RF_bus_reg_dataout_1024_port, regs(1023) =>
                           DataPath_RF_bus_reg_dataout_1023_port, regs(1022) =>
                           DataPath_RF_bus_reg_dataout_1022_port, regs(1021) =>
                           DataPath_RF_bus_reg_dataout_1021_port, regs(1020) =>
                           DataPath_RF_bus_reg_dataout_1020_port, regs(1019) =>
                           DataPath_RF_bus_reg_dataout_1019_port, regs(1018) =>
                           DataPath_RF_bus_reg_dataout_1018_port, regs(1017) =>
                           DataPath_RF_bus_reg_dataout_1017_port, regs(1016) =>
                           DataPath_RF_bus_reg_dataout_1016_port, regs(1015) =>
                           DataPath_RF_bus_reg_dataout_1015_port, regs(1014) =>
                           DataPath_RF_bus_reg_dataout_1014_port, regs(1013) =>
                           DataPath_RF_bus_reg_dataout_1013_port, regs(1012) =>
                           DataPath_RF_bus_reg_dataout_1012_port, regs(1011) =>
                           DataPath_RF_bus_reg_dataout_1011_port, regs(1010) =>
                           DataPath_RF_bus_reg_dataout_1010_port, regs(1009) =>
                           DataPath_RF_bus_reg_dataout_1009_port, regs(1008) =>
                           DataPath_RF_bus_reg_dataout_1008_port, regs(1007) =>
                           DataPath_RF_bus_reg_dataout_1007_port, regs(1006) =>
                           DataPath_RF_bus_reg_dataout_1006_port, regs(1005) =>
                           DataPath_RF_bus_reg_dataout_1005_port, regs(1004) =>
                           DataPath_RF_bus_reg_dataout_1004_port, regs(1003) =>
                           DataPath_RF_bus_reg_dataout_1003_port, regs(1002) =>
                           DataPath_RF_bus_reg_dataout_1002_port, regs(1001) =>
                           DataPath_RF_bus_reg_dataout_1001_port, regs(1000) =>
                           DataPath_RF_bus_reg_dataout_1000_port, regs(999) => 
                           DataPath_RF_bus_reg_dataout_999_port, regs(998) => 
                           DataPath_RF_bus_reg_dataout_998_port, regs(997) => 
                           DataPath_RF_bus_reg_dataout_997_port, regs(996) => 
                           DataPath_RF_bus_reg_dataout_996_port, regs(995) => 
                           DataPath_RF_bus_reg_dataout_995_port, regs(994) => 
                           DataPath_RF_bus_reg_dataout_994_port, regs(993) => 
                           DataPath_RF_bus_reg_dataout_993_port, regs(992) => 
                           DataPath_RF_bus_reg_dataout_992_port, regs(991) => 
                           DataPath_RF_bus_reg_dataout_991_port, regs(990) => 
                           DataPath_RF_bus_reg_dataout_990_port, regs(989) => 
                           DataPath_RF_bus_reg_dataout_989_port, regs(988) => 
                           DataPath_RF_bus_reg_dataout_988_port, regs(987) => 
                           DataPath_RF_bus_reg_dataout_987_port, regs(986) => 
                           DataPath_RF_bus_reg_dataout_986_port, regs(985) => 
                           DataPath_RF_bus_reg_dataout_985_port, regs(984) => 
                           DataPath_RF_bus_reg_dataout_984_port, regs(983) => 
                           DataPath_RF_bus_reg_dataout_983_port, regs(982) => 
                           DataPath_RF_bus_reg_dataout_982_port, regs(981) => 
                           DataPath_RF_bus_reg_dataout_981_port, regs(980) => 
                           DataPath_RF_bus_reg_dataout_980_port, regs(979) => 
                           DataPath_RF_bus_reg_dataout_979_port, regs(978) => 
                           DataPath_RF_bus_reg_dataout_978_port, regs(977) => 
                           DataPath_RF_bus_reg_dataout_977_port, regs(976) => 
                           DataPath_RF_bus_reg_dataout_976_port, regs(975) => 
                           DataPath_RF_bus_reg_dataout_975_port, regs(974) => 
                           DataPath_RF_bus_reg_dataout_974_port, regs(973) => 
                           DataPath_RF_bus_reg_dataout_973_port, regs(972) => 
                           DataPath_RF_bus_reg_dataout_972_port, regs(971) => 
                           DataPath_RF_bus_reg_dataout_971_port, regs(970) => 
                           DataPath_RF_bus_reg_dataout_970_port, regs(969) => 
                           DataPath_RF_bus_reg_dataout_969_port, regs(968) => 
                           DataPath_RF_bus_reg_dataout_968_port, regs(967) => 
                           DataPath_RF_bus_reg_dataout_967_port, regs(966) => 
                           DataPath_RF_bus_reg_dataout_966_port, regs(965) => 
                           DataPath_RF_bus_reg_dataout_965_port, regs(964) => 
                           DataPath_RF_bus_reg_dataout_964_port, regs(963) => 
                           DataPath_RF_bus_reg_dataout_963_port, regs(962) => 
                           DataPath_RF_bus_reg_dataout_962_port, regs(961) => 
                           DataPath_RF_bus_reg_dataout_961_port, regs(960) => 
                           DataPath_RF_bus_reg_dataout_960_port, regs(959) => 
                           DataPath_RF_bus_reg_dataout_959_port, regs(958) => 
                           DataPath_RF_bus_reg_dataout_958_port, regs(957) => 
                           DataPath_RF_bus_reg_dataout_957_port, regs(956) => 
                           DataPath_RF_bus_reg_dataout_956_port, regs(955) => 
                           DataPath_RF_bus_reg_dataout_955_port, regs(954) => 
                           DataPath_RF_bus_reg_dataout_954_port, regs(953) => 
                           DataPath_RF_bus_reg_dataout_953_port, regs(952) => 
                           DataPath_RF_bus_reg_dataout_952_port, regs(951) => 
                           DataPath_RF_bus_reg_dataout_951_port, regs(950) => 
                           DataPath_RF_bus_reg_dataout_950_port, regs(949) => 
                           DataPath_RF_bus_reg_dataout_949_port, regs(948) => 
                           DataPath_RF_bus_reg_dataout_948_port, regs(947) => 
                           DataPath_RF_bus_reg_dataout_947_port, regs(946) => 
                           DataPath_RF_bus_reg_dataout_946_port, regs(945) => 
                           DataPath_RF_bus_reg_dataout_945_port, regs(944) => 
                           DataPath_RF_bus_reg_dataout_944_port, regs(943) => 
                           DataPath_RF_bus_reg_dataout_943_port, regs(942) => 
                           DataPath_RF_bus_reg_dataout_942_port, regs(941) => 
                           DataPath_RF_bus_reg_dataout_941_port, regs(940) => 
                           DataPath_RF_bus_reg_dataout_940_port, regs(939) => 
                           DataPath_RF_bus_reg_dataout_939_port, regs(938) => 
                           DataPath_RF_bus_reg_dataout_938_port, regs(937) => 
                           DataPath_RF_bus_reg_dataout_937_port, regs(936) => 
                           DataPath_RF_bus_reg_dataout_936_port, regs(935) => 
                           DataPath_RF_bus_reg_dataout_935_port, regs(934) => 
                           DataPath_RF_bus_reg_dataout_934_port, regs(933) => 
                           DataPath_RF_bus_reg_dataout_933_port, regs(932) => 
                           DataPath_RF_bus_reg_dataout_932_port, regs(931) => 
                           DataPath_RF_bus_reg_dataout_931_port, regs(930) => 
                           DataPath_RF_bus_reg_dataout_930_port, regs(929) => 
                           DataPath_RF_bus_reg_dataout_929_port, regs(928) => 
                           DataPath_RF_bus_reg_dataout_928_port, regs(927) => 
                           DataPath_RF_bus_reg_dataout_927_port, regs(926) => 
                           DataPath_RF_bus_reg_dataout_926_port, regs(925) => 
                           DataPath_RF_bus_reg_dataout_925_port, regs(924) => 
                           DataPath_RF_bus_reg_dataout_924_port, regs(923) => 
                           DataPath_RF_bus_reg_dataout_923_port, regs(922) => 
                           DataPath_RF_bus_reg_dataout_922_port, regs(921) => 
                           DataPath_RF_bus_reg_dataout_921_port, regs(920) => 
                           DataPath_RF_bus_reg_dataout_920_port, regs(919) => 
                           DataPath_RF_bus_reg_dataout_919_port, regs(918) => 
                           DataPath_RF_bus_reg_dataout_918_port, regs(917) => 
                           DataPath_RF_bus_reg_dataout_917_port, regs(916) => 
                           DataPath_RF_bus_reg_dataout_916_port, regs(915) => 
                           DataPath_RF_bus_reg_dataout_915_port, regs(914) => 
                           DataPath_RF_bus_reg_dataout_914_port, regs(913) => 
                           DataPath_RF_bus_reg_dataout_913_port, regs(912) => 
                           DataPath_RF_bus_reg_dataout_912_port, regs(911) => 
                           DataPath_RF_bus_reg_dataout_911_port, regs(910) => 
                           DataPath_RF_bus_reg_dataout_910_port, regs(909) => 
                           DataPath_RF_bus_reg_dataout_909_port, regs(908) => 
                           DataPath_RF_bus_reg_dataout_908_port, regs(907) => 
                           DataPath_RF_bus_reg_dataout_907_port, regs(906) => 
                           DataPath_RF_bus_reg_dataout_906_port, regs(905) => 
                           DataPath_RF_bus_reg_dataout_905_port, regs(904) => 
                           DataPath_RF_bus_reg_dataout_904_port, regs(903) => 
                           DataPath_RF_bus_reg_dataout_903_port, regs(902) => 
                           DataPath_RF_bus_reg_dataout_902_port, regs(901) => 
                           DataPath_RF_bus_reg_dataout_901_port, regs(900) => 
                           DataPath_RF_bus_reg_dataout_900_port, regs(899) => 
                           DataPath_RF_bus_reg_dataout_899_port, regs(898) => 
                           DataPath_RF_bus_reg_dataout_898_port, regs(897) => 
                           DataPath_RF_bus_reg_dataout_897_port, regs(896) => 
                           DataPath_RF_bus_reg_dataout_896_port, regs(895) => 
                           DataPath_RF_bus_reg_dataout_895_port, regs(894) => 
                           DataPath_RF_bus_reg_dataout_894_port, regs(893) => 
                           DataPath_RF_bus_reg_dataout_893_port, regs(892) => 
                           DataPath_RF_bus_reg_dataout_892_port, regs(891) => 
                           DataPath_RF_bus_reg_dataout_891_port, regs(890) => 
                           DataPath_RF_bus_reg_dataout_890_port, regs(889) => 
                           DataPath_RF_bus_reg_dataout_889_port, regs(888) => 
                           DataPath_RF_bus_reg_dataout_888_port, regs(887) => 
                           DataPath_RF_bus_reg_dataout_887_port, regs(886) => 
                           DataPath_RF_bus_reg_dataout_886_port, regs(885) => 
                           DataPath_RF_bus_reg_dataout_885_port, regs(884) => 
                           DataPath_RF_bus_reg_dataout_884_port, regs(883) => 
                           DataPath_RF_bus_reg_dataout_883_port, regs(882) => 
                           DataPath_RF_bus_reg_dataout_882_port, regs(881) => 
                           DataPath_RF_bus_reg_dataout_881_port, regs(880) => 
                           DataPath_RF_bus_reg_dataout_880_port, regs(879) => 
                           DataPath_RF_bus_reg_dataout_879_port, regs(878) => 
                           DataPath_RF_bus_reg_dataout_878_port, regs(877) => 
                           DataPath_RF_bus_reg_dataout_877_port, regs(876) => 
                           DataPath_RF_bus_reg_dataout_876_port, regs(875) => 
                           DataPath_RF_bus_reg_dataout_875_port, regs(874) => 
                           DataPath_RF_bus_reg_dataout_874_port, regs(873) => 
                           DataPath_RF_bus_reg_dataout_873_port, regs(872) => 
                           DataPath_RF_bus_reg_dataout_872_port, regs(871) => 
                           DataPath_RF_bus_reg_dataout_871_port, regs(870) => 
                           DataPath_RF_bus_reg_dataout_870_port, regs(869) => 
                           DataPath_RF_bus_reg_dataout_869_port, regs(868) => 
                           DataPath_RF_bus_reg_dataout_868_port, regs(867) => 
                           DataPath_RF_bus_reg_dataout_867_port, regs(866) => 
                           DataPath_RF_bus_reg_dataout_866_port, regs(865) => 
                           DataPath_RF_bus_reg_dataout_865_port, regs(864) => 
                           DataPath_RF_bus_reg_dataout_864_port, regs(863) => 
                           DataPath_RF_bus_reg_dataout_863_port, regs(862) => 
                           DataPath_RF_bus_reg_dataout_862_port, regs(861) => 
                           DataPath_RF_bus_reg_dataout_861_port, regs(860) => 
                           DataPath_RF_bus_reg_dataout_860_port, regs(859) => 
                           DataPath_RF_bus_reg_dataout_859_port, regs(858) => 
                           DataPath_RF_bus_reg_dataout_858_port, regs(857) => 
                           DataPath_RF_bus_reg_dataout_857_port, regs(856) => 
                           DataPath_RF_bus_reg_dataout_856_port, regs(855) => 
                           DataPath_RF_bus_reg_dataout_855_port, regs(854) => 
                           DataPath_RF_bus_reg_dataout_854_port, regs(853) => 
                           DataPath_RF_bus_reg_dataout_853_port, regs(852) => 
                           DataPath_RF_bus_reg_dataout_852_port, regs(851) => 
                           DataPath_RF_bus_reg_dataout_851_port, regs(850) => 
                           DataPath_RF_bus_reg_dataout_850_port, regs(849) => 
                           DataPath_RF_bus_reg_dataout_849_port, regs(848) => 
                           DataPath_RF_bus_reg_dataout_848_port, regs(847) => 
                           DataPath_RF_bus_reg_dataout_847_port, regs(846) => 
                           DataPath_RF_bus_reg_dataout_846_port, regs(845) => 
                           DataPath_RF_bus_reg_dataout_845_port, regs(844) => 
                           DataPath_RF_bus_reg_dataout_844_port, regs(843) => 
                           DataPath_RF_bus_reg_dataout_843_port, regs(842) => 
                           DataPath_RF_bus_reg_dataout_842_port, regs(841) => 
                           DataPath_RF_bus_reg_dataout_841_port, regs(840) => 
                           DataPath_RF_bus_reg_dataout_840_port, regs(839) => 
                           DataPath_RF_bus_reg_dataout_839_port, regs(838) => 
                           DataPath_RF_bus_reg_dataout_838_port, regs(837) => 
                           DataPath_RF_bus_reg_dataout_837_port, regs(836) => 
                           DataPath_RF_bus_reg_dataout_836_port, regs(835) => 
                           DataPath_RF_bus_reg_dataout_835_port, regs(834) => 
                           DataPath_RF_bus_reg_dataout_834_port, regs(833) => 
                           DataPath_RF_bus_reg_dataout_833_port, regs(832) => 
                           DataPath_RF_bus_reg_dataout_832_port, regs(831) => 
                           DataPath_RF_bus_reg_dataout_831_port, regs(830) => 
                           DataPath_RF_bus_reg_dataout_830_port, regs(829) => 
                           DataPath_RF_bus_reg_dataout_829_port, regs(828) => 
                           DataPath_RF_bus_reg_dataout_828_port, regs(827) => 
                           DataPath_RF_bus_reg_dataout_827_port, regs(826) => 
                           DataPath_RF_bus_reg_dataout_826_port, regs(825) => 
                           DataPath_RF_bus_reg_dataout_825_port, regs(824) => 
                           DataPath_RF_bus_reg_dataout_824_port, regs(823) => 
                           DataPath_RF_bus_reg_dataout_823_port, regs(822) => 
                           DataPath_RF_bus_reg_dataout_822_port, regs(821) => 
                           DataPath_RF_bus_reg_dataout_821_port, regs(820) => 
                           DataPath_RF_bus_reg_dataout_820_port, regs(819) => 
                           DataPath_RF_bus_reg_dataout_819_port, regs(818) => 
                           DataPath_RF_bus_reg_dataout_818_port, regs(817) => 
                           DataPath_RF_bus_reg_dataout_817_port, regs(816) => 
                           DataPath_RF_bus_reg_dataout_816_port, regs(815) => 
                           DataPath_RF_bus_reg_dataout_815_port, regs(814) => 
                           DataPath_RF_bus_reg_dataout_814_port, regs(813) => 
                           DataPath_RF_bus_reg_dataout_813_port, regs(812) => 
                           DataPath_RF_bus_reg_dataout_812_port, regs(811) => 
                           DataPath_RF_bus_reg_dataout_811_port, regs(810) => 
                           DataPath_RF_bus_reg_dataout_810_port, regs(809) => 
                           DataPath_RF_bus_reg_dataout_809_port, regs(808) => 
                           DataPath_RF_bus_reg_dataout_808_port, regs(807) => 
                           DataPath_RF_bus_reg_dataout_807_port, regs(806) => 
                           DataPath_RF_bus_reg_dataout_806_port, regs(805) => 
                           DataPath_RF_bus_reg_dataout_805_port, regs(804) => 
                           DataPath_RF_bus_reg_dataout_804_port, regs(803) => 
                           DataPath_RF_bus_reg_dataout_803_port, regs(802) => 
                           DataPath_RF_bus_reg_dataout_802_port, regs(801) => 
                           DataPath_RF_bus_reg_dataout_801_port, regs(800) => 
                           DataPath_RF_bus_reg_dataout_800_port, regs(799) => 
                           DataPath_RF_bus_reg_dataout_799_port, regs(798) => 
                           DataPath_RF_bus_reg_dataout_798_port, regs(797) => 
                           DataPath_RF_bus_reg_dataout_797_port, regs(796) => 
                           DataPath_RF_bus_reg_dataout_796_port, regs(795) => 
                           DataPath_RF_bus_reg_dataout_795_port, regs(794) => 
                           DataPath_RF_bus_reg_dataout_794_port, regs(793) => 
                           DataPath_RF_bus_reg_dataout_793_port, regs(792) => 
                           DataPath_RF_bus_reg_dataout_792_port, regs(791) => 
                           DataPath_RF_bus_reg_dataout_791_port, regs(790) => 
                           DataPath_RF_bus_reg_dataout_790_port, regs(789) => 
                           DataPath_RF_bus_reg_dataout_789_port, regs(788) => 
                           DataPath_RF_bus_reg_dataout_788_port, regs(787) => 
                           DataPath_RF_bus_reg_dataout_787_port, regs(786) => 
                           DataPath_RF_bus_reg_dataout_786_port, regs(785) => 
                           DataPath_RF_bus_reg_dataout_785_port, regs(784) => 
                           DataPath_RF_bus_reg_dataout_784_port, regs(783) => 
                           DataPath_RF_bus_reg_dataout_783_port, regs(782) => 
                           DataPath_RF_bus_reg_dataout_782_port, regs(781) => 
                           DataPath_RF_bus_reg_dataout_781_port, regs(780) => 
                           DataPath_RF_bus_reg_dataout_780_port, regs(779) => 
                           DataPath_RF_bus_reg_dataout_779_port, regs(778) => 
                           DataPath_RF_bus_reg_dataout_778_port, regs(777) => 
                           DataPath_RF_bus_reg_dataout_777_port, regs(776) => 
                           DataPath_RF_bus_reg_dataout_776_port, regs(775) => 
                           DataPath_RF_bus_reg_dataout_775_port, regs(774) => 
                           DataPath_RF_bus_reg_dataout_774_port, regs(773) => 
                           DataPath_RF_bus_reg_dataout_773_port, regs(772) => 
                           DataPath_RF_bus_reg_dataout_772_port, regs(771) => 
                           DataPath_RF_bus_reg_dataout_771_port, regs(770) => 
                           DataPath_RF_bus_reg_dataout_770_port, regs(769) => 
                           DataPath_RF_bus_reg_dataout_769_port, regs(768) => 
                           DataPath_RF_bus_reg_dataout_768_port, regs(767) => 
                           DataPath_RF_bus_reg_dataout_767_port, regs(766) => 
                           DataPath_RF_bus_reg_dataout_766_port, regs(765) => 
                           DataPath_RF_bus_reg_dataout_765_port, regs(764) => 
                           DataPath_RF_bus_reg_dataout_764_port, regs(763) => 
                           DataPath_RF_bus_reg_dataout_763_port, regs(762) => 
                           DataPath_RF_bus_reg_dataout_762_port, regs(761) => 
                           DataPath_RF_bus_reg_dataout_761_port, regs(760) => 
                           DataPath_RF_bus_reg_dataout_760_port, regs(759) => 
                           DataPath_RF_bus_reg_dataout_759_port, regs(758) => 
                           DataPath_RF_bus_reg_dataout_758_port, regs(757) => 
                           DataPath_RF_bus_reg_dataout_757_port, regs(756) => 
                           DataPath_RF_bus_reg_dataout_756_port, regs(755) => 
                           DataPath_RF_bus_reg_dataout_755_port, regs(754) => 
                           DataPath_RF_bus_reg_dataout_754_port, regs(753) => 
                           DataPath_RF_bus_reg_dataout_753_port, regs(752) => 
                           DataPath_RF_bus_reg_dataout_752_port, regs(751) => 
                           DataPath_RF_bus_reg_dataout_751_port, regs(750) => 
                           DataPath_RF_bus_reg_dataout_750_port, regs(749) => 
                           DataPath_RF_bus_reg_dataout_749_port, regs(748) => 
                           DataPath_RF_bus_reg_dataout_748_port, regs(747) => 
                           DataPath_RF_bus_reg_dataout_747_port, regs(746) => 
                           DataPath_RF_bus_reg_dataout_746_port, regs(745) => 
                           DataPath_RF_bus_reg_dataout_745_port, regs(744) => 
                           DataPath_RF_bus_reg_dataout_744_port, regs(743) => 
                           DataPath_RF_bus_reg_dataout_743_port, regs(742) => 
                           DataPath_RF_bus_reg_dataout_742_port, regs(741) => 
                           DataPath_RF_bus_reg_dataout_741_port, regs(740) => 
                           DataPath_RF_bus_reg_dataout_740_port, regs(739) => 
                           DataPath_RF_bus_reg_dataout_739_port, regs(738) => 
                           DataPath_RF_bus_reg_dataout_738_port, regs(737) => 
                           DataPath_RF_bus_reg_dataout_737_port, regs(736) => 
                           DataPath_RF_bus_reg_dataout_736_port, regs(735) => 
                           DataPath_RF_bus_reg_dataout_735_port, regs(734) => 
                           DataPath_RF_bus_reg_dataout_734_port, regs(733) => 
                           DataPath_RF_bus_reg_dataout_733_port, regs(732) => 
                           DataPath_RF_bus_reg_dataout_732_port, regs(731) => 
                           DataPath_RF_bus_reg_dataout_731_port, regs(730) => 
                           DataPath_RF_bus_reg_dataout_730_port, regs(729) => 
                           DataPath_RF_bus_reg_dataout_729_port, regs(728) => 
                           DataPath_RF_bus_reg_dataout_728_port, regs(727) => 
                           DataPath_RF_bus_reg_dataout_727_port, regs(726) => 
                           DataPath_RF_bus_reg_dataout_726_port, regs(725) => 
                           DataPath_RF_bus_reg_dataout_725_port, regs(724) => 
                           DataPath_RF_bus_reg_dataout_724_port, regs(723) => 
                           DataPath_RF_bus_reg_dataout_723_port, regs(722) => 
                           DataPath_RF_bus_reg_dataout_722_port, regs(721) => 
                           DataPath_RF_bus_reg_dataout_721_port, regs(720) => 
                           DataPath_RF_bus_reg_dataout_720_port, regs(719) => 
                           DataPath_RF_bus_reg_dataout_719_port, regs(718) => 
                           DataPath_RF_bus_reg_dataout_718_port, regs(717) => 
                           DataPath_RF_bus_reg_dataout_717_port, regs(716) => 
                           DataPath_RF_bus_reg_dataout_716_port, regs(715) => 
                           DataPath_RF_bus_reg_dataout_715_port, regs(714) => 
                           DataPath_RF_bus_reg_dataout_714_port, regs(713) => 
                           DataPath_RF_bus_reg_dataout_713_port, regs(712) => 
                           DataPath_RF_bus_reg_dataout_712_port, regs(711) => 
                           DataPath_RF_bus_reg_dataout_711_port, regs(710) => 
                           DataPath_RF_bus_reg_dataout_710_port, regs(709) => 
                           DataPath_RF_bus_reg_dataout_709_port, regs(708) => 
                           DataPath_RF_bus_reg_dataout_708_port, regs(707) => 
                           DataPath_RF_bus_reg_dataout_707_port, regs(706) => 
                           DataPath_RF_bus_reg_dataout_706_port, regs(705) => 
                           DataPath_RF_bus_reg_dataout_705_port, regs(704) => 
                           DataPath_RF_bus_reg_dataout_704_port, regs(703) => 
                           DataPath_RF_bus_reg_dataout_703_port, regs(702) => 
                           DataPath_RF_bus_reg_dataout_702_port, regs(701) => 
                           DataPath_RF_bus_reg_dataout_701_port, regs(700) => 
                           DataPath_RF_bus_reg_dataout_700_port, regs(699) => 
                           DataPath_RF_bus_reg_dataout_699_port, regs(698) => 
                           DataPath_RF_bus_reg_dataout_698_port, regs(697) => 
                           DataPath_RF_bus_reg_dataout_697_port, regs(696) => 
                           DataPath_RF_bus_reg_dataout_696_port, regs(695) => 
                           DataPath_RF_bus_reg_dataout_695_port, regs(694) => 
                           DataPath_RF_bus_reg_dataout_694_port, regs(693) => 
                           DataPath_RF_bus_reg_dataout_693_port, regs(692) => 
                           DataPath_RF_bus_reg_dataout_692_port, regs(691) => 
                           DataPath_RF_bus_reg_dataout_691_port, regs(690) => 
                           DataPath_RF_bus_reg_dataout_690_port, regs(689) => 
                           DataPath_RF_bus_reg_dataout_689_port, regs(688) => 
                           DataPath_RF_bus_reg_dataout_688_port, regs(687) => 
                           DataPath_RF_bus_reg_dataout_687_port, regs(686) => 
                           DataPath_RF_bus_reg_dataout_686_port, regs(685) => 
                           DataPath_RF_bus_reg_dataout_685_port, regs(684) => 
                           DataPath_RF_bus_reg_dataout_684_port, regs(683) => 
                           DataPath_RF_bus_reg_dataout_683_port, regs(682) => 
                           DataPath_RF_bus_reg_dataout_682_port, regs(681) => 
                           DataPath_RF_bus_reg_dataout_681_port, regs(680) => 
                           DataPath_RF_bus_reg_dataout_680_port, regs(679) => 
                           DataPath_RF_bus_reg_dataout_679_port, regs(678) => 
                           DataPath_RF_bus_reg_dataout_678_port, regs(677) => 
                           DataPath_RF_bus_reg_dataout_677_port, regs(676) => 
                           DataPath_RF_bus_reg_dataout_676_port, regs(675) => 
                           DataPath_RF_bus_reg_dataout_675_port, regs(674) => 
                           DataPath_RF_bus_reg_dataout_674_port, regs(673) => 
                           DataPath_RF_bus_reg_dataout_673_port, regs(672) => 
                           DataPath_RF_bus_reg_dataout_672_port, regs(671) => 
                           DataPath_RF_bus_reg_dataout_671_port, regs(670) => 
                           DataPath_RF_bus_reg_dataout_670_port, regs(669) => 
                           DataPath_RF_bus_reg_dataout_669_port, regs(668) => 
                           DataPath_RF_bus_reg_dataout_668_port, regs(667) => 
                           DataPath_RF_bus_reg_dataout_667_port, regs(666) => 
                           DataPath_RF_bus_reg_dataout_666_port, regs(665) => 
                           DataPath_RF_bus_reg_dataout_665_port, regs(664) => 
                           DataPath_RF_bus_reg_dataout_664_port, regs(663) => 
                           DataPath_RF_bus_reg_dataout_663_port, regs(662) => 
                           DataPath_RF_bus_reg_dataout_662_port, regs(661) => 
                           DataPath_RF_bus_reg_dataout_661_port, regs(660) => 
                           DataPath_RF_bus_reg_dataout_660_port, regs(659) => 
                           DataPath_RF_bus_reg_dataout_659_port, regs(658) => 
                           DataPath_RF_bus_reg_dataout_658_port, regs(657) => 
                           DataPath_RF_bus_reg_dataout_657_port, regs(656) => 
                           DataPath_RF_bus_reg_dataout_656_port, regs(655) => 
                           DataPath_RF_bus_reg_dataout_655_port, regs(654) => 
                           DataPath_RF_bus_reg_dataout_654_port, regs(653) => 
                           DataPath_RF_bus_reg_dataout_653_port, regs(652) => 
                           DataPath_RF_bus_reg_dataout_652_port, regs(651) => 
                           DataPath_RF_bus_reg_dataout_651_port, regs(650) => 
                           DataPath_RF_bus_reg_dataout_650_port, regs(649) => 
                           DataPath_RF_bus_reg_dataout_649_port, regs(648) => 
                           DataPath_RF_bus_reg_dataout_648_port, regs(647) => 
                           DataPath_RF_bus_reg_dataout_647_port, regs(646) => 
                           DataPath_RF_bus_reg_dataout_646_port, regs(645) => 
                           DataPath_RF_bus_reg_dataout_645_port, regs(644) => 
                           DataPath_RF_bus_reg_dataout_644_port, regs(643) => 
                           DataPath_RF_bus_reg_dataout_643_port, regs(642) => 
                           DataPath_RF_bus_reg_dataout_642_port, regs(641) => 
                           DataPath_RF_bus_reg_dataout_641_port, regs(640) => 
                           DataPath_RF_bus_reg_dataout_640_port, regs(639) => 
                           DataPath_RF_bus_reg_dataout_639_port, regs(638) => 
                           DataPath_RF_bus_reg_dataout_638_port, regs(637) => 
                           DataPath_RF_bus_reg_dataout_637_port, regs(636) => 
                           DataPath_RF_bus_reg_dataout_636_port, regs(635) => 
                           DataPath_RF_bus_reg_dataout_635_port, regs(634) => 
                           DataPath_RF_bus_reg_dataout_634_port, regs(633) => 
                           DataPath_RF_bus_reg_dataout_633_port, regs(632) => 
                           DataPath_RF_bus_reg_dataout_632_port, regs(631) => 
                           DataPath_RF_bus_reg_dataout_631_port, regs(630) => 
                           DataPath_RF_bus_reg_dataout_630_port, regs(629) => 
                           DataPath_RF_bus_reg_dataout_629_port, regs(628) => 
                           DataPath_RF_bus_reg_dataout_628_port, regs(627) => 
                           DataPath_RF_bus_reg_dataout_627_port, regs(626) => 
                           DataPath_RF_bus_reg_dataout_626_port, regs(625) => 
                           DataPath_RF_bus_reg_dataout_625_port, regs(624) => 
                           DataPath_RF_bus_reg_dataout_624_port, regs(623) => 
                           DataPath_RF_bus_reg_dataout_623_port, regs(622) => 
                           DataPath_RF_bus_reg_dataout_622_port, regs(621) => 
                           DataPath_RF_bus_reg_dataout_621_port, regs(620) => 
                           DataPath_RF_bus_reg_dataout_620_port, regs(619) => 
                           DataPath_RF_bus_reg_dataout_619_port, regs(618) => 
                           DataPath_RF_bus_reg_dataout_618_port, regs(617) => 
                           DataPath_RF_bus_reg_dataout_617_port, regs(616) => 
                           DataPath_RF_bus_reg_dataout_616_port, regs(615) => 
                           DataPath_RF_bus_reg_dataout_615_port, regs(614) => 
                           DataPath_RF_bus_reg_dataout_614_port, regs(613) => 
                           DataPath_RF_bus_reg_dataout_613_port, regs(612) => 
                           DataPath_RF_bus_reg_dataout_612_port, regs(611) => 
                           DataPath_RF_bus_reg_dataout_611_port, regs(610) => 
                           DataPath_RF_bus_reg_dataout_610_port, regs(609) => 
                           DataPath_RF_bus_reg_dataout_609_port, regs(608) => 
                           DataPath_RF_bus_reg_dataout_608_port, regs(607) => 
                           DataPath_RF_bus_reg_dataout_607_port, regs(606) => 
                           DataPath_RF_bus_reg_dataout_606_port, regs(605) => 
                           DataPath_RF_bus_reg_dataout_605_port, regs(604) => 
                           DataPath_RF_bus_reg_dataout_604_port, regs(603) => 
                           DataPath_RF_bus_reg_dataout_603_port, regs(602) => 
                           DataPath_RF_bus_reg_dataout_602_port, regs(601) => 
                           DataPath_RF_bus_reg_dataout_601_port, regs(600) => 
                           DataPath_RF_bus_reg_dataout_600_port, regs(599) => 
                           DataPath_RF_bus_reg_dataout_599_port, regs(598) => 
                           DataPath_RF_bus_reg_dataout_598_port, regs(597) => 
                           DataPath_RF_bus_reg_dataout_597_port, regs(596) => 
                           DataPath_RF_bus_reg_dataout_596_port, regs(595) => 
                           DataPath_RF_bus_reg_dataout_595_port, regs(594) => 
                           DataPath_RF_bus_reg_dataout_594_port, regs(593) => 
                           DataPath_RF_bus_reg_dataout_593_port, regs(592) => 
                           DataPath_RF_bus_reg_dataout_592_port, regs(591) => 
                           DataPath_RF_bus_reg_dataout_591_port, regs(590) => 
                           DataPath_RF_bus_reg_dataout_590_port, regs(589) => 
                           DataPath_RF_bus_reg_dataout_589_port, regs(588) => 
                           DataPath_RF_bus_reg_dataout_588_port, regs(587) => 
                           DataPath_RF_bus_reg_dataout_587_port, regs(586) => 
                           DataPath_RF_bus_reg_dataout_586_port, regs(585) => 
                           DataPath_RF_bus_reg_dataout_585_port, regs(584) => 
                           DataPath_RF_bus_reg_dataout_584_port, regs(583) => 
                           DataPath_RF_bus_reg_dataout_583_port, regs(582) => 
                           DataPath_RF_bus_reg_dataout_582_port, regs(581) => 
                           DataPath_RF_bus_reg_dataout_581_port, regs(580) => 
                           DataPath_RF_bus_reg_dataout_580_port, regs(579) => 
                           DataPath_RF_bus_reg_dataout_579_port, regs(578) => 
                           DataPath_RF_bus_reg_dataout_578_port, regs(577) => 
                           DataPath_RF_bus_reg_dataout_577_port, regs(576) => 
                           DataPath_RF_bus_reg_dataout_576_port, regs(575) => 
                           DataPath_RF_bus_reg_dataout_575_port, regs(574) => 
                           DataPath_RF_bus_reg_dataout_574_port, regs(573) => 
                           DataPath_RF_bus_reg_dataout_573_port, regs(572) => 
                           DataPath_RF_bus_reg_dataout_572_port, regs(571) => 
                           DataPath_RF_bus_reg_dataout_571_port, regs(570) => 
                           DataPath_RF_bus_reg_dataout_570_port, regs(569) => 
                           DataPath_RF_bus_reg_dataout_569_port, regs(568) => 
                           DataPath_RF_bus_reg_dataout_568_port, regs(567) => 
                           DataPath_RF_bus_reg_dataout_567_port, regs(566) => 
                           DataPath_RF_bus_reg_dataout_566_port, regs(565) => 
                           DataPath_RF_bus_reg_dataout_565_port, regs(564) => 
                           DataPath_RF_bus_reg_dataout_564_port, regs(563) => 
                           DataPath_RF_bus_reg_dataout_563_port, regs(562) => 
                           DataPath_RF_bus_reg_dataout_562_port, regs(561) => 
                           DataPath_RF_bus_reg_dataout_561_port, regs(560) => 
                           DataPath_RF_bus_reg_dataout_560_port, regs(559) => 
                           DataPath_RF_bus_reg_dataout_559_port, regs(558) => 
                           DataPath_RF_bus_reg_dataout_558_port, regs(557) => 
                           DataPath_RF_bus_reg_dataout_557_port, regs(556) => 
                           DataPath_RF_bus_reg_dataout_556_port, regs(555) => 
                           DataPath_RF_bus_reg_dataout_555_port, regs(554) => 
                           DataPath_RF_bus_reg_dataout_554_port, regs(553) => 
                           DataPath_RF_bus_reg_dataout_553_port, regs(552) => 
                           DataPath_RF_bus_reg_dataout_552_port, regs(551) => 
                           DataPath_RF_bus_reg_dataout_551_port, regs(550) => 
                           DataPath_RF_bus_reg_dataout_550_port, regs(549) => 
                           DataPath_RF_bus_reg_dataout_549_port, regs(548) => 
                           DataPath_RF_bus_reg_dataout_548_port, regs(547) => 
                           DataPath_RF_bus_reg_dataout_547_port, regs(546) => 
                           DataPath_RF_bus_reg_dataout_546_port, regs(545) => 
                           DataPath_RF_bus_reg_dataout_545_port, regs(544) => 
                           DataPath_RF_bus_reg_dataout_544_port, regs(543) => 
                           DataPath_RF_bus_reg_dataout_543_port, regs(542) => 
                           DataPath_RF_bus_reg_dataout_542_port, regs(541) => 
                           DataPath_RF_bus_reg_dataout_541_port, regs(540) => 
                           DataPath_RF_bus_reg_dataout_540_port, regs(539) => 
                           DataPath_RF_bus_reg_dataout_539_port, regs(538) => 
                           DataPath_RF_bus_reg_dataout_538_port, regs(537) => 
                           DataPath_RF_bus_reg_dataout_537_port, regs(536) => 
                           DataPath_RF_bus_reg_dataout_536_port, regs(535) => 
                           DataPath_RF_bus_reg_dataout_535_port, regs(534) => 
                           DataPath_RF_bus_reg_dataout_534_port, regs(533) => 
                           DataPath_RF_bus_reg_dataout_533_port, regs(532) => 
                           DataPath_RF_bus_reg_dataout_532_port, regs(531) => 
                           DataPath_RF_bus_reg_dataout_531_port, regs(530) => 
                           DataPath_RF_bus_reg_dataout_530_port, regs(529) => 
                           DataPath_RF_bus_reg_dataout_529_port, regs(528) => 
                           DataPath_RF_bus_reg_dataout_528_port, regs(527) => 
                           DataPath_RF_bus_reg_dataout_527_port, regs(526) => 
                           DataPath_RF_bus_reg_dataout_526_port, regs(525) => 
                           DataPath_RF_bus_reg_dataout_525_port, regs(524) => 
                           DataPath_RF_bus_reg_dataout_524_port, regs(523) => 
                           DataPath_RF_bus_reg_dataout_523_port, regs(522) => 
                           DataPath_RF_bus_reg_dataout_522_port, regs(521) => 
                           DataPath_RF_bus_reg_dataout_521_port, regs(520) => 
                           DataPath_RF_bus_reg_dataout_520_port, regs(519) => 
                           DataPath_RF_bus_reg_dataout_519_port, regs(518) => 
                           DataPath_RF_bus_reg_dataout_518_port, regs(517) => 
                           DataPath_RF_bus_reg_dataout_517_port, regs(516) => 
                           DataPath_RF_bus_reg_dataout_516_port, regs(515) => 
                           DataPath_RF_bus_reg_dataout_515_port, regs(514) => 
                           DataPath_RF_bus_reg_dataout_514_port, regs(513) => 
                           DataPath_RF_bus_reg_dataout_513_port, regs(512) => 
                           DataPath_RF_bus_reg_dataout_512_port, regs(511) => 
                           DataPath_RF_bus_reg_dataout_511_port, regs(510) => 
                           DataPath_RF_bus_reg_dataout_510_port, regs(509) => 
                           DataPath_RF_bus_reg_dataout_509_port, regs(508) => 
                           DataPath_RF_bus_reg_dataout_508_port, regs(507) => 
                           DataPath_RF_bus_reg_dataout_507_port, regs(506) => 
                           DataPath_RF_bus_reg_dataout_506_port, regs(505) => 
                           DataPath_RF_bus_reg_dataout_505_port, regs(504) => 
                           DataPath_RF_bus_reg_dataout_504_port, regs(503) => 
                           DataPath_RF_bus_reg_dataout_503_port, regs(502) => 
                           DataPath_RF_bus_reg_dataout_502_port, regs(501) => 
                           DataPath_RF_bus_reg_dataout_501_port, regs(500) => 
                           DataPath_RF_bus_reg_dataout_500_port, regs(499) => 
                           DataPath_RF_bus_reg_dataout_499_port, regs(498) => 
                           DataPath_RF_bus_reg_dataout_498_port, regs(497) => 
                           DataPath_RF_bus_reg_dataout_497_port, regs(496) => 
                           DataPath_RF_bus_reg_dataout_496_port, regs(495) => 
                           DataPath_RF_bus_reg_dataout_495_port, regs(494) => 
                           DataPath_RF_bus_reg_dataout_494_port, regs(493) => 
                           DataPath_RF_bus_reg_dataout_493_port, regs(492) => 
                           DataPath_RF_bus_reg_dataout_492_port, regs(491) => 
                           DataPath_RF_bus_reg_dataout_491_port, regs(490) => 
                           DataPath_RF_bus_reg_dataout_490_port, regs(489) => 
                           DataPath_RF_bus_reg_dataout_489_port, regs(488) => 
                           DataPath_RF_bus_reg_dataout_488_port, regs(487) => 
                           DataPath_RF_bus_reg_dataout_487_port, regs(486) => 
                           DataPath_RF_bus_reg_dataout_486_port, regs(485) => 
                           DataPath_RF_bus_reg_dataout_485_port, regs(484) => 
                           DataPath_RF_bus_reg_dataout_484_port, regs(483) => 
                           DataPath_RF_bus_reg_dataout_483_port, regs(482) => 
                           DataPath_RF_bus_reg_dataout_482_port, regs(481) => 
                           DataPath_RF_bus_reg_dataout_481_port, regs(480) => 
                           DataPath_RF_bus_reg_dataout_480_port, regs(479) => 
                           DataPath_RF_bus_reg_dataout_479_port, regs(478) => 
                           DataPath_RF_bus_reg_dataout_478_port, regs(477) => 
                           DataPath_RF_bus_reg_dataout_477_port, regs(476) => 
                           DataPath_RF_bus_reg_dataout_476_port, regs(475) => 
                           DataPath_RF_bus_reg_dataout_475_port, regs(474) => 
                           DataPath_RF_bus_reg_dataout_474_port, regs(473) => 
                           DataPath_RF_bus_reg_dataout_473_port, regs(472) => 
                           DataPath_RF_bus_reg_dataout_472_port, regs(471) => 
                           DataPath_RF_bus_reg_dataout_471_port, regs(470) => 
                           DataPath_RF_bus_reg_dataout_470_port, regs(469) => 
                           DataPath_RF_bus_reg_dataout_469_port, regs(468) => 
                           DataPath_RF_bus_reg_dataout_468_port, regs(467) => 
                           DataPath_RF_bus_reg_dataout_467_port, regs(466) => 
                           DataPath_RF_bus_reg_dataout_466_port, regs(465) => 
                           DataPath_RF_bus_reg_dataout_465_port, regs(464) => 
                           DataPath_RF_bus_reg_dataout_464_port, regs(463) => 
                           DataPath_RF_bus_reg_dataout_463_port, regs(462) => 
                           DataPath_RF_bus_reg_dataout_462_port, regs(461) => 
                           DataPath_RF_bus_reg_dataout_461_port, regs(460) => 
                           DataPath_RF_bus_reg_dataout_460_port, regs(459) => 
                           DataPath_RF_bus_reg_dataout_459_port, regs(458) => 
                           DataPath_RF_bus_reg_dataout_458_port, regs(457) => 
                           DataPath_RF_bus_reg_dataout_457_port, regs(456) => 
                           DataPath_RF_bus_reg_dataout_456_port, regs(455) => 
                           DataPath_RF_bus_reg_dataout_455_port, regs(454) => 
                           DataPath_RF_bus_reg_dataout_454_port, regs(453) => 
                           DataPath_RF_bus_reg_dataout_453_port, regs(452) => 
                           DataPath_RF_bus_reg_dataout_452_port, regs(451) => 
                           DataPath_RF_bus_reg_dataout_451_port, regs(450) => 
                           DataPath_RF_bus_reg_dataout_450_port, regs(449) => 
                           DataPath_RF_bus_reg_dataout_449_port, regs(448) => 
                           DataPath_RF_bus_reg_dataout_448_port, regs(447) => 
                           DataPath_RF_bus_reg_dataout_447_port, regs(446) => 
                           DataPath_RF_bus_reg_dataout_446_port, regs(445) => 
                           DataPath_RF_bus_reg_dataout_445_port, regs(444) => 
                           DataPath_RF_bus_reg_dataout_444_port, regs(443) => 
                           DataPath_RF_bus_reg_dataout_443_port, regs(442) => 
                           DataPath_RF_bus_reg_dataout_442_port, regs(441) => 
                           DataPath_RF_bus_reg_dataout_441_port, regs(440) => 
                           DataPath_RF_bus_reg_dataout_440_port, regs(439) => 
                           DataPath_RF_bus_reg_dataout_439_port, regs(438) => 
                           DataPath_RF_bus_reg_dataout_438_port, regs(437) => 
                           DataPath_RF_bus_reg_dataout_437_port, regs(436) => 
                           DataPath_RF_bus_reg_dataout_436_port, regs(435) => 
                           DataPath_RF_bus_reg_dataout_435_port, regs(434) => 
                           DataPath_RF_bus_reg_dataout_434_port, regs(433) => 
                           DataPath_RF_bus_reg_dataout_433_port, regs(432) => 
                           DataPath_RF_bus_reg_dataout_432_port, regs(431) => 
                           DataPath_RF_bus_reg_dataout_431_port, regs(430) => 
                           DataPath_RF_bus_reg_dataout_430_port, regs(429) => 
                           DataPath_RF_bus_reg_dataout_429_port, regs(428) => 
                           DataPath_RF_bus_reg_dataout_428_port, regs(427) => 
                           DataPath_RF_bus_reg_dataout_427_port, regs(426) => 
                           DataPath_RF_bus_reg_dataout_426_port, regs(425) => 
                           DataPath_RF_bus_reg_dataout_425_port, regs(424) => 
                           DataPath_RF_bus_reg_dataout_424_port, regs(423) => 
                           DataPath_RF_bus_reg_dataout_423_port, regs(422) => 
                           DataPath_RF_bus_reg_dataout_422_port, regs(421) => 
                           DataPath_RF_bus_reg_dataout_421_port, regs(420) => 
                           DataPath_RF_bus_reg_dataout_420_port, regs(419) => 
                           DataPath_RF_bus_reg_dataout_419_port, regs(418) => 
                           DataPath_RF_bus_reg_dataout_418_port, regs(417) => 
                           DataPath_RF_bus_reg_dataout_417_port, regs(416) => 
                           DataPath_RF_bus_reg_dataout_416_port, regs(415) => 
                           DataPath_RF_bus_reg_dataout_415_port, regs(414) => 
                           DataPath_RF_bus_reg_dataout_414_port, regs(413) => 
                           DataPath_RF_bus_reg_dataout_413_port, regs(412) => 
                           DataPath_RF_bus_reg_dataout_412_port, regs(411) => 
                           DataPath_RF_bus_reg_dataout_411_port, regs(410) => 
                           DataPath_RF_bus_reg_dataout_410_port, regs(409) => 
                           DataPath_RF_bus_reg_dataout_409_port, regs(408) => 
                           DataPath_RF_bus_reg_dataout_408_port, regs(407) => 
                           DataPath_RF_bus_reg_dataout_407_port, regs(406) => 
                           DataPath_RF_bus_reg_dataout_406_port, regs(405) => 
                           DataPath_RF_bus_reg_dataout_405_port, regs(404) => 
                           DataPath_RF_bus_reg_dataout_404_port, regs(403) => 
                           DataPath_RF_bus_reg_dataout_403_port, regs(402) => 
                           DataPath_RF_bus_reg_dataout_402_port, regs(401) => 
                           DataPath_RF_bus_reg_dataout_401_port, regs(400) => 
                           DataPath_RF_bus_reg_dataout_400_port, regs(399) => 
                           DataPath_RF_bus_reg_dataout_399_port, regs(398) => 
                           DataPath_RF_bus_reg_dataout_398_port, regs(397) => 
                           DataPath_RF_bus_reg_dataout_397_port, regs(396) => 
                           DataPath_RF_bus_reg_dataout_396_port, regs(395) => 
                           DataPath_RF_bus_reg_dataout_395_port, regs(394) => 
                           DataPath_RF_bus_reg_dataout_394_port, regs(393) => 
                           DataPath_RF_bus_reg_dataout_393_port, regs(392) => 
                           DataPath_RF_bus_reg_dataout_392_port, regs(391) => 
                           DataPath_RF_bus_reg_dataout_391_port, regs(390) => 
                           DataPath_RF_bus_reg_dataout_390_port, regs(389) => 
                           DataPath_RF_bus_reg_dataout_389_port, regs(388) => 
                           DataPath_RF_bus_reg_dataout_388_port, regs(387) => 
                           DataPath_RF_bus_reg_dataout_387_port, regs(386) => 
                           DataPath_RF_bus_reg_dataout_386_port, regs(385) => 
                           DataPath_RF_bus_reg_dataout_385_port, regs(384) => 
                           DataPath_RF_bus_reg_dataout_384_port, regs(383) => 
                           DataPath_RF_bus_reg_dataout_383_port, regs(382) => 
                           DataPath_RF_bus_reg_dataout_382_port, regs(381) => 
                           DataPath_RF_bus_reg_dataout_381_port, regs(380) => 
                           DataPath_RF_bus_reg_dataout_380_port, regs(379) => 
                           DataPath_RF_bus_reg_dataout_379_port, regs(378) => 
                           DataPath_RF_bus_reg_dataout_378_port, regs(377) => 
                           DataPath_RF_bus_reg_dataout_377_port, regs(376) => 
                           DataPath_RF_bus_reg_dataout_376_port, regs(375) => 
                           DataPath_RF_bus_reg_dataout_375_port, regs(374) => 
                           DataPath_RF_bus_reg_dataout_374_port, regs(373) => 
                           DataPath_RF_bus_reg_dataout_373_port, regs(372) => 
                           DataPath_RF_bus_reg_dataout_372_port, regs(371) => 
                           DataPath_RF_bus_reg_dataout_371_port, regs(370) => 
                           DataPath_RF_bus_reg_dataout_370_port, regs(369) => 
                           DataPath_RF_bus_reg_dataout_369_port, regs(368) => 
                           DataPath_RF_bus_reg_dataout_368_port, regs(367) => 
                           DataPath_RF_bus_reg_dataout_367_port, regs(366) => 
                           DataPath_RF_bus_reg_dataout_366_port, regs(365) => 
                           DataPath_RF_bus_reg_dataout_365_port, regs(364) => 
                           DataPath_RF_bus_reg_dataout_364_port, regs(363) => 
                           DataPath_RF_bus_reg_dataout_363_port, regs(362) => 
                           DataPath_RF_bus_reg_dataout_362_port, regs(361) => 
                           DataPath_RF_bus_reg_dataout_361_port, regs(360) => 
                           DataPath_RF_bus_reg_dataout_360_port, regs(359) => 
                           DataPath_RF_bus_reg_dataout_359_port, regs(358) => 
                           DataPath_RF_bus_reg_dataout_358_port, regs(357) => 
                           DataPath_RF_bus_reg_dataout_357_port, regs(356) => 
                           DataPath_RF_bus_reg_dataout_356_port, regs(355) => 
                           DataPath_RF_bus_reg_dataout_355_port, regs(354) => 
                           DataPath_RF_bus_reg_dataout_354_port, regs(353) => 
                           DataPath_RF_bus_reg_dataout_353_port, regs(352) => 
                           DataPath_RF_bus_reg_dataout_352_port, regs(351) => 
                           DataPath_RF_bus_reg_dataout_351_port, regs(350) => 
                           DataPath_RF_bus_reg_dataout_350_port, regs(349) => 
                           DataPath_RF_bus_reg_dataout_349_port, regs(348) => 
                           DataPath_RF_bus_reg_dataout_348_port, regs(347) => 
                           DataPath_RF_bus_reg_dataout_347_port, regs(346) => 
                           DataPath_RF_bus_reg_dataout_346_port, regs(345) => 
                           DataPath_RF_bus_reg_dataout_345_port, regs(344) => 
                           DataPath_RF_bus_reg_dataout_344_port, regs(343) => 
                           DataPath_RF_bus_reg_dataout_343_port, regs(342) => 
                           DataPath_RF_bus_reg_dataout_342_port, regs(341) => 
                           DataPath_RF_bus_reg_dataout_341_port, regs(340) => 
                           DataPath_RF_bus_reg_dataout_340_port, regs(339) => 
                           DataPath_RF_bus_reg_dataout_339_port, regs(338) => 
                           DataPath_RF_bus_reg_dataout_338_port, regs(337) => 
                           DataPath_RF_bus_reg_dataout_337_port, regs(336) => 
                           DataPath_RF_bus_reg_dataout_336_port, regs(335) => 
                           DataPath_RF_bus_reg_dataout_335_port, regs(334) => 
                           DataPath_RF_bus_reg_dataout_334_port, regs(333) => 
                           DataPath_RF_bus_reg_dataout_333_port, regs(332) => 
                           DataPath_RF_bus_reg_dataout_332_port, regs(331) => 
                           DataPath_RF_bus_reg_dataout_331_port, regs(330) => 
                           DataPath_RF_bus_reg_dataout_330_port, regs(329) => 
                           DataPath_RF_bus_reg_dataout_329_port, regs(328) => 
                           DataPath_RF_bus_reg_dataout_328_port, regs(327) => 
                           DataPath_RF_bus_reg_dataout_327_port, regs(326) => 
                           DataPath_RF_bus_reg_dataout_326_port, regs(325) => 
                           DataPath_RF_bus_reg_dataout_325_port, regs(324) => 
                           DataPath_RF_bus_reg_dataout_324_port, regs(323) => 
                           DataPath_RF_bus_reg_dataout_323_port, regs(322) => 
                           DataPath_RF_bus_reg_dataout_322_port, regs(321) => 
                           DataPath_RF_bus_reg_dataout_321_port, regs(320) => 
                           DataPath_RF_bus_reg_dataout_320_port, regs(319) => 
                           DataPath_RF_bus_reg_dataout_319_port, regs(318) => 
                           DataPath_RF_bus_reg_dataout_318_port, regs(317) => 
                           DataPath_RF_bus_reg_dataout_317_port, regs(316) => 
                           DataPath_RF_bus_reg_dataout_316_port, regs(315) => 
                           DataPath_RF_bus_reg_dataout_315_port, regs(314) => 
                           DataPath_RF_bus_reg_dataout_314_port, regs(313) => 
                           DataPath_RF_bus_reg_dataout_313_port, regs(312) => 
                           DataPath_RF_bus_reg_dataout_312_port, regs(311) => 
                           DataPath_RF_bus_reg_dataout_311_port, regs(310) => 
                           DataPath_RF_bus_reg_dataout_310_port, regs(309) => 
                           DataPath_RF_bus_reg_dataout_309_port, regs(308) => 
                           DataPath_RF_bus_reg_dataout_308_port, regs(307) => 
                           DataPath_RF_bus_reg_dataout_307_port, regs(306) => 
                           DataPath_RF_bus_reg_dataout_306_port, regs(305) => 
                           DataPath_RF_bus_reg_dataout_305_port, regs(304) => 
                           DataPath_RF_bus_reg_dataout_304_port, regs(303) => 
                           DataPath_RF_bus_reg_dataout_303_port, regs(302) => 
                           DataPath_RF_bus_reg_dataout_302_port, regs(301) => 
                           DataPath_RF_bus_reg_dataout_301_port, regs(300) => 
                           DataPath_RF_bus_reg_dataout_300_port, regs(299) => 
                           DataPath_RF_bus_reg_dataout_299_port, regs(298) => 
                           DataPath_RF_bus_reg_dataout_298_port, regs(297) => 
                           DataPath_RF_bus_reg_dataout_297_port, regs(296) => 
                           DataPath_RF_bus_reg_dataout_296_port, regs(295) => 
                           DataPath_RF_bus_reg_dataout_295_port, regs(294) => 
                           DataPath_RF_bus_reg_dataout_294_port, regs(293) => 
                           DataPath_RF_bus_reg_dataout_293_port, regs(292) => 
                           DataPath_RF_bus_reg_dataout_292_port, regs(291) => 
                           DataPath_RF_bus_reg_dataout_291_port, regs(290) => 
                           DataPath_RF_bus_reg_dataout_290_port, regs(289) => 
                           DataPath_RF_bus_reg_dataout_289_port, regs(288) => 
                           DataPath_RF_bus_reg_dataout_288_port, regs(287) => 
                           DataPath_RF_bus_reg_dataout_287_port, regs(286) => 
                           DataPath_RF_bus_reg_dataout_286_port, regs(285) => 
                           DataPath_RF_bus_reg_dataout_285_port, regs(284) => 
                           DataPath_RF_bus_reg_dataout_284_port, regs(283) => 
                           DataPath_RF_bus_reg_dataout_283_port, regs(282) => 
                           DataPath_RF_bus_reg_dataout_282_port, regs(281) => 
                           DataPath_RF_bus_reg_dataout_281_port, regs(280) => 
                           DataPath_RF_bus_reg_dataout_280_port, regs(279) => 
                           DataPath_RF_bus_reg_dataout_279_port, regs(278) => 
                           DataPath_RF_bus_reg_dataout_278_port, regs(277) => 
                           DataPath_RF_bus_reg_dataout_277_port, regs(276) => 
                           DataPath_RF_bus_reg_dataout_276_port, regs(275) => 
                           DataPath_RF_bus_reg_dataout_275_port, regs(274) => 
                           DataPath_RF_bus_reg_dataout_274_port, regs(273) => 
                           DataPath_RF_bus_reg_dataout_273_port, regs(272) => 
                           DataPath_RF_bus_reg_dataout_272_port, regs(271) => 
                           DataPath_RF_bus_reg_dataout_271_port, regs(270) => 
                           DataPath_RF_bus_reg_dataout_270_port, regs(269) => 
                           DataPath_RF_bus_reg_dataout_269_port, regs(268) => 
                           DataPath_RF_bus_reg_dataout_268_port, regs(267) => 
                           DataPath_RF_bus_reg_dataout_267_port, regs(266) => 
                           DataPath_RF_bus_reg_dataout_266_port, regs(265) => 
                           DataPath_RF_bus_reg_dataout_265_port, regs(264) => 
                           DataPath_RF_bus_reg_dataout_264_port, regs(263) => 
                           DataPath_RF_bus_reg_dataout_263_port, regs(262) => 
                           DataPath_RF_bus_reg_dataout_262_port, regs(261) => 
                           DataPath_RF_bus_reg_dataout_261_port, regs(260) => 
                           DataPath_RF_bus_reg_dataout_260_port, regs(259) => 
                           DataPath_RF_bus_reg_dataout_259_port, regs(258) => 
                           DataPath_RF_bus_reg_dataout_258_port, regs(257) => 
                           DataPath_RF_bus_reg_dataout_257_port, regs(256) => 
                           DataPath_RF_bus_reg_dataout_256_port, regs(255) => 
                           DataPath_RF_bus_reg_dataout_255_port, regs(254) => 
                           DataPath_RF_bus_reg_dataout_254_port, regs(253) => 
                           DataPath_RF_bus_reg_dataout_253_port, regs(252) => 
                           DataPath_RF_bus_reg_dataout_252_port, regs(251) => 
                           DataPath_RF_bus_reg_dataout_251_port, regs(250) => 
                           DataPath_RF_bus_reg_dataout_250_port, regs(249) => 
                           DataPath_RF_bus_reg_dataout_249_port, regs(248) => 
                           DataPath_RF_bus_reg_dataout_248_port, regs(247) => 
                           DataPath_RF_bus_reg_dataout_247_port, regs(246) => 
                           DataPath_RF_bus_reg_dataout_246_port, regs(245) => 
                           DataPath_RF_bus_reg_dataout_245_port, regs(244) => 
                           DataPath_RF_bus_reg_dataout_244_port, regs(243) => 
                           DataPath_RF_bus_reg_dataout_243_port, regs(242) => 
                           DataPath_RF_bus_reg_dataout_242_port, regs(241) => 
                           DataPath_RF_bus_reg_dataout_241_port, regs(240) => 
                           DataPath_RF_bus_reg_dataout_240_port, regs(239) => 
                           DataPath_RF_bus_reg_dataout_239_port, regs(238) => 
                           DataPath_RF_bus_reg_dataout_238_port, regs(237) => 
                           DataPath_RF_bus_reg_dataout_237_port, regs(236) => 
                           DataPath_RF_bus_reg_dataout_236_port, regs(235) => 
                           DataPath_RF_bus_reg_dataout_235_port, regs(234) => 
                           DataPath_RF_bus_reg_dataout_234_port, regs(233) => 
                           DataPath_RF_bus_reg_dataout_233_port, regs(232) => 
                           DataPath_RF_bus_reg_dataout_232_port, regs(231) => 
                           DataPath_RF_bus_reg_dataout_231_port, regs(230) => 
                           DataPath_RF_bus_reg_dataout_230_port, regs(229) => 
                           DataPath_RF_bus_reg_dataout_229_port, regs(228) => 
                           DataPath_RF_bus_reg_dataout_228_port, regs(227) => 
                           DataPath_RF_bus_reg_dataout_227_port, regs(226) => 
                           DataPath_RF_bus_reg_dataout_226_port, regs(225) => 
                           DataPath_RF_bus_reg_dataout_225_port, regs(224) => 
                           DataPath_RF_bus_reg_dataout_224_port, regs(223) => 
                           DataPath_RF_bus_reg_dataout_223_port, regs(222) => 
                           DataPath_RF_bus_reg_dataout_222_port, regs(221) => 
                           DataPath_RF_bus_reg_dataout_221_port, regs(220) => 
                           DataPath_RF_bus_reg_dataout_220_port, regs(219) => 
                           DataPath_RF_bus_reg_dataout_219_port, regs(218) => 
                           DataPath_RF_bus_reg_dataout_218_port, regs(217) => 
                           DataPath_RF_bus_reg_dataout_217_port, regs(216) => 
                           DataPath_RF_bus_reg_dataout_216_port, regs(215) => 
                           DataPath_RF_bus_reg_dataout_215_port, regs(214) => 
                           DataPath_RF_bus_reg_dataout_214_port, regs(213) => 
                           DataPath_RF_bus_reg_dataout_213_port, regs(212) => 
                           DataPath_RF_bus_reg_dataout_212_port, regs(211) => 
                           DataPath_RF_bus_reg_dataout_211_port, regs(210) => 
                           DataPath_RF_bus_reg_dataout_210_port, regs(209) => 
                           DataPath_RF_bus_reg_dataout_209_port, regs(208) => 
                           DataPath_RF_bus_reg_dataout_208_port, regs(207) => 
                           DataPath_RF_bus_reg_dataout_207_port, regs(206) => 
                           DataPath_RF_bus_reg_dataout_206_port, regs(205) => 
                           DataPath_RF_bus_reg_dataout_205_port, regs(204) => 
                           DataPath_RF_bus_reg_dataout_204_port, regs(203) => 
                           DataPath_RF_bus_reg_dataout_203_port, regs(202) => 
                           DataPath_RF_bus_reg_dataout_202_port, regs(201) => 
                           DataPath_RF_bus_reg_dataout_201_port, regs(200) => 
                           DataPath_RF_bus_reg_dataout_200_port, regs(199) => 
                           DataPath_RF_bus_reg_dataout_199_port, regs(198) => 
                           DataPath_RF_bus_reg_dataout_198_port, regs(197) => 
                           DataPath_RF_bus_reg_dataout_197_port, regs(196) => 
                           DataPath_RF_bus_reg_dataout_196_port, regs(195) => 
                           DataPath_RF_bus_reg_dataout_195_port, regs(194) => 
                           DataPath_RF_bus_reg_dataout_194_port, regs(193) => 
                           DataPath_RF_bus_reg_dataout_193_port, regs(192) => 
                           DataPath_RF_bus_reg_dataout_192_port, regs(191) => 
                           DataPath_RF_bus_reg_dataout_191_port, regs(190) => 
                           DataPath_RF_bus_reg_dataout_190_port, regs(189) => 
                           DataPath_RF_bus_reg_dataout_189_port, regs(188) => 
                           DataPath_RF_bus_reg_dataout_188_port, regs(187) => 
                           DataPath_RF_bus_reg_dataout_187_port, regs(186) => 
                           DataPath_RF_bus_reg_dataout_186_port, regs(185) => 
                           DataPath_RF_bus_reg_dataout_185_port, regs(184) => 
                           DataPath_RF_bus_reg_dataout_184_port, regs(183) => 
                           DataPath_RF_bus_reg_dataout_183_port, regs(182) => 
                           DataPath_RF_bus_reg_dataout_182_port, regs(181) => 
                           DataPath_RF_bus_reg_dataout_181_port, regs(180) => 
                           DataPath_RF_bus_reg_dataout_180_port, regs(179) => 
                           DataPath_RF_bus_reg_dataout_179_port, regs(178) => 
                           DataPath_RF_bus_reg_dataout_178_port, regs(177) => 
                           DataPath_RF_bus_reg_dataout_177_port, regs(176) => 
                           DataPath_RF_bus_reg_dataout_176_port, regs(175) => 
                           DataPath_RF_bus_reg_dataout_175_port, regs(174) => 
                           DataPath_RF_bus_reg_dataout_174_port, regs(173) => 
                           DataPath_RF_bus_reg_dataout_173_port, regs(172) => 
                           DataPath_RF_bus_reg_dataout_172_port, regs(171) => 
                           DataPath_RF_bus_reg_dataout_171_port, regs(170) => 
                           DataPath_RF_bus_reg_dataout_170_port, regs(169) => 
                           DataPath_RF_bus_reg_dataout_169_port, regs(168) => 
                           DataPath_RF_bus_reg_dataout_168_port, regs(167) => 
                           DataPath_RF_bus_reg_dataout_167_port, regs(166) => 
                           DataPath_RF_bus_reg_dataout_166_port, regs(165) => 
                           DataPath_RF_bus_reg_dataout_165_port, regs(164) => 
                           DataPath_RF_bus_reg_dataout_164_port, regs(163) => 
                           DataPath_RF_bus_reg_dataout_163_port, regs(162) => 
                           DataPath_RF_bus_reg_dataout_162_port, regs(161) => 
                           DataPath_RF_bus_reg_dataout_161_port, regs(160) => 
                           DataPath_RF_bus_reg_dataout_160_port, regs(159) => 
                           DataPath_RF_bus_reg_dataout_159_port, regs(158) => 
                           DataPath_RF_bus_reg_dataout_158_port, regs(157) => 
                           DataPath_RF_bus_reg_dataout_157_port, regs(156) => 
                           DataPath_RF_bus_reg_dataout_156_port, regs(155) => 
                           DataPath_RF_bus_reg_dataout_155_port, regs(154) => 
                           DataPath_RF_bus_reg_dataout_154_port, regs(153) => 
                           DataPath_RF_bus_reg_dataout_153_port, regs(152) => 
                           DataPath_RF_bus_reg_dataout_152_port, regs(151) => 
                           DataPath_RF_bus_reg_dataout_151_port, regs(150) => 
                           DataPath_RF_bus_reg_dataout_150_port, regs(149) => 
                           DataPath_RF_bus_reg_dataout_149_port, regs(148) => 
                           DataPath_RF_bus_reg_dataout_148_port, regs(147) => 
                           DataPath_RF_bus_reg_dataout_147_port, regs(146) => 
                           DataPath_RF_bus_reg_dataout_146_port, regs(145) => 
                           DataPath_RF_bus_reg_dataout_145_port, regs(144) => 
                           DataPath_RF_bus_reg_dataout_144_port, regs(143) => 
                           DataPath_RF_bus_reg_dataout_143_port, regs(142) => 
                           DataPath_RF_bus_reg_dataout_142_port, regs(141) => 
                           DataPath_RF_bus_reg_dataout_141_port, regs(140) => 
                           DataPath_RF_bus_reg_dataout_140_port, regs(139) => 
                           DataPath_RF_bus_reg_dataout_139_port, regs(138) => 
                           DataPath_RF_bus_reg_dataout_138_port, regs(137) => 
                           DataPath_RF_bus_reg_dataout_137_port, regs(136) => 
                           DataPath_RF_bus_reg_dataout_136_port, regs(135) => 
                           DataPath_RF_bus_reg_dataout_135_port, regs(134) => 
                           DataPath_RF_bus_reg_dataout_134_port, regs(133) => 
                           DataPath_RF_bus_reg_dataout_133_port, regs(132) => 
                           DataPath_RF_bus_reg_dataout_132_port, regs(131) => 
                           DataPath_RF_bus_reg_dataout_131_port, regs(130) => 
                           DataPath_RF_bus_reg_dataout_130_port, regs(129) => 
                           DataPath_RF_bus_reg_dataout_129_port, regs(128) => 
                           DataPath_RF_bus_reg_dataout_128_port, regs(127) => 
                           DataPath_RF_bus_reg_dataout_127_port, regs(126) => 
                           DataPath_RF_bus_reg_dataout_126_port, regs(125) => 
                           DataPath_RF_bus_reg_dataout_125_port, regs(124) => 
                           DataPath_RF_bus_reg_dataout_124_port, regs(123) => 
                           DataPath_RF_bus_reg_dataout_123_port, regs(122) => 
                           DataPath_RF_bus_reg_dataout_122_port, regs(121) => 
                           DataPath_RF_bus_reg_dataout_121_port, regs(120) => 
                           DataPath_RF_bus_reg_dataout_120_port, regs(119) => 
                           DataPath_RF_bus_reg_dataout_119_port, regs(118) => 
                           DataPath_RF_bus_reg_dataout_118_port, regs(117) => 
                           DataPath_RF_bus_reg_dataout_117_port, regs(116) => 
                           DataPath_RF_bus_reg_dataout_116_port, regs(115) => 
                           DataPath_RF_bus_reg_dataout_115_port, regs(114) => 
                           DataPath_RF_bus_reg_dataout_114_port, regs(113) => 
                           DataPath_RF_bus_reg_dataout_113_port, regs(112) => 
                           DataPath_RF_bus_reg_dataout_112_port, regs(111) => 
                           DataPath_RF_bus_reg_dataout_111_port, regs(110) => 
                           DataPath_RF_bus_reg_dataout_110_port, regs(109) => 
                           DataPath_RF_bus_reg_dataout_109_port, regs(108) => 
                           DataPath_RF_bus_reg_dataout_108_port, regs(107) => 
                           DataPath_RF_bus_reg_dataout_107_port, regs(106) => 
                           DataPath_RF_bus_reg_dataout_106_port, regs(105) => 
                           DataPath_RF_bus_reg_dataout_105_port, regs(104) => 
                           DataPath_RF_bus_reg_dataout_104_port, regs(103) => 
                           DataPath_RF_bus_reg_dataout_103_port, regs(102) => 
                           DataPath_RF_bus_reg_dataout_102_port, regs(101) => 
                           DataPath_RF_bus_reg_dataout_101_port, regs(100) => 
                           DataPath_RF_bus_reg_dataout_100_port, regs(99) => 
                           DataPath_RF_bus_reg_dataout_99_port, regs(98) => 
                           DataPath_RF_bus_reg_dataout_98_port, regs(97) => 
                           DataPath_RF_bus_reg_dataout_97_port, regs(96) => 
                           DataPath_RF_bus_reg_dataout_96_port, regs(95) => 
                           DataPath_RF_bus_reg_dataout_95_port, regs(94) => 
                           DataPath_RF_bus_reg_dataout_94_port, regs(93) => 
                           DataPath_RF_bus_reg_dataout_93_port, regs(92) => 
                           DataPath_RF_bus_reg_dataout_92_port, regs(91) => 
                           DataPath_RF_bus_reg_dataout_91_port, regs(90) => 
                           DataPath_RF_bus_reg_dataout_90_port, regs(89) => 
                           DataPath_RF_bus_reg_dataout_89_port, regs(88) => 
                           DataPath_RF_bus_reg_dataout_88_port, regs(87) => 
                           DataPath_RF_bus_reg_dataout_87_port, regs(86) => 
                           DataPath_RF_bus_reg_dataout_86_port, regs(85) => 
                           DataPath_RF_bus_reg_dataout_85_port, regs(84) => 
                           DataPath_RF_bus_reg_dataout_84_port, regs(83) => 
                           DataPath_RF_bus_reg_dataout_83_port, regs(82) => 
                           DataPath_RF_bus_reg_dataout_82_port, regs(81) => 
                           DataPath_RF_bus_reg_dataout_81_port, regs(80) => 
                           DataPath_RF_bus_reg_dataout_80_port, regs(79) => 
                           DataPath_RF_bus_reg_dataout_79_port, regs(78) => 
                           DataPath_RF_bus_reg_dataout_78_port, regs(77) => 
                           DataPath_RF_bus_reg_dataout_77_port, regs(76) => 
                           DataPath_RF_bus_reg_dataout_76_port, regs(75) => 
                           DataPath_RF_bus_reg_dataout_75_port, regs(74) => 
                           DataPath_RF_bus_reg_dataout_74_port, regs(73) => 
                           DataPath_RF_bus_reg_dataout_73_port, regs(72) => 
                           DataPath_RF_bus_reg_dataout_72_port, regs(71) => 
                           DataPath_RF_bus_reg_dataout_71_port, regs(70) => 
                           DataPath_RF_bus_reg_dataout_70_port, regs(69) => 
                           DataPath_RF_bus_reg_dataout_69_port, regs(68) => 
                           DataPath_RF_bus_reg_dataout_68_port, regs(67) => 
                           DataPath_RF_bus_reg_dataout_67_port, regs(66) => 
                           DataPath_RF_bus_reg_dataout_66_port, regs(65) => 
                           DataPath_RF_bus_reg_dataout_65_port, regs(64) => 
                           DataPath_RF_bus_reg_dataout_64_port, regs(63) => 
                           DataPath_RF_bus_reg_dataout_63_port, regs(62) => 
                           DataPath_RF_bus_reg_dataout_62_port, regs(61) => 
                           DataPath_RF_bus_reg_dataout_61_port, regs(60) => 
                           DataPath_RF_bus_reg_dataout_60_port, regs(59) => 
                           DataPath_RF_bus_reg_dataout_59_port, regs(58) => 
                           DataPath_RF_bus_reg_dataout_58_port, regs(57) => 
                           DataPath_RF_bus_reg_dataout_57_port, regs(56) => 
                           DataPath_RF_bus_reg_dataout_56_port, regs(55) => 
                           DataPath_RF_bus_reg_dataout_55_port, regs(54) => 
                           DataPath_RF_bus_reg_dataout_54_port, regs(53) => 
                           DataPath_RF_bus_reg_dataout_53_port, regs(52) => 
                           DataPath_RF_bus_reg_dataout_52_port, regs(51) => 
                           DataPath_RF_bus_reg_dataout_51_port, regs(50) => 
                           DataPath_RF_bus_reg_dataout_50_port, regs(49) => 
                           DataPath_RF_bus_reg_dataout_49_port, regs(48) => 
                           DataPath_RF_bus_reg_dataout_48_port, regs(47) => 
                           DataPath_RF_bus_reg_dataout_47_port, regs(46) => 
                           DataPath_RF_bus_reg_dataout_46_port, regs(45) => 
                           DataPath_RF_bus_reg_dataout_45_port, regs(44) => 
                           DataPath_RF_bus_reg_dataout_44_port, regs(43) => 
                           DataPath_RF_bus_reg_dataout_43_port, regs(42) => 
                           DataPath_RF_bus_reg_dataout_42_port, regs(41) => 
                           DataPath_RF_bus_reg_dataout_41_port, regs(40) => 
                           DataPath_RF_bus_reg_dataout_40_port, regs(39) => 
                           DataPath_RF_bus_reg_dataout_39_port, regs(38) => 
                           DataPath_RF_bus_reg_dataout_38_port, regs(37) => 
                           DataPath_RF_bus_reg_dataout_37_port, regs(36) => 
                           DataPath_RF_bus_reg_dataout_36_port, regs(35) => 
                           DataPath_RF_bus_reg_dataout_35_port, regs(34) => 
                           DataPath_RF_bus_reg_dataout_34_port, regs(33) => 
                           DataPath_RF_bus_reg_dataout_33_port, regs(32) => 
                           DataPath_RF_bus_reg_dataout_32_port, regs(31) => 
                           DataPath_RF_bus_reg_dataout_31_port, regs(30) => 
                           DataPath_RF_bus_reg_dataout_30_port, regs(29) => 
                           DataPath_RF_bus_reg_dataout_29_port, regs(28) => 
                           DataPath_RF_bus_reg_dataout_28_port, regs(27) => 
                           DataPath_RF_bus_reg_dataout_27_port, regs(26) => 
                           DataPath_RF_bus_reg_dataout_26_port, regs(25) => 
                           DataPath_RF_bus_reg_dataout_25_port, regs(24) => 
                           DataPath_RF_bus_reg_dataout_24_port, regs(23) => 
                           DataPath_RF_bus_reg_dataout_23_port, regs(22) => 
                           DataPath_RF_bus_reg_dataout_22_port, regs(21) => 
                           DataPath_RF_bus_reg_dataout_21_port, regs(20) => 
                           DataPath_RF_bus_reg_dataout_20_port, regs(19) => 
                           DataPath_RF_bus_reg_dataout_19_port, regs(18) => 
                           DataPath_RF_bus_reg_dataout_18_port, regs(17) => 
                           DataPath_RF_bus_reg_dataout_17_port, regs(16) => 
                           DataPath_RF_bus_reg_dataout_16_port, regs(15) => 
                           DataPath_RF_bus_reg_dataout_15_port, regs(14) => 
                           DataPath_RF_bus_reg_dataout_14_port, regs(13) => 
                           DataPath_RF_bus_reg_dataout_13_port, regs(12) => 
                           DataPath_RF_bus_reg_dataout_12_port, regs(11) => 
                           DataPath_RF_bus_reg_dataout_11_port, regs(10) => 
                           DataPath_RF_bus_reg_dataout_10_port, regs(9) => 
                           DataPath_RF_bus_reg_dataout_9_port, regs(8) => 
                           DataPath_RF_bus_reg_dataout_8_port, regs(7) => 
                           DataPath_RF_bus_reg_dataout_7_port, regs(6) => 
                           DataPath_RF_bus_reg_dataout_6_port, regs(5) => 
                           DataPath_RF_bus_reg_dataout_5_port, regs(4) => 
                           DataPath_RF_bus_reg_dataout_4_port, regs(3) => 
                           DataPath_RF_bus_reg_dataout_3_port, regs(2) => 
                           DataPath_RF_bus_reg_dataout_2_port, regs(1) => 
                           DataPath_RF_bus_reg_dataout_1_port, regs(0) => 
                           DataPath_RF_bus_reg_dataout_0_port, win(4) => n8564,
                           win(3) => n11814, win(2) => n8554, win(1) => 
                           DataPath_RF_c_win_1_port, win(0) => 
                           DataPath_RF_c_win_0_port, curr_proc_regs(767) => 
                           DataPath_RF_bus_selected_win_data_767_port, 
                           curr_proc_regs(766) => 
                           DataPath_RF_bus_selected_win_data_766_port, 
                           curr_proc_regs(765) => 
                           DataPath_RF_bus_selected_win_data_765_port, 
                           curr_proc_regs(764) => 
                           DataPath_RF_bus_selected_win_data_764_port, 
                           curr_proc_regs(763) => 
                           DataPath_RF_bus_selected_win_data_763_port, 
                           curr_proc_regs(762) => 
                           DataPath_RF_bus_selected_win_data_762_port, 
                           curr_proc_regs(761) => 
                           DataPath_RF_bus_selected_win_data_761_port, 
                           curr_proc_regs(760) => 
                           DataPath_RF_bus_selected_win_data_760_port, 
                           curr_proc_regs(759) => 
                           DataPath_RF_bus_selected_win_data_759_port, 
                           curr_proc_regs(758) => 
                           DataPath_RF_bus_selected_win_data_758_port, 
                           curr_proc_regs(757) => 
                           DataPath_RF_bus_selected_win_data_757_port, 
                           curr_proc_regs(756) => 
                           DataPath_RF_bus_selected_win_data_756_port, 
                           curr_proc_regs(755) => 
                           DataPath_RF_bus_selected_win_data_755_port, 
                           curr_proc_regs(754) => 
                           DataPath_RF_bus_selected_win_data_754_port, 
                           curr_proc_regs(753) => 
                           DataPath_RF_bus_selected_win_data_753_port, 
                           curr_proc_regs(752) => 
                           DataPath_RF_bus_selected_win_data_752_port, 
                           curr_proc_regs(751) => 
                           DataPath_RF_bus_selected_win_data_751_port, 
                           curr_proc_regs(750) => 
                           DataPath_RF_bus_selected_win_data_750_port, 
                           curr_proc_regs(749) => 
                           DataPath_RF_bus_selected_win_data_749_port, 
                           curr_proc_regs(748) => 
                           DataPath_RF_bus_selected_win_data_748_port, 
                           curr_proc_regs(747) => 
                           DataPath_RF_bus_selected_win_data_747_port, 
                           curr_proc_regs(746) => 
                           DataPath_RF_bus_selected_win_data_746_port, 
                           curr_proc_regs(745) => 
                           DataPath_RF_bus_selected_win_data_745_port, 
                           curr_proc_regs(744) => 
                           DataPath_RF_bus_selected_win_data_744_port, 
                           curr_proc_regs(743) => 
                           DataPath_RF_bus_selected_win_data_743_port, 
                           curr_proc_regs(742) => 
                           DataPath_RF_bus_selected_win_data_742_port, 
                           curr_proc_regs(741) => 
                           DataPath_RF_bus_selected_win_data_741_port, 
                           curr_proc_regs(740) => 
                           DataPath_RF_bus_selected_win_data_740_port, 
                           curr_proc_regs(739) => 
                           DataPath_RF_bus_selected_win_data_739_port, 
                           curr_proc_regs(738) => 
                           DataPath_RF_bus_selected_win_data_738_port, 
                           curr_proc_regs(737) => 
                           DataPath_RF_bus_selected_win_data_737_port, 
                           curr_proc_regs(736) => 
                           DataPath_RF_bus_selected_win_data_736_port, 
                           curr_proc_regs(735) => 
                           DataPath_RF_bus_selected_win_data_735_port, 
                           curr_proc_regs(734) => 
                           DataPath_RF_bus_selected_win_data_734_port, 
                           curr_proc_regs(733) => 
                           DataPath_RF_bus_selected_win_data_733_port, 
                           curr_proc_regs(732) => 
                           DataPath_RF_bus_selected_win_data_732_port, 
                           curr_proc_regs(731) => 
                           DataPath_RF_bus_selected_win_data_731_port, 
                           curr_proc_regs(730) => 
                           DataPath_RF_bus_selected_win_data_730_port, 
                           curr_proc_regs(729) => 
                           DataPath_RF_bus_selected_win_data_729_port, 
                           curr_proc_regs(728) => 
                           DataPath_RF_bus_selected_win_data_728_port, 
                           curr_proc_regs(727) => 
                           DataPath_RF_bus_selected_win_data_727_port, 
                           curr_proc_regs(726) => 
                           DataPath_RF_bus_selected_win_data_726_port, 
                           curr_proc_regs(725) => 
                           DataPath_RF_bus_selected_win_data_725_port, 
                           curr_proc_regs(724) => 
                           DataPath_RF_bus_selected_win_data_724_port, 
                           curr_proc_regs(723) => 
                           DataPath_RF_bus_selected_win_data_723_port, 
                           curr_proc_regs(722) => 
                           DataPath_RF_bus_selected_win_data_722_port, 
                           curr_proc_regs(721) => 
                           DataPath_RF_bus_selected_win_data_721_port, 
                           curr_proc_regs(720) => 
                           DataPath_RF_bus_selected_win_data_720_port, 
                           curr_proc_regs(719) => 
                           DataPath_RF_bus_selected_win_data_719_port, 
                           curr_proc_regs(718) => 
                           DataPath_RF_bus_selected_win_data_718_port, 
                           curr_proc_regs(717) => 
                           DataPath_RF_bus_selected_win_data_717_port, 
                           curr_proc_regs(716) => 
                           DataPath_RF_bus_selected_win_data_716_port, 
                           curr_proc_regs(715) => 
                           DataPath_RF_bus_selected_win_data_715_port, 
                           curr_proc_regs(714) => 
                           DataPath_RF_bus_selected_win_data_714_port, 
                           curr_proc_regs(713) => 
                           DataPath_RF_bus_selected_win_data_713_port, 
                           curr_proc_regs(712) => 
                           DataPath_RF_bus_selected_win_data_712_port, 
                           curr_proc_regs(711) => 
                           DataPath_RF_bus_selected_win_data_711_port, 
                           curr_proc_regs(710) => 
                           DataPath_RF_bus_selected_win_data_710_port, 
                           curr_proc_regs(709) => 
                           DataPath_RF_bus_selected_win_data_709_port, 
                           curr_proc_regs(708) => 
                           DataPath_RF_bus_selected_win_data_708_port, 
                           curr_proc_regs(707) => 
                           DataPath_RF_bus_selected_win_data_707_port, 
                           curr_proc_regs(706) => 
                           DataPath_RF_bus_selected_win_data_706_port, 
                           curr_proc_regs(705) => 
                           DataPath_RF_bus_selected_win_data_705_port, 
                           curr_proc_regs(704) => 
                           DataPath_RF_bus_selected_win_data_704_port, 
                           curr_proc_regs(703) => 
                           DataPath_RF_bus_selected_win_data_703_port, 
                           curr_proc_regs(702) => 
                           DataPath_RF_bus_selected_win_data_702_port, 
                           curr_proc_regs(701) => 
                           DataPath_RF_bus_selected_win_data_701_port, 
                           curr_proc_regs(700) => 
                           DataPath_RF_bus_selected_win_data_700_port, 
                           curr_proc_regs(699) => 
                           DataPath_RF_bus_selected_win_data_699_port, 
                           curr_proc_regs(698) => 
                           DataPath_RF_bus_selected_win_data_698_port, 
                           curr_proc_regs(697) => 
                           DataPath_RF_bus_selected_win_data_697_port, 
                           curr_proc_regs(696) => 
                           DataPath_RF_bus_selected_win_data_696_port, 
                           curr_proc_regs(695) => 
                           DataPath_RF_bus_selected_win_data_695_port, 
                           curr_proc_regs(694) => 
                           DataPath_RF_bus_selected_win_data_694_port, 
                           curr_proc_regs(693) => 
                           DataPath_RF_bus_selected_win_data_693_port, 
                           curr_proc_regs(692) => 
                           DataPath_RF_bus_selected_win_data_692_port, 
                           curr_proc_regs(691) => 
                           DataPath_RF_bus_selected_win_data_691_port, 
                           curr_proc_regs(690) => 
                           DataPath_RF_bus_selected_win_data_690_port, 
                           curr_proc_regs(689) => 
                           DataPath_RF_bus_selected_win_data_689_port, 
                           curr_proc_regs(688) => 
                           DataPath_RF_bus_selected_win_data_688_port, 
                           curr_proc_regs(687) => 
                           DataPath_RF_bus_selected_win_data_687_port, 
                           curr_proc_regs(686) => 
                           DataPath_RF_bus_selected_win_data_686_port, 
                           curr_proc_regs(685) => 
                           DataPath_RF_bus_selected_win_data_685_port, 
                           curr_proc_regs(684) => 
                           DataPath_RF_bus_selected_win_data_684_port, 
                           curr_proc_regs(683) => 
                           DataPath_RF_bus_selected_win_data_683_port, 
                           curr_proc_regs(682) => 
                           DataPath_RF_bus_selected_win_data_682_port, 
                           curr_proc_regs(681) => 
                           DataPath_RF_bus_selected_win_data_681_port, 
                           curr_proc_regs(680) => 
                           DataPath_RF_bus_selected_win_data_680_port, 
                           curr_proc_regs(679) => 
                           DataPath_RF_bus_selected_win_data_679_port, 
                           curr_proc_regs(678) => 
                           DataPath_RF_bus_selected_win_data_678_port, 
                           curr_proc_regs(677) => 
                           DataPath_RF_bus_selected_win_data_677_port, 
                           curr_proc_regs(676) => 
                           DataPath_RF_bus_selected_win_data_676_port, 
                           curr_proc_regs(675) => 
                           DataPath_RF_bus_selected_win_data_675_port, 
                           curr_proc_regs(674) => 
                           DataPath_RF_bus_selected_win_data_674_port, 
                           curr_proc_regs(673) => 
                           DataPath_RF_bus_selected_win_data_673_port, 
                           curr_proc_regs(672) => 
                           DataPath_RF_bus_selected_win_data_672_port, 
                           curr_proc_regs(671) => 
                           DataPath_RF_bus_selected_win_data_671_port, 
                           curr_proc_regs(670) => 
                           DataPath_RF_bus_selected_win_data_670_port, 
                           curr_proc_regs(669) => 
                           DataPath_RF_bus_selected_win_data_669_port, 
                           curr_proc_regs(668) => 
                           DataPath_RF_bus_selected_win_data_668_port, 
                           curr_proc_regs(667) => 
                           DataPath_RF_bus_selected_win_data_667_port, 
                           curr_proc_regs(666) => 
                           DataPath_RF_bus_selected_win_data_666_port, 
                           curr_proc_regs(665) => 
                           DataPath_RF_bus_selected_win_data_665_port, 
                           curr_proc_regs(664) => 
                           DataPath_RF_bus_selected_win_data_664_port, 
                           curr_proc_regs(663) => 
                           DataPath_RF_bus_selected_win_data_663_port, 
                           curr_proc_regs(662) => 
                           DataPath_RF_bus_selected_win_data_662_port, 
                           curr_proc_regs(661) => 
                           DataPath_RF_bus_selected_win_data_661_port, 
                           curr_proc_regs(660) => 
                           DataPath_RF_bus_selected_win_data_660_port, 
                           curr_proc_regs(659) => 
                           DataPath_RF_bus_selected_win_data_659_port, 
                           curr_proc_regs(658) => 
                           DataPath_RF_bus_selected_win_data_658_port, 
                           curr_proc_regs(657) => 
                           DataPath_RF_bus_selected_win_data_657_port, 
                           curr_proc_regs(656) => 
                           DataPath_RF_bus_selected_win_data_656_port, 
                           curr_proc_regs(655) => 
                           DataPath_RF_bus_selected_win_data_655_port, 
                           curr_proc_regs(654) => 
                           DataPath_RF_bus_selected_win_data_654_port, 
                           curr_proc_regs(653) => 
                           DataPath_RF_bus_selected_win_data_653_port, 
                           curr_proc_regs(652) => 
                           DataPath_RF_bus_selected_win_data_652_port, 
                           curr_proc_regs(651) => 
                           DataPath_RF_bus_selected_win_data_651_port, 
                           curr_proc_regs(650) => 
                           DataPath_RF_bus_selected_win_data_650_port, 
                           curr_proc_regs(649) => 
                           DataPath_RF_bus_selected_win_data_649_port, 
                           curr_proc_regs(648) => 
                           DataPath_RF_bus_selected_win_data_648_port, 
                           curr_proc_regs(647) => 
                           DataPath_RF_bus_selected_win_data_647_port, 
                           curr_proc_regs(646) => 
                           DataPath_RF_bus_selected_win_data_646_port, 
                           curr_proc_regs(645) => 
                           DataPath_RF_bus_selected_win_data_645_port, 
                           curr_proc_regs(644) => 
                           DataPath_RF_bus_selected_win_data_644_port, 
                           curr_proc_regs(643) => 
                           DataPath_RF_bus_selected_win_data_643_port, 
                           curr_proc_regs(642) => 
                           DataPath_RF_bus_selected_win_data_642_port, 
                           curr_proc_regs(641) => 
                           DataPath_RF_bus_selected_win_data_641_port, 
                           curr_proc_regs(640) => 
                           DataPath_RF_bus_selected_win_data_640_port, 
                           curr_proc_regs(639) => 
                           DataPath_RF_bus_selected_win_data_639_port, 
                           curr_proc_regs(638) => 
                           DataPath_RF_bus_selected_win_data_638_port, 
                           curr_proc_regs(637) => 
                           DataPath_RF_bus_selected_win_data_637_port, 
                           curr_proc_regs(636) => 
                           DataPath_RF_bus_selected_win_data_636_port, 
                           curr_proc_regs(635) => 
                           DataPath_RF_bus_selected_win_data_635_port, 
                           curr_proc_regs(634) => 
                           DataPath_RF_bus_selected_win_data_634_port, 
                           curr_proc_regs(633) => 
                           DataPath_RF_bus_selected_win_data_633_port, 
                           curr_proc_regs(632) => 
                           DataPath_RF_bus_selected_win_data_632_port, 
                           curr_proc_regs(631) => 
                           DataPath_RF_bus_selected_win_data_631_port, 
                           curr_proc_regs(630) => 
                           DataPath_RF_bus_selected_win_data_630_port, 
                           curr_proc_regs(629) => 
                           DataPath_RF_bus_selected_win_data_629_port, 
                           curr_proc_regs(628) => 
                           DataPath_RF_bus_selected_win_data_628_port, 
                           curr_proc_regs(627) => 
                           DataPath_RF_bus_selected_win_data_627_port, 
                           curr_proc_regs(626) => 
                           DataPath_RF_bus_selected_win_data_626_port, 
                           curr_proc_regs(625) => 
                           DataPath_RF_bus_selected_win_data_625_port, 
                           curr_proc_regs(624) => 
                           DataPath_RF_bus_selected_win_data_624_port, 
                           curr_proc_regs(623) => 
                           DataPath_RF_bus_selected_win_data_623_port, 
                           curr_proc_regs(622) => 
                           DataPath_RF_bus_selected_win_data_622_port, 
                           curr_proc_regs(621) => 
                           DataPath_RF_bus_selected_win_data_621_port, 
                           curr_proc_regs(620) => 
                           DataPath_RF_bus_selected_win_data_620_port, 
                           curr_proc_regs(619) => 
                           DataPath_RF_bus_selected_win_data_619_port, 
                           curr_proc_regs(618) => 
                           DataPath_RF_bus_selected_win_data_618_port, 
                           curr_proc_regs(617) => 
                           DataPath_RF_bus_selected_win_data_617_port, 
                           curr_proc_regs(616) => 
                           DataPath_RF_bus_selected_win_data_616_port, 
                           curr_proc_regs(615) => 
                           DataPath_RF_bus_selected_win_data_615_port, 
                           curr_proc_regs(614) => 
                           DataPath_RF_bus_selected_win_data_614_port, 
                           curr_proc_regs(613) => 
                           DataPath_RF_bus_selected_win_data_613_port, 
                           curr_proc_regs(612) => 
                           DataPath_RF_bus_selected_win_data_612_port, 
                           curr_proc_regs(611) => 
                           DataPath_RF_bus_selected_win_data_611_port, 
                           curr_proc_regs(610) => 
                           DataPath_RF_bus_selected_win_data_610_port, 
                           curr_proc_regs(609) => 
                           DataPath_RF_bus_selected_win_data_609_port, 
                           curr_proc_regs(608) => 
                           DataPath_RF_bus_selected_win_data_608_port, 
                           curr_proc_regs(607) => 
                           DataPath_RF_bus_selected_win_data_607_port, 
                           curr_proc_regs(606) => 
                           DataPath_RF_bus_selected_win_data_606_port, 
                           curr_proc_regs(605) => 
                           DataPath_RF_bus_selected_win_data_605_port, 
                           curr_proc_regs(604) => 
                           DataPath_RF_bus_selected_win_data_604_port, 
                           curr_proc_regs(603) => 
                           DataPath_RF_bus_selected_win_data_603_port, 
                           curr_proc_regs(602) => 
                           DataPath_RF_bus_selected_win_data_602_port, 
                           curr_proc_regs(601) => 
                           DataPath_RF_bus_selected_win_data_601_port, 
                           curr_proc_regs(600) => 
                           DataPath_RF_bus_selected_win_data_600_port, 
                           curr_proc_regs(599) => 
                           DataPath_RF_bus_selected_win_data_599_port, 
                           curr_proc_regs(598) => 
                           DataPath_RF_bus_selected_win_data_598_port, 
                           curr_proc_regs(597) => 
                           DataPath_RF_bus_selected_win_data_597_port, 
                           curr_proc_regs(596) => 
                           DataPath_RF_bus_selected_win_data_596_port, 
                           curr_proc_regs(595) => 
                           DataPath_RF_bus_selected_win_data_595_port, 
                           curr_proc_regs(594) => 
                           DataPath_RF_bus_selected_win_data_594_port, 
                           curr_proc_regs(593) => 
                           DataPath_RF_bus_selected_win_data_593_port, 
                           curr_proc_regs(592) => 
                           DataPath_RF_bus_selected_win_data_592_port, 
                           curr_proc_regs(591) => 
                           DataPath_RF_bus_selected_win_data_591_port, 
                           curr_proc_regs(590) => 
                           DataPath_RF_bus_selected_win_data_590_port, 
                           curr_proc_regs(589) => 
                           DataPath_RF_bus_selected_win_data_589_port, 
                           curr_proc_regs(588) => 
                           DataPath_RF_bus_selected_win_data_588_port, 
                           curr_proc_regs(587) => 
                           DataPath_RF_bus_selected_win_data_587_port, 
                           curr_proc_regs(586) => 
                           DataPath_RF_bus_selected_win_data_586_port, 
                           curr_proc_regs(585) => 
                           DataPath_RF_bus_selected_win_data_585_port, 
                           curr_proc_regs(584) => 
                           DataPath_RF_bus_selected_win_data_584_port, 
                           curr_proc_regs(583) => 
                           DataPath_RF_bus_selected_win_data_583_port, 
                           curr_proc_regs(582) => 
                           DataPath_RF_bus_selected_win_data_582_port, 
                           curr_proc_regs(581) => 
                           DataPath_RF_bus_selected_win_data_581_port, 
                           curr_proc_regs(580) => 
                           DataPath_RF_bus_selected_win_data_580_port, 
                           curr_proc_regs(579) => 
                           DataPath_RF_bus_selected_win_data_579_port, 
                           curr_proc_regs(578) => 
                           DataPath_RF_bus_selected_win_data_578_port, 
                           curr_proc_regs(577) => 
                           DataPath_RF_bus_selected_win_data_577_port, 
                           curr_proc_regs(576) => 
                           DataPath_RF_bus_selected_win_data_576_port, 
                           curr_proc_regs(575) => 
                           DataPath_RF_bus_selected_win_data_575_port, 
                           curr_proc_regs(574) => 
                           DataPath_RF_bus_selected_win_data_574_port, 
                           curr_proc_regs(573) => 
                           DataPath_RF_bus_selected_win_data_573_port, 
                           curr_proc_regs(572) => 
                           DataPath_RF_bus_selected_win_data_572_port, 
                           curr_proc_regs(571) => 
                           DataPath_RF_bus_selected_win_data_571_port, 
                           curr_proc_regs(570) => 
                           DataPath_RF_bus_selected_win_data_570_port, 
                           curr_proc_regs(569) => 
                           DataPath_RF_bus_selected_win_data_569_port, 
                           curr_proc_regs(568) => 
                           DataPath_RF_bus_selected_win_data_568_port, 
                           curr_proc_regs(567) => 
                           DataPath_RF_bus_selected_win_data_567_port, 
                           curr_proc_regs(566) => 
                           DataPath_RF_bus_selected_win_data_566_port, 
                           curr_proc_regs(565) => 
                           DataPath_RF_bus_selected_win_data_565_port, 
                           curr_proc_regs(564) => 
                           DataPath_RF_bus_selected_win_data_564_port, 
                           curr_proc_regs(563) => 
                           DataPath_RF_bus_selected_win_data_563_port, 
                           curr_proc_regs(562) => 
                           DataPath_RF_bus_selected_win_data_562_port, 
                           curr_proc_regs(561) => 
                           DataPath_RF_bus_selected_win_data_561_port, 
                           curr_proc_regs(560) => 
                           DataPath_RF_bus_selected_win_data_560_port, 
                           curr_proc_regs(559) => 
                           DataPath_RF_bus_selected_win_data_559_port, 
                           curr_proc_regs(558) => 
                           DataPath_RF_bus_selected_win_data_558_port, 
                           curr_proc_regs(557) => 
                           DataPath_RF_bus_selected_win_data_557_port, 
                           curr_proc_regs(556) => 
                           DataPath_RF_bus_selected_win_data_556_port, 
                           curr_proc_regs(555) => 
                           DataPath_RF_bus_selected_win_data_555_port, 
                           curr_proc_regs(554) => 
                           DataPath_RF_bus_selected_win_data_554_port, 
                           curr_proc_regs(553) => 
                           DataPath_RF_bus_selected_win_data_553_port, 
                           curr_proc_regs(552) => 
                           DataPath_RF_bus_selected_win_data_552_port, 
                           curr_proc_regs(551) => 
                           DataPath_RF_bus_selected_win_data_551_port, 
                           curr_proc_regs(550) => 
                           DataPath_RF_bus_selected_win_data_550_port, 
                           curr_proc_regs(549) => 
                           DataPath_RF_bus_selected_win_data_549_port, 
                           curr_proc_regs(548) => 
                           DataPath_RF_bus_selected_win_data_548_port, 
                           curr_proc_regs(547) => 
                           DataPath_RF_bus_selected_win_data_547_port, 
                           curr_proc_regs(546) => 
                           DataPath_RF_bus_selected_win_data_546_port, 
                           curr_proc_regs(545) => 
                           DataPath_RF_bus_selected_win_data_545_port, 
                           curr_proc_regs(544) => 
                           DataPath_RF_bus_selected_win_data_544_port, 
                           curr_proc_regs(543) => 
                           DataPath_RF_bus_selected_win_data_543_port, 
                           curr_proc_regs(542) => 
                           DataPath_RF_bus_selected_win_data_542_port, 
                           curr_proc_regs(541) => 
                           DataPath_RF_bus_selected_win_data_541_port, 
                           curr_proc_regs(540) => 
                           DataPath_RF_bus_selected_win_data_540_port, 
                           curr_proc_regs(539) => 
                           DataPath_RF_bus_selected_win_data_539_port, 
                           curr_proc_regs(538) => 
                           DataPath_RF_bus_selected_win_data_538_port, 
                           curr_proc_regs(537) => 
                           DataPath_RF_bus_selected_win_data_537_port, 
                           curr_proc_regs(536) => 
                           DataPath_RF_bus_selected_win_data_536_port, 
                           curr_proc_regs(535) => 
                           DataPath_RF_bus_selected_win_data_535_port, 
                           curr_proc_regs(534) => 
                           DataPath_RF_bus_selected_win_data_534_port, 
                           curr_proc_regs(533) => 
                           DataPath_RF_bus_selected_win_data_533_port, 
                           curr_proc_regs(532) => 
                           DataPath_RF_bus_selected_win_data_532_port, 
                           curr_proc_regs(531) => 
                           DataPath_RF_bus_selected_win_data_531_port, 
                           curr_proc_regs(530) => 
                           DataPath_RF_bus_selected_win_data_530_port, 
                           curr_proc_regs(529) => 
                           DataPath_RF_bus_selected_win_data_529_port, 
                           curr_proc_regs(528) => 
                           DataPath_RF_bus_selected_win_data_528_port, 
                           curr_proc_regs(527) => 
                           DataPath_RF_bus_selected_win_data_527_port, 
                           curr_proc_regs(526) => 
                           DataPath_RF_bus_selected_win_data_526_port, 
                           curr_proc_regs(525) => 
                           DataPath_RF_bus_selected_win_data_525_port, 
                           curr_proc_regs(524) => 
                           DataPath_RF_bus_selected_win_data_524_port, 
                           curr_proc_regs(523) => 
                           DataPath_RF_bus_selected_win_data_523_port, 
                           curr_proc_regs(522) => 
                           DataPath_RF_bus_selected_win_data_522_port, 
                           curr_proc_regs(521) => 
                           DataPath_RF_bus_selected_win_data_521_port, 
                           curr_proc_regs(520) => 
                           DataPath_RF_bus_selected_win_data_520_port, 
                           curr_proc_regs(519) => 
                           DataPath_RF_bus_selected_win_data_519_port, 
                           curr_proc_regs(518) => 
                           DataPath_RF_bus_selected_win_data_518_port, 
                           curr_proc_regs(517) => 
                           DataPath_RF_bus_selected_win_data_517_port, 
                           curr_proc_regs(516) => 
                           DataPath_RF_bus_selected_win_data_516_port, 
                           curr_proc_regs(515) => 
                           DataPath_RF_bus_selected_win_data_515_port, 
                           curr_proc_regs(514) => 
                           DataPath_RF_bus_selected_win_data_514_port, 
                           curr_proc_regs(513) => 
                           DataPath_RF_bus_selected_win_data_513_port, 
                           curr_proc_regs(512) => 
                           DataPath_RF_bus_selected_win_data_512_port, 
                           curr_proc_regs(511) => 
                           DataPath_RF_bus_selected_win_data_511_port, 
                           curr_proc_regs(510) => 
                           DataPath_RF_bus_selected_win_data_510_port, 
                           curr_proc_regs(509) => 
                           DataPath_RF_bus_selected_win_data_509_port, 
                           curr_proc_regs(508) => 
                           DataPath_RF_bus_selected_win_data_508_port, 
                           curr_proc_regs(507) => 
                           DataPath_RF_bus_selected_win_data_507_port, 
                           curr_proc_regs(506) => 
                           DataPath_RF_bus_selected_win_data_506_port, 
                           curr_proc_regs(505) => 
                           DataPath_RF_bus_selected_win_data_505_port, 
                           curr_proc_regs(504) => 
                           DataPath_RF_bus_selected_win_data_504_port, 
                           curr_proc_regs(503) => 
                           DataPath_RF_bus_selected_win_data_503_port, 
                           curr_proc_regs(502) => 
                           DataPath_RF_bus_selected_win_data_502_port, 
                           curr_proc_regs(501) => 
                           DataPath_RF_bus_selected_win_data_501_port, 
                           curr_proc_regs(500) => 
                           DataPath_RF_bus_selected_win_data_500_port, 
                           curr_proc_regs(499) => 
                           DataPath_RF_bus_selected_win_data_499_port, 
                           curr_proc_regs(498) => 
                           DataPath_RF_bus_selected_win_data_498_port, 
                           curr_proc_regs(497) => 
                           DataPath_RF_bus_selected_win_data_497_port, 
                           curr_proc_regs(496) => 
                           DataPath_RF_bus_selected_win_data_496_port, 
                           curr_proc_regs(495) => 
                           DataPath_RF_bus_selected_win_data_495_port, 
                           curr_proc_regs(494) => 
                           DataPath_RF_bus_selected_win_data_494_port, 
                           curr_proc_regs(493) => 
                           DataPath_RF_bus_selected_win_data_493_port, 
                           curr_proc_regs(492) => 
                           DataPath_RF_bus_selected_win_data_492_port, 
                           curr_proc_regs(491) => 
                           DataPath_RF_bus_selected_win_data_491_port, 
                           curr_proc_regs(490) => 
                           DataPath_RF_bus_selected_win_data_490_port, 
                           curr_proc_regs(489) => 
                           DataPath_RF_bus_selected_win_data_489_port, 
                           curr_proc_regs(488) => 
                           DataPath_RF_bus_selected_win_data_488_port, 
                           curr_proc_regs(487) => 
                           DataPath_RF_bus_selected_win_data_487_port, 
                           curr_proc_regs(486) => 
                           DataPath_RF_bus_selected_win_data_486_port, 
                           curr_proc_regs(485) => 
                           DataPath_RF_bus_selected_win_data_485_port, 
                           curr_proc_regs(484) => 
                           DataPath_RF_bus_selected_win_data_484_port, 
                           curr_proc_regs(483) => 
                           DataPath_RF_bus_selected_win_data_483_port, 
                           curr_proc_regs(482) => 
                           DataPath_RF_bus_selected_win_data_482_port, 
                           curr_proc_regs(481) => 
                           DataPath_RF_bus_selected_win_data_481_port, 
                           curr_proc_regs(480) => 
                           DataPath_RF_bus_selected_win_data_480_port, 
                           curr_proc_regs(479) => 
                           DataPath_RF_bus_selected_win_data_479_port, 
                           curr_proc_regs(478) => 
                           DataPath_RF_bus_selected_win_data_478_port, 
                           curr_proc_regs(477) => 
                           DataPath_RF_bus_selected_win_data_477_port, 
                           curr_proc_regs(476) => 
                           DataPath_RF_bus_selected_win_data_476_port, 
                           curr_proc_regs(475) => 
                           DataPath_RF_bus_selected_win_data_475_port, 
                           curr_proc_regs(474) => 
                           DataPath_RF_bus_selected_win_data_474_port, 
                           curr_proc_regs(473) => 
                           DataPath_RF_bus_selected_win_data_473_port, 
                           curr_proc_regs(472) => 
                           DataPath_RF_bus_selected_win_data_472_port, 
                           curr_proc_regs(471) => 
                           DataPath_RF_bus_selected_win_data_471_port, 
                           curr_proc_regs(470) => 
                           DataPath_RF_bus_selected_win_data_470_port, 
                           curr_proc_regs(469) => 
                           DataPath_RF_bus_selected_win_data_469_port, 
                           curr_proc_regs(468) => 
                           DataPath_RF_bus_selected_win_data_468_port, 
                           curr_proc_regs(467) => 
                           DataPath_RF_bus_selected_win_data_467_port, 
                           curr_proc_regs(466) => 
                           DataPath_RF_bus_selected_win_data_466_port, 
                           curr_proc_regs(465) => 
                           DataPath_RF_bus_selected_win_data_465_port, 
                           curr_proc_regs(464) => 
                           DataPath_RF_bus_selected_win_data_464_port, 
                           curr_proc_regs(463) => 
                           DataPath_RF_bus_selected_win_data_463_port, 
                           curr_proc_regs(462) => 
                           DataPath_RF_bus_selected_win_data_462_port, 
                           curr_proc_regs(461) => 
                           DataPath_RF_bus_selected_win_data_461_port, 
                           curr_proc_regs(460) => 
                           DataPath_RF_bus_selected_win_data_460_port, 
                           curr_proc_regs(459) => 
                           DataPath_RF_bus_selected_win_data_459_port, 
                           curr_proc_regs(458) => 
                           DataPath_RF_bus_selected_win_data_458_port, 
                           curr_proc_regs(457) => 
                           DataPath_RF_bus_selected_win_data_457_port, 
                           curr_proc_regs(456) => 
                           DataPath_RF_bus_selected_win_data_456_port, 
                           curr_proc_regs(455) => 
                           DataPath_RF_bus_selected_win_data_455_port, 
                           curr_proc_regs(454) => 
                           DataPath_RF_bus_selected_win_data_454_port, 
                           curr_proc_regs(453) => 
                           DataPath_RF_bus_selected_win_data_453_port, 
                           curr_proc_regs(452) => 
                           DataPath_RF_bus_selected_win_data_452_port, 
                           curr_proc_regs(451) => 
                           DataPath_RF_bus_selected_win_data_451_port, 
                           curr_proc_regs(450) => 
                           DataPath_RF_bus_selected_win_data_450_port, 
                           curr_proc_regs(449) => 
                           DataPath_RF_bus_selected_win_data_449_port, 
                           curr_proc_regs(448) => 
                           DataPath_RF_bus_selected_win_data_448_port, 
                           curr_proc_regs(447) => 
                           DataPath_RF_bus_selected_win_data_447_port, 
                           curr_proc_regs(446) => 
                           DataPath_RF_bus_selected_win_data_446_port, 
                           curr_proc_regs(445) => 
                           DataPath_RF_bus_selected_win_data_445_port, 
                           curr_proc_regs(444) => 
                           DataPath_RF_bus_selected_win_data_444_port, 
                           curr_proc_regs(443) => 
                           DataPath_RF_bus_selected_win_data_443_port, 
                           curr_proc_regs(442) => 
                           DataPath_RF_bus_selected_win_data_442_port, 
                           curr_proc_regs(441) => 
                           DataPath_RF_bus_selected_win_data_441_port, 
                           curr_proc_regs(440) => 
                           DataPath_RF_bus_selected_win_data_440_port, 
                           curr_proc_regs(439) => 
                           DataPath_RF_bus_selected_win_data_439_port, 
                           curr_proc_regs(438) => 
                           DataPath_RF_bus_selected_win_data_438_port, 
                           curr_proc_regs(437) => 
                           DataPath_RF_bus_selected_win_data_437_port, 
                           curr_proc_regs(436) => 
                           DataPath_RF_bus_selected_win_data_436_port, 
                           curr_proc_regs(435) => 
                           DataPath_RF_bus_selected_win_data_435_port, 
                           curr_proc_regs(434) => 
                           DataPath_RF_bus_selected_win_data_434_port, 
                           curr_proc_regs(433) => 
                           DataPath_RF_bus_selected_win_data_433_port, 
                           curr_proc_regs(432) => 
                           DataPath_RF_bus_selected_win_data_432_port, 
                           curr_proc_regs(431) => 
                           DataPath_RF_bus_selected_win_data_431_port, 
                           curr_proc_regs(430) => 
                           DataPath_RF_bus_selected_win_data_430_port, 
                           curr_proc_regs(429) => 
                           DataPath_RF_bus_selected_win_data_429_port, 
                           curr_proc_regs(428) => 
                           DataPath_RF_bus_selected_win_data_428_port, 
                           curr_proc_regs(427) => 
                           DataPath_RF_bus_selected_win_data_427_port, 
                           curr_proc_regs(426) => 
                           DataPath_RF_bus_selected_win_data_426_port, 
                           curr_proc_regs(425) => 
                           DataPath_RF_bus_selected_win_data_425_port, 
                           curr_proc_regs(424) => 
                           DataPath_RF_bus_selected_win_data_424_port, 
                           curr_proc_regs(423) => 
                           DataPath_RF_bus_selected_win_data_423_port, 
                           curr_proc_regs(422) => 
                           DataPath_RF_bus_selected_win_data_422_port, 
                           curr_proc_regs(421) => 
                           DataPath_RF_bus_selected_win_data_421_port, 
                           curr_proc_regs(420) => 
                           DataPath_RF_bus_selected_win_data_420_port, 
                           curr_proc_regs(419) => 
                           DataPath_RF_bus_selected_win_data_419_port, 
                           curr_proc_regs(418) => 
                           DataPath_RF_bus_selected_win_data_418_port, 
                           curr_proc_regs(417) => 
                           DataPath_RF_bus_selected_win_data_417_port, 
                           curr_proc_regs(416) => 
                           DataPath_RF_bus_selected_win_data_416_port, 
                           curr_proc_regs(415) => 
                           DataPath_RF_bus_selected_win_data_415_port, 
                           curr_proc_regs(414) => 
                           DataPath_RF_bus_selected_win_data_414_port, 
                           curr_proc_regs(413) => 
                           DataPath_RF_bus_selected_win_data_413_port, 
                           curr_proc_regs(412) => 
                           DataPath_RF_bus_selected_win_data_412_port, 
                           curr_proc_regs(411) => 
                           DataPath_RF_bus_selected_win_data_411_port, 
                           curr_proc_regs(410) => 
                           DataPath_RF_bus_selected_win_data_410_port, 
                           curr_proc_regs(409) => 
                           DataPath_RF_bus_selected_win_data_409_port, 
                           curr_proc_regs(408) => 
                           DataPath_RF_bus_selected_win_data_408_port, 
                           curr_proc_regs(407) => 
                           DataPath_RF_bus_selected_win_data_407_port, 
                           curr_proc_regs(406) => 
                           DataPath_RF_bus_selected_win_data_406_port, 
                           curr_proc_regs(405) => 
                           DataPath_RF_bus_selected_win_data_405_port, 
                           curr_proc_regs(404) => 
                           DataPath_RF_bus_selected_win_data_404_port, 
                           curr_proc_regs(403) => 
                           DataPath_RF_bus_selected_win_data_403_port, 
                           curr_proc_regs(402) => 
                           DataPath_RF_bus_selected_win_data_402_port, 
                           curr_proc_regs(401) => 
                           DataPath_RF_bus_selected_win_data_401_port, 
                           curr_proc_regs(400) => 
                           DataPath_RF_bus_selected_win_data_400_port, 
                           curr_proc_regs(399) => 
                           DataPath_RF_bus_selected_win_data_399_port, 
                           curr_proc_regs(398) => 
                           DataPath_RF_bus_selected_win_data_398_port, 
                           curr_proc_regs(397) => 
                           DataPath_RF_bus_selected_win_data_397_port, 
                           curr_proc_regs(396) => 
                           DataPath_RF_bus_selected_win_data_396_port, 
                           curr_proc_regs(395) => 
                           DataPath_RF_bus_selected_win_data_395_port, 
                           curr_proc_regs(394) => 
                           DataPath_RF_bus_selected_win_data_394_port, 
                           curr_proc_regs(393) => 
                           DataPath_RF_bus_selected_win_data_393_port, 
                           curr_proc_regs(392) => 
                           DataPath_RF_bus_selected_win_data_392_port, 
                           curr_proc_regs(391) => 
                           DataPath_RF_bus_selected_win_data_391_port, 
                           curr_proc_regs(390) => 
                           DataPath_RF_bus_selected_win_data_390_port, 
                           curr_proc_regs(389) => 
                           DataPath_RF_bus_selected_win_data_389_port, 
                           curr_proc_regs(388) => 
                           DataPath_RF_bus_selected_win_data_388_port, 
                           curr_proc_regs(387) => 
                           DataPath_RF_bus_selected_win_data_387_port, 
                           curr_proc_regs(386) => 
                           DataPath_RF_bus_selected_win_data_386_port, 
                           curr_proc_regs(385) => 
                           DataPath_RF_bus_selected_win_data_385_port, 
                           curr_proc_regs(384) => 
                           DataPath_RF_bus_selected_win_data_384_port, 
                           curr_proc_regs(383) => 
                           DataPath_RF_bus_selected_win_data_383_port, 
                           curr_proc_regs(382) => 
                           DataPath_RF_bus_selected_win_data_382_port, 
                           curr_proc_regs(381) => 
                           DataPath_RF_bus_selected_win_data_381_port, 
                           curr_proc_regs(380) => 
                           DataPath_RF_bus_selected_win_data_380_port, 
                           curr_proc_regs(379) => 
                           DataPath_RF_bus_selected_win_data_379_port, 
                           curr_proc_regs(378) => 
                           DataPath_RF_bus_selected_win_data_378_port, 
                           curr_proc_regs(377) => 
                           DataPath_RF_bus_selected_win_data_377_port, 
                           curr_proc_regs(376) => 
                           DataPath_RF_bus_selected_win_data_376_port, 
                           curr_proc_regs(375) => 
                           DataPath_RF_bus_selected_win_data_375_port, 
                           curr_proc_regs(374) => 
                           DataPath_RF_bus_selected_win_data_374_port, 
                           curr_proc_regs(373) => 
                           DataPath_RF_bus_selected_win_data_373_port, 
                           curr_proc_regs(372) => 
                           DataPath_RF_bus_selected_win_data_372_port, 
                           curr_proc_regs(371) => 
                           DataPath_RF_bus_selected_win_data_371_port, 
                           curr_proc_regs(370) => 
                           DataPath_RF_bus_selected_win_data_370_port, 
                           curr_proc_regs(369) => 
                           DataPath_RF_bus_selected_win_data_369_port, 
                           curr_proc_regs(368) => 
                           DataPath_RF_bus_selected_win_data_368_port, 
                           curr_proc_regs(367) => 
                           DataPath_RF_bus_selected_win_data_367_port, 
                           curr_proc_regs(366) => 
                           DataPath_RF_bus_selected_win_data_366_port, 
                           curr_proc_regs(365) => 
                           DataPath_RF_bus_selected_win_data_365_port, 
                           curr_proc_regs(364) => 
                           DataPath_RF_bus_selected_win_data_364_port, 
                           curr_proc_regs(363) => 
                           DataPath_RF_bus_selected_win_data_363_port, 
                           curr_proc_regs(362) => 
                           DataPath_RF_bus_selected_win_data_362_port, 
                           curr_proc_regs(361) => 
                           DataPath_RF_bus_selected_win_data_361_port, 
                           curr_proc_regs(360) => 
                           DataPath_RF_bus_selected_win_data_360_port, 
                           curr_proc_regs(359) => 
                           DataPath_RF_bus_selected_win_data_359_port, 
                           curr_proc_regs(358) => 
                           DataPath_RF_bus_selected_win_data_358_port, 
                           curr_proc_regs(357) => 
                           DataPath_RF_bus_selected_win_data_357_port, 
                           curr_proc_regs(356) => 
                           DataPath_RF_bus_selected_win_data_356_port, 
                           curr_proc_regs(355) => 
                           DataPath_RF_bus_selected_win_data_355_port, 
                           curr_proc_regs(354) => 
                           DataPath_RF_bus_selected_win_data_354_port, 
                           curr_proc_regs(353) => 
                           DataPath_RF_bus_selected_win_data_353_port, 
                           curr_proc_regs(352) => 
                           DataPath_RF_bus_selected_win_data_352_port, 
                           curr_proc_regs(351) => 
                           DataPath_RF_bus_selected_win_data_351_port, 
                           curr_proc_regs(350) => 
                           DataPath_RF_bus_selected_win_data_350_port, 
                           curr_proc_regs(349) => 
                           DataPath_RF_bus_selected_win_data_349_port, 
                           curr_proc_regs(348) => 
                           DataPath_RF_bus_selected_win_data_348_port, 
                           curr_proc_regs(347) => 
                           DataPath_RF_bus_selected_win_data_347_port, 
                           curr_proc_regs(346) => 
                           DataPath_RF_bus_selected_win_data_346_port, 
                           curr_proc_regs(345) => 
                           DataPath_RF_bus_selected_win_data_345_port, 
                           curr_proc_regs(344) => 
                           DataPath_RF_bus_selected_win_data_344_port, 
                           curr_proc_regs(343) => 
                           DataPath_RF_bus_selected_win_data_343_port, 
                           curr_proc_regs(342) => 
                           DataPath_RF_bus_selected_win_data_342_port, 
                           curr_proc_regs(341) => 
                           DataPath_RF_bus_selected_win_data_341_port, 
                           curr_proc_regs(340) => 
                           DataPath_RF_bus_selected_win_data_340_port, 
                           curr_proc_regs(339) => 
                           DataPath_RF_bus_selected_win_data_339_port, 
                           curr_proc_regs(338) => 
                           DataPath_RF_bus_selected_win_data_338_port, 
                           curr_proc_regs(337) => 
                           DataPath_RF_bus_selected_win_data_337_port, 
                           curr_proc_regs(336) => 
                           DataPath_RF_bus_selected_win_data_336_port, 
                           curr_proc_regs(335) => 
                           DataPath_RF_bus_selected_win_data_335_port, 
                           curr_proc_regs(334) => 
                           DataPath_RF_bus_selected_win_data_334_port, 
                           curr_proc_regs(333) => 
                           DataPath_RF_bus_selected_win_data_333_port, 
                           curr_proc_regs(332) => 
                           DataPath_RF_bus_selected_win_data_332_port, 
                           curr_proc_regs(331) => 
                           DataPath_RF_bus_selected_win_data_331_port, 
                           curr_proc_regs(330) => 
                           DataPath_RF_bus_selected_win_data_330_port, 
                           curr_proc_regs(329) => 
                           DataPath_RF_bus_selected_win_data_329_port, 
                           curr_proc_regs(328) => 
                           DataPath_RF_bus_selected_win_data_328_port, 
                           curr_proc_regs(327) => 
                           DataPath_RF_bus_selected_win_data_327_port, 
                           curr_proc_regs(326) => 
                           DataPath_RF_bus_selected_win_data_326_port, 
                           curr_proc_regs(325) => 
                           DataPath_RF_bus_selected_win_data_325_port, 
                           curr_proc_regs(324) => 
                           DataPath_RF_bus_selected_win_data_324_port, 
                           curr_proc_regs(323) => 
                           DataPath_RF_bus_selected_win_data_323_port, 
                           curr_proc_regs(322) => 
                           DataPath_RF_bus_selected_win_data_322_port, 
                           curr_proc_regs(321) => 
                           DataPath_RF_bus_selected_win_data_321_port, 
                           curr_proc_regs(320) => 
                           DataPath_RF_bus_selected_win_data_320_port, 
                           curr_proc_regs(319) => 
                           DataPath_RF_bus_selected_win_data_319_port, 
                           curr_proc_regs(318) => 
                           DataPath_RF_bus_selected_win_data_318_port, 
                           curr_proc_regs(317) => 
                           DataPath_RF_bus_selected_win_data_317_port, 
                           curr_proc_regs(316) => 
                           DataPath_RF_bus_selected_win_data_316_port, 
                           curr_proc_regs(315) => 
                           DataPath_RF_bus_selected_win_data_315_port, 
                           curr_proc_regs(314) => 
                           DataPath_RF_bus_selected_win_data_314_port, 
                           curr_proc_regs(313) => 
                           DataPath_RF_bus_selected_win_data_313_port, 
                           curr_proc_regs(312) => 
                           DataPath_RF_bus_selected_win_data_312_port, 
                           curr_proc_regs(311) => 
                           DataPath_RF_bus_selected_win_data_311_port, 
                           curr_proc_regs(310) => 
                           DataPath_RF_bus_selected_win_data_310_port, 
                           curr_proc_regs(309) => 
                           DataPath_RF_bus_selected_win_data_309_port, 
                           curr_proc_regs(308) => 
                           DataPath_RF_bus_selected_win_data_308_port, 
                           curr_proc_regs(307) => 
                           DataPath_RF_bus_selected_win_data_307_port, 
                           curr_proc_regs(306) => 
                           DataPath_RF_bus_selected_win_data_306_port, 
                           curr_proc_regs(305) => 
                           DataPath_RF_bus_selected_win_data_305_port, 
                           curr_proc_regs(304) => 
                           DataPath_RF_bus_selected_win_data_304_port, 
                           curr_proc_regs(303) => 
                           DataPath_RF_bus_selected_win_data_303_port, 
                           curr_proc_regs(302) => 
                           DataPath_RF_bus_selected_win_data_302_port, 
                           curr_proc_regs(301) => 
                           DataPath_RF_bus_selected_win_data_301_port, 
                           curr_proc_regs(300) => 
                           DataPath_RF_bus_selected_win_data_300_port, 
                           curr_proc_regs(299) => 
                           DataPath_RF_bus_selected_win_data_299_port, 
                           curr_proc_regs(298) => 
                           DataPath_RF_bus_selected_win_data_298_port, 
                           curr_proc_regs(297) => 
                           DataPath_RF_bus_selected_win_data_297_port, 
                           curr_proc_regs(296) => 
                           DataPath_RF_bus_selected_win_data_296_port, 
                           curr_proc_regs(295) => 
                           DataPath_RF_bus_selected_win_data_295_port, 
                           curr_proc_regs(294) => 
                           DataPath_RF_bus_selected_win_data_294_port, 
                           curr_proc_regs(293) => 
                           DataPath_RF_bus_selected_win_data_293_port, 
                           curr_proc_regs(292) => 
                           DataPath_RF_bus_selected_win_data_292_port, 
                           curr_proc_regs(291) => 
                           DataPath_RF_bus_selected_win_data_291_port, 
                           curr_proc_regs(290) => 
                           DataPath_RF_bus_selected_win_data_290_port, 
                           curr_proc_regs(289) => 
                           DataPath_RF_bus_selected_win_data_289_port, 
                           curr_proc_regs(288) => 
                           DataPath_RF_bus_selected_win_data_288_port, 
                           curr_proc_regs(287) => 
                           DataPath_RF_bus_selected_win_data_287_port, 
                           curr_proc_regs(286) => 
                           DataPath_RF_bus_selected_win_data_286_port, 
                           curr_proc_regs(285) => 
                           DataPath_RF_bus_selected_win_data_285_port, 
                           curr_proc_regs(284) => 
                           DataPath_RF_bus_selected_win_data_284_port, 
                           curr_proc_regs(283) => 
                           DataPath_RF_bus_selected_win_data_283_port, 
                           curr_proc_regs(282) => 
                           DataPath_RF_bus_selected_win_data_282_port, 
                           curr_proc_regs(281) => 
                           DataPath_RF_bus_selected_win_data_281_port, 
                           curr_proc_regs(280) => 
                           DataPath_RF_bus_selected_win_data_280_port, 
                           curr_proc_regs(279) => 
                           DataPath_RF_bus_selected_win_data_279_port, 
                           curr_proc_regs(278) => 
                           DataPath_RF_bus_selected_win_data_278_port, 
                           curr_proc_regs(277) => 
                           DataPath_RF_bus_selected_win_data_277_port, 
                           curr_proc_regs(276) => 
                           DataPath_RF_bus_selected_win_data_276_port, 
                           curr_proc_regs(275) => 
                           DataPath_RF_bus_selected_win_data_275_port, 
                           curr_proc_regs(274) => 
                           DataPath_RF_bus_selected_win_data_274_port, 
                           curr_proc_regs(273) => 
                           DataPath_RF_bus_selected_win_data_273_port, 
                           curr_proc_regs(272) => 
                           DataPath_RF_bus_selected_win_data_272_port, 
                           curr_proc_regs(271) => 
                           DataPath_RF_bus_selected_win_data_271_port, 
                           curr_proc_regs(270) => 
                           DataPath_RF_bus_selected_win_data_270_port, 
                           curr_proc_regs(269) => 
                           DataPath_RF_bus_selected_win_data_269_port, 
                           curr_proc_regs(268) => 
                           DataPath_RF_bus_selected_win_data_268_port, 
                           curr_proc_regs(267) => 
                           DataPath_RF_bus_selected_win_data_267_port, 
                           curr_proc_regs(266) => 
                           DataPath_RF_bus_selected_win_data_266_port, 
                           curr_proc_regs(265) => 
                           DataPath_RF_bus_selected_win_data_265_port, 
                           curr_proc_regs(264) => 
                           DataPath_RF_bus_selected_win_data_264_port, 
                           curr_proc_regs(263) => 
                           DataPath_RF_bus_selected_win_data_263_port, 
                           curr_proc_regs(262) => 
                           DataPath_RF_bus_selected_win_data_262_port, 
                           curr_proc_regs(261) => 
                           DataPath_RF_bus_selected_win_data_261_port, 
                           curr_proc_regs(260) => 
                           DataPath_RF_bus_selected_win_data_260_port, 
                           curr_proc_regs(259) => 
                           DataPath_RF_bus_selected_win_data_259_port, 
                           curr_proc_regs(258) => 
                           DataPath_RF_bus_selected_win_data_258_port, 
                           curr_proc_regs(257) => 
                           DataPath_RF_bus_selected_win_data_257_port, 
                           curr_proc_regs(256) => 
                           DataPath_RF_bus_selected_win_data_256_port, 
                           curr_proc_regs(255) => 
                           DataPath_RF_bus_selected_win_data_255_port, 
                           curr_proc_regs(254) => 
                           DataPath_RF_bus_selected_win_data_254_port, 
                           curr_proc_regs(253) => 
                           DataPath_RF_bus_selected_win_data_253_port, 
                           curr_proc_regs(252) => 
                           DataPath_RF_bus_selected_win_data_252_port, 
                           curr_proc_regs(251) => 
                           DataPath_RF_bus_selected_win_data_251_port, 
                           curr_proc_regs(250) => 
                           DataPath_RF_bus_selected_win_data_250_port, 
                           curr_proc_regs(249) => 
                           DataPath_RF_bus_selected_win_data_249_port, 
                           curr_proc_regs(248) => 
                           DataPath_RF_bus_selected_win_data_248_port, 
                           curr_proc_regs(247) => 
                           DataPath_RF_bus_selected_win_data_247_port, 
                           curr_proc_regs(246) => 
                           DataPath_RF_bus_selected_win_data_246_port, 
                           curr_proc_regs(245) => 
                           DataPath_RF_bus_selected_win_data_245_port, 
                           curr_proc_regs(244) => 
                           DataPath_RF_bus_selected_win_data_244_port, 
                           curr_proc_regs(243) => 
                           DataPath_RF_bus_selected_win_data_243_port, 
                           curr_proc_regs(242) => 
                           DataPath_RF_bus_selected_win_data_242_port, 
                           curr_proc_regs(241) => 
                           DataPath_RF_bus_selected_win_data_241_port, 
                           curr_proc_regs(240) => 
                           DataPath_RF_bus_selected_win_data_240_port, 
                           curr_proc_regs(239) => 
                           DataPath_RF_bus_selected_win_data_239_port, 
                           curr_proc_regs(238) => 
                           DataPath_RF_bus_selected_win_data_238_port, 
                           curr_proc_regs(237) => 
                           DataPath_RF_bus_selected_win_data_237_port, 
                           curr_proc_regs(236) => 
                           DataPath_RF_bus_selected_win_data_236_port, 
                           curr_proc_regs(235) => 
                           DataPath_RF_bus_selected_win_data_235_port, 
                           curr_proc_regs(234) => 
                           DataPath_RF_bus_selected_win_data_234_port, 
                           curr_proc_regs(233) => 
                           DataPath_RF_bus_selected_win_data_233_port, 
                           curr_proc_regs(232) => 
                           DataPath_RF_bus_selected_win_data_232_port, 
                           curr_proc_regs(231) => 
                           DataPath_RF_bus_selected_win_data_231_port, 
                           curr_proc_regs(230) => 
                           DataPath_RF_bus_selected_win_data_230_port, 
                           curr_proc_regs(229) => 
                           DataPath_RF_bus_selected_win_data_229_port, 
                           curr_proc_regs(228) => 
                           DataPath_RF_bus_selected_win_data_228_port, 
                           curr_proc_regs(227) => 
                           DataPath_RF_bus_selected_win_data_227_port, 
                           curr_proc_regs(226) => 
                           DataPath_RF_bus_selected_win_data_226_port, 
                           curr_proc_regs(225) => 
                           DataPath_RF_bus_selected_win_data_225_port, 
                           curr_proc_regs(224) => 
                           DataPath_RF_bus_selected_win_data_224_port, 
                           curr_proc_regs(223) => 
                           DataPath_RF_bus_selected_win_data_223_port, 
                           curr_proc_regs(222) => 
                           DataPath_RF_bus_selected_win_data_222_port, 
                           curr_proc_regs(221) => 
                           DataPath_RF_bus_selected_win_data_221_port, 
                           curr_proc_regs(220) => 
                           DataPath_RF_bus_selected_win_data_220_port, 
                           curr_proc_regs(219) => 
                           DataPath_RF_bus_selected_win_data_219_port, 
                           curr_proc_regs(218) => 
                           DataPath_RF_bus_selected_win_data_218_port, 
                           curr_proc_regs(217) => 
                           DataPath_RF_bus_selected_win_data_217_port, 
                           curr_proc_regs(216) => 
                           DataPath_RF_bus_selected_win_data_216_port, 
                           curr_proc_regs(215) => 
                           DataPath_RF_bus_selected_win_data_215_port, 
                           curr_proc_regs(214) => 
                           DataPath_RF_bus_selected_win_data_214_port, 
                           curr_proc_regs(213) => 
                           DataPath_RF_bus_selected_win_data_213_port, 
                           curr_proc_regs(212) => 
                           DataPath_RF_bus_selected_win_data_212_port, 
                           curr_proc_regs(211) => 
                           DataPath_RF_bus_selected_win_data_211_port, 
                           curr_proc_regs(210) => 
                           DataPath_RF_bus_selected_win_data_210_port, 
                           curr_proc_regs(209) => 
                           DataPath_RF_bus_selected_win_data_209_port, 
                           curr_proc_regs(208) => 
                           DataPath_RF_bus_selected_win_data_208_port, 
                           curr_proc_regs(207) => 
                           DataPath_RF_bus_selected_win_data_207_port, 
                           curr_proc_regs(206) => 
                           DataPath_RF_bus_selected_win_data_206_port, 
                           curr_proc_regs(205) => 
                           DataPath_RF_bus_selected_win_data_205_port, 
                           curr_proc_regs(204) => 
                           DataPath_RF_bus_selected_win_data_204_port, 
                           curr_proc_regs(203) => 
                           DataPath_RF_bus_selected_win_data_203_port, 
                           curr_proc_regs(202) => 
                           DataPath_RF_bus_selected_win_data_202_port, 
                           curr_proc_regs(201) => 
                           DataPath_RF_bus_selected_win_data_201_port, 
                           curr_proc_regs(200) => 
                           DataPath_RF_bus_selected_win_data_200_port, 
                           curr_proc_regs(199) => 
                           DataPath_RF_bus_selected_win_data_199_port, 
                           curr_proc_regs(198) => 
                           DataPath_RF_bus_selected_win_data_198_port, 
                           curr_proc_regs(197) => 
                           DataPath_RF_bus_selected_win_data_197_port, 
                           curr_proc_regs(196) => 
                           DataPath_RF_bus_selected_win_data_196_port, 
                           curr_proc_regs(195) => 
                           DataPath_RF_bus_selected_win_data_195_port, 
                           curr_proc_regs(194) => 
                           DataPath_RF_bus_selected_win_data_194_port, 
                           curr_proc_regs(193) => 
                           DataPath_RF_bus_selected_win_data_193_port, 
                           curr_proc_regs(192) => 
                           DataPath_RF_bus_selected_win_data_192_port, 
                           curr_proc_regs(191) => 
                           DataPath_RF_bus_selected_win_data_191_port, 
                           curr_proc_regs(190) => 
                           DataPath_RF_bus_selected_win_data_190_port, 
                           curr_proc_regs(189) => 
                           DataPath_RF_bus_selected_win_data_189_port, 
                           curr_proc_regs(188) => 
                           DataPath_RF_bus_selected_win_data_188_port, 
                           curr_proc_regs(187) => 
                           DataPath_RF_bus_selected_win_data_187_port, 
                           curr_proc_regs(186) => 
                           DataPath_RF_bus_selected_win_data_186_port, 
                           curr_proc_regs(185) => 
                           DataPath_RF_bus_selected_win_data_185_port, 
                           curr_proc_regs(184) => 
                           DataPath_RF_bus_selected_win_data_184_port, 
                           curr_proc_regs(183) => 
                           DataPath_RF_bus_selected_win_data_183_port, 
                           curr_proc_regs(182) => 
                           DataPath_RF_bus_selected_win_data_182_port, 
                           curr_proc_regs(181) => 
                           DataPath_RF_bus_selected_win_data_181_port, 
                           curr_proc_regs(180) => 
                           DataPath_RF_bus_selected_win_data_180_port, 
                           curr_proc_regs(179) => 
                           DataPath_RF_bus_selected_win_data_179_port, 
                           curr_proc_regs(178) => 
                           DataPath_RF_bus_selected_win_data_178_port, 
                           curr_proc_regs(177) => 
                           DataPath_RF_bus_selected_win_data_177_port, 
                           curr_proc_regs(176) => 
                           DataPath_RF_bus_selected_win_data_176_port, 
                           curr_proc_regs(175) => 
                           DataPath_RF_bus_selected_win_data_175_port, 
                           curr_proc_regs(174) => 
                           DataPath_RF_bus_selected_win_data_174_port, 
                           curr_proc_regs(173) => 
                           DataPath_RF_bus_selected_win_data_173_port, 
                           curr_proc_regs(172) => 
                           DataPath_RF_bus_selected_win_data_172_port, 
                           curr_proc_regs(171) => 
                           DataPath_RF_bus_selected_win_data_171_port, 
                           curr_proc_regs(170) => 
                           DataPath_RF_bus_selected_win_data_170_port, 
                           curr_proc_regs(169) => 
                           DataPath_RF_bus_selected_win_data_169_port, 
                           curr_proc_regs(168) => 
                           DataPath_RF_bus_selected_win_data_168_port, 
                           curr_proc_regs(167) => 
                           DataPath_RF_bus_selected_win_data_167_port, 
                           curr_proc_regs(166) => 
                           DataPath_RF_bus_selected_win_data_166_port, 
                           curr_proc_regs(165) => 
                           DataPath_RF_bus_selected_win_data_165_port, 
                           curr_proc_regs(164) => 
                           DataPath_RF_bus_selected_win_data_164_port, 
                           curr_proc_regs(163) => 
                           DataPath_RF_bus_selected_win_data_163_port, 
                           curr_proc_regs(162) => 
                           DataPath_RF_bus_selected_win_data_162_port, 
                           curr_proc_regs(161) => 
                           DataPath_RF_bus_selected_win_data_161_port, 
                           curr_proc_regs(160) => 
                           DataPath_RF_bus_selected_win_data_160_port, 
                           curr_proc_regs(159) => 
                           DataPath_RF_bus_selected_win_data_159_port, 
                           curr_proc_regs(158) => 
                           DataPath_RF_bus_selected_win_data_158_port, 
                           curr_proc_regs(157) => 
                           DataPath_RF_bus_selected_win_data_157_port, 
                           curr_proc_regs(156) => 
                           DataPath_RF_bus_selected_win_data_156_port, 
                           curr_proc_regs(155) => 
                           DataPath_RF_bus_selected_win_data_155_port, 
                           curr_proc_regs(154) => 
                           DataPath_RF_bus_selected_win_data_154_port, 
                           curr_proc_regs(153) => 
                           DataPath_RF_bus_selected_win_data_153_port, 
                           curr_proc_regs(152) => 
                           DataPath_RF_bus_selected_win_data_152_port, 
                           curr_proc_regs(151) => 
                           DataPath_RF_bus_selected_win_data_151_port, 
                           curr_proc_regs(150) => 
                           DataPath_RF_bus_selected_win_data_150_port, 
                           curr_proc_regs(149) => 
                           DataPath_RF_bus_selected_win_data_149_port, 
                           curr_proc_regs(148) => 
                           DataPath_RF_bus_selected_win_data_148_port, 
                           curr_proc_regs(147) => 
                           DataPath_RF_bus_selected_win_data_147_port, 
                           curr_proc_regs(146) => 
                           DataPath_RF_bus_selected_win_data_146_port, 
                           curr_proc_regs(145) => 
                           DataPath_RF_bus_selected_win_data_145_port, 
                           curr_proc_regs(144) => 
                           DataPath_RF_bus_selected_win_data_144_port, 
                           curr_proc_regs(143) => 
                           DataPath_RF_bus_selected_win_data_143_port, 
                           curr_proc_regs(142) => 
                           DataPath_RF_bus_selected_win_data_142_port, 
                           curr_proc_regs(141) => 
                           DataPath_RF_bus_selected_win_data_141_port, 
                           curr_proc_regs(140) => 
                           DataPath_RF_bus_selected_win_data_140_port, 
                           curr_proc_regs(139) => 
                           DataPath_RF_bus_selected_win_data_139_port, 
                           curr_proc_regs(138) => 
                           DataPath_RF_bus_selected_win_data_138_port, 
                           curr_proc_regs(137) => 
                           DataPath_RF_bus_selected_win_data_137_port, 
                           curr_proc_regs(136) => 
                           DataPath_RF_bus_selected_win_data_136_port, 
                           curr_proc_regs(135) => 
                           DataPath_RF_bus_selected_win_data_135_port, 
                           curr_proc_regs(134) => 
                           DataPath_RF_bus_selected_win_data_134_port, 
                           curr_proc_regs(133) => 
                           DataPath_RF_bus_selected_win_data_133_port, 
                           curr_proc_regs(132) => 
                           DataPath_RF_bus_selected_win_data_132_port, 
                           curr_proc_regs(131) => 
                           DataPath_RF_bus_selected_win_data_131_port, 
                           curr_proc_regs(130) => 
                           DataPath_RF_bus_selected_win_data_130_port, 
                           curr_proc_regs(129) => 
                           DataPath_RF_bus_selected_win_data_129_port, 
                           curr_proc_regs(128) => 
                           DataPath_RF_bus_selected_win_data_128_port, 
                           curr_proc_regs(127) => 
                           DataPath_RF_bus_selected_win_data_127_port, 
                           curr_proc_regs(126) => 
                           DataPath_RF_bus_selected_win_data_126_port, 
                           curr_proc_regs(125) => 
                           DataPath_RF_bus_selected_win_data_125_port, 
                           curr_proc_regs(124) => 
                           DataPath_RF_bus_selected_win_data_124_port, 
                           curr_proc_regs(123) => 
                           DataPath_RF_bus_selected_win_data_123_port, 
                           curr_proc_regs(122) => 
                           DataPath_RF_bus_selected_win_data_122_port, 
                           curr_proc_regs(121) => 
                           DataPath_RF_bus_selected_win_data_121_port, 
                           curr_proc_regs(120) => 
                           DataPath_RF_bus_selected_win_data_120_port, 
                           curr_proc_regs(119) => 
                           DataPath_RF_bus_selected_win_data_119_port, 
                           curr_proc_regs(118) => 
                           DataPath_RF_bus_selected_win_data_118_port, 
                           curr_proc_regs(117) => 
                           DataPath_RF_bus_selected_win_data_117_port, 
                           curr_proc_regs(116) => 
                           DataPath_RF_bus_selected_win_data_116_port, 
                           curr_proc_regs(115) => 
                           DataPath_RF_bus_selected_win_data_115_port, 
                           curr_proc_regs(114) => 
                           DataPath_RF_bus_selected_win_data_114_port, 
                           curr_proc_regs(113) => 
                           DataPath_RF_bus_selected_win_data_113_port, 
                           curr_proc_regs(112) => 
                           DataPath_RF_bus_selected_win_data_112_port, 
                           curr_proc_regs(111) => 
                           DataPath_RF_bus_selected_win_data_111_port, 
                           curr_proc_regs(110) => 
                           DataPath_RF_bus_selected_win_data_110_port, 
                           curr_proc_regs(109) => 
                           DataPath_RF_bus_selected_win_data_109_port, 
                           curr_proc_regs(108) => 
                           DataPath_RF_bus_selected_win_data_108_port, 
                           curr_proc_regs(107) => 
                           DataPath_RF_bus_selected_win_data_107_port, 
                           curr_proc_regs(106) => 
                           DataPath_RF_bus_selected_win_data_106_port, 
                           curr_proc_regs(105) => 
                           DataPath_RF_bus_selected_win_data_105_port, 
                           curr_proc_regs(104) => 
                           DataPath_RF_bus_selected_win_data_104_port, 
                           curr_proc_regs(103) => 
                           DataPath_RF_bus_selected_win_data_103_port, 
                           curr_proc_regs(102) => 
                           DataPath_RF_bus_selected_win_data_102_port, 
                           curr_proc_regs(101) => 
                           DataPath_RF_bus_selected_win_data_101_port, 
                           curr_proc_regs(100) => 
                           DataPath_RF_bus_selected_win_data_100_port, 
                           curr_proc_regs(99) => 
                           DataPath_RF_bus_selected_win_data_99_port, 
                           curr_proc_regs(98) => 
                           DataPath_RF_bus_selected_win_data_98_port, 
                           curr_proc_regs(97) => 
                           DataPath_RF_bus_selected_win_data_97_port, 
                           curr_proc_regs(96) => 
                           DataPath_RF_bus_selected_win_data_96_port, 
                           curr_proc_regs(95) => 
                           DataPath_RF_bus_selected_win_data_95_port, 
                           curr_proc_regs(94) => 
                           DataPath_RF_bus_selected_win_data_94_port, 
                           curr_proc_regs(93) => 
                           DataPath_RF_bus_selected_win_data_93_port, 
                           curr_proc_regs(92) => 
                           DataPath_RF_bus_selected_win_data_92_port, 
                           curr_proc_regs(91) => 
                           DataPath_RF_bus_selected_win_data_91_port, 
                           curr_proc_regs(90) => 
                           DataPath_RF_bus_selected_win_data_90_port, 
                           curr_proc_regs(89) => 
                           DataPath_RF_bus_selected_win_data_89_port, 
                           curr_proc_regs(88) => 
                           DataPath_RF_bus_selected_win_data_88_port, 
                           curr_proc_regs(87) => 
                           DataPath_RF_bus_selected_win_data_87_port, 
                           curr_proc_regs(86) => 
                           DataPath_RF_bus_selected_win_data_86_port, 
                           curr_proc_regs(85) => 
                           DataPath_RF_bus_selected_win_data_85_port, 
                           curr_proc_regs(84) => 
                           DataPath_RF_bus_selected_win_data_84_port, 
                           curr_proc_regs(83) => 
                           DataPath_RF_bus_selected_win_data_83_port, 
                           curr_proc_regs(82) => 
                           DataPath_RF_bus_selected_win_data_82_port, 
                           curr_proc_regs(81) => 
                           DataPath_RF_bus_selected_win_data_81_port, 
                           curr_proc_regs(80) => 
                           DataPath_RF_bus_selected_win_data_80_port, 
                           curr_proc_regs(79) => 
                           DataPath_RF_bus_selected_win_data_79_port, 
                           curr_proc_regs(78) => 
                           DataPath_RF_bus_selected_win_data_78_port, 
                           curr_proc_regs(77) => 
                           DataPath_RF_bus_selected_win_data_77_port, 
                           curr_proc_regs(76) => 
                           DataPath_RF_bus_selected_win_data_76_port, 
                           curr_proc_regs(75) => 
                           DataPath_RF_bus_selected_win_data_75_port, 
                           curr_proc_regs(74) => 
                           DataPath_RF_bus_selected_win_data_74_port, 
                           curr_proc_regs(73) => 
                           DataPath_RF_bus_selected_win_data_73_port, 
                           curr_proc_regs(72) => 
                           DataPath_RF_bus_selected_win_data_72_port, 
                           curr_proc_regs(71) => 
                           DataPath_RF_bus_selected_win_data_71_port, 
                           curr_proc_regs(70) => 
                           DataPath_RF_bus_selected_win_data_70_port, 
                           curr_proc_regs(69) => 
                           DataPath_RF_bus_selected_win_data_69_port, 
                           curr_proc_regs(68) => 
                           DataPath_RF_bus_selected_win_data_68_port, 
                           curr_proc_regs(67) => 
                           DataPath_RF_bus_selected_win_data_67_port, 
                           curr_proc_regs(66) => 
                           DataPath_RF_bus_selected_win_data_66_port, 
                           curr_proc_regs(65) => 
                           DataPath_RF_bus_selected_win_data_65_port, 
                           curr_proc_regs(64) => 
                           DataPath_RF_bus_selected_win_data_64_port, 
                           curr_proc_regs(63) => 
                           DataPath_RF_bus_selected_win_data_63_port, 
                           curr_proc_regs(62) => 
                           DataPath_RF_bus_selected_win_data_62_port, 
                           curr_proc_regs(61) => 
                           DataPath_RF_bus_selected_win_data_61_port, 
                           curr_proc_regs(60) => 
                           DataPath_RF_bus_selected_win_data_60_port, 
                           curr_proc_regs(59) => 
                           DataPath_RF_bus_selected_win_data_59_port, 
                           curr_proc_regs(58) => 
                           DataPath_RF_bus_selected_win_data_58_port, 
                           curr_proc_regs(57) => 
                           DataPath_RF_bus_selected_win_data_57_port, 
                           curr_proc_regs(56) => 
                           DataPath_RF_bus_selected_win_data_56_port, 
                           curr_proc_regs(55) => 
                           DataPath_RF_bus_selected_win_data_55_port, 
                           curr_proc_regs(54) => 
                           DataPath_RF_bus_selected_win_data_54_port, 
                           curr_proc_regs(53) => 
                           DataPath_RF_bus_selected_win_data_53_port, 
                           curr_proc_regs(52) => 
                           DataPath_RF_bus_selected_win_data_52_port, 
                           curr_proc_regs(51) => 
                           DataPath_RF_bus_selected_win_data_51_port, 
                           curr_proc_regs(50) => 
                           DataPath_RF_bus_selected_win_data_50_port, 
                           curr_proc_regs(49) => 
                           DataPath_RF_bus_selected_win_data_49_port, 
                           curr_proc_regs(48) => 
                           DataPath_RF_bus_selected_win_data_48_port, 
                           curr_proc_regs(47) => 
                           DataPath_RF_bus_selected_win_data_47_port, 
                           curr_proc_regs(46) => 
                           DataPath_RF_bus_selected_win_data_46_port, 
                           curr_proc_regs(45) => 
                           DataPath_RF_bus_selected_win_data_45_port, 
                           curr_proc_regs(44) => 
                           DataPath_RF_bus_selected_win_data_44_port, 
                           curr_proc_regs(43) => 
                           DataPath_RF_bus_selected_win_data_43_port, 
                           curr_proc_regs(42) => 
                           DataPath_RF_bus_selected_win_data_42_port, 
                           curr_proc_regs(41) => 
                           DataPath_RF_bus_selected_win_data_41_port, 
                           curr_proc_regs(40) => 
                           DataPath_RF_bus_selected_win_data_40_port, 
                           curr_proc_regs(39) => 
                           DataPath_RF_bus_selected_win_data_39_port, 
                           curr_proc_regs(38) => 
                           DataPath_RF_bus_selected_win_data_38_port, 
                           curr_proc_regs(37) => 
                           DataPath_RF_bus_selected_win_data_37_port, 
                           curr_proc_regs(36) => 
                           DataPath_RF_bus_selected_win_data_36_port, 
                           curr_proc_regs(35) => 
                           DataPath_RF_bus_selected_win_data_35_port, 
                           curr_proc_regs(34) => 
                           DataPath_RF_bus_selected_win_data_34_port, 
                           curr_proc_regs(33) => 
                           DataPath_RF_bus_selected_win_data_33_port, 
                           curr_proc_regs(32) => 
                           DataPath_RF_bus_selected_win_data_32_port, 
                           curr_proc_regs(31) => 
                           DataPath_RF_bus_selected_win_data_31_port, 
                           curr_proc_regs(30) => 
                           DataPath_RF_bus_selected_win_data_30_port, 
                           curr_proc_regs(29) => 
                           DataPath_RF_bus_selected_win_data_29_port, 
                           curr_proc_regs(28) => 
                           DataPath_RF_bus_selected_win_data_28_port, 
                           curr_proc_regs(27) => 
                           DataPath_RF_bus_selected_win_data_27_port, 
                           curr_proc_regs(26) => 
                           DataPath_RF_bus_selected_win_data_26_port, 
                           curr_proc_regs(25) => 
                           DataPath_RF_bus_selected_win_data_25_port, 
                           curr_proc_regs(24) => 
                           DataPath_RF_bus_selected_win_data_24_port, 
                           curr_proc_regs(23) => 
                           DataPath_RF_bus_selected_win_data_23_port, 
                           curr_proc_regs(22) => 
                           DataPath_RF_bus_selected_win_data_22_port, 
                           curr_proc_regs(21) => 
                           DataPath_RF_bus_selected_win_data_21_port, 
                           curr_proc_regs(20) => 
                           DataPath_RF_bus_selected_win_data_20_port, 
                           curr_proc_regs(19) => 
                           DataPath_RF_bus_selected_win_data_19_port, 
                           curr_proc_regs(18) => 
                           DataPath_RF_bus_selected_win_data_18_port, 
                           curr_proc_regs(17) => 
                           DataPath_RF_bus_selected_win_data_17_port, 
                           curr_proc_regs(16) => 
                           DataPath_RF_bus_selected_win_data_16_port, 
                           curr_proc_regs(15) => 
                           DataPath_RF_bus_selected_win_data_15_port, 
                           curr_proc_regs(14) => 
                           DataPath_RF_bus_selected_win_data_14_port, 
                           curr_proc_regs(13) => 
                           DataPath_RF_bus_selected_win_data_13_port, 
                           curr_proc_regs(12) => 
                           DataPath_RF_bus_selected_win_data_12_port, 
                           curr_proc_regs(11) => 
                           DataPath_RF_bus_selected_win_data_11_port, 
                           curr_proc_regs(10) => 
                           DataPath_RF_bus_selected_win_data_10_port, 
                           curr_proc_regs(9) => 
                           DataPath_RF_bus_selected_win_data_9_port, 
                           curr_proc_regs(8) => 
                           DataPath_RF_bus_selected_win_data_8_port, 
                           curr_proc_regs(7) => 
                           DataPath_RF_bus_selected_win_data_7_port, 
                           curr_proc_regs(6) => 
                           DataPath_RF_bus_selected_win_data_6_port, 
                           curr_proc_regs(5) => 
                           DataPath_RF_bus_selected_win_data_5_port, 
                           curr_proc_regs(4) => 
                           DataPath_RF_bus_selected_win_data_4_port, 
                           curr_proc_regs(3) => 
                           DataPath_RF_bus_selected_win_data_3_port, 
                           curr_proc_regs(2) => 
                           DataPath_RF_bus_selected_win_data_2_port, 
                           curr_proc_regs(1) => 
                           DataPath_RF_bus_selected_win_data_1_port, 
                           curr_proc_regs(0) => 
                           DataPath_RF_bus_selected_win_data_0_port);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_6_inst : DFF_X1 port map( D => 
                           n7159, CK => CLK, Q => DECODEhw_i_tickcounter_6_port
                           , QN => n_1065);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_8_inst : DFF_X1 port map( D => 
                           n7157, CK => CLK, Q => DECODEhw_i_tickcounter_8_port
                           , QN => n_1066);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_10_inst : DFF_X1 port map( D => 
                           n7155, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_10_port, QN => n_1067);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_12_inst : DFF_X1 port map( D => 
                           n7153, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_12_port, QN => n8265);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_13_inst : DFF_X1 port map( D => 
                           n7152, CK => CLK, Q => n_1068, QN => n554);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_14_inst : DFF_X1 port map( D => 
                           n7151, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_14_port, QN => n_1069);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_15_inst : DFF_X1 port map( D => 
                           n7150, CK => CLK, Q => n_1070, QN => n556);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_16_inst : DFF_X1 port map( D => 
                           n7149, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_16_port, QN => n_1071);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_17_inst : DFF_X1 port map( D => 
                           n7148, CK => CLK, Q => n_1072, QN => n558);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_18_inst : DFF_X1 port map( D => 
                           n7147, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_18_port, QN => n_1073);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_19_inst : DFF_X1 port map( D => 
                           n7146, CK => CLK, Q => n_1074, QN => n560);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_20_inst : DFF_X1 port map( D => 
                           n7145, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_20_port, QN => n_1075);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_21_inst : DFF_X1 port map( D => 
                           n7144, CK => CLK, Q => n_1076, QN => n562);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_22_inst : DFF_X1 port map( D => 
                           n7143, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_22_port, QN => n_1077);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_23_inst : DFF_X1 port map( D => 
                           n7142, CK => CLK, Q => n_1078, QN => n564);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_24_inst : DFF_X1 port map( D => 
                           n7141, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_24_port, QN => n_1079);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_25_inst : DFF_X1 port map( D => 
                           n7140, CK => CLK, Q => n_1080, QN => n566);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_26_inst : DFF_X1 port map( D => 
                           n7139, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_26_port, QN => n_1081);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_27_inst : DFF_X1 port map( D => 
                           n7138, CK => CLK, Q => n_1082, QN => n568);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_28_inst : DFF_X1 port map( D => 
                           n7137, CK => CLK, Q => n_1083, QN => n569);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_29_inst : DFF_X1 port map( D => 
                           n3160, CK => CLK, Q => n_1084, QN => 
                           DECODEhw_i_tickcounter_29_port);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_30_inst : DFF_X1 port map( D => 
                           n7136, CK => CLK, Q => n_1085, QN => n570);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_31_inst : DFF_X1 port map( D => 
                           n7166, CK => CLK, Q => 
                           DECODEhw_i_tickcounter_31_port, QN => n_1086);
   DataPath_RF_BLOCKi_72_Q_reg_0_inst : DFF_X1 port map( D => n5788, CK => CLK,
                           Q => n_1087, QN => 
                           DataPath_RF_bus_reg_dataout_2048_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_31_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N35, Q => i_RD2_31_port
                           );
   DataPath_REG_B_Q_reg_31_inst : DFF_X1 port map( D => n2732, CK => CLK, Q => 
                           n8297, QN => DataPath_i_PIPLIN_B_31_port);
   DataPath_REG_ME_Q_reg_31_inst : DFF_X1 port map( D => n2700, CK => CLK, Q =>
                           n_1088, QN => DataPath_i_REG_ME_DATA_DATAMEM_31_port
                           );
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_7_inst : DFF_X1 port map( D => n2202, CK =>
                           CLK, Q => n_1089, QN => 
                           DataPath_i_REG_LDSTR_OUT_7_port);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_31_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N35, Q => i_RD1_31_port
                           );
   IR_reg_25_inst : DFFR_X1 port map( D => n7124, CK => CLK, RN => n8582, Q => 
                           n8305, QN => n169);
   IR_reg_23_inst : DFFR_X1 port map( D => n7125, CK => CLK, RN => n8571, Q => 
                           n_1090, QN => n170);
   IR_reg_20_inst : DFFR_X1 port map( D => n7127, CK => CLK, RN => n8578, Q => 
                           n_1091, QN => n172);
   IR_reg_19_inst : DFFR_X1 port map( D => n7128, CK => CLK, RN => n8574, Q => 
                           n_1092, QN => n173);
   IR_reg_18_inst : DFFR_X1 port map( D => n7129, CK => CLK, RN => n8580, Q => 
                           n8287, QN => n174);
   IR_reg_17_inst : DFFR_X1 port map( D => n7130, CK => CLK, RN => n8577, Q => 
                           n_1093, QN => n175);
   IR_reg_16_inst : DFFR_X1 port map( D => n7131, CK => CLK, RN => n8576, Q => 
                           n_1094, QN => n176);
   IR_reg_15_inst : DFFR_X1 port map( D => n7132, CK => CLK, RN => n8570, Q => 
                           n8210, QN => n177);
   IR_reg_14_inst : DFFR_X1 port map( D => n7133, CK => CLK, RN => n8570, Q => 
                           n8282, QN => n178);
   IR_reg_9_inst : DFFR_X1 port map( D => n7134, CK => CLK, RN => n8570, Q => 
                           IR_9_port, QN => n8241);
   IR_reg_8_inst : DFFR_X1 port map( D => n7135, CK => CLK, RN => n8570, Q => 
                           IR_8_port, QN => n8238);
   IR_reg_0_inst : DFFR_X1 port map( D => n34, CK => CLK, RN => n8570, Q => 
                           n8309, QN => n193);
   IR_reg_2_inst : DFFR_X1 port map( D => n36, CK => CLK, RN => n8570, Q => 
                           IR_2_port, QN => n8224);
   IR_reg_3_inst : DFFR_X1 port map( D => n37, CK => CLK, RN => n8570, Q => 
                           IR_3_port, QN => n8226);
   IR_reg_4_inst : DFFR_X1 port map( D => n38, CK => CLK, RN => n8570, Q => 
                           IR_4_port, QN => n8190);
   IR_reg_5_inst : DFFR_X1 port map( D => n39, CK => CLK, RN => n8570, Q => 
                           IR_5_port, QN => n8198);
   IR_reg_7_inst : DFFR_X1 port map( D => n41, CK => CLK, RN => n8571, Q => 
                           IR_7_port, QN => n8234);
   IR_reg_10_inst : DFFS_X1 port map( D => n2886, CK => CLK, SN => n8572, Q => 
                           n8233, QN => IR_10_port);
   IR_reg_11_inst : DFFR_X1 port map( D => n42, CK => CLK, RN => n8571, Q => 
                           n8280, QN => n180);
   IR_reg_12_inst : DFFR_X1 port map( D => n43, CK => CLK, RN => n8582, Q => 
                           n8196, QN => n179);
   IR_reg_13_inst : DFFS_X1 port map( D => n2883, CK => CLK, SN => n8570, Q => 
                           n8199, QN => IR_13_port);
   IR_reg_21_inst : DFFS_X1 port map( D => n2878, CK => CLK, SN => n8580, Q => 
                           n8232, QN => IR_21_port);
   IR_reg_24_inst : DFFS_X1 port map( D => n2875, CK => CLK, SN => n8573, Q => 
                           n8231, QN => IR_24_port);
   IR_reg_28_inst : DFFS_X1 port map( D => n7121, CK => CLK, SN => n8571, Q => 
                           n8195, QN => n163);
   DataPath_WRB1_Q_reg_0_inst : DFF_X1 port map( D => n2865, CK => CLK, Q => 
                           n_1095, QN => DataPath_i_PIPLIN_WRB1_0_port);
   DataPath_WRB2_Q_reg_0_inst : DFF_X1 port map( D => n2766, CK => CLK, Q => 
                           n_1096, QN => DataPath_i_PIPLIN_WRB2_0_port);
   DataPath_WRB3_Q_reg_0_inst : DFF_X1 port map( D => n355, CK => CLK, Q => 
                           i_ADD_WB_0_port, QN => n523);
   CU_I_CW_ID_reg_MEM_EN_inst : DLL_X1 port map( D => CU_I_CW_IF_MEM_EN_port, 
                           GN => n2867, Q => CU_I_CW_ID_MEM_EN_port);
   CU_I_CW_EX_reg_MEM_EN_inst : DFF_X1 port map( D => n365, CK => CLK, Q => 
                           CU_I_CW_EX_MEM_EN_port, QN => n_1097);
   CU_I_CW_MEM_reg_MEM_EN_inst : DFF_X1 port map( D => n7099, CK => CLK, Q => 
                           CU_I_CW_MEM_MEM_EN_port, QN => n_1098);
   CU_I_aluOpcode1_reg_0_inst : DFF_X1 port map( D => n7095, CK => CLK, Q => 
                           i_ALU_OP_0_port, QN => n8292);
   CU_I_setcmp_1_reg_1_inst : DFF_X1 port map( D => n7089, CK => CLK, Q => 
                           i_SEL_LGET_1_port, QN => n8283);
   CU_I_i_FILL_delay_reg : DFF_X1 port map( D => CU_I_N317, CK => CLK, Q => 
                           CU_I_i_FILL_delay, QN => n_1099);
   DataPath_RF_PUSH_ADDRGEN_curr_state_reg_0_inst : DFF_X1 port map( D => n7069
                           , CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_state_0_port, QN => 
                           n_1100);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_1_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N47, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, QN => 
                           n_1101);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_2_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N48, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, QN => 
                           n_1102);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_3_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N49, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, QN => 
                           n_1103);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_4_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N50, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, QN => 
                           n_1104);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_5_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N51, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, QN => 
                           n_1105);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_6_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N52, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, QN => 
                           n_1106);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_7_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N53, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, QN => 
                           n_1107);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_8_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N54, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, QN => 
                           n_1108);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_9_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N55, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, QN => 
                           n_1109);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_10_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N56, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, QN => 
                           n_1110);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_11_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N57, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, QN => 
                           n_1111);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_12_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N58, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, QN => 
                           n_1112);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_13_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N59, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, QN => 
                           n_1113);
   DataPath_RF_POP_ADDRGEN_curr_state_reg_1_inst : DFF_X1 port map( D => n7062,
                           CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_state_1_port, QN => 
                           n_1114);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_1_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N47, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_1_port, QN => 
                           n_1115);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_2_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N48, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_2_port, QN => 
                           n_1116);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_3_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N49, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_3_port, QN => 
                           n_1117);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_4_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N50, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_4_port, QN => 
                           n_1118);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_5_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N51, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_5_port, QN => 
                           n_1119);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_6_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N52, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_6_port, QN => 
                           n_1120);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_7_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N53, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_7_port, QN => 
                           n_1121);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_9_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N55, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_9_port, QN => 
                           n_1122);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_10_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N56, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_10_port, QN => 
                           n_1123);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_11_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N57, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_11_port, QN => 
                           n_1124);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_12_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N58, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_12_port, QN => 
                           n_1125);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_13_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N59, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_13_port, QN => 
                           n_1126);
   CU_I_CW_ID_reg_RF_RD1_EN_inst : DLL_X1 port map( D => CU_I_CW_RF_RD1_EN_port
                           , GN => n2867, Q => i_RF1);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_0_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N4, Q => i_RD1_0_port);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_1_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N5, Q => i_RD1_1_port);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_2_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N6, Q => i_RD1_2_port);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_3_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N7, Q => i_RD1_3_port);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_4_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N8, Q => i_RD1_4_port);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_5_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N9, Q => i_RD1_5_port);
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_6_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N10, Q => i_RD1_6_port)
                           ;
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_7_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N11, Q => i_RD1_7_port)
                           ;
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_8_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N12, Q => i_RD1_8_port)
                           ;
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_9_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N13, Q => i_RD1_9_port)
                           ;
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_10_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N14, Q => i_RD1_10_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_11_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N15, Q => i_RD1_11_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_12_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N16, Q => i_RD1_12_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_13_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N17, Q => i_RD1_13_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_14_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N18, Q => i_RD1_14_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_15_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N19, Q => i_RD1_15_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_16_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N20, Q => i_RD1_16_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_17_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N21, Q => i_RD1_17_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_18_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N22, Q => i_RD1_18_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_19_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N23, Q => i_RD1_19_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_20_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N24, Q => i_RD1_20_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_21_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N25, Q => i_RD1_21_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_22_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N26, Q => i_RD1_22_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_23_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N27, Q => i_RD1_23_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_24_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N28, Q => i_RD1_24_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_25_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N29, Q => i_RD1_25_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_26_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N30, Q => i_RD1_26_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_27_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N31, Q => i_RD1_27_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_28_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N32, Q => i_RD1_28_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_29_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N33, Q => i_RD1_29_port
                           );
   DataPath_RF_RDPORT0_OUTLATCH_q_mem_reg_30_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT0_OUTLATCH_N34, Q => i_RD1_30_port
                           );
   CU_I_CW_ID_reg_RF_RD2_EN_inst : DLL_X1 port map( D => CU_I_CW_RF_RD2_EN_port
                           , GN => n8458, Q => i_RF2);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_0_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N4, Q => i_RD2_0_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_1_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N5, Q => i_RD2_1_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_2_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N6, Q => i_RD2_2_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_3_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N7, Q => i_RD2_3_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_4_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N8, Q => i_RD2_4_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_5_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N9, Q => i_RD2_5_port);
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_6_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N10, Q => i_RD2_6_port)
                           ;
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_7_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N11, Q => i_RD2_7_port)
                           ;
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_8_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N12, Q => i_RD2_8_port)
                           ;
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_9_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N13, Q => i_RD2_9_port)
                           ;
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_10_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N14, Q => i_RD2_10_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_11_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N15, Q => i_RD2_11_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_12_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N16, Q => i_RD2_12_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_13_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N17, Q => i_RD2_13_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_14_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N18, Q => i_RD2_14_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_15_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N19, Q => i_RD2_15_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_16_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N20, Q => i_RD2_16_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_17_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N21, Q => i_RD2_17_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_18_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N22, Q => i_RD2_18_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_19_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N23, Q => i_RD2_19_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_20_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N24, Q => i_RD2_20_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_21_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N25, Q => i_RD2_21_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_22_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N26, Q => i_RD2_22_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_23_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N27, Q => i_RD2_23_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_24_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N28, Q => i_RD2_24_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_25_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N29, Q => i_RD2_25_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_26_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N30, Q => i_RD2_26_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_27_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N31, Q => i_RD2_27_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_28_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N32, Q => i_RD2_28_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_29_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N33, Q => i_RD2_29_port
                           );
   DataPath_RF_RDPORT1_OUTLATCH_q_mem_reg_30_inst : DLH_X1 port map( G => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3, D => 
                           DataPath_RF_RDPORT1_OUTLATCH_N34, Q => i_RD2_30_port
                           );
   CU_I_CW_ID_reg_SEL_CMPB_inst : DLL_X1 port map( D => CU_I_CW_SEL_CMPB_port, 
                           GN => n8458, Q => i_SEL_CMPB);
   CU_I_CW_ID_reg_UNSIGNED_ID_inst : DLL_X1 port map( D => 
                           CU_I_CW_UNSIGNED_ID_port, GN => n8458, Q => 
                           CU_I_CW_ID_UNSIGNED_ID_port);
   CU_I_CW_ID_reg_NPC_SEL_inst : DLL_X1 port map( D => CU_I_CW_NPC_SEL_port, GN
                           => n2867, Q => i_NPC_SEL);
   PC_reg_0_inst : DFFR_X1 port map( D => n7061, CK => CLK, RN => n8571, Q => 
                           IRAM_ADDRESS_0_port, QN => n211);
   PC_reg_1_inst : DFFR_X1 port map( D => n7060, CK => CLK, RN => n8571, Q => 
                           IRAM_ADDRESS_1_port, QN => n_1127);
   PC_reg_2_inst : DFFR_X1 port map( D => n7059, CK => CLK, RN => n8571, Q => 
                           IRAM_ADDRESS_2_port, QN => n_1128);
   PC_reg_3_inst : DFFR_X1 port map( D => n7058, CK => CLK, RN => n8571, Q => 
                           IRAM_ADDRESS_3_port, QN => n8321);
   PC_reg_5_inst : DFFR_X1 port map( D => n7056, CK => CLK, RN => n8570, Q => 
                           IRAM_ADDRESS_5_port, QN => n207);
   PC_reg_6_inst : DFFR_X1 port map( D => n7055, CK => CLK, RN => n8578, Q => 
                           IRAM_ADDRESS_6_port, QN => n8307);
   PC_reg_7_inst : DFFR_X1 port map( D => n7054, CK => CLK, RN => n8579, Q => 
                           IRAM_ADDRESS_7_port, QN => n8284);
   PC_reg_8_inst : DFFR_X1 port map( D => n7053, CK => CLK, RN => n8572, Q => 
                           IRAM_ADDRESS_8_port, QN => n206);
   PC_reg_9_inst : DFFR_X1 port map( D => n7052, CK => CLK, RN => n8577, Q => 
                           IRAM_ADDRESS_9_port, QN => n205);
   PC_reg_12_inst : DFFR_X1 port map( D => n7049, CK => CLK, RN => n8571, Q => 
                           IRAM_ADDRESS_12_port, QN => n8311);
   PC_reg_13_inst : DFFR_X1 port map( D => n7048, CK => CLK, RN => n8576, Q => 
                           IRAM_ADDRESS_13_port, QN => n8290);
   PC_reg_14_inst : DFFR_X1 port map( D => n7047, CK => CLK, RN => n8577, Q => 
                           IRAM_ADDRESS_14_port, QN => n8279);
   PC_reg_15_inst : DFFR_X1 port map( D => n7046, CK => CLK, RN => n8570, Q => 
                           IRAM_ADDRESS_15_port, QN => n8300);
   PC_reg_16_inst : DFFR_X1 port map( D => n7045, CK => CLK, RN => n8571, Q => 
                           IRAM_ADDRESS_16_port, QN => n_1129);
   PC_reg_17_inst : DFFR_X1 port map( D => n7044, CK => CLK, RN => n8574, Q => 
                           IRAM_ADDRESS_17_port, QN => n_1130);
   PC_reg_18_inst : DFFR_X1 port map( D => n7043, CK => CLK, RN => n8573, Q => 
                           IRAM_ADDRESS_18_port, QN => n8322);
   PC_reg_19_inst : DFFR_X1 port map( D => n7042, CK => CLK, RN => n8578, Q => 
                           IRAM_ADDRESS_19_port, QN => n_1131);
   PC_reg_20_inst : DFFR_X1 port map( D => n7041, CK => CLK, RN => n8573, Q => 
                           IRAM_ADDRESS_20_port, QN => n_1132);
   PC_reg_21_inst : DFFR_X1 port map( D => n7040, CK => CLK, RN => n8575, Q => 
                           IRAM_ADDRESS_21_port, QN => n8275);
   PC_reg_22_inst : DFFR_X1 port map( D => n7039, CK => CLK, RN => n8571, Q => 
                           IRAM_ADDRESS_22_port, QN => n8274);
   PC_reg_24_inst : DFFR_X1 port map( D => n7037, CK => CLK, RN => n8577, Q => 
                           IRAM_ADDRESS_24_port, QN => n7611);
   PC_reg_25_inst : DFFR_X1 port map( D => n7036, CK => CLK, RN => n8571, Q => 
                           IRAM_ADDRESS_25_port, QN => n_1133);
   PC_reg_26_inst : DFFR_X1 port map( D => n7035, CK => CLK, RN => n8571, Q => 
                           IRAM_ADDRESS_26_port, QN => n8323);
   PC_reg_27_inst : DFFR_X1 port map( D => n7034, CK => CLK, RN => n8573, Q => 
                           IRAM_ADDRESS_27_port, QN => n_1134);
   CU_I_CW_ID_reg_HAZARD_TABLE_WR1_inst : DLL_X1 port map( D => n6692, GN => 
                           n8458, Q => n461);
   CU_I_CW_ID_reg_MUXA_SEL_inst : DLL_X1 port map( D => CU_I_CW_MUXA_SEL_port, 
                           GN => n8458, Q => CU_I_CW_ID_MUXA_SEL_port);
   CU_I_CW_EX_reg_MUXA_SEL_inst : DFF_X1 port map( D => n7085, CK => CLK, Q => 
                           n8225, QN => n460);
   CU_I_CW_ID_reg_MUXB_SEL_inst : DLL_X1 port map( D => CU_I_CW_MUXB_SEL_port, 
                           GN => n2867, Q => CU_I_CW_ID_MUXB_SEL_port);
   CU_I_CW_ID_reg_DRAM_WE_inst : DLL_X1 port map( D => n143, GN => n8458, Q => 
                           CU_I_CW_ID_DRAM_WE_port);
   CU_I_CW_EX_reg_DRAM_WE_inst : DFF_X1 port map( D => n364, CK => CLK, Q => 
                           CU_I_CW_EX_DRAM_WE_port, QN => n_1135);
   CU_I_CW_MEM_reg_DRAM_WE_inst : DFF_X1 port map( D => n7118, CK => CLK, Q => 
                           i_DATAMEM_WM, QN => DRAM_READNOTWRITE);
   CU_I_CW_ID_reg_DRAM_RE_inst : DLL_X1 port map( D => CU_I_CW_WB_MUX_SEL_port,
                           GN => n8458, Q => CU_I_CW_ID_DRAM_RE_port);
   CU_I_CW_EX_reg_DRAM_RE_inst : DFF_X1 port map( D => n368, CK => CLK, Q => 
                           CU_I_CW_EX_DRAM_RE_port, QN => n_1136);
   CU_I_CW_ID_reg_DATA_SIZE_1_inst : DLL_X1 port map( D => 
                           CU_I_CW_DATA_SIZE_1_port, GN => n2867, Q => 
                           CU_I_CW_ID_DATA_SIZE_1_port);
   CU_I_CW_EX_reg_DATA_SIZE_1_inst : DFF_X1 port map( D => n367, CK => CLK, Q 
                           => CU_I_CW_EX_DATA_SIZE_1_port, QN => n_1137);
   CU_I_CW_MEM_reg_DATA_SIZE_1_inst : DFF_X1 port map( D => n7097, CK => CLK, Q
                           => DATA_SIZE_1_port, QN => n376);
   CU_I_CW_ID_reg_DATA_SIZE_0_inst : DLL_X1 port map( D => 
                           CU_I_CW_DATA_SIZE_0_port, GN => n8458, Q => 
                           CU_I_CW_ID_DATA_SIZE_0_port);
   CU_I_CW_EX_reg_DATA_SIZE_0_inst : DFF_X1 port map( D => n366, CK => CLK, Q 
                           => CU_I_CW_EX_DATA_SIZE_0_port, QN => n_1138);
   CU_I_CW_MEM_reg_DATA_SIZE_0_inst : DFF_X1 port map( D => n7098, CK => CLK, Q
                           => DATA_SIZE_0_port, QN => n375);
   CU_I_CW_ID_reg_WB_MUX_SEL_inst : DLL_X1 port map( D => 
                           CU_I_CW_WB_MUX_SEL_port, GN => n8458, Q => 
                           CU_I_CW_ID_WB_MUX_SEL_port);
   CU_I_CW_WB_reg_WB_MUX_SEL_inst : DFF_X1 port map( D => CU_I_N305, CK => CLK,
                           Q => i_S3, QN => n_1139);
   CU_I_CW_ID_reg_WB_EN_inst : DLL_X1 port map( D => CU_I_CW_IF_WB_EN_port, GN 
                           => n8458, Q => CU_I_CW_ID_WB_EN_port);
   CU_I_CW_WB_reg_WB_EN_inst : DFF_X1 port map( D => CU_I_N304, CK => CLK, Q =>
                           i_WF, QN => n8306);
   CU_I_CW_ID_reg_EX_EN_inst : DLL_X1 port map( D => CU_I_CW_IF_MEM_EN_port, GN
                           => n8458, Q => CU_I_CW_ID_EX_EN_port);
   CU_I_CW_EX_reg_EX_EN_inst : DFF_X1 port map( D => n2767, CK => CLK, Q => 
                           n8301, QN => CU_I_CW_EX_EX_EN_port);
   CU_I_CW_ID_reg_ID_EN_inst : DLL_X1 port map( D => CU_I_CW_IF_MEM_EN_port, GN
                           => n8458, Q => CU_I_CW_ID_ID_EN_port);
   DataPath_REG_IN2_Q_reg_20_inst : DFF_X1 port map( D => n7021, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_20_port, QN => n_1140);
   DataPath_REG_IN2_Q_reg_14_inst : DFF_X1 port map( D => n7022, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_14_port, QN => n_1141);
   DataPath_REG_IN2_Q_reg_13_inst : DFF_X1 port map( D => n7023, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_13_port, QN => n8316);
   DataPath_REG_IN2_Q_reg_12_inst : DFF_X1 port map( D => n7024, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_12_port, QN => n8326);
   DataPath_REG_IN2_Q_reg_10_inst : DFF_X1 port map( D => n7025, CK => CLK, Q 
                           => DataPath_i_PIPLIN_IN2_10_port, QN => n8315);
   DataPath_REG_IN2_Q_reg_4_inst : DFF_X1 port map( D => n7027, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_4_port, QN => n_1142);
   DataPath_REG_IN2_Q_reg_3_inst : DFF_X1 port map( D => n7028, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_3_port, QN => n_1143);
   DataPath_REG_IN2_Q_reg_1_inst : DFF_X1 port map( D => n7029, CK => CLK, Q =>
                           DataPath_i_PIPLIN_IN2_1_port, QN => n_1144);
   DataPath_REG_B_Q_reg_20_inst : DFF_X1 port map( D => n7075, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_20_port, QN => n_1145);
   DataPath_REG_ME_Q_reg_20_inst : DFF_X1 port map( D => n2711, CK => CLK, Q =>
                           n_1146, QN => DataPath_i_REG_ME_DATA_DATAMEM_20_port
                           );
   DataPath_REG_B_Q_reg_14_inst : DFF_X1 port map( D => n7076, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_14_port, QN => n_1147);
   DataPath_REG_ME_Q_reg_14_inst : DFF_X1 port map( D => n2717, CK => CLK, Q =>
                           n_1148, QN => DataPath_i_REG_ME_DATA_DATAMEM_14_port
                           );
   DataPath_REG_ME_Q_reg_13_inst : DFF_X1 port map( D => n2718, CK => CLK, Q =>
                           n_1149, QN => DataPath_i_REG_ME_DATA_DATAMEM_13_port
                           );
   DataPath_REG_B_Q_reg_12_inst : DFF_X1 port map( D => n7078, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_12_port, QN => n_1150);
   DataPath_REG_ME_Q_reg_12_inst : DFF_X1 port map( D => n2719, CK => CLK, Q =>
                           n_1151, QN => DataPath_i_REG_ME_DATA_DATAMEM_12_port
                           );
   DataPath_REG_B_Q_reg_10_inst : DFF_X1 port map( D => n7079, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_10_port, QN => n_1152);
   DataPath_REG_ME_Q_reg_10_inst : DFF_X1 port map( D => n2721, CK => CLK, Q =>
                           n_1153, QN => DataPath_i_REG_ME_DATA_DATAMEM_10_port
                           );
   DataPath_REG_ME_Q_reg_6_inst : DFF_X1 port map( D => n2725, CK => CLK, Q => 
                           n_1154, QN => DataPath_i_REG_ME_DATA_DATAMEM_6_port)
                           ;
   DataPath_REG_B_Q_reg_4_inst : DFF_X1 port map( D => n7081, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_4_port, QN => n_1155);
   DataPath_REG_ME_Q_reg_4_inst : DFF_X1 port map( D => n2727, CK => CLK, Q => 
                           n_1156, QN => DataPath_i_REG_ME_DATA_DATAMEM_4_port)
                           ;
   DataPath_REG_B_Q_reg_3_inst : DFF_X1 port map( D => n7082, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_3_port, QN => n_1157);
   DataPath_REG_ME_Q_reg_3_inst : DFF_X1 port map( D => n2728, CK => CLK, Q => 
                           n_1158, QN => DataPath_i_REG_ME_DATA_DATAMEM_3_port)
                           ;
   DataPath_REG_CMP_Q_reg_1_inst : DFF_X1 port map( D => n7116, CK => CLK, Q =>
                           n_1159, QN => n493);
   DataPath_REG_CMP_Q_reg_0_inst : DFF_X1 port map( D => n7117, CK => CLK, Q =>
                           n8319, QN => n492);
   DataPath_REG_A_Q_reg_20_inst : DFF_X1 port map( D => n6728, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_20_port, QN => n_1160);
   DataPath_REG_A_Q_reg_14_inst : DFF_X1 port map( D => n6729, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_14_port, QN => n_1161);
   DataPath_REG_A_Q_reg_13_inst : DFF_X1 port map( D => n6730, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_13_port, QN => n_1162);
   DataPath_REG_A_Q_reg_12_inst : DFF_X1 port map( D => n6731, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_12_port, QN => n7692);
   DataPath_REG_A_Q_reg_10_inst : DFF_X1 port map( D => n6732, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_10_port, QN => n_1163);
   DataPath_REG_A_Q_reg_8_inst : DFF_X1 port map( D => n6733, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_8_port, QN => n_1164);
   DataPath_REG_A_Q_reg_3_inst : DFF_X1 port map( D => n6734, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_3_port, QN => n_1165);
   DataPath_REG_A_Q_reg_1_inst : DFF_X1 port map( D => n6735, CK => CLK, Q => 
                           DataPath_i_PIPLIN_A_1_port, QN => n_1166);
   DataPath_REG_A_Q_reg_0_inst : DFF_X1 port map( D => n3261, CK => CLK, Q => 
                           n_1167, QN => DataPath_i_PIPLIN_A_0_port);
   DataPath_REG_A_Q_reg_2_inst : DFF_X1 port map( D => n3260, CK => CLK, Q => 
                           n_1168, QN => DataPath_i_PIPLIN_A_2_port);
   DataPath_REG_A_Q_reg_4_inst : DFF_X1 port map( D => n3259, CK => CLK, Q => 
                           n_1169, QN => DataPath_i_PIPLIN_A_4_port);
   DataPath_REG_A_Q_reg_5_inst : DFF_X1 port map( D => n3258, CK => CLK, Q => 
                           n_1170, QN => DataPath_i_PIPLIN_A_5_port);
   DataPath_REG_A_Q_reg_6_inst : DFF_X1 port map( D => n3257, CK => CLK, Q => 
                           n_1171, QN => DataPath_i_PIPLIN_A_6_port);
   DataPath_REG_A_Q_reg_7_inst : DFF_X1 port map( D => n3256, CK => CLK, Q => 
                           n_1172, QN => DataPath_i_PIPLIN_A_7_port);
   DataPath_REG_A_Q_reg_9_inst : DFF_X1 port map( D => n3255, CK => CLK, Q => 
                           n_1173, QN => DataPath_i_PIPLIN_A_9_port);
   DataPath_REG_A_Q_reg_11_inst : DFF_X1 port map( D => n3254, CK => CLK, Q => 
                           n_1174, QN => DataPath_i_PIPLIN_A_11_port);
   DataPath_REG_A_Q_reg_15_inst : DFF_X1 port map( D => n3253, CK => CLK, Q => 
                           n_1175, QN => DataPath_i_PIPLIN_A_15_port);
   DataPath_REG_A_Q_reg_16_inst : DFF_X1 port map( D => n3252, CK => CLK, Q => 
                           n_1176, QN => DataPath_i_PIPLIN_A_16_port);
   DataPath_REG_A_Q_reg_17_inst : DFF_X1 port map( D => n3251, CK => CLK, Q => 
                           n_1177, QN => DataPath_i_PIPLIN_A_17_port);
   DataPath_REG_A_Q_reg_18_inst : DFF_X1 port map( D => n3250, CK => CLK, Q => 
                           n_1178, QN => DataPath_i_PIPLIN_A_18_port);
   DataPath_REG_A_Q_reg_19_inst : DFF_X1 port map( D => n3249, CK => CLK, Q => 
                           n_1179, QN => DataPath_i_PIPLIN_A_19_port);
   DataPath_REG_A_Q_reg_21_inst : DFF_X1 port map( D => n3248, CK => CLK, Q => 
                           n_1180, QN => DataPath_i_PIPLIN_A_21_port);
   DataPath_REG_A_Q_reg_22_inst : DFF_X1 port map( D => n3247, CK => CLK, Q => 
                           n_1181, QN => DataPath_i_PIPLIN_A_22_port);
   DataPath_REG_A_Q_reg_23_inst : DFF_X1 port map( D => n3246, CK => CLK, Q => 
                           n_1182, QN => DataPath_i_PIPLIN_A_23_port);
   DataPath_REG_A_Q_reg_24_inst : DFF_X1 port map( D => n3245, CK => CLK, Q => 
                           n_1183, QN => DataPath_i_PIPLIN_A_24_port);
   DataPath_REG_A_Q_reg_25_inst : DFF_X1 port map( D => n3244, CK => CLK, Q => 
                           n_1184, QN => DataPath_i_PIPLIN_A_25_port);
   DataPath_REG_A_Q_reg_26_inst : DFF_X1 port map( D => n3243, CK => CLK, Q => 
                           n_1185, QN => DataPath_i_PIPLIN_A_26_port);
   DataPath_REG_A_Q_reg_27_inst : DFF_X1 port map( D => n3242, CK => CLK, Q => 
                           n_1186, QN => DataPath_i_PIPLIN_A_27_port);
   DataPath_REG_A_Q_reg_28_inst : DFF_X1 port map( D => n3241, CK => CLK, Q => 
                           n_1187, QN => DataPath_i_PIPLIN_A_28_port);
   DataPath_REG_A_Q_reg_29_inst : DFF_X1 port map( D => n3240, CK => CLK, Q => 
                           n_1188, QN => DataPath_i_PIPLIN_A_29_port);
   DataPath_REG_A_Q_reg_31_inst : DFF_X1 port map( D => n3238, CK => CLK, Q => 
                           n_1189, QN => DataPath_i_PIPLIN_A_31_port);
   DataPath_WRB1_Q_reg_1_inst : DFF_X1 port map( D => n2864, CK => CLK, Q => 
                           n_1190, QN => DataPath_i_PIPLIN_WRB1_1_port);
   DataPath_WRB2_Q_reg_1_inst : DFF_X1 port map( D => n2765, CK => CLK, Q => 
                           n_1191, QN => DataPath_i_PIPLIN_WRB2_1_port);
   DataPath_WRB3_Q_reg_1_inst : DFF_X1 port map( D => n356, CK => CLK, Q => 
                           i_ADD_WB_1_port, QN => n8276);
   DataPath_WRB1_Q_reg_2_inst : DFF_X1 port map( D => n2863, CK => CLK, Q => 
                           n_1192, QN => DataPath_i_PIPLIN_WRB1_2_port);
   DataPath_WRB2_Q_reg_2_inst : DFF_X1 port map( D => n2764, CK => CLK, Q => 
                           n_1193, QN => DataPath_i_PIPLIN_WRB2_2_port);
   DataPath_WRB3_Q_reg_2_inst : DFF_X1 port map( D => n357, CK => CLK, Q => 
                           i_ADD_WB_2_port, QN => n525);
   DataPath_WRB1_Q_reg_3_inst : DFF_X1 port map( D => n2862, CK => CLK, Q => 
                           n_1194, QN => DataPath_i_PIPLIN_WRB1_3_port);
   DataPath_WRB2_Q_reg_3_inst : DFF_X1 port map( D => n2763, CK => CLK, Q => 
                           n_1195, QN => DataPath_i_PIPLIN_WRB2_3_port);
   DataPath_WRB3_Q_reg_3_inst : DFF_X1 port map( D => n358, CK => CLK, Q => 
                           i_ADD_WB_3_port, QN => n_1196);
   DataPath_WRB1_Q_reg_4_inst : DFF_X1 port map( D => n2861, CK => CLK, Q => 
                           n_1197, QN => DataPath_i_PIPLIN_WRB1_4_port);
   DataPath_WRB2_Q_reg_4_inst : DFF_X1 port map( D => n2762, CK => CLK, Q => 
                           n_1198, QN => DataPath_i_PIPLIN_WRB2_4_port);
   DataPath_WRB3_Q_reg_4_inst : DFF_X1 port map( D => n359, CK => CLK, Q => 
                           i_ADD_WB_4_port, QN => n8209);
   DataPath_REG_IN1_Q_reg_0_inst : DFF_X1 port map( D => n2859, CK => CLK, Q =>
                           n8262, QN => DataPath_i_PIPLIN_IN1_0_port);
   DataPath_REG_IN1_Q_reg_2_inst : DFF_X1 port map( D => n2854, CK => CLK, Q =>
                           n_1199, QN => DataPath_i_PIPLIN_IN1_2_port);
   DataPath_REG_IN1_Q_reg_4_inst : DFF_X1 port map( D => n2852, CK => CLK, Q =>
                           n8259, QN => DataPath_i_PIPLIN_IN1_4_port);
   DataPath_REG_IN1_Q_reg_5_inst : DFF_X1 port map( D => n2851, CK => CLK, Q =>
                           n8258, QN => DataPath_i_PIPLIN_IN1_5_port);
   DataPath_REG_IN1_Q_reg_6_inst : DFF_X1 port map( D => n2850, CK => CLK, Q =>
                           n8263, QN => DataPath_i_PIPLIN_IN1_6_port);
   DataPath_REG_IN1_Q_reg_7_inst : DFF_X1 port map( D => n2849, CK => CLK, Q =>
                           n8264, QN => DataPath_i_PIPLIN_IN1_7_port);
   DataPath_REG_IN1_Q_reg_9_inst : DFF_X1 port map( D => n2847, CK => CLK, Q =>
                           n8261, QN => DataPath_i_PIPLIN_IN1_9_port);
   DataPath_REG_IN1_Q_reg_11_inst : DFF_X1 port map( D => n2845, CK => CLK, Q 
                           => n8260, QN => DataPath_i_PIPLIN_IN1_11_port);
   DataPath_REG_IN1_Q_reg_15_inst : DFF_X1 port map( D => n2840, CK => CLK, Q 
                           => n8257, QN => DataPath_i_PIPLIN_IN1_15_port);
   DataPath_REG_B_Q_reg_0_inst : DFF_X1 port map( D => n2755, CK => CLK, Q => 
                           n8235, QN => DataPath_i_PIPLIN_B_0_port);
   DataPath_REG_ME_Q_reg_0_inst : DFF_X1 port map( D => n2731, CK => CLK, Q => 
                           n_1200, QN => DataPath_i_REG_ME_DATA_DATAMEM_0_port)
                           ;
   DataPath_REG_B_Q_reg_1_inst : DFF_X1 port map( D => n2754, CK => CLK, Q => 
                           n8268, QN => DataPath_i_PIPLIN_B_1_port);
   DataPath_REG_ME_Q_reg_1_inst : DFF_X1 port map( D => n2730, CK => CLK, Q => 
                           n_1201, QN => DataPath_i_REG_ME_DATA_DATAMEM_1_port)
                           ;
   DataPath_REG_B_Q_reg_2_inst : DFF_X1 port map( D => n2753, CK => CLK, Q => 
                           n8244, QN => DataPath_i_PIPLIN_B_2_port);
   DataPath_REG_ME_Q_reg_2_inst : DFF_X1 port map( D => n2729, CK => CLK, Q => 
                           n_1202, QN => DataPath_i_REG_ME_DATA_DATAMEM_2_port)
                           ;
   DataPath_REG_B_Q_reg_5_inst : DFF_X1 port map( D => n2752, CK => CLK, Q => 
                           n_1203, QN => DataPath_i_PIPLIN_B_5_port);
   DataPath_REG_ME_Q_reg_5_inst : DFF_X1 port map( D => n2726, CK => CLK, Q => 
                           n_1204, QN => DataPath_i_REG_ME_DATA_DATAMEM_5_port)
                           ;
   DataPath_REG_B_Q_reg_7_inst : DFF_X1 port map( D => n2751, CK => CLK, Q => 
                           n8245, QN => DataPath_i_PIPLIN_B_7_port);
   DataPath_REG_ME_Q_reg_7_inst : DFF_X1 port map( D => n2724, CK => CLK, Q => 
                           n_1205, QN => DataPath_i_REG_ME_DATA_DATAMEM_7_port)
                           ;
   DataPath_REG_B_Q_reg_8_inst : DFF_X1 port map( D => n2750, CK => CLK, Q => 
                           n8247, QN => DataPath_i_PIPLIN_B_8_port);
   DataPath_REG_ME_Q_reg_8_inst : DFF_X1 port map( D => n2723, CK => CLK, Q => 
                           n_1206, QN => DataPath_i_REG_ME_DATA_DATAMEM_8_port)
                           ;
   DataPath_REG_B_Q_reg_9_inst : DFF_X1 port map( D => n2749, CK => CLK, Q => 
                           n8246, QN => DataPath_i_PIPLIN_B_9_port);
   DataPath_REG_ME_Q_reg_9_inst : DFF_X1 port map( D => n2722, CK => CLK, Q => 
                           n_1207, QN => DataPath_i_REG_ME_DATA_DATAMEM_9_port)
                           ;
   DataPath_REG_B_Q_reg_11_inst : DFF_X1 port map( D => n2748, CK => CLK, Q => 
                           n8248, QN => DataPath_i_PIPLIN_B_11_port);
   DataPath_REG_ME_Q_reg_11_inst : DFF_X1 port map( D => n2720, CK => CLK, Q =>
                           n_1208, QN => DataPath_i_REG_ME_DATA_DATAMEM_11_port
                           );
   DataPath_REG_B_Q_reg_15_inst : DFF_X1 port map( D => n2747, CK => CLK, Q => 
                           n8249, QN => DataPath_i_PIPLIN_B_15_port);
   DataPath_REG_ME_Q_reg_15_inst : DFF_X1 port map( D => n2716, CK => CLK, Q =>
                           n_1209, QN => DataPath_i_REG_ME_DATA_DATAMEM_15_port
                           );
   DataPath_REG_B_Q_reg_16_inst : DFF_X1 port map( D => n2746, CK => CLK, Q => 
                           n8251, QN => DataPath_i_PIPLIN_B_16_port);
   DataPath_REG_ME_Q_reg_16_inst : DFF_X1 port map( D => n2715, CK => CLK, Q =>
                           n_1210, QN => DataPath_i_REG_ME_DATA_DATAMEM_16_port
                           );
   DataPath_REG_B_Q_reg_17_inst : DFF_X1 port map( D => n2745, CK => CLK, Q => 
                           n8250, QN => DataPath_i_PIPLIN_B_17_port);
   DataPath_REG_ME_Q_reg_17_inst : DFF_X1 port map( D => n2714, CK => CLK, Q =>
                           n_1211, QN => DataPath_i_REG_ME_DATA_DATAMEM_17_port
                           );
   DataPath_REG_B_Q_reg_18_inst : DFF_X1 port map( D => n2744, CK => CLK, Q => 
                           n8253, QN => DataPath_i_PIPLIN_B_18_port);
   DataPath_REG_ME_Q_reg_18_inst : DFF_X1 port map( D => n2713, CK => CLK, Q =>
                           n_1212, QN => DataPath_i_REG_ME_DATA_DATAMEM_18_port
                           );
   DataPath_REG_B_Q_reg_19_inst : DFF_X1 port map( D => n2743, CK => CLK, Q => 
                           n8252, QN => DataPath_i_PIPLIN_B_19_port);
   DataPath_REG_ME_Q_reg_19_inst : DFF_X1 port map( D => n2712, CK => CLK, Q =>
                           n_1213, QN => DataPath_i_REG_ME_DATA_DATAMEM_19_port
                           );
   DataPath_REG_ME_Q_reg_21_inst : DFF_X1 port map( D => n2710, CK => CLK, Q =>
                           n_1214, QN => DataPath_i_REG_ME_DATA_DATAMEM_21_port
                           );
   DataPath_REG_B_Q_reg_22_inst : DFF_X1 port map( D => n2741, CK => CLK, Q => 
                           n8254, QN => DataPath_i_PIPLIN_B_22_port);
   DataPath_REG_ME_Q_reg_22_inst : DFF_X1 port map( D => n2709, CK => CLK, Q =>
                           n_1215, QN => DataPath_i_REG_ME_DATA_DATAMEM_22_port
                           );
   DataPath_REG_ME_Q_reg_23_inst : DFF_X1 port map( D => n2708, CK => CLK, Q =>
                           n_1216, QN => DataPath_i_REG_ME_DATA_DATAMEM_23_port
                           );
   DataPath_REG_B_Q_reg_24_inst : DFF_X1 port map( D => n2739, CK => CLK, Q => 
                           n8255, QN => DataPath_i_PIPLIN_B_24_port);
   DataPath_REG_ME_Q_reg_24_inst : DFF_X1 port map( D => n2707, CK => CLK, Q =>
                           n_1217, QN => DataPath_i_REG_ME_DATA_DATAMEM_24_port
                           );
   DataPath_REG_B_Q_reg_25_inst : DFF_X1 port map( D => n2738, CK => CLK, Q => 
                           n8201, QN => DataPath_i_PIPLIN_B_25_port);
   DataPath_REG_ME_Q_reg_25_inst : DFF_X1 port map( D => n2706, CK => CLK, Q =>
                           n_1218, QN => DataPath_i_REG_ME_DATA_DATAMEM_25_port
                           );
   DataPath_REG_B_Q_reg_26_inst : DFF_X1 port map( D => n2737, CK => CLK, Q => 
                           n8256, QN => DataPath_i_PIPLIN_B_26_port);
   DataPath_REG_ME_Q_reg_26_inst : DFF_X1 port map( D => n2705, CK => CLK, Q =>
                           n_1219, QN => DataPath_i_REG_ME_DATA_DATAMEM_26_port
                           );
   DataPath_REG_B_Q_reg_27_inst : DFF_X1 port map( D => n2736, CK => CLK, Q => 
                           n8288, QN => DataPath_i_PIPLIN_B_27_port);
   DataPath_REG_ME_Q_reg_27_inst : DFF_X1 port map( D => n2704, CK => CLK, Q =>
                           n_1220, QN => DataPath_i_REG_ME_DATA_DATAMEM_27_port
                           );
   DataPath_REG_B_Q_reg_28_inst : DFF_X1 port map( D => n2735, CK => CLK, Q => 
                           n8299, QN => DataPath_i_PIPLIN_B_28_port);
   DataPath_REG_ME_Q_reg_28_inst : DFF_X1 port map( D => n2703, CK => CLK, Q =>
                           n_1221, QN => DataPath_i_REG_ME_DATA_DATAMEM_28_port
                           );
   DataPath_REG_B_Q_reg_29_inst : DFF_X1 port map( D => n2734, CK => CLK, Q => 
                           n8243, QN => DataPath_i_PIPLIN_B_29_port);
   DataPath_REG_ME_Q_reg_29_inst : DFF_X1 port map( D => n2702, CK => CLK, Q =>
                           n_1222, QN => DataPath_i_REG_ME_DATA_DATAMEM_29_port
                           );
   DataPath_REG_B_Q_reg_30_inst : DFF_X1 port map( D => n2733, CK => CLK, Q => 
                           n8298, QN => DataPath_i_PIPLIN_B_30_port);
   DataPath_REG_ME_Q_reg_30_inst : DFF_X1 port map( D => n2701, CK => CLK, Q =>
                           n_1223, QN => DataPath_i_REG_ME_DATA_DATAMEM_30_port
                           );
   DataPath_REG_IN2_Q_reg_0_inst : DFF_X1 port map( D => n2387, CK => CLK, Q =>
                           n_1224, QN => DataPath_i_PIPLIN_IN2_0_port);
   DataPath_REG_IN2_Q_reg_2_inst : DFF_X1 port map( D => n2384, CK => CLK, Q =>
                           n_1225, QN => DataPath_i_PIPLIN_IN2_2_port);
   DataPath_REG_IN2_Q_reg_7_inst : DFF_X1 port map( D => n2377, CK => CLK, Q =>
                           n_1226, QN => DataPath_i_PIPLIN_IN2_7_port);
   DataPath_REG_IN2_Q_reg_8_inst : DFF_X1 port map( D => n2375, CK => CLK, Q =>
                           n_1227, QN => DataPath_i_PIPLIN_IN2_8_port);
   DataPath_REG_IN2_Q_reg_9_inst : DFF_X1 port map( D => n2373, CK => CLK, Q =>
                           n_1228, QN => DataPath_i_PIPLIN_IN2_9_port);
   DataPath_REG_IN2_Q_reg_11_inst : DFF_X1 port map( D => n2370, CK => CLK, Q 
                           => n_1229, QN => DataPath_i_PIPLIN_IN2_11_port);
   DataPath_REG_IN2_Q_reg_15_inst : DFF_X1 port map( D => n2365, CK => CLK, Q 
                           => n_1230, QN => DataPath_i_PIPLIN_IN2_15_port);
   DataPath_REG_IN2_Q_reg_16_inst : DFF_X1 port map( D => n2363, CK => CLK, Q 
                           => n_1231, QN => DataPath_i_PIPLIN_IN2_16_port);
   DataPath_REG_IN2_Q_reg_17_inst : DFF_X1 port map( D => n2361, CK => CLK, Q 
                           => n_1232, QN => DataPath_i_PIPLIN_IN2_17_port);
   DataPath_REG_IN2_Q_reg_18_inst : DFF_X1 port map( D => n2359, CK => CLK, Q 
                           => n_1233, QN => DataPath_i_PIPLIN_IN2_18_port);
   DataPath_REG_IN2_Q_reg_19_inst : DFF_X1 port map( D => n2357, CK => CLK, Q 
                           => n_1234, QN => DataPath_i_PIPLIN_IN2_19_port);
   DataPath_REG_IN2_Q_reg_21_inst : DFF_X1 port map( D => n2352, CK => CLK, Q 
                           => n_1235, QN => DataPath_i_PIPLIN_IN2_21_port);
   DataPath_REG_IN2_Q_reg_22_inst : DFF_X1 port map( D => n2350, CK => CLK, Q 
                           => n_1236, QN => DataPath_i_PIPLIN_IN2_22_port);
   DataPath_REG_IN2_Q_reg_23_inst : DFF_X1 port map( D => n2348, CK => CLK, Q 
                           => n_1237, QN => DataPath_i_PIPLIN_IN2_23_port);
   DataPath_REG_IN2_Q_reg_24_inst : DFF_X1 port map( D => n2346, CK => CLK, Q 
                           => n_1238, QN => DataPath_i_PIPLIN_IN2_24_port);
   DataPath_REG_IN2_Q_reg_25_inst : DFF_X1 port map( D => n2344, CK => CLK, Q 
                           => n_1239, QN => DataPath_i_PIPLIN_IN2_25_port);
   DataPath_REG_IN2_Q_reg_26_inst : DFF_X1 port map( D => n2342, CK => CLK, Q 
                           => n_1240, QN => DataPath_i_PIPLIN_IN2_26_port);
   DataPath_REG_IN2_Q_reg_27_inst : DFF_X1 port map( D => n2340, CK => CLK, Q 
                           => n_1241, QN => DataPath_i_PIPLIN_IN2_27_port);
   DataPath_REG_IN2_Q_reg_28_inst : DFF_X1 port map( D => n2338, CK => CLK, Q 
                           => n_1242, QN => DataPath_i_PIPLIN_IN2_28_port);
   DataPath_REG_IN2_Q_reg_29_inst : DFF_X1 port map( D => n2336, CK => CLK, Q 
                           => n_1243, QN => DataPath_i_PIPLIN_IN2_29_port);
   DataPath_REG_IN2_Q_reg_30_inst : DFF_X1 port map( D => n2334, CK => CLK, Q 
                           => n_1244, QN => DataPath_i_PIPLIN_IN2_30_port);
   DataPath_REG_IN2_Q_reg_31_inst : DFF_X1 port map( D => n2332, CK => CLK, Q 
                           => n_1245, QN => DataPath_i_PIPLIN_IN2_31_port);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_7_inst : DFF_X1 port map( D => n6952, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_199_port
                           , QN => n766);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_7_inst : DFF_X1 port map( D => n6888, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_135_port
                           , QN => n702);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_7_inst : DFF_X1 port map( D => n6856, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_103_port
                           , QN => n670);
   CU_I_setcmp_1_reg_0_inst : DFF_X1 port map( D => n7090, CK => CLK, Q => 
                           i_SEL_LGET_0_port, QN => n8332);
   CU_I_aluOpcode1_reg_4_inst : DFF_X1 port map( D => n7091, CK => CLK, Q => 
                           i_ALU_OP_4_port, QN => n8189);
   CU_I_aluOpcode1_reg_3_inst : DFF_X1 port map( D => n7092, CK => CLK, Q => 
                           i_ALU_OP_3_port, QN => n8197);
   CU_I_aluOpcode1_reg_1_inst : DFF_X1 port map( D => n7094, CK => CLK, Q => 
                           i_ALU_OP_1_port, QN => n_1246);
   DataPath_REG_MEM_ALUOUT_Q_reg_31_inst : DFF_X1 port map( D => n1116, CK => 
                           CLK, Q => n_1247, QN => 
                           DataPath_i_REG_MEM_ALUOUT_31_port);
   DataPath_REG_ALU_OUT_Q_reg_7_inst : DFF_X1 port map( D => n1998, CK => CLK, 
                           Q => n_1248, QN => DRAM_ADDRESS_7_port);
   DataPath_REG_MEM_ALUOUT_Q_reg_7_inst : DFF_X1 port map( D => n1142, CK => 
                           CLK, Q => n_1249, QN => 
                           DataPath_i_REG_MEM_ALUOUT_7_port);
   DataPath_REG_ALU_OUT_Q_reg_6_inst : DFF_X1 port map( D => n7016, CK => CLK, 
                           Q => DRAM_ADDRESS_6_port, QN => n497);
   DataPath_REG_MEM_ALUOUT_Q_reg_6_inst : DFF_X1 port map( D => n1143, CK => 
                           CLK, Q => n_1250, QN => 
                           DataPath_i_REG_MEM_ALUOUT_6_port);
   DataPath_REG_ALU_OUT_Q_reg_0_inst : DFF_X1 port map( D => n7020, CK => CLK, 
                           Q => n8278, QN => n494);
   DataPath_REG_MEM_ALUOUT_Q_reg_0_inst : DFF_X1 port map( D => n1149, CK => 
                           CLK, Q => n_1251, QN => 
                           DataPath_i_REG_MEM_ALUOUT_0_port);
   DataPath_REG_ALU_OUT_Q_reg_17_inst : DFF_X1 port map( D => n7006, CK => CLK,
                           Q => DRAM_ADDRESS_17_port, QN => n8331);
   DataPath_REG_MEM_ALUOUT_Q_reg_17_inst : DFF_X1 port map( D => n1132, CK => 
                           CLK, Q => n_1252, QN => 
                           DataPath_i_REG_MEM_ALUOUT_17_port);
   DataPath_REG_ALU_OUT_Q_reg_13_inst : DFF_X1 port map( D => n7010, CK => CLK,
                           Q => DRAM_ADDRESS_13_port, QN => n8330);
   DataPath_REG_MEM_ALUOUT_Q_reg_13_inst : DFF_X1 port map( D => n1136, CK => 
                           CLK, Q => n_1253, QN => 
                           DataPath_i_REG_MEM_ALUOUT_13_port);
   DataPath_REG_ALU_OUT_Q_reg_9_inst : DFF_X1 port map( D => n7014, CK => CLK, 
                           Q => DRAM_ADDRESS_9_port, QN => n8318);
   DataPath_REG_MEM_ALUOUT_Q_reg_9_inst : DFF_X1 port map( D => n1140, CK => 
                           CLK, Q => n_1254, QN => 
                           DataPath_i_REG_MEM_ALUOUT_9_port);
   DataPath_REG_ALU_OUT_Q_reg_5_inst : DFF_X1 port map( D => n7017, CK => CLK, 
                           Q => DRAM_ADDRESS_5_port, QN => n8317);
   DataPath_REG_MEM_ALUOUT_Q_reg_5_inst : DFF_X1 port map( D => n1144, CK => 
                           CLK, Q => n_1255, QN => 
                           DataPath_i_REG_MEM_ALUOUT_5_port);
   DataPath_REG_ALU_OUT_Q_reg_1_inst : DFF_X1 port map( D => n7019, CK => CLK, 
                           Q => n8285, QN => n495);
   DataPath_REG_MEM_ALUOUT_Q_reg_1_inst : DFF_X1 port map( D => n1148, CK => 
                           CLK, Q => n_1256, QN => 
                           DataPath_i_REG_MEM_ALUOUT_1_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_23_inst : DFF_X1 port map( D => n2186, CK 
                           => CLK, Q => n_1257, QN => 
                           DataPath_i_REG_LDSTR_OUT_23_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_31_inst : DFF_X1 port map( D => n2178, CK 
                           => CLK, Q => n_1258, QN => 
                           DataPath_i_REG_LDSTR_OUT_31_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_31_inst : DFF_X1 port map( D => n6768, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_63_port,
                           QN => n630);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_31_inst : DFF_X1 port map( D => n6800, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_95_port,
                           QN => n662);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_31_inst : DFF_X1 port map( D => n6832, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_127_port
                           , QN => n694);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_31_inst : DFF_X1 port map( D => n6864, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_159_port
                           , QN => n726);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_31_inst : DFF_X1 port map( D => n6896, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_191_port
                           , QN => n758);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_31_inst : DFF_X1 port map( D => n6928, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_223_port
                           , QN => n790);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_31_inst : DFF_X1 port map( D => n6960, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_255_port
                           , QN => n822);
   DataPath_RF_BLOCKi_8_Q_reg_31_inst : DFF_X1 port map( D => n3154, CK => CLK,
                           Q => n_1259, QN => 
                           DataPath_RF_bus_reg_dataout_31_port);
   DataPath_RF_BLOCKi_9_Q_reg_31_inst : DFF_X1 port map( D => n3379, CK => CLK,
                           Q => n_1260, QN => 
                           DataPath_RF_bus_reg_dataout_63_port);
   DataPath_RF_BLOCKi_10_Q_reg_31_inst : DFF_X1 port map( D => n3417, CK => CLK
                           , Q => n_1261, QN => 
                           DataPath_RF_bus_reg_dataout_95_port);
   DataPath_RF_BLOCKi_11_Q_reg_31_inst : DFF_X1 port map( D => n3455, CK => CLK
                           , Q => n_1262, QN => 
                           DataPath_RF_bus_reg_dataout_127_port);
   DataPath_RF_BLOCKi_12_Q_reg_31_inst : DFF_X1 port map( D => n3493, CK => CLK
                           , Q => n_1263, QN => 
                           DataPath_RF_bus_reg_dataout_159_port);
   DataPath_RF_BLOCKi_13_Q_reg_31_inst : DFF_X1 port map( D => n3531, CK => CLK
                           , Q => n_1264, QN => 
                           DataPath_RF_bus_reg_dataout_191_port);
   DataPath_RF_BLOCKi_14_Q_reg_31_inst : DFF_X1 port map( D => n3569, CK => CLK
                           , Q => n_1265, QN => 
                           DataPath_RF_bus_reg_dataout_223_port);
   DataPath_RF_BLOCKi_15_Q_reg_31_inst : DFF_X1 port map( D => n3607, CK => CLK
                           , Q => n_1266, QN => 
                           DataPath_RF_bus_reg_dataout_255_port);
   DataPath_RF_BLOCKi_16_Q_reg_31_inst : DFF_X1 port map( D => n3645, CK => CLK
                           , Q => n_1267, QN => 
                           DataPath_RF_bus_reg_dataout_287_port);
   DataPath_RF_BLOCKi_17_Q_reg_31_inst : DFF_X1 port map( D => n3682, CK => CLK
                           , Q => n_1268, QN => 
                           DataPath_RF_bus_reg_dataout_319_port);
   DataPath_RF_BLOCKi_18_Q_reg_31_inst : DFF_X1 port map( D => n3719, CK => CLK
                           , Q => n_1269, QN => 
                           DataPath_RF_bus_reg_dataout_351_port);
   DataPath_RF_BLOCKi_19_Q_reg_31_inst : DFF_X1 port map( D => n3756, CK => CLK
                           , Q => n_1270, QN => 
                           DataPath_RF_bus_reg_dataout_383_port);
   DataPath_RF_BLOCKi_20_Q_reg_31_inst : DFF_X1 port map( D => n3791, CK => CLK
                           , Q => n_1271, QN => 
                           DataPath_RF_bus_reg_dataout_415_port);
   DataPath_RF_BLOCKi_21_Q_reg_31_inst : DFF_X1 port map( D => n3826, CK => CLK
                           , Q => n_1272, QN => 
                           DataPath_RF_bus_reg_dataout_447_port);
   DataPath_RF_BLOCKi_22_Q_reg_31_inst : DFF_X1 port map( D => n3861, CK => CLK
                           , Q => n_1273, QN => 
                           DataPath_RF_bus_reg_dataout_479_port);
   DataPath_RF_BLOCKi_23_Q_reg_31_inst : DFF_X1 port map( D => n3896, CK => CLK
                           , Q => n_1274, QN => 
                           DataPath_RF_bus_reg_dataout_511_port);
   DataPath_RF_BLOCKi_24_Q_reg_31_inst : DFF_X1 port map( D => n3964, CK => CLK
                           , Q => n_1275, QN => 
                           DataPath_RF_bus_reg_dataout_543_port);
   DataPath_RF_BLOCKi_25_Q_reg_31_inst : DFF_X1 port map( D => n4032, CK => CLK
                           , Q => n_1276, QN => 
                           DataPath_RF_bus_reg_dataout_575_port);
   DataPath_RF_BLOCKi_26_Q_reg_31_inst : DFF_X1 port map( D => n4067, CK => CLK
                           , Q => n_1277, QN => 
                           DataPath_RF_bus_reg_dataout_607_port);
   DataPath_RF_BLOCKi_27_Q_reg_31_inst : DFF_X1 port map( D => n4102, CK => CLK
                           , Q => n_1278, QN => 
                           DataPath_RF_bus_reg_dataout_639_port);
   DataPath_RF_BLOCKi_28_Q_reg_31_inst : DFF_X1 port map( D => n4137, CK => CLK
                           , Q => n_1279, QN => 
                           DataPath_RF_bus_reg_dataout_671_port);
   DataPath_RF_BLOCKi_29_Q_reg_31_inst : DFF_X1 port map( D => n4172, CK => CLK
                           , Q => n_1280, QN => 
                           DataPath_RF_bus_reg_dataout_703_port);
   DataPath_RF_BLOCKi_30_Q_reg_31_inst : DFF_X1 port map( D => n4207, CK => CLK
                           , Q => n_1281, QN => 
                           DataPath_RF_bus_reg_dataout_735_port);
   DataPath_RF_BLOCKi_31_Q_reg_31_inst : DFF_X1 port map( D => n4242, CK => CLK
                           , Q => n_1282, QN => 
                           DataPath_RF_bus_reg_dataout_767_port);
   DataPath_RF_BLOCKi_32_Q_reg_31_inst : DFF_X1 port map( D => n4277, CK => CLK
                           , Q => n_1283, QN => 
                           DataPath_RF_bus_reg_dataout_799_port);
   DataPath_RF_BLOCKi_33_Q_reg_31_inst : DFF_X1 port map( D => n4312, CK => CLK
                           , Q => n_1284, QN => 
                           DataPath_RF_bus_reg_dataout_831_port);
   DataPath_RF_BLOCKi_34_Q_reg_31_inst : DFF_X1 port map( D => n4347, CK => CLK
                           , Q => n_1285, QN => 
                           DataPath_RF_bus_reg_dataout_863_port);
   DataPath_RF_BLOCKi_35_Q_reg_31_inst : DFF_X1 port map( D => n4382, CK => CLK
                           , Q => n_1286, QN => 
                           DataPath_RF_bus_reg_dataout_895_port);
   DataPath_RF_BLOCKi_36_Q_reg_31_inst : DFF_X1 port map( D => n4417, CK => CLK
                           , Q => n_1287, QN => 
                           DataPath_RF_bus_reg_dataout_927_port);
   DataPath_RF_BLOCKi_37_Q_reg_31_inst : DFF_X1 port map( D => n4452, CK => CLK
                           , Q => n_1288, QN => 
                           DataPath_RF_bus_reg_dataout_959_port);
   DataPath_RF_BLOCKi_38_Q_reg_31_inst : DFF_X1 port map( D => n4487, CK => CLK
                           , Q => n_1289, QN => 
                           DataPath_RF_bus_reg_dataout_991_port);
   DataPath_RF_BLOCKi_39_Q_reg_31_inst : DFF_X1 port map( D => n4522, CK => CLK
                           , Q => n_1290, QN => 
                           DataPath_RF_bus_reg_dataout_1023_port);
   DataPath_RF_BLOCKi_40_Q_reg_31_inst : DFF_X1 port map( D => n4557, CK => CLK
                           , Q => n_1291, QN => 
                           DataPath_RF_bus_reg_dataout_1055_port);
   DataPath_RF_BLOCKi_41_Q_reg_31_inst : DFF_X1 port map( D => n4625, CK => CLK
                           , Q => n_1292, QN => 
                           DataPath_RF_bus_reg_dataout_1087_port);
   DataPath_RF_BLOCKi_42_Q_reg_31_inst : DFF_X1 port map( D => n4660, CK => CLK
                           , Q => n_1293, QN => 
                           DataPath_RF_bus_reg_dataout_1119_port);
   DataPath_RF_BLOCKi_43_Q_reg_31_inst : DFF_X1 port map( D => n4695, CK => CLK
                           , Q => n_1294, QN => 
                           DataPath_RF_bus_reg_dataout_1151_port);
   DataPath_RF_BLOCKi_44_Q_reg_31_inst : DFF_X1 port map( D => n4730, CK => CLK
                           , Q => n_1295, QN => 
                           DataPath_RF_bus_reg_dataout_1183_port);
   DataPath_RF_BLOCKi_45_Q_reg_31_inst : DFF_X1 port map( D => n4765, CK => CLK
                           , Q => n_1296, QN => 
                           DataPath_RF_bus_reg_dataout_1215_port);
   DataPath_RF_BLOCKi_46_Q_reg_31_inst : DFF_X1 port map( D => n4800, CK => CLK
                           , Q => n_1297, QN => 
                           DataPath_RF_bus_reg_dataout_1247_port);
   DataPath_RF_BLOCKi_47_Q_reg_31_inst : DFF_X1 port map( D => n4835, CK => CLK
                           , Q => n_1298, QN => 
                           DataPath_RF_bus_reg_dataout_1279_port);
   DataPath_RF_BLOCKi_48_Q_reg_31_inst : DFF_X1 port map( D => n4870, CK => CLK
                           , Q => n_1299, QN => 
                           DataPath_RF_bus_reg_dataout_1311_port);
   DataPath_RF_BLOCKi_49_Q_reg_31_inst : DFF_X1 port map( D => n4905, CK => CLK
                           , Q => n_1300, QN => 
                           DataPath_RF_bus_reg_dataout_1343_port);
   DataPath_RF_BLOCKi_50_Q_reg_31_inst : DFF_X1 port map( D => n4940, CK => CLK
                           , Q => n_1301, QN => 
                           DataPath_RF_bus_reg_dataout_1375_port);
   DataPath_RF_BLOCKi_51_Q_reg_31_inst : DFF_X1 port map( D => n4975, CK => CLK
                           , Q => n_1302, QN => 
                           DataPath_RF_bus_reg_dataout_1407_port);
   DataPath_RF_BLOCKi_52_Q_reg_31_inst : DFF_X1 port map( D => n5010, CK => CLK
                           , Q => n_1303, QN => 
                           DataPath_RF_bus_reg_dataout_1439_port);
   DataPath_RF_BLOCKi_53_Q_reg_31_inst : DFF_X1 port map( D => n5045, CK => CLK
                           , Q => n_1304, QN => 
                           DataPath_RF_bus_reg_dataout_1471_port);
   DataPath_RF_BLOCKi_54_Q_reg_31_inst : DFF_X1 port map( D => n5080, CK => CLK
                           , Q => n_1305, QN => 
                           DataPath_RF_bus_reg_dataout_1503_port);
   DataPath_RF_BLOCKi_55_Q_reg_31_inst : DFF_X1 port map( D => n5115, CK => CLK
                           , Q => n_1306, QN => 
                           DataPath_RF_bus_reg_dataout_1535_port);
   DataPath_RF_BLOCKi_56_Q_reg_31_inst : DFF_X1 port map( D => n5150, CK => CLK
                           , Q => n_1307, QN => 
                           DataPath_RF_bus_reg_dataout_1567_port);
   DataPath_RF_BLOCKi_57_Q_reg_31_inst : DFF_X1 port map( D => n5217, CK => CLK
                           , Q => n_1308, QN => 
                           DataPath_RF_bus_reg_dataout_1599_port);
   DataPath_RF_BLOCKi_58_Q_reg_31_inst : DFF_X1 port map( D => n5253, CK => CLK
                           , Q => n_1309, QN => 
                           DataPath_RF_bus_reg_dataout_1631_port);
   DataPath_RF_BLOCKi_59_Q_reg_31_inst : DFF_X1 port map( D => n5288, CK => CLK
                           , Q => n_1310, QN => 
                           DataPath_RF_bus_reg_dataout_1663_port);
   DataPath_RF_BLOCKi_60_Q_reg_31_inst : DFF_X1 port map( D => n5323, CK => CLK
                           , Q => n_1311, QN => 
                           DataPath_RF_bus_reg_dataout_1695_port);
   DataPath_RF_BLOCKi_61_Q_reg_31_inst : DFF_X1 port map( D => n5358, CK => CLK
                           , Q => n_1312, QN => 
                           DataPath_RF_bus_reg_dataout_1727_port);
   DataPath_RF_BLOCKi_62_Q_reg_31_inst : DFF_X1 port map( D => n5393, CK => CLK
                           , Q => n_1313, QN => 
                           DataPath_RF_bus_reg_dataout_1759_port);
   DataPath_RF_BLOCKi_63_Q_reg_31_inst : DFF_X1 port map( D => n5428, CK => CLK
                           , Q => n_1314, QN => 
                           DataPath_RF_bus_reg_dataout_1791_port);
   DataPath_RF_BLOCKi_64_Q_reg_31_inst : DFF_X1 port map( D => n5463, CK => CLK
                           , Q => n_1315, QN => 
                           DataPath_RF_bus_reg_dataout_1823_port);
   DataPath_RF_BLOCKi_65_Q_reg_31_inst : DFF_X1 port map( D => n5498, CK => CLK
                           , Q => n_1316, QN => 
                           DataPath_RF_bus_reg_dataout_1855_port);
   DataPath_RF_BLOCKi_66_Q_reg_31_inst : DFF_X1 port map( D => n5533, CK => CLK
                           , Q => n_1317, QN => 
                           DataPath_RF_bus_reg_dataout_1887_port);
   DataPath_RF_BLOCKi_67_Q_reg_31_inst : DFF_X1 port map( D => n5568, CK => CLK
                           , Q => n_1318, QN => 
                           DataPath_RF_bus_reg_dataout_1919_port);
   DataPath_RF_BLOCKi_68_Q_reg_31_inst : DFF_X1 port map( D => n5607, CK => CLK
                           , Q => n_1319, QN => 
                           DataPath_RF_bus_reg_dataout_1951_port);
   DataPath_RF_BLOCKi_69_Q_reg_31_inst : DFF_X1 port map( D => n5644, CK => CLK
                           , Q => n_1320, QN => 
                           DataPath_RF_bus_reg_dataout_1983_port);
   DataPath_RF_BLOCKi_70_Q_reg_31_inst : DFF_X1 port map( D => n5681, CK => CLK
                           , Q => n_1321, QN => 
                           DataPath_RF_bus_reg_dataout_2015_port);
   DataPath_RF_BLOCKi_71_Q_reg_31_inst : DFF_X1 port map( D => n5718, CK => CLK
                           , Q => n_1322, QN => 
                           DataPath_RF_bus_reg_dataout_2047_port);
   DataPath_RF_BLOCKi_83_Q_reg_31_inst : DFF_X1 port map( D => n914, CK => CLK,
                           Q => n_1323, QN => 
                           DataPath_RF_bus_reg_dataout_2431_port);
   DataPath_RF_BLOCKi_84_Q_reg_31_inst : DFF_X1 port map( D => n968, CK => CLK,
                           Q => n_1324, QN => 
                           DataPath_RF_bus_reg_dataout_2463_port);
   DataPath_RF_BLOCKi_85_Q_reg_31_inst : DFF_X1 port map( D => n1005, CK => CLK
                           , Q => n_1325, QN => 
                           DataPath_RF_bus_reg_dataout_2495_port);
   DataPath_RF_BLOCKi_86_Q_reg_31_inst : DFF_X1 port map( D => n1042, CK => CLK
                           , Q => n_1326, QN => 
                           DataPath_RF_bus_reg_dataout_2527_port);
   DataPath_RF_BLOCKi_87_Q_reg_31_inst : DFF_X1 port map( D => n1079, CK => CLK
                           , Q => n_1327, QN => 
                           DataPath_RF_bus_reg_dataout_2559_port);
   DataPath_RF_BLOCKi_72_Q_reg_31_inst : DFF_X1 port map( D => n5755, CK => CLK
                           , Q => n_1328, QN => 
                           DataPath_RF_bus_reg_dataout_2079_port);
   DataPath_RF_BLOCKi_73_Q_reg_31_inst : DFF_X1 port map( D => n5794, CK => CLK
                           , Q => n_1329, QN => 
                           DataPath_RF_bus_reg_dataout_2111_port);
   DataPath_RF_BLOCKi_74_Q_reg_31_inst : DFF_X1 port map( D => n5830, CK => CLK
                           , Q => n_1330, QN => 
                           DataPath_RF_bus_reg_dataout_2143_port);
   DataPath_RF_BLOCKi_75_Q_reg_31_inst : DFF_X1 port map( D => n5866, CK => CLK
                           , Q => n_1331, QN => 
                           DataPath_RF_bus_reg_dataout_2175_port);
   DataPath_RF_BLOCKi_76_Q_reg_31_inst : DFF_X1 port map( D => n5902, CK => CLK
                           , Q => n_1332, QN => 
                           DataPath_RF_bus_reg_dataout_2207_port);
   DataPath_RF_BLOCKi_77_Q_reg_31_inst : DFF_X1 port map( D => n5938, CK => CLK
                           , Q => n_1333, QN => 
                           DataPath_RF_bus_reg_dataout_2239_port);
   DataPath_RF_BLOCKi_78_Q_reg_31_inst : DFF_X1 port map( D => n5974, CK => CLK
                           , Q => n_1334, QN => 
                           DataPath_RF_bus_reg_dataout_2271_port);
   DataPath_RF_BLOCKi_79_Q_reg_31_inst : DFF_X1 port map( D => n6010, CK => CLK
                           , Q => n_1335, QN => 
                           DataPath_RF_bus_reg_dataout_2303_port);
   DataPath_RF_BLOCKi_80_Q_reg_31_inst : DFF_X1 port map( D => n6047, CK => CLK
                           , Q => n_1336, QN => 
                           DataPath_RF_bus_reg_dataout_2335_port);
   DataPath_RF_BLOCKi_81_Q_reg_31_inst : DFF_X1 port map( D => n6083, CK => CLK
                           , Q => n_1337, QN => 
                           DataPath_RF_bus_reg_dataout_2367_port);
   DataPath_RF_BLOCKi_82_Q_reg_31_inst : DFF_X1 port map( D => n6119, CK => CLK
                           , Q => n_1338, QN => 
                           DataPath_RF_bus_reg_dataout_2399_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_15_inst : DFF_X1 port map( D => n2194, CK 
                           => CLK, Q => n_1339, QN => 
                           DataPath_i_REG_LDSTR_OUT_15_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_17_inst : DFF_X1 port map( D => n2192, CK 
                           => CLK, Q => n_1340, QN => 
                           DataPath_i_REG_LDSTR_OUT_17_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_17_inst : DFF_X1 port map( D => n6782, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_49_port,
                           QN => n616);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_17_inst : DFF_X1 port map( D => n6814, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_81_port,
                           QN => n648);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_17_inst : DFF_X1 port map( D => n6846, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_113_port
                           , QN => n680);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_17_inst : DFF_X1 port map( D => n6878, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_145_port
                           , QN => n712);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_17_inst : DFF_X1 port map( D => n6910, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_177_port
                           , QN => n744);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_17_inst : DFF_X1 port map( D => n6942, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_209_port
                           , QN => n776);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_17_inst : DFF_X1 port map( D => n6974, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_241_port
                           , QN => n808);
   DataPath_RF_BLOCKi_8_Q_reg_17_inst : DFF_X1 port map( D => n3338, CK => CLK,
                           Q => n_1341, QN => 
                           DataPath_RF_bus_reg_dataout_17_port);
   DataPath_RF_BLOCKi_9_Q_reg_17_inst : DFF_X1 port map( D => n3395, CK => CLK,
                           Q => n_1342, QN => 
                           DataPath_RF_bus_reg_dataout_49_port);
   DataPath_RF_BLOCKi_10_Q_reg_17_inst : DFF_X1 port map( D => n3433, CK => CLK
                           , Q => n_1343, QN => 
                           DataPath_RF_bus_reg_dataout_81_port);
   DataPath_RF_BLOCKi_11_Q_reg_17_inst : DFF_X1 port map( D => n3471, CK => CLK
                           , Q => n_1344, QN => 
                           DataPath_RF_bus_reg_dataout_113_port);
   DataPath_RF_BLOCKi_12_Q_reg_17_inst : DFF_X1 port map( D => n3509, CK => CLK
                           , Q => n_1345, QN => 
                           DataPath_RF_bus_reg_dataout_145_port);
   DataPath_RF_BLOCKi_13_Q_reg_17_inst : DFF_X1 port map( D => n3547, CK => CLK
                           , Q => n_1346, QN => 
                           DataPath_RF_bus_reg_dataout_177_port);
   DataPath_RF_BLOCKi_14_Q_reg_17_inst : DFF_X1 port map( D => n3585, CK => CLK
                           , Q => n_1347, QN => 
                           DataPath_RF_bus_reg_dataout_209_port);
   DataPath_RF_BLOCKi_15_Q_reg_17_inst : DFF_X1 port map( D => n3623, CK => CLK
                           , Q => n_1348, QN => 
                           DataPath_RF_bus_reg_dataout_241_port);
   DataPath_RF_BLOCKi_16_Q_reg_17_inst : DFF_X1 port map( D => n3661, CK => CLK
                           , Q => n_1349, QN => 
                           DataPath_RF_bus_reg_dataout_273_port);
   DataPath_RF_BLOCKi_17_Q_reg_17_inst : DFF_X1 port map( D => n3698, CK => CLK
                           , Q => n_1350, QN => 
                           DataPath_RF_bus_reg_dataout_305_port);
   DataPath_RF_BLOCKi_18_Q_reg_17_inst : DFF_X1 port map( D => n3735, CK => CLK
                           , Q => n_1351, QN => 
                           DataPath_RF_bus_reg_dataout_337_port);
   DataPath_RF_BLOCKi_19_Q_reg_17_inst : DFF_X1 port map( D => n3772, CK => CLK
                           , Q => n_1352, QN => 
                           DataPath_RF_bus_reg_dataout_369_port);
   DataPath_RF_BLOCKi_20_Q_reg_17_inst : DFF_X1 port map( D => n3807, CK => CLK
                           , Q => n_1353, QN => 
                           DataPath_RF_bus_reg_dataout_401_port);
   DataPath_RF_BLOCKi_21_Q_reg_17_inst : DFF_X1 port map( D => n3842, CK => CLK
                           , Q => n_1354, QN => 
                           DataPath_RF_bus_reg_dataout_433_port);
   DataPath_RF_BLOCKi_22_Q_reg_17_inst : DFF_X1 port map( D => n3877, CK => CLK
                           , Q => n_1355, QN => 
                           DataPath_RF_bus_reg_dataout_465_port);
   DataPath_RF_BLOCKi_23_Q_reg_17_inst : DFF_X1 port map( D => n3926, CK => CLK
                           , Q => n_1356, QN => 
                           DataPath_RF_bus_reg_dataout_497_port);
   DataPath_RF_BLOCKi_24_Q_reg_17_inst : DFF_X1 port map( D => n3994, CK => CLK
                           , Q => n_1357, QN => 
                           DataPath_RF_bus_reg_dataout_529_port);
   DataPath_RF_BLOCKi_25_Q_reg_17_inst : DFF_X1 port map( D => n4048, CK => CLK
                           , Q => n_1358, QN => 
                           DataPath_RF_bus_reg_dataout_561_port);
   DataPath_RF_BLOCKi_26_Q_reg_17_inst : DFF_X1 port map( D => n4083, CK => CLK
                           , Q => n_1359, QN => 
                           DataPath_RF_bus_reg_dataout_593_port);
   DataPath_RF_BLOCKi_27_Q_reg_17_inst : DFF_X1 port map( D => n4118, CK => CLK
                           , Q => n_1360, QN => 
                           DataPath_RF_bus_reg_dataout_625_port);
   DataPath_RF_BLOCKi_28_Q_reg_17_inst : DFF_X1 port map( D => n4153, CK => CLK
                           , Q => n_1361, QN => 
                           DataPath_RF_bus_reg_dataout_657_port);
   DataPath_RF_BLOCKi_29_Q_reg_17_inst : DFF_X1 port map( D => n4188, CK => CLK
                           , Q => n_1362, QN => 
                           DataPath_RF_bus_reg_dataout_689_port);
   DataPath_RF_BLOCKi_30_Q_reg_17_inst : DFF_X1 port map( D => n4223, CK => CLK
                           , Q => n_1363, QN => 
                           DataPath_RF_bus_reg_dataout_721_port);
   DataPath_RF_BLOCKi_31_Q_reg_17_inst : DFF_X1 port map( D => n4258, CK => CLK
                           , Q => n_1364, QN => 
                           DataPath_RF_bus_reg_dataout_753_port);
   DataPath_RF_BLOCKi_32_Q_reg_17_inst : DFF_X1 port map( D => n4293, CK => CLK
                           , Q => n_1365, QN => 
                           DataPath_RF_bus_reg_dataout_785_port);
   DataPath_RF_BLOCKi_33_Q_reg_17_inst : DFF_X1 port map( D => n4328, CK => CLK
                           , Q => n_1366, QN => 
                           DataPath_RF_bus_reg_dataout_817_port);
   DataPath_RF_BLOCKi_34_Q_reg_17_inst : DFF_X1 port map( D => n4363, CK => CLK
                           , Q => n_1367, QN => 
                           DataPath_RF_bus_reg_dataout_849_port);
   DataPath_RF_BLOCKi_35_Q_reg_17_inst : DFF_X1 port map( D => n4398, CK => CLK
                           , Q => n_1368, QN => 
                           DataPath_RF_bus_reg_dataout_881_port);
   DataPath_RF_BLOCKi_36_Q_reg_17_inst : DFF_X1 port map( D => n4433, CK => CLK
                           , Q => n_1369, QN => 
                           DataPath_RF_bus_reg_dataout_913_port);
   DataPath_RF_BLOCKi_37_Q_reg_17_inst : DFF_X1 port map( D => n4468, CK => CLK
                           , Q => n_1370, QN => 
                           DataPath_RF_bus_reg_dataout_945_port);
   DataPath_RF_BLOCKi_38_Q_reg_17_inst : DFF_X1 port map( D => n4503, CK => CLK
                           , Q => n_1371, QN => 
                           DataPath_RF_bus_reg_dataout_977_port);
   DataPath_RF_BLOCKi_39_Q_reg_17_inst : DFF_X1 port map( D => n4538, CK => CLK
                           , Q => n_1372, QN => 
                           DataPath_RF_bus_reg_dataout_1009_port);
   DataPath_RF_BLOCKi_40_Q_reg_17_inst : DFF_X1 port map( D => n4587, CK => CLK
                           , Q => n_1373, QN => 
                           DataPath_RF_bus_reg_dataout_1041_port);
   DataPath_RF_BLOCKi_41_Q_reg_17_inst : DFF_X1 port map( D => n4641, CK => CLK
                           , Q => n_1374, QN => 
                           DataPath_RF_bus_reg_dataout_1073_port);
   DataPath_RF_BLOCKi_42_Q_reg_17_inst : DFF_X1 port map( D => n4676, CK => CLK
                           , Q => n_1375, QN => 
                           DataPath_RF_bus_reg_dataout_1105_port);
   DataPath_RF_BLOCKi_43_Q_reg_17_inst : DFF_X1 port map( D => n4711, CK => CLK
                           , Q => n_1376, QN => 
                           DataPath_RF_bus_reg_dataout_1137_port);
   DataPath_RF_BLOCKi_44_Q_reg_17_inst : DFF_X1 port map( D => n4746, CK => CLK
                           , Q => n_1377, QN => 
                           DataPath_RF_bus_reg_dataout_1169_port);
   DataPath_RF_BLOCKi_45_Q_reg_17_inst : DFF_X1 port map( D => n4781, CK => CLK
                           , Q => n_1378, QN => 
                           DataPath_RF_bus_reg_dataout_1201_port);
   DataPath_RF_BLOCKi_46_Q_reg_17_inst : DFF_X1 port map( D => n4816, CK => CLK
                           , Q => n_1379, QN => 
                           DataPath_RF_bus_reg_dataout_1233_port);
   DataPath_RF_BLOCKi_47_Q_reg_17_inst : DFF_X1 port map( D => n4851, CK => CLK
                           , Q => n_1380, QN => 
                           DataPath_RF_bus_reg_dataout_1265_port);
   DataPath_RF_BLOCKi_48_Q_reg_17_inst : DFF_X1 port map( D => n4886, CK => CLK
                           , Q => n_1381, QN => 
                           DataPath_RF_bus_reg_dataout_1297_port);
   DataPath_RF_BLOCKi_49_Q_reg_17_inst : DFF_X1 port map( D => n4921, CK => CLK
                           , Q => n_1382, QN => 
                           DataPath_RF_bus_reg_dataout_1329_port);
   DataPath_RF_BLOCKi_50_Q_reg_17_inst : DFF_X1 port map( D => n4956, CK => CLK
                           , Q => n_1383, QN => 
                           DataPath_RF_bus_reg_dataout_1361_port);
   DataPath_RF_BLOCKi_51_Q_reg_17_inst : DFF_X1 port map( D => n4991, CK => CLK
                           , Q => n_1384, QN => 
                           DataPath_RF_bus_reg_dataout_1393_port);
   DataPath_RF_BLOCKi_52_Q_reg_17_inst : DFF_X1 port map( D => n5026, CK => CLK
                           , Q => n_1385, QN => 
                           DataPath_RF_bus_reg_dataout_1425_port);
   DataPath_RF_BLOCKi_53_Q_reg_17_inst : DFF_X1 port map( D => n5061, CK => CLK
                           , Q => n_1386, QN => 
                           DataPath_RF_bus_reg_dataout_1457_port);
   DataPath_RF_BLOCKi_54_Q_reg_17_inst : DFF_X1 port map( D => n5096, CK => CLK
                           , Q => n_1387, QN => 
                           DataPath_RF_bus_reg_dataout_1489_port);
   DataPath_RF_BLOCKi_55_Q_reg_17_inst : DFF_X1 port map( D => n5131, CK => CLK
                           , Q => n_1388, QN => 
                           DataPath_RF_bus_reg_dataout_1521_port);
   DataPath_RF_BLOCKi_56_Q_reg_17_inst : DFF_X1 port map( D => n5180, CK => CLK
                           , Q => n_1389, QN => 
                           DataPath_RF_bus_reg_dataout_1553_port);
   DataPath_RF_BLOCKi_57_Q_reg_17_inst : DFF_X1 port map( D => n5233, CK => CLK
                           , Q => n_1390, QN => 
                           DataPath_RF_bus_reg_dataout_1585_port);
   DataPath_RF_BLOCKi_58_Q_reg_17_inst : DFF_X1 port map( D => n5269, CK => CLK
                           , Q => n_1391, QN => 
                           DataPath_RF_bus_reg_dataout_1617_port);
   DataPath_RF_BLOCKi_59_Q_reg_17_inst : DFF_X1 port map( D => n5304, CK => CLK
                           , Q => n_1392, QN => 
                           DataPath_RF_bus_reg_dataout_1649_port);
   DataPath_RF_BLOCKi_60_Q_reg_17_inst : DFF_X1 port map( D => n5339, CK => CLK
                           , Q => n_1393, QN => 
                           DataPath_RF_bus_reg_dataout_1681_port);
   DataPath_RF_BLOCKi_61_Q_reg_17_inst : DFF_X1 port map( D => n5374, CK => CLK
                           , Q => n_1394, QN => 
                           DataPath_RF_bus_reg_dataout_1713_port);
   DataPath_RF_BLOCKi_62_Q_reg_17_inst : DFF_X1 port map( D => n5409, CK => CLK
                           , Q => n_1395, QN => 
                           DataPath_RF_bus_reg_dataout_1745_port);
   DataPath_RF_BLOCKi_63_Q_reg_17_inst : DFF_X1 port map( D => n5444, CK => CLK
                           , Q => n_1396, QN => 
                           DataPath_RF_bus_reg_dataout_1777_port);
   DataPath_RF_BLOCKi_64_Q_reg_17_inst : DFF_X1 port map( D => n5479, CK => CLK
                           , Q => n_1397, QN => 
                           DataPath_RF_bus_reg_dataout_1809_port);
   DataPath_RF_BLOCKi_65_Q_reg_17_inst : DFF_X1 port map( D => n5514, CK => CLK
                           , Q => n_1398, QN => 
                           DataPath_RF_bus_reg_dataout_1841_port);
   DataPath_RF_BLOCKi_66_Q_reg_17_inst : DFF_X1 port map( D => n5549, CK => CLK
                           , Q => n_1399, QN => 
                           DataPath_RF_bus_reg_dataout_1873_port);
   DataPath_RF_BLOCKi_67_Q_reg_17_inst : DFF_X1 port map( D => n5584, CK => CLK
                           , Q => n_1400, QN => 
                           DataPath_RF_bus_reg_dataout_1905_port);
   DataPath_RF_BLOCKi_68_Q_reg_17_inst : DFF_X1 port map( D => n5623, CK => CLK
                           , Q => n_1401, QN => 
                           DataPath_RF_bus_reg_dataout_1937_port);
   DataPath_RF_BLOCKi_69_Q_reg_17_inst : DFF_X1 port map( D => n5660, CK => CLK
                           , Q => n_1402, QN => 
                           DataPath_RF_bus_reg_dataout_1969_port);
   DataPath_RF_BLOCKi_70_Q_reg_17_inst : DFF_X1 port map( D => n5697, CK => CLK
                           , Q => n_1403, QN => 
                           DataPath_RF_bus_reg_dataout_2001_port);
   DataPath_RF_BLOCKi_71_Q_reg_17_inst : DFF_X1 port map( D => n5734, CK => CLK
                           , Q => n_1404, QN => 
                           DataPath_RF_bus_reg_dataout_2033_port);
   DataPath_RF_BLOCKi_83_Q_reg_17_inst : DFF_X1 port map( D => n944, CK => CLK,
                           Q => n_1405, QN => 
                           DataPath_RF_bus_reg_dataout_2417_port);
   DataPath_RF_BLOCKi_84_Q_reg_17_inst : DFF_X1 port map( D => n984, CK => CLK,
                           Q => n_1406, QN => 
                           DataPath_RF_bus_reg_dataout_2449_port);
   DataPath_RF_BLOCKi_85_Q_reg_17_inst : DFF_X1 port map( D => n1021, CK => CLK
                           , Q => n_1407, QN => 
                           DataPath_RF_bus_reg_dataout_2481_port);
   DataPath_RF_BLOCKi_86_Q_reg_17_inst : DFF_X1 port map( D => n1058, CK => CLK
                           , Q => n_1408, QN => 
                           DataPath_RF_bus_reg_dataout_2513_port);
   DataPath_RF_BLOCKi_87_Q_reg_17_inst : DFF_X1 port map( D => n1095, CK => CLK
                           , Q => n_1409, QN => 
                           DataPath_RF_bus_reg_dataout_2545_port);
   DataPath_RF_BLOCKi_72_Q_reg_17_inst : DFF_X1 port map( D => n5771, CK => CLK
                           , Q => n_1410, QN => 
                           DataPath_RF_bus_reg_dataout_2065_port);
   DataPath_RF_BLOCKi_73_Q_reg_17_inst : DFF_X1 port map( D => n5810, CK => CLK
                           , Q => n_1411, QN => 
                           DataPath_RF_bus_reg_dataout_2097_port);
   DataPath_RF_BLOCKi_74_Q_reg_17_inst : DFF_X1 port map( D => n5846, CK => CLK
                           , Q => n_1412, QN => 
                           DataPath_RF_bus_reg_dataout_2129_port);
   DataPath_RF_BLOCKi_75_Q_reg_17_inst : DFF_X1 port map( D => n5882, CK => CLK
                           , Q => n_1413, QN => 
                           DataPath_RF_bus_reg_dataout_2161_port);
   DataPath_RF_BLOCKi_76_Q_reg_17_inst : DFF_X1 port map( D => n5918, CK => CLK
                           , Q => n_1414, QN => 
                           DataPath_RF_bus_reg_dataout_2193_port);
   DataPath_RF_BLOCKi_77_Q_reg_17_inst : DFF_X1 port map( D => n5954, CK => CLK
                           , Q => n_1415, QN => 
                           DataPath_RF_bus_reg_dataout_2225_port);
   DataPath_RF_BLOCKi_78_Q_reg_17_inst : DFF_X1 port map( D => n5990, CK => CLK
                           , Q => n_1416, QN => 
                           DataPath_RF_bus_reg_dataout_2257_port);
   DataPath_RF_BLOCKi_79_Q_reg_17_inst : DFF_X1 port map( D => n6026, CK => CLK
                           , Q => n_1417, QN => 
                           DataPath_RF_bus_reg_dataout_2289_port);
   DataPath_RF_BLOCKi_80_Q_reg_17_inst : DFF_X1 port map( D => n6063, CK => CLK
                           , Q => n_1418, QN => 
                           DataPath_RF_bus_reg_dataout_2321_port);
   DataPath_RF_BLOCKi_81_Q_reg_17_inst : DFF_X1 port map( D => n6099, CK => CLK
                           , Q => n_1419, QN => 
                           DataPath_RF_bus_reg_dataout_2353_port);
   DataPath_RF_BLOCKi_82_Q_reg_17_inst : DFF_X1 port map( D => n6133, CK => CLK
                           , Q => n_1420, QN => 
                           DataPath_RF_bus_reg_dataout_2385_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_25_inst : DFF_X1 port map( D => n2184, CK 
                           => CLK, Q => n_1421, QN => 
                           DataPath_i_REG_LDSTR_OUT_25_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_9_inst : DFF_X1 port map( D => n2200, CK =>
                           CLK, Q => n_1422, QN => 
                           DataPath_i_REG_LDSTR_OUT_9_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_9_inst : DFF_X1 port map( D => n6790, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_41_port,
                           QN => n608);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_9_inst : DFF_X1 port map( D => n6822, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_73_port,
                           QN => n640);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_9_inst : DFF_X1 port map( D => n6854, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_105_port
                           , QN => n672);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_9_inst : DFF_X1 port map( D => n6886, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_137_port
                           , QN => n704);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_9_inst : DFF_X1 port map( D => n6918, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_169_port
                           , QN => n736);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_9_inst : DFF_X1 port map( D => n6950, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_201_port
                           , QN => n768);
   DataPath_RF_BLOCKi_8_Q_reg_9_inst : DFF_X1 port map( D => n3354, CK => CLK, 
                           Q => n_1423, QN => 
                           DataPath_RF_bus_reg_dataout_9_port);
   DataPath_RF_BLOCKi_9_Q_reg_9_inst : DFF_X1 port map( D => n3403, CK => CLK, 
                           Q => n_1424, QN => 
                           DataPath_RF_bus_reg_dataout_41_port);
   DataPath_RF_BLOCKi_10_Q_reg_9_inst : DFF_X1 port map( D => n3441, CK => CLK,
                           Q => n_1425, QN => 
                           DataPath_RF_bus_reg_dataout_73_port);
   DataPath_RF_BLOCKi_11_Q_reg_9_inst : DFF_X1 port map( D => n3479, CK => CLK,
                           Q => n_1426, QN => 
                           DataPath_RF_bus_reg_dataout_105_port);
   DataPath_RF_BLOCKi_12_Q_reg_9_inst : DFF_X1 port map( D => n3517, CK => CLK,
                           Q => n_1427, QN => 
                           DataPath_RF_bus_reg_dataout_137_port);
   DataPath_RF_BLOCKi_13_Q_reg_9_inst : DFF_X1 port map( D => n3555, CK => CLK,
                           Q => n_1428, QN => 
                           DataPath_RF_bus_reg_dataout_169_port);
   DataPath_RF_BLOCKi_14_Q_reg_9_inst : DFF_X1 port map( D => n3593, CK => CLK,
                           Q => n_1429, QN => 
                           DataPath_RF_bus_reg_dataout_201_port);
   DataPath_RF_BLOCKi_15_Q_reg_9_inst : DFF_X1 port map( D => n3631, CK => CLK,
                           Q => n_1430, QN => 
                           DataPath_RF_bus_reg_dataout_233_port);
   DataPath_RF_BLOCKi_16_Q_reg_9_inst : DFF_X1 port map( D => n3669, CK => CLK,
                           Q => n_1431, QN => 
                           DataPath_RF_bus_reg_dataout_265_port);
   DataPath_RF_BLOCKi_17_Q_reg_9_inst : DFF_X1 port map( D => n3706, CK => CLK,
                           Q => n_1432, QN => 
                           DataPath_RF_bus_reg_dataout_297_port);
   DataPath_RF_BLOCKi_18_Q_reg_9_inst : DFF_X1 port map( D => n3743, CK => CLK,
                           Q => n_1433, QN => 
                           DataPath_RF_bus_reg_dataout_329_port);
   DataPath_RF_BLOCKi_19_Q_reg_9_inst : DFF_X1 port map( D => n3780, CK => CLK,
                           Q => n_1434, QN => 
                           DataPath_RF_bus_reg_dataout_361_port);
   DataPath_RF_BLOCKi_20_Q_reg_9_inst : DFF_X1 port map( D => n3815, CK => CLK,
                           Q => n_1435, QN => 
                           DataPath_RF_bus_reg_dataout_393_port);
   DataPath_RF_BLOCKi_21_Q_reg_9_inst : DFF_X1 port map( D => n3850, CK => CLK,
                           Q => n_1436, QN => 
                           DataPath_RF_bus_reg_dataout_425_port);
   DataPath_RF_BLOCKi_22_Q_reg_9_inst : DFF_X1 port map( D => n3885, CK => CLK,
                           Q => n_1437, QN => 
                           DataPath_RF_bus_reg_dataout_457_port);
   DataPath_RF_BLOCKi_23_Q_reg_9_inst : DFF_X1 port map( D => n3942, CK => CLK,
                           Q => n_1438, QN => 
                           DataPath_RF_bus_reg_dataout_489_port);
   DataPath_RF_BLOCKi_24_Q_reg_9_inst : DFF_X1 port map( D => n4010, CK => CLK,
                           Q => n_1439, QN => 
                           DataPath_RF_bus_reg_dataout_521_port);
   DataPath_RF_BLOCKi_25_Q_reg_9_inst : DFF_X1 port map( D => n4056, CK => CLK,
                           Q => n_1440, QN => 
                           DataPath_RF_bus_reg_dataout_553_port);
   DataPath_RF_BLOCKi_26_Q_reg_9_inst : DFF_X1 port map( D => n4091, CK => CLK,
                           Q => n_1441, QN => 
                           DataPath_RF_bus_reg_dataout_585_port);
   DataPath_RF_BLOCKi_27_Q_reg_9_inst : DFF_X1 port map( D => n4126, CK => CLK,
                           Q => n_1442, QN => 
                           DataPath_RF_bus_reg_dataout_617_port);
   DataPath_RF_BLOCKi_28_Q_reg_9_inst : DFF_X1 port map( D => n4161, CK => CLK,
                           Q => n_1443, QN => 
                           DataPath_RF_bus_reg_dataout_649_port);
   DataPath_RF_BLOCKi_29_Q_reg_9_inst : DFF_X1 port map( D => n4196, CK => CLK,
                           Q => n_1444, QN => 
                           DataPath_RF_bus_reg_dataout_681_port);
   DataPath_RF_BLOCKi_30_Q_reg_9_inst : DFF_X1 port map( D => n4231, CK => CLK,
                           Q => n_1445, QN => 
                           DataPath_RF_bus_reg_dataout_713_port);
   DataPath_RF_BLOCKi_31_Q_reg_9_inst : DFF_X1 port map( D => n4266, CK => CLK,
                           Q => n_1446, QN => 
                           DataPath_RF_bus_reg_dataout_745_port);
   DataPath_RF_BLOCKi_32_Q_reg_9_inst : DFF_X1 port map( D => n4301, CK => CLK,
                           Q => n_1447, QN => 
                           DataPath_RF_bus_reg_dataout_777_port);
   DataPath_RF_BLOCKi_33_Q_reg_9_inst : DFF_X1 port map( D => n4336, CK => CLK,
                           Q => n_1448, QN => 
                           DataPath_RF_bus_reg_dataout_809_port);
   DataPath_RF_BLOCKi_34_Q_reg_9_inst : DFF_X1 port map( D => n4371, CK => CLK,
                           Q => n_1449, QN => 
                           DataPath_RF_bus_reg_dataout_841_port);
   DataPath_RF_BLOCKi_35_Q_reg_9_inst : DFF_X1 port map( D => n4406, CK => CLK,
                           Q => n_1450, QN => 
                           DataPath_RF_bus_reg_dataout_873_port);
   DataPath_RF_BLOCKi_36_Q_reg_9_inst : DFF_X1 port map( D => n4441, CK => CLK,
                           Q => n_1451, QN => 
                           DataPath_RF_bus_reg_dataout_905_port);
   DataPath_RF_BLOCKi_37_Q_reg_9_inst : DFF_X1 port map( D => n4476, CK => CLK,
                           Q => n_1452, QN => 
                           DataPath_RF_bus_reg_dataout_937_port);
   DataPath_RF_BLOCKi_38_Q_reg_9_inst : DFF_X1 port map( D => n4511, CK => CLK,
                           Q => n_1453, QN => 
                           DataPath_RF_bus_reg_dataout_969_port);
   DataPath_RF_BLOCKi_39_Q_reg_9_inst : DFF_X1 port map( D => n4546, CK => CLK,
                           Q => n_1454, QN => 
                           DataPath_RF_bus_reg_dataout_1001_port);
   DataPath_RF_BLOCKi_40_Q_reg_9_inst : DFF_X1 port map( D => n4603, CK => CLK,
                           Q => n_1455, QN => 
                           DataPath_RF_bus_reg_dataout_1033_port);
   DataPath_RF_BLOCKi_41_Q_reg_9_inst : DFF_X1 port map( D => n4649, CK => CLK,
                           Q => n_1456, QN => 
                           DataPath_RF_bus_reg_dataout_1065_port);
   DataPath_RF_BLOCKi_42_Q_reg_9_inst : DFF_X1 port map( D => n4684, CK => CLK,
                           Q => n_1457, QN => 
                           DataPath_RF_bus_reg_dataout_1097_port);
   DataPath_RF_BLOCKi_43_Q_reg_9_inst : DFF_X1 port map( D => n4719, CK => CLK,
                           Q => n_1458, QN => 
                           DataPath_RF_bus_reg_dataout_1129_port);
   DataPath_RF_BLOCKi_44_Q_reg_9_inst : DFF_X1 port map( D => n4754, CK => CLK,
                           Q => n_1459, QN => 
                           DataPath_RF_bus_reg_dataout_1161_port);
   DataPath_RF_BLOCKi_45_Q_reg_9_inst : DFF_X1 port map( D => n4789, CK => CLK,
                           Q => n_1460, QN => 
                           DataPath_RF_bus_reg_dataout_1193_port);
   DataPath_RF_BLOCKi_46_Q_reg_9_inst : DFF_X1 port map( D => n4824, CK => CLK,
                           Q => n_1461, QN => 
                           DataPath_RF_bus_reg_dataout_1225_port);
   DataPath_RF_BLOCKi_47_Q_reg_9_inst : DFF_X1 port map( D => n4859, CK => CLK,
                           Q => n_1462, QN => 
                           DataPath_RF_bus_reg_dataout_1257_port);
   DataPath_RF_BLOCKi_48_Q_reg_9_inst : DFF_X1 port map( D => n4894, CK => CLK,
                           Q => n_1463, QN => 
                           DataPath_RF_bus_reg_dataout_1289_port);
   DataPath_RF_BLOCKi_49_Q_reg_9_inst : DFF_X1 port map( D => n4929, CK => CLK,
                           Q => n_1464, QN => 
                           DataPath_RF_bus_reg_dataout_1321_port);
   DataPath_RF_BLOCKi_50_Q_reg_9_inst : DFF_X1 port map( D => n4964, CK => CLK,
                           Q => n_1465, QN => 
                           DataPath_RF_bus_reg_dataout_1353_port);
   DataPath_RF_BLOCKi_51_Q_reg_9_inst : DFF_X1 port map( D => n4999, CK => CLK,
                           Q => n_1466, QN => 
                           DataPath_RF_bus_reg_dataout_1385_port);
   DataPath_RF_BLOCKi_52_Q_reg_9_inst : DFF_X1 port map( D => n5034, CK => CLK,
                           Q => n_1467, QN => 
                           DataPath_RF_bus_reg_dataout_1417_port);
   DataPath_RF_BLOCKi_53_Q_reg_9_inst : DFF_X1 port map( D => n5069, CK => CLK,
                           Q => n_1468, QN => 
                           DataPath_RF_bus_reg_dataout_1449_port);
   DataPath_RF_BLOCKi_54_Q_reg_9_inst : DFF_X1 port map( D => n5104, CK => CLK,
                           Q => n_1469, QN => 
                           DataPath_RF_bus_reg_dataout_1481_port);
   DataPath_RF_BLOCKi_55_Q_reg_9_inst : DFF_X1 port map( D => n5139, CK => CLK,
                           Q => n_1470, QN => 
                           DataPath_RF_bus_reg_dataout_1513_port);
   DataPath_RF_BLOCKi_56_Q_reg_9_inst : DFF_X1 port map( D => n5196, CK => CLK,
                           Q => n_1471, QN => 
                           DataPath_RF_bus_reg_dataout_1545_port);
   DataPath_RF_BLOCKi_57_Q_reg_9_inst : DFF_X1 port map( D => n5241, CK => CLK,
                           Q => n_1472, QN => 
                           DataPath_RF_bus_reg_dataout_1577_port);
   DataPath_RF_BLOCKi_58_Q_reg_9_inst : DFF_X1 port map( D => n5277, CK => CLK,
                           Q => n_1473, QN => 
                           DataPath_RF_bus_reg_dataout_1609_port);
   DataPath_RF_BLOCKi_59_Q_reg_9_inst : DFF_X1 port map( D => n5312, CK => CLK,
                           Q => n_1474, QN => 
                           DataPath_RF_bus_reg_dataout_1641_port);
   DataPath_RF_BLOCKi_60_Q_reg_9_inst : DFF_X1 port map( D => n5347, CK => CLK,
                           Q => n_1475, QN => 
                           DataPath_RF_bus_reg_dataout_1673_port);
   DataPath_RF_BLOCKi_61_Q_reg_9_inst : DFF_X1 port map( D => n5382, CK => CLK,
                           Q => n_1476, QN => 
                           DataPath_RF_bus_reg_dataout_1705_port);
   DataPath_RF_BLOCKi_62_Q_reg_9_inst : DFF_X1 port map( D => n5417, CK => CLK,
                           Q => n_1477, QN => 
                           DataPath_RF_bus_reg_dataout_1737_port);
   DataPath_RF_BLOCKi_63_Q_reg_9_inst : DFF_X1 port map( D => n5452, CK => CLK,
                           Q => n_1478, QN => 
                           DataPath_RF_bus_reg_dataout_1769_port);
   DataPath_RF_BLOCKi_64_Q_reg_9_inst : DFF_X1 port map( D => n5487, CK => CLK,
                           Q => n_1479, QN => 
                           DataPath_RF_bus_reg_dataout_1801_port);
   DataPath_RF_BLOCKi_65_Q_reg_9_inst : DFF_X1 port map( D => n5522, CK => CLK,
                           Q => n_1480, QN => 
                           DataPath_RF_bus_reg_dataout_1833_port);
   DataPath_RF_BLOCKi_66_Q_reg_9_inst : DFF_X1 port map( D => n5557, CK => CLK,
                           Q => n_1481, QN => 
                           DataPath_RF_bus_reg_dataout_1865_port);
   DataPath_RF_BLOCKi_67_Q_reg_9_inst : DFF_X1 port map( D => n5592, CK => CLK,
                           Q => n_1482, QN => 
                           DataPath_RF_bus_reg_dataout_1897_port);
   DataPath_RF_BLOCKi_68_Q_reg_9_inst : DFF_X1 port map( D => n5631, CK => CLK,
                           Q => n_1483, QN => 
                           DataPath_RF_bus_reg_dataout_1929_port);
   DataPath_RF_BLOCKi_69_Q_reg_9_inst : DFF_X1 port map( D => n5668, CK => CLK,
                           Q => n_1484, QN => 
                           DataPath_RF_bus_reg_dataout_1961_port);
   DataPath_RF_BLOCKi_70_Q_reg_9_inst : DFF_X1 port map( D => n5705, CK => CLK,
                           Q => n_1485, QN => 
                           DataPath_RF_bus_reg_dataout_1993_port);
   DataPath_RF_BLOCKi_71_Q_reg_9_inst : DFF_X1 port map( D => n5742, CK => CLK,
                           Q => n_1486, QN => 
                           DataPath_RF_bus_reg_dataout_2025_port);
   DataPath_RF_BLOCKi_82_Q_reg_9_inst : DFF_X1 port map( D => n894, CK => CLK, 
                           Q => n_1487, QN => 
                           DataPath_RF_bus_reg_dataout_2377_port);
   DataPath_RF_BLOCKi_83_Q_reg_9_inst : DFF_X1 port map( D => n954, CK => CLK, 
                           Q => n_1488, QN => 
                           DataPath_RF_bus_reg_dataout_2409_port);
   DataPath_RF_BLOCKi_84_Q_reg_9_inst : DFF_X1 port map( D => n992, CK => CLK, 
                           Q => n_1489, QN => 
                           DataPath_RF_bus_reg_dataout_2441_port);
   DataPath_RF_BLOCKi_85_Q_reg_9_inst : DFF_X1 port map( D => n1029, CK => CLK,
                           Q => n_1490, QN => 
                           DataPath_RF_bus_reg_dataout_2473_port);
   DataPath_RF_BLOCKi_86_Q_reg_9_inst : DFF_X1 port map( D => n1066, CK => CLK,
                           Q => n_1491, QN => 
                           DataPath_RF_bus_reg_dataout_2505_port);
   DataPath_RF_BLOCKi_87_Q_reg_9_inst : DFF_X1 port map( D => n1103, CK => CLK,
                           Q => n_1492, QN => 
                           DataPath_RF_bus_reg_dataout_2537_port);
   DataPath_RF_BLOCKi_72_Q_reg_9_inst : DFF_X1 port map( D => n5779, CK => CLK,
                           Q => n_1493, QN => 
                           DataPath_RF_bus_reg_dataout_2057_port);
   DataPath_RF_BLOCKi_73_Q_reg_9_inst : DFF_X1 port map( D => n5818, CK => CLK,
                           Q => n_1494, QN => 
                           DataPath_RF_bus_reg_dataout_2089_port);
   DataPath_RF_BLOCKi_74_Q_reg_9_inst : DFF_X1 port map( D => n5854, CK => CLK,
                           Q => n_1495, QN => 
                           DataPath_RF_bus_reg_dataout_2121_port);
   DataPath_RF_BLOCKi_75_Q_reg_9_inst : DFF_X1 port map( D => n5890, CK => CLK,
                           Q => n_1496, QN => 
                           DataPath_RF_bus_reg_dataout_2153_port);
   DataPath_RF_BLOCKi_76_Q_reg_9_inst : DFF_X1 port map( D => n5926, CK => CLK,
                           Q => n_1497, QN => 
                           DataPath_RF_bus_reg_dataout_2185_port);
   DataPath_RF_BLOCKi_77_Q_reg_9_inst : DFF_X1 port map( D => n5962, CK => CLK,
                           Q => n_1498, QN => 
                           DataPath_RF_bus_reg_dataout_2217_port);
   DataPath_RF_BLOCKi_78_Q_reg_9_inst : DFF_X1 port map( D => n5998, CK => CLK,
                           Q => n_1499, QN => 
                           DataPath_RF_bus_reg_dataout_2249_port);
   DataPath_RF_BLOCKi_79_Q_reg_9_inst : DFF_X1 port map( D => n6034, CK => CLK,
                           Q => n_1500, QN => 
                           DataPath_RF_bus_reg_dataout_2281_port);
   DataPath_RF_BLOCKi_80_Q_reg_9_inst : DFF_X1 port map( D => n6071, CK => CLK,
                           Q => n_1501, QN => 
                           DataPath_RF_bus_reg_dataout_2313_port);
   DataPath_RF_BLOCKi_81_Q_reg_9_inst : DFF_X1 port map( D => n6107, CK => CLK,
                           Q => n_1502, QN => 
                           DataPath_RF_bus_reg_dataout_2345_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_1_inst : DFF_X1 port map( D => n2208, CK =>
                           CLK, Q => n_1503, QN => 
                           DataPath_i_REG_LDSTR_OUT_1_port);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_1_inst : DFF_X1 port map( D => n6862, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_97_port,
                           QN => n664);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_1_inst : DFF_X1 port map( D => n6894, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_129_port
                           , QN => n696);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_1_inst : DFF_X1 port map( D => n6958, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_193_port
                           , QN => n760);
   DataPath_RF_BLOCKi_8_Q_reg_1_inst : DFF_X1 port map( D => n3370, CK => CLK, 
                           Q => n_1504, QN => 
                           DataPath_RF_bus_reg_dataout_1_port);
   DataPath_RF_BLOCKi_9_Q_reg_1_inst : DFF_X1 port map( D => n3411, CK => CLK, 
                           Q => n_1505, QN => 
                           DataPath_RF_bus_reg_dataout_33_port);
   DataPath_RF_BLOCKi_10_Q_reg_1_inst : DFF_X1 port map( D => n3449, CK => CLK,
                           Q => n_1506, QN => 
                           DataPath_RF_bus_reg_dataout_65_port);
   DataPath_RF_BLOCKi_11_Q_reg_1_inst : DFF_X1 port map( D => n3487, CK => CLK,
                           Q => n_1507, QN => 
                           DataPath_RF_bus_reg_dataout_97_port);
   DataPath_RF_BLOCKi_12_Q_reg_1_inst : DFF_X1 port map( D => n3525, CK => CLK,
                           Q => n_1508, QN => 
                           DataPath_RF_bus_reg_dataout_129_port);
   DataPath_RF_BLOCKi_13_Q_reg_1_inst : DFF_X1 port map( D => n3563, CK => CLK,
                           Q => n_1509, QN => 
                           DataPath_RF_bus_reg_dataout_161_port);
   DataPath_RF_BLOCKi_14_Q_reg_1_inst : DFF_X1 port map( D => n3601, CK => CLK,
                           Q => n_1510, QN => 
                           DataPath_RF_bus_reg_dataout_193_port);
   DataPath_RF_BLOCKi_15_Q_reg_1_inst : DFF_X1 port map( D => n3639, CK => CLK,
                           Q => n_1511, QN => 
                           DataPath_RF_bus_reg_dataout_225_port);
   DataPath_RF_BLOCKi_16_Q_reg_1_inst : DFF_X1 port map( D => n3677, CK => CLK,
                           Q => n_1512, QN => 
                           DataPath_RF_bus_reg_dataout_257_port);
   DataPath_RF_BLOCKi_17_Q_reg_1_inst : DFF_X1 port map( D => n3714, CK => CLK,
                           Q => n_1513, QN => 
                           DataPath_RF_bus_reg_dataout_289_port);
   DataPath_RF_BLOCKi_18_Q_reg_1_inst : DFF_X1 port map( D => n3751, CK => CLK,
                           Q => n_1514, QN => 
                           DataPath_RF_bus_reg_dataout_321_port);
   DataPath_RF_BLOCKi_19_Q_reg_1_inst : DFF_X1 port map( D => n3788, CK => CLK,
                           Q => n_1515, QN => 
                           DataPath_RF_bus_reg_dataout_353_port);
   DataPath_RF_BLOCKi_20_Q_reg_1_inst : DFF_X1 port map( D => n3823, CK => CLK,
                           Q => n_1516, QN => 
                           DataPath_RF_bus_reg_dataout_385_port);
   DataPath_RF_BLOCKi_21_Q_reg_1_inst : DFF_X1 port map( D => n3858, CK => CLK,
                           Q => n_1517, QN => 
                           DataPath_RF_bus_reg_dataout_417_port);
   DataPath_RF_BLOCKi_22_Q_reg_1_inst : DFF_X1 port map( D => n3893, CK => CLK,
                           Q => n_1518, QN => 
                           DataPath_RF_bus_reg_dataout_449_port);
   DataPath_RF_BLOCKi_23_Q_reg_1_inst : DFF_X1 port map( D => n3958, CK => CLK,
                           Q => n_1519, QN => 
                           DataPath_RF_bus_reg_dataout_481_port);
   DataPath_RF_BLOCKi_24_Q_reg_1_inst : DFF_X1 port map( D => n4026, CK => CLK,
                           Q => n_1520, QN => 
                           DataPath_RF_bus_reg_dataout_513_port);
   DataPath_RF_BLOCKi_25_Q_reg_1_inst : DFF_X1 port map( D => n4064, CK => CLK,
                           Q => n_1521, QN => 
                           DataPath_RF_bus_reg_dataout_545_port);
   DataPath_RF_BLOCKi_26_Q_reg_1_inst : DFF_X1 port map( D => n4099, CK => CLK,
                           Q => n_1522, QN => 
                           DataPath_RF_bus_reg_dataout_577_port);
   DataPath_RF_BLOCKi_27_Q_reg_1_inst : DFF_X1 port map( D => n4134, CK => CLK,
                           Q => n_1523, QN => 
                           DataPath_RF_bus_reg_dataout_609_port);
   DataPath_RF_BLOCKi_28_Q_reg_1_inst : DFF_X1 port map( D => n4169, CK => CLK,
                           Q => n_1524, QN => 
                           DataPath_RF_bus_reg_dataout_641_port);
   DataPath_RF_BLOCKi_29_Q_reg_1_inst : DFF_X1 port map( D => n4204, CK => CLK,
                           Q => n_1525, QN => 
                           DataPath_RF_bus_reg_dataout_673_port);
   DataPath_RF_BLOCKi_30_Q_reg_1_inst : DFF_X1 port map( D => n4239, CK => CLK,
                           Q => n_1526, QN => 
                           DataPath_RF_bus_reg_dataout_705_port);
   DataPath_RF_BLOCKi_31_Q_reg_1_inst : DFF_X1 port map( D => n4274, CK => CLK,
                           Q => n_1527, QN => 
                           DataPath_RF_bus_reg_dataout_737_port);
   DataPath_RF_BLOCKi_32_Q_reg_1_inst : DFF_X1 port map( D => n4309, CK => CLK,
                           Q => n_1528, QN => 
                           DataPath_RF_bus_reg_dataout_769_port);
   DataPath_RF_BLOCKi_33_Q_reg_1_inst : DFF_X1 port map( D => n4344, CK => CLK,
                           Q => n_1529, QN => 
                           DataPath_RF_bus_reg_dataout_801_port);
   DataPath_RF_BLOCKi_34_Q_reg_1_inst : DFF_X1 port map( D => n4379, CK => CLK,
                           Q => n_1530, QN => 
                           DataPath_RF_bus_reg_dataout_833_port);
   DataPath_RF_BLOCKi_35_Q_reg_1_inst : DFF_X1 port map( D => n4414, CK => CLK,
                           Q => n_1531, QN => 
                           DataPath_RF_bus_reg_dataout_865_port);
   DataPath_RF_BLOCKi_36_Q_reg_1_inst : DFF_X1 port map( D => n4449, CK => CLK,
                           Q => n_1532, QN => 
                           DataPath_RF_bus_reg_dataout_897_port);
   DataPath_RF_BLOCKi_37_Q_reg_1_inst : DFF_X1 port map( D => n4484, CK => CLK,
                           Q => n_1533, QN => 
                           DataPath_RF_bus_reg_dataout_929_port);
   DataPath_RF_BLOCKi_38_Q_reg_1_inst : DFF_X1 port map( D => n4519, CK => CLK,
                           Q => n_1534, QN => 
                           DataPath_RF_bus_reg_dataout_961_port);
   DataPath_RF_BLOCKi_39_Q_reg_1_inst : DFF_X1 port map( D => n4554, CK => CLK,
                           Q => n_1535, QN => 
                           DataPath_RF_bus_reg_dataout_993_port);
   DataPath_RF_BLOCKi_40_Q_reg_1_inst : DFF_X1 port map( D => n4619, CK => CLK,
                           Q => n_1536, QN => 
                           DataPath_RF_bus_reg_dataout_1025_port);
   DataPath_RF_BLOCKi_41_Q_reg_1_inst : DFF_X1 port map( D => n4657, CK => CLK,
                           Q => n_1537, QN => 
                           DataPath_RF_bus_reg_dataout_1057_port);
   DataPath_RF_BLOCKi_42_Q_reg_1_inst : DFF_X1 port map( D => n4692, CK => CLK,
                           Q => n_1538, QN => 
                           DataPath_RF_bus_reg_dataout_1089_port);
   DataPath_RF_BLOCKi_43_Q_reg_1_inst : DFF_X1 port map( D => n4727, CK => CLK,
                           Q => n_1539, QN => 
                           DataPath_RF_bus_reg_dataout_1121_port);
   DataPath_RF_BLOCKi_44_Q_reg_1_inst : DFF_X1 port map( D => n4762, CK => CLK,
                           Q => n_1540, QN => 
                           DataPath_RF_bus_reg_dataout_1153_port);
   DataPath_RF_BLOCKi_45_Q_reg_1_inst : DFF_X1 port map( D => n4797, CK => CLK,
                           Q => n_1541, QN => 
                           DataPath_RF_bus_reg_dataout_1185_port);
   DataPath_RF_BLOCKi_46_Q_reg_1_inst : DFF_X1 port map( D => n4832, CK => CLK,
                           Q => n_1542, QN => 
                           DataPath_RF_bus_reg_dataout_1217_port);
   DataPath_RF_BLOCKi_47_Q_reg_1_inst : DFF_X1 port map( D => n4867, CK => CLK,
                           Q => n_1543, QN => 
                           DataPath_RF_bus_reg_dataout_1249_port);
   DataPath_RF_BLOCKi_48_Q_reg_1_inst : DFF_X1 port map( D => n4902, CK => CLK,
                           Q => n_1544, QN => 
                           DataPath_RF_bus_reg_dataout_1281_port);
   DataPath_RF_BLOCKi_49_Q_reg_1_inst : DFF_X1 port map( D => n4937, CK => CLK,
                           Q => n_1545, QN => 
                           DataPath_RF_bus_reg_dataout_1313_port);
   DataPath_RF_BLOCKi_50_Q_reg_1_inst : DFF_X1 port map( D => n4972, CK => CLK,
                           Q => n_1546, QN => 
                           DataPath_RF_bus_reg_dataout_1345_port);
   DataPath_RF_BLOCKi_51_Q_reg_1_inst : DFF_X1 port map( D => n5007, CK => CLK,
                           Q => n_1547, QN => 
                           DataPath_RF_bus_reg_dataout_1377_port);
   DataPath_RF_BLOCKi_52_Q_reg_1_inst : DFF_X1 port map( D => n5042, CK => CLK,
                           Q => n_1548, QN => 
                           DataPath_RF_bus_reg_dataout_1409_port);
   DataPath_RF_BLOCKi_53_Q_reg_1_inst : DFF_X1 port map( D => n5077, CK => CLK,
                           Q => n_1549, QN => 
                           DataPath_RF_bus_reg_dataout_1441_port);
   DataPath_RF_BLOCKi_54_Q_reg_1_inst : DFF_X1 port map( D => n5112, CK => CLK,
                           Q => n_1550, QN => 
                           DataPath_RF_bus_reg_dataout_1473_port);
   DataPath_RF_BLOCKi_55_Q_reg_1_inst : DFF_X1 port map( D => n5147, CK => CLK,
                           Q => n_1551, QN => 
                           DataPath_RF_bus_reg_dataout_1505_port);
   DataPath_RF_BLOCKi_56_Q_reg_1_inst : DFF_X1 port map( D => n5212, CK => CLK,
                           Q => n_1552, QN => 
                           DataPath_RF_bus_reg_dataout_1537_port);
   DataPath_RF_BLOCKi_57_Q_reg_1_inst : DFF_X1 port map( D => n5249, CK => CLK,
                           Q => n_1553, QN => 
                           DataPath_RF_bus_reg_dataout_1569_port);
   DataPath_RF_BLOCKi_58_Q_reg_1_inst : DFF_X1 port map( D => n5285, CK => CLK,
                           Q => n_1554, QN => 
                           DataPath_RF_bus_reg_dataout_1601_port);
   DataPath_RF_BLOCKi_59_Q_reg_1_inst : DFF_X1 port map( D => n5320, CK => CLK,
                           Q => n_1555, QN => 
                           DataPath_RF_bus_reg_dataout_1633_port);
   DataPath_RF_BLOCKi_60_Q_reg_1_inst : DFF_X1 port map( D => n5355, CK => CLK,
                           Q => n_1556, QN => 
                           DataPath_RF_bus_reg_dataout_1665_port);
   DataPath_RF_BLOCKi_61_Q_reg_1_inst : DFF_X1 port map( D => n5390, CK => CLK,
                           Q => n_1557, QN => 
                           DataPath_RF_bus_reg_dataout_1697_port);
   DataPath_RF_BLOCKi_62_Q_reg_1_inst : DFF_X1 port map( D => n5425, CK => CLK,
                           Q => n_1558, QN => 
                           DataPath_RF_bus_reg_dataout_1729_port);
   DataPath_RF_BLOCKi_63_Q_reg_1_inst : DFF_X1 port map( D => n5460, CK => CLK,
                           Q => n_1559, QN => 
                           DataPath_RF_bus_reg_dataout_1761_port);
   DataPath_RF_BLOCKi_64_Q_reg_1_inst : DFF_X1 port map( D => n5495, CK => CLK,
                           Q => n_1560, QN => 
                           DataPath_RF_bus_reg_dataout_1793_port);
   DataPath_RF_BLOCKi_65_Q_reg_1_inst : DFF_X1 port map( D => n5530, CK => CLK,
                           Q => n_1561, QN => 
                           DataPath_RF_bus_reg_dataout_1825_port);
   DataPath_RF_BLOCKi_66_Q_reg_1_inst : DFF_X1 port map( D => n5565, CK => CLK,
                           Q => n_1562, QN => 
                           DataPath_RF_bus_reg_dataout_1857_port);
   DataPath_RF_BLOCKi_67_Q_reg_1_inst : DFF_X1 port map( D => n5600, CK => CLK,
                           Q => n_1563, QN => 
                           DataPath_RF_bus_reg_dataout_1889_port);
   DataPath_RF_BLOCKi_68_Q_reg_1_inst : DFF_X1 port map( D => n5639, CK => CLK,
                           Q => n_1564, QN => 
                           DataPath_RF_bus_reg_dataout_1921_port);
   DataPath_RF_BLOCKi_69_Q_reg_1_inst : DFF_X1 port map( D => n5676, CK => CLK,
                           Q => n_1565, QN => 
                           DataPath_RF_bus_reg_dataout_1953_port);
   DataPath_RF_BLOCKi_70_Q_reg_1_inst : DFF_X1 port map( D => n5713, CK => CLK,
                           Q => n_1566, QN => 
                           DataPath_RF_bus_reg_dataout_1985_port);
   DataPath_RF_BLOCKi_71_Q_reg_1_inst : DFF_X1 port map( D => n5750, CK => CLK,
                           Q => n_1567, QN => 
                           DataPath_RF_bus_reg_dataout_2017_port);
   DataPath_RF_BLOCKi_82_Q_reg_1_inst : DFF_X1 port map( D => n910, CK => CLK, 
                           Q => n_1568, QN => 
                           DataPath_RF_bus_reg_dataout_2369_port);
   DataPath_RF_BLOCKi_83_Q_reg_1_inst : DFF_X1 port map( D => n962, CK => CLK, 
                           Q => n_1569, QN => 
                           DataPath_RF_bus_reg_dataout_2401_port);
   DataPath_RF_BLOCKi_84_Q_reg_1_inst : DFF_X1 port map( D => n1000, CK => CLK,
                           Q => n_1570, QN => 
                           DataPath_RF_bus_reg_dataout_2433_port);
   DataPath_RF_BLOCKi_85_Q_reg_1_inst : DFF_X1 port map( D => n1037, CK => CLK,
                           Q => n_1571, QN => 
                           DataPath_RF_bus_reg_dataout_2465_port);
   DataPath_RF_BLOCKi_86_Q_reg_1_inst : DFF_X1 port map( D => n1074, CK => CLK,
                           Q => n_1572, QN => 
                           DataPath_RF_bus_reg_dataout_2497_port);
   DataPath_RF_BLOCKi_87_Q_reg_1_inst : DFF_X1 port map( D => n1111, CK => CLK,
                           Q => n_1573, QN => 
                           DataPath_RF_bus_reg_dataout_2529_port);
   DataPath_RF_BLOCKi_72_Q_reg_1_inst : DFF_X1 port map( D => n5787, CK => CLK,
                           Q => n_1574, QN => 
                           DataPath_RF_bus_reg_dataout_2049_port);
   DataPath_RF_BLOCKi_73_Q_reg_1_inst : DFF_X1 port map( D => n5826, CK => CLK,
                           Q => n_1575, QN => 
                           DataPath_RF_bus_reg_dataout_2081_port);
   DataPath_RF_BLOCKi_74_Q_reg_1_inst : DFF_X1 port map( D => n5862, CK => CLK,
                           Q => n_1576, QN => 
                           DataPath_RF_bus_reg_dataout_2113_port);
   DataPath_RF_BLOCKi_75_Q_reg_1_inst : DFF_X1 port map( D => n5898, CK => CLK,
                           Q => n_1577, QN => 
                           DataPath_RF_bus_reg_dataout_2145_port);
   DataPath_RF_BLOCKi_76_Q_reg_1_inst : DFF_X1 port map( D => n5934, CK => CLK,
                           Q => n_1578, QN => 
                           DataPath_RF_bus_reg_dataout_2177_port);
   DataPath_RF_BLOCKi_77_Q_reg_1_inst : DFF_X1 port map( D => n5970, CK => CLK,
                           Q => n_1579, QN => 
                           DataPath_RF_bus_reg_dataout_2209_port);
   DataPath_RF_BLOCKi_78_Q_reg_1_inst : DFF_X1 port map( D => n6006, CK => CLK,
                           Q => n_1580, QN => 
                           DataPath_RF_bus_reg_dataout_2241_port);
   DataPath_RF_BLOCKi_79_Q_reg_1_inst : DFF_X1 port map( D => n6042, CK => CLK,
                           Q => n_1581, QN => 
                           DataPath_RF_bus_reg_dataout_2273_port);
   DataPath_RF_BLOCKi_80_Q_reg_1_inst : DFF_X1 port map( D => n6079, CK => CLK,
                           Q => n_1582, QN => 
                           DataPath_RF_bus_reg_dataout_2305_port);
   DataPath_RF_BLOCKi_81_Q_reg_1_inst : DFF_X1 port map( D => n6115, CK => CLK,
                           Q => n_1583, QN => 
                           DataPath_RF_bus_reg_dataout_2337_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_14_inst : DFF_X1 port map( D => n2195, CK 
                           => CLK, Q => n_1584, QN => 
                           DataPath_i_REG_LDSTR_OUT_14_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_22_inst : DFF_X1 port map( D => n2187, CK 
                           => CLK, Q => n_1585, QN => 
                           DataPath_i_REG_LDSTR_OUT_22_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_30_inst : DFF_X1 port map( D => n2179, CK 
                           => CLK, Q => n_1586, QN => 
                           DataPath_i_REG_LDSTR_OUT_30_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_6_inst : DFF_X1 port map( D => n2203, CK =>
                           CLK, Q => n_1587, QN => 
                           DataPath_i_REG_LDSTR_OUT_6_port);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_6_inst : DFF_X1 port map( D => n6857, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_102_port
                           , QN => n669);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_6_inst : DFF_X1 port map( D => n6889, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_134_port
                           , QN => n701);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_6_inst : DFF_X1 port map( D => n6953, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_198_port
                           , QN => n765);
   DataPath_RF_BLOCKi_8_Q_reg_6_inst : DFF_X1 port map( D => n3360, CK => CLK, 
                           Q => n_1588, QN => 
                           DataPath_RF_bus_reg_dataout_6_port);
   DataPath_RF_BLOCKi_9_Q_reg_6_inst : DFF_X1 port map( D => n3406, CK => CLK, 
                           Q => n_1589, QN => 
                           DataPath_RF_bus_reg_dataout_38_port);
   DataPath_RF_BLOCKi_10_Q_reg_6_inst : DFF_X1 port map( D => n3444, CK => CLK,
                           Q => n_1590, QN => 
                           DataPath_RF_bus_reg_dataout_70_port);
   DataPath_RF_BLOCKi_11_Q_reg_6_inst : DFF_X1 port map( D => n3482, CK => CLK,
                           Q => n_1591, QN => 
                           DataPath_RF_bus_reg_dataout_102_port);
   DataPath_RF_BLOCKi_12_Q_reg_6_inst : DFF_X1 port map( D => n3520, CK => CLK,
                           Q => n_1592, QN => 
                           DataPath_RF_bus_reg_dataout_134_port);
   DataPath_RF_BLOCKi_13_Q_reg_6_inst : DFF_X1 port map( D => n3558, CK => CLK,
                           Q => n_1593, QN => 
                           DataPath_RF_bus_reg_dataout_166_port);
   DataPath_RF_BLOCKi_14_Q_reg_6_inst : DFF_X1 port map( D => n3596, CK => CLK,
                           Q => n_1594, QN => 
                           DataPath_RF_bus_reg_dataout_198_port);
   DataPath_RF_BLOCKi_15_Q_reg_6_inst : DFF_X1 port map( D => n3634, CK => CLK,
                           Q => n_1595, QN => 
                           DataPath_RF_bus_reg_dataout_230_port);
   DataPath_RF_BLOCKi_16_Q_reg_6_inst : DFF_X1 port map( D => n3672, CK => CLK,
                           Q => n_1596, QN => 
                           DataPath_RF_bus_reg_dataout_262_port);
   DataPath_RF_BLOCKi_17_Q_reg_6_inst : DFF_X1 port map( D => n3709, CK => CLK,
                           Q => n_1597, QN => 
                           DataPath_RF_bus_reg_dataout_294_port);
   DataPath_RF_BLOCKi_18_Q_reg_6_inst : DFF_X1 port map( D => n3746, CK => CLK,
                           Q => n_1598, QN => 
                           DataPath_RF_bus_reg_dataout_326_port);
   DataPath_RF_BLOCKi_19_Q_reg_6_inst : DFF_X1 port map( D => n3783, CK => CLK,
                           Q => n_1599, QN => 
                           DataPath_RF_bus_reg_dataout_358_port);
   DataPath_RF_BLOCKi_20_Q_reg_6_inst : DFF_X1 port map( D => n3818, CK => CLK,
                           Q => n_1600, QN => 
                           DataPath_RF_bus_reg_dataout_390_port);
   DataPath_RF_BLOCKi_21_Q_reg_6_inst : DFF_X1 port map( D => n3853, CK => CLK,
                           Q => n_1601, QN => 
                           DataPath_RF_bus_reg_dataout_422_port);
   DataPath_RF_BLOCKi_22_Q_reg_6_inst : DFF_X1 port map( D => n3888, CK => CLK,
                           Q => n_1602, QN => 
                           DataPath_RF_bus_reg_dataout_454_port);
   DataPath_RF_BLOCKi_23_Q_reg_6_inst : DFF_X1 port map( D => n3948, CK => CLK,
                           Q => n_1603, QN => 
                           DataPath_RF_bus_reg_dataout_486_port);
   DataPath_RF_BLOCKi_24_Q_reg_6_inst : DFF_X1 port map( D => n4016, CK => CLK,
                           Q => n_1604, QN => 
                           DataPath_RF_bus_reg_dataout_518_port);
   DataPath_RF_BLOCKi_25_Q_reg_6_inst : DFF_X1 port map( D => n4059, CK => CLK,
                           Q => n_1605, QN => 
                           DataPath_RF_bus_reg_dataout_550_port);
   DataPath_RF_BLOCKi_26_Q_reg_6_inst : DFF_X1 port map( D => n4094, CK => CLK,
                           Q => n_1606, QN => 
                           DataPath_RF_bus_reg_dataout_582_port);
   DataPath_RF_BLOCKi_27_Q_reg_6_inst : DFF_X1 port map( D => n4129, CK => CLK,
                           Q => n_1607, QN => 
                           DataPath_RF_bus_reg_dataout_614_port);
   DataPath_RF_BLOCKi_28_Q_reg_6_inst : DFF_X1 port map( D => n4164, CK => CLK,
                           Q => n_1608, QN => 
                           DataPath_RF_bus_reg_dataout_646_port);
   DataPath_RF_BLOCKi_29_Q_reg_6_inst : DFF_X1 port map( D => n4199, CK => CLK,
                           Q => n_1609, QN => 
                           DataPath_RF_bus_reg_dataout_678_port);
   DataPath_RF_BLOCKi_30_Q_reg_6_inst : DFF_X1 port map( D => n4234, CK => CLK,
                           Q => n_1610, QN => 
                           DataPath_RF_bus_reg_dataout_710_port);
   DataPath_RF_BLOCKi_31_Q_reg_6_inst : DFF_X1 port map( D => n4269, CK => CLK,
                           Q => n_1611, QN => 
                           DataPath_RF_bus_reg_dataout_742_port);
   DataPath_RF_BLOCKi_32_Q_reg_6_inst : DFF_X1 port map( D => n4304, CK => CLK,
                           Q => n_1612, QN => 
                           DataPath_RF_bus_reg_dataout_774_port);
   DataPath_RF_BLOCKi_33_Q_reg_6_inst : DFF_X1 port map( D => n4339, CK => CLK,
                           Q => n_1613, QN => 
                           DataPath_RF_bus_reg_dataout_806_port);
   DataPath_RF_BLOCKi_34_Q_reg_6_inst : DFF_X1 port map( D => n4374, CK => CLK,
                           Q => n_1614, QN => 
                           DataPath_RF_bus_reg_dataout_838_port);
   DataPath_RF_BLOCKi_35_Q_reg_6_inst : DFF_X1 port map( D => n4409, CK => CLK,
                           Q => n_1615, QN => 
                           DataPath_RF_bus_reg_dataout_870_port);
   DataPath_RF_BLOCKi_36_Q_reg_6_inst : DFF_X1 port map( D => n4444, CK => CLK,
                           Q => n_1616, QN => 
                           DataPath_RF_bus_reg_dataout_902_port);
   DataPath_RF_BLOCKi_37_Q_reg_6_inst : DFF_X1 port map( D => n4479, CK => CLK,
                           Q => n_1617, QN => 
                           DataPath_RF_bus_reg_dataout_934_port);
   DataPath_RF_BLOCKi_38_Q_reg_6_inst : DFF_X1 port map( D => n4514, CK => CLK,
                           Q => n_1618, QN => 
                           DataPath_RF_bus_reg_dataout_966_port);
   DataPath_RF_BLOCKi_39_Q_reg_6_inst : DFF_X1 port map( D => n4549, CK => CLK,
                           Q => n_1619, QN => 
                           DataPath_RF_bus_reg_dataout_998_port);
   DataPath_RF_BLOCKi_40_Q_reg_6_inst : DFF_X1 port map( D => n4609, CK => CLK,
                           Q => n_1620, QN => 
                           DataPath_RF_bus_reg_dataout_1030_port);
   DataPath_RF_BLOCKi_41_Q_reg_6_inst : DFF_X1 port map( D => n4652, CK => CLK,
                           Q => n_1621, QN => 
                           DataPath_RF_bus_reg_dataout_1062_port);
   DataPath_RF_BLOCKi_42_Q_reg_6_inst : DFF_X1 port map( D => n4687, CK => CLK,
                           Q => n_1622, QN => 
                           DataPath_RF_bus_reg_dataout_1094_port);
   DataPath_RF_BLOCKi_43_Q_reg_6_inst : DFF_X1 port map( D => n4722, CK => CLK,
                           Q => n_1623, QN => 
                           DataPath_RF_bus_reg_dataout_1126_port);
   DataPath_RF_BLOCKi_44_Q_reg_6_inst : DFF_X1 port map( D => n4757, CK => CLK,
                           Q => n_1624, QN => 
                           DataPath_RF_bus_reg_dataout_1158_port);
   DataPath_RF_BLOCKi_45_Q_reg_6_inst : DFF_X1 port map( D => n4792, CK => CLK,
                           Q => n_1625, QN => 
                           DataPath_RF_bus_reg_dataout_1190_port);
   DataPath_RF_BLOCKi_46_Q_reg_6_inst : DFF_X1 port map( D => n4827, CK => CLK,
                           Q => n_1626, QN => 
                           DataPath_RF_bus_reg_dataout_1222_port);
   DataPath_RF_BLOCKi_47_Q_reg_6_inst : DFF_X1 port map( D => n4862, CK => CLK,
                           Q => n_1627, QN => 
                           DataPath_RF_bus_reg_dataout_1254_port);
   DataPath_RF_BLOCKi_48_Q_reg_6_inst : DFF_X1 port map( D => n4897, CK => CLK,
                           Q => n_1628, QN => 
                           DataPath_RF_bus_reg_dataout_1286_port);
   DataPath_RF_BLOCKi_49_Q_reg_6_inst : DFF_X1 port map( D => n4932, CK => CLK,
                           Q => n_1629, QN => 
                           DataPath_RF_bus_reg_dataout_1318_port);
   DataPath_RF_BLOCKi_50_Q_reg_6_inst : DFF_X1 port map( D => n4967, CK => CLK,
                           Q => n_1630, QN => 
                           DataPath_RF_bus_reg_dataout_1350_port);
   DataPath_RF_BLOCKi_51_Q_reg_6_inst : DFF_X1 port map( D => n5002, CK => CLK,
                           Q => n_1631, QN => 
                           DataPath_RF_bus_reg_dataout_1382_port);
   DataPath_RF_BLOCKi_52_Q_reg_6_inst : DFF_X1 port map( D => n5037, CK => CLK,
                           Q => n_1632, QN => 
                           DataPath_RF_bus_reg_dataout_1414_port);
   DataPath_RF_BLOCKi_53_Q_reg_6_inst : DFF_X1 port map( D => n5072, CK => CLK,
                           Q => n_1633, QN => 
                           DataPath_RF_bus_reg_dataout_1446_port);
   DataPath_RF_BLOCKi_54_Q_reg_6_inst : DFF_X1 port map( D => n5107, CK => CLK,
                           Q => n_1634, QN => 
                           DataPath_RF_bus_reg_dataout_1478_port);
   DataPath_RF_BLOCKi_55_Q_reg_6_inst : DFF_X1 port map( D => n5142, CK => CLK,
                           Q => n_1635, QN => 
                           DataPath_RF_bus_reg_dataout_1510_port);
   DataPath_RF_BLOCKi_56_Q_reg_6_inst : DFF_X1 port map( D => n5202, CK => CLK,
                           Q => n_1636, QN => 
                           DataPath_RF_bus_reg_dataout_1542_port);
   DataPath_RF_BLOCKi_57_Q_reg_6_inst : DFF_X1 port map( D => n5244, CK => CLK,
                           Q => n_1637, QN => 
                           DataPath_RF_bus_reg_dataout_1574_port);
   DataPath_RF_BLOCKi_58_Q_reg_6_inst : DFF_X1 port map( D => n5280, CK => CLK,
                           Q => n_1638, QN => 
                           DataPath_RF_bus_reg_dataout_1606_port);
   DataPath_RF_BLOCKi_59_Q_reg_6_inst : DFF_X1 port map( D => n5315, CK => CLK,
                           Q => n_1639, QN => 
                           DataPath_RF_bus_reg_dataout_1638_port);
   DataPath_RF_BLOCKi_60_Q_reg_6_inst : DFF_X1 port map( D => n5350, CK => CLK,
                           Q => n_1640, QN => 
                           DataPath_RF_bus_reg_dataout_1670_port);
   DataPath_RF_BLOCKi_61_Q_reg_6_inst : DFF_X1 port map( D => n5385, CK => CLK,
                           Q => n_1641, QN => 
                           DataPath_RF_bus_reg_dataout_1702_port);
   DataPath_RF_BLOCKi_62_Q_reg_6_inst : DFF_X1 port map( D => n5420, CK => CLK,
                           Q => n_1642, QN => 
                           DataPath_RF_bus_reg_dataout_1734_port);
   DataPath_RF_BLOCKi_63_Q_reg_6_inst : DFF_X1 port map( D => n5455, CK => CLK,
                           Q => n_1643, QN => 
                           DataPath_RF_bus_reg_dataout_1766_port);
   DataPath_RF_BLOCKi_64_Q_reg_6_inst : DFF_X1 port map( D => n5490, CK => CLK,
                           Q => n_1644, QN => 
                           DataPath_RF_bus_reg_dataout_1798_port);
   DataPath_RF_BLOCKi_65_Q_reg_6_inst : DFF_X1 port map( D => n5525, CK => CLK,
                           Q => n_1645, QN => 
                           DataPath_RF_bus_reg_dataout_1830_port);
   DataPath_RF_BLOCKi_66_Q_reg_6_inst : DFF_X1 port map( D => n5560, CK => CLK,
                           Q => n_1646, QN => 
                           DataPath_RF_bus_reg_dataout_1862_port);
   DataPath_RF_BLOCKi_67_Q_reg_6_inst : DFF_X1 port map( D => n5595, CK => CLK,
                           Q => n_1647, QN => 
                           DataPath_RF_bus_reg_dataout_1894_port);
   DataPath_RF_BLOCKi_68_Q_reg_6_inst : DFF_X1 port map( D => n5634, CK => CLK,
                           Q => n_1648, QN => 
                           DataPath_RF_bus_reg_dataout_1926_port);
   DataPath_RF_BLOCKi_69_Q_reg_6_inst : DFF_X1 port map( D => n5671, CK => CLK,
                           Q => n_1649, QN => 
                           DataPath_RF_bus_reg_dataout_1958_port);
   DataPath_RF_BLOCKi_70_Q_reg_6_inst : DFF_X1 port map( D => n5708, CK => CLK,
                           Q => n_1650, QN => 
                           DataPath_RF_bus_reg_dataout_1990_port);
   DataPath_RF_BLOCKi_71_Q_reg_6_inst : DFF_X1 port map( D => n5745, CK => CLK,
                           Q => n_1651, QN => 
                           DataPath_RF_bus_reg_dataout_2022_port);
   DataPath_RF_BLOCKi_82_Q_reg_6_inst : DFF_X1 port map( D => n900, CK => CLK, 
                           Q => n_1652, QN => 
                           DataPath_RF_bus_reg_dataout_2374_port);
   DataPath_RF_BLOCKi_83_Q_reg_6_inst : DFF_X1 port map( D => n957, CK => CLK, 
                           Q => n_1653, QN => 
                           DataPath_RF_bus_reg_dataout_2406_port);
   DataPath_RF_BLOCKi_84_Q_reg_6_inst : DFF_X1 port map( D => n995, CK => CLK, 
                           Q => n_1654, QN => 
                           DataPath_RF_bus_reg_dataout_2438_port);
   DataPath_RF_BLOCKi_85_Q_reg_6_inst : DFF_X1 port map( D => n1032, CK => CLK,
                           Q => n_1655, QN => 
                           DataPath_RF_bus_reg_dataout_2470_port);
   DataPath_RF_BLOCKi_86_Q_reg_6_inst : DFF_X1 port map( D => n1069, CK => CLK,
                           Q => n_1656, QN => 
                           DataPath_RF_bus_reg_dataout_2502_port);
   DataPath_RF_BLOCKi_87_Q_reg_6_inst : DFF_X1 port map( D => n1106, CK => CLK,
                           Q => n_1657, QN => 
                           DataPath_RF_bus_reg_dataout_2534_port);
   DataPath_RF_BLOCKi_72_Q_reg_6_inst : DFF_X1 port map( D => n5782, CK => CLK,
                           Q => n_1658, QN => 
                           DataPath_RF_bus_reg_dataout_2054_port);
   DataPath_RF_BLOCKi_73_Q_reg_6_inst : DFF_X1 port map( D => n5821, CK => CLK,
                           Q => n_1659, QN => 
                           DataPath_RF_bus_reg_dataout_2086_port);
   DataPath_RF_BLOCKi_74_Q_reg_6_inst : DFF_X1 port map( D => n5857, CK => CLK,
                           Q => n_1660, QN => 
                           DataPath_RF_bus_reg_dataout_2118_port);
   DataPath_RF_BLOCKi_75_Q_reg_6_inst : DFF_X1 port map( D => n5893, CK => CLK,
                           Q => n_1661, QN => 
                           DataPath_RF_bus_reg_dataout_2150_port);
   DataPath_RF_BLOCKi_76_Q_reg_6_inst : DFF_X1 port map( D => n5929, CK => CLK,
                           Q => n_1662, QN => 
                           DataPath_RF_bus_reg_dataout_2182_port);
   DataPath_RF_BLOCKi_77_Q_reg_6_inst : DFF_X1 port map( D => n5965, CK => CLK,
                           Q => n_1663, QN => 
                           DataPath_RF_bus_reg_dataout_2214_port);
   DataPath_RF_BLOCKi_78_Q_reg_6_inst : DFF_X1 port map( D => n6001, CK => CLK,
                           Q => n_1664, QN => 
                           DataPath_RF_bus_reg_dataout_2246_port);
   DataPath_RF_BLOCKi_79_Q_reg_6_inst : DFF_X1 port map( D => n6037, CK => CLK,
                           Q => n_1665, QN => 
                           DataPath_RF_bus_reg_dataout_2278_port);
   DataPath_RF_BLOCKi_80_Q_reg_6_inst : DFF_X1 port map( D => n6074, CK => CLK,
                           Q => n_1666, QN => 
                           DataPath_RF_bus_reg_dataout_2310_port);
   DataPath_RF_BLOCKi_81_Q_reg_6_inst : DFF_X1 port map( D => n6110, CK => CLK,
                           Q => n_1667, QN => 
                           DataPath_RF_bus_reg_dataout_2342_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_13_inst : DFF_X1 port map( D => n2196, CK 
                           => CLK, Q => n_1668, QN => 
                           DataPath_i_REG_LDSTR_OUT_13_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_13_inst : DFF_X1 port map( D => n6786, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_45_port,
                           QN => n612);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_13_inst : DFF_X1 port map( D => n6818, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_77_port,
                           QN => n644);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_13_inst : DFF_X1 port map( D => n6850, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_109_port
                           , QN => n676);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_13_inst : DFF_X1 port map( D => n6882, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_141_port
                           , QN => n708);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_13_inst : DFF_X1 port map( D => n6914, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_173_port
                           , QN => n740);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_13_inst : DFF_X1 port map( D => n6946, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_205_port
                           , QN => n772);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_13_inst : DFF_X1 port map( D => n6978, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_237_port
                           , QN => n804);
   DataPath_RF_BLOCKi_8_Q_reg_13_inst : DFF_X1 port map( D => n3346, CK => CLK,
                           Q => n_1669, QN => 
                           DataPath_RF_bus_reg_dataout_13_port);
   DataPath_RF_BLOCKi_9_Q_reg_13_inst : DFF_X1 port map( D => n3399, CK => CLK,
                           Q => n_1670, QN => 
                           DataPath_RF_bus_reg_dataout_45_port);
   DataPath_RF_BLOCKi_10_Q_reg_13_inst : DFF_X1 port map( D => n3437, CK => CLK
                           , Q => n_1671, QN => 
                           DataPath_RF_bus_reg_dataout_77_port);
   DataPath_RF_BLOCKi_11_Q_reg_13_inst : DFF_X1 port map( D => n3475, CK => CLK
                           , Q => n_1672, QN => 
                           DataPath_RF_bus_reg_dataout_109_port);
   DataPath_RF_BLOCKi_12_Q_reg_13_inst : DFF_X1 port map( D => n3513, CK => CLK
                           , Q => n_1673, QN => 
                           DataPath_RF_bus_reg_dataout_141_port);
   DataPath_RF_BLOCKi_13_Q_reg_13_inst : DFF_X1 port map( D => n3551, CK => CLK
                           , Q => n_1674, QN => 
                           DataPath_RF_bus_reg_dataout_173_port);
   DataPath_RF_BLOCKi_14_Q_reg_13_inst : DFF_X1 port map( D => n3589, CK => CLK
                           , Q => n_1675, QN => 
                           DataPath_RF_bus_reg_dataout_205_port);
   DataPath_RF_BLOCKi_15_Q_reg_13_inst : DFF_X1 port map( D => n3627, CK => CLK
                           , Q => n_1676, QN => 
                           DataPath_RF_bus_reg_dataout_237_port);
   DataPath_RF_BLOCKi_16_Q_reg_13_inst : DFF_X1 port map( D => n3665, CK => CLK
                           , Q => n_1677, QN => 
                           DataPath_RF_bus_reg_dataout_269_port);
   DataPath_RF_BLOCKi_17_Q_reg_13_inst : DFF_X1 port map( D => n3702, CK => CLK
                           , Q => n_1678, QN => 
                           DataPath_RF_bus_reg_dataout_301_port);
   DataPath_RF_BLOCKi_18_Q_reg_13_inst : DFF_X1 port map( D => n3739, CK => CLK
                           , Q => n_1679, QN => 
                           DataPath_RF_bus_reg_dataout_333_port);
   DataPath_RF_BLOCKi_19_Q_reg_13_inst : DFF_X1 port map( D => n3776, CK => CLK
                           , Q => n_1680, QN => 
                           DataPath_RF_bus_reg_dataout_365_port);
   DataPath_RF_BLOCKi_20_Q_reg_13_inst : DFF_X1 port map( D => n3811, CK => CLK
                           , Q => n_1681, QN => 
                           DataPath_RF_bus_reg_dataout_397_port);
   DataPath_RF_BLOCKi_21_Q_reg_13_inst : DFF_X1 port map( D => n3846, CK => CLK
                           , Q => n_1682, QN => 
                           DataPath_RF_bus_reg_dataout_429_port);
   DataPath_RF_BLOCKi_22_Q_reg_13_inst : DFF_X1 port map( D => n3881, CK => CLK
                           , Q => n_1683, QN => 
                           DataPath_RF_bus_reg_dataout_461_port);
   DataPath_RF_BLOCKi_23_Q_reg_13_inst : DFF_X1 port map( D => n3934, CK => CLK
                           , Q => n_1684, QN => 
                           DataPath_RF_bus_reg_dataout_493_port);
   DataPath_RF_BLOCKi_24_Q_reg_13_inst : DFF_X1 port map( D => n4002, CK => CLK
                           , Q => n_1685, QN => 
                           DataPath_RF_bus_reg_dataout_525_port);
   DataPath_RF_BLOCKi_25_Q_reg_13_inst : DFF_X1 port map( D => n4052, CK => CLK
                           , Q => n_1686, QN => 
                           DataPath_RF_bus_reg_dataout_557_port);
   DataPath_RF_BLOCKi_26_Q_reg_13_inst : DFF_X1 port map( D => n4087, CK => CLK
                           , Q => n_1687, QN => 
                           DataPath_RF_bus_reg_dataout_589_port);
   DataPath_RF_BLOCKi_27_Q_reg_13_inst : DFF_X1 port map( D => n4122, CK => CLK
                           , Q => n_1688, QN => 
                           DataPath_RF_bus_reg_dataout_621_port);
   DataPath_RF_BLOCKi_28_Q_reg_13_inst : DFF_X1 port map( D => n4157, CK => CLK
                           , Q => n_1689, QN => 
                           DataPath_RF_bus_reg_dataout_653_port);
   DataPath_RF_BLOCKi_29_Q_reg_13_inst : DFF_X1 port map( D => n4192, CK => CLK
                           , Q => n_1690, QN => 
                           DataPath_RF_bus_reg_dataout_685_port);
   DataPath_RF_BLOCKi_30_Q_reg_13_inst : DFF_X1 port map( D => n4227, CK => CLK
                           , Q => n_1691, QN => 
                           DataPath_RF_bus_reg_dataout_717_port);
   DataPath_RF_BLOCKi_31_Q_reg_13_inst : DFF_X1 port map( D => n4262, CK => CLK
                           , Q => n_1692, QN => 
                           DataPath_RF_bus_reg_dataout_749_port);
   DataPath_RF_BLOCKi_32_Q_reg_13_inst : DFF_X1 port map( D => n4297, CK => CLK
                           , Q => n_1693, QN => 
                           DataPath_RF_bus_reg_dataout_781_port);
   DataPath_RF_BLOCKi_33_Q_reg_13_inst : DFF_X1 port map( D => n4332, CK => CLK
                           , Q => n_1694, QN => 
                           DataPath_RF_bus_reg_dataout_813_port);
   DataPath_RF_BLOCKi_34_Q_reg_13_inst : DFF_X1 port map( D => n4367, CK => CLK
                           , Q => n_1695, QN => 
                           DataPath_RF_bus_reg_dataout_845_port);
   DataPath_RF_BLOCKi_35_Q_reg_13_inst : DFF_X1 port map( D => n4402, CK => CLK
                           , Q => n_1696, QN => 
                           DataPath_RF_bus_reg_dataout_877_port);
   DataPath_RF_BLOCKi_36_Q_reg_13_inst : DFF_X1 port map( D => n4437, CK => CLK
                           , Q => n_1697, QN => 
                           DataPath_RF_bus_reg_dataout_909_port);
   DataPath_RF_BLOCKi_37_Q_reg_13_inst : DFF_X1 port map( D => n4472, CK => CLK
                           , Q => n_1698, QN => 
                           DataPath_RF_bus_reg_dataout_941_port);
   DataPath_RF_BLOCKi_38_Q_reg_13_inst : DFF_X1 port map( D => n4507, CK => CLK
                           , Q => n_1699, QN => 
                           DataPath_RF_bus_reg_dataout_973_port);
   DataPath_RF_BLOCKi_39_Q_reg_13_inst : DFF_X1 port map( D => n4542, CK => CLK
                           , Q => n_1700, QN => 
                           DataPath_RF_bus_reg_dataout_1005_port);
   DataPath_RF_BLOCKi_40_Q_reg_13_inst : DFF_X1 port map( D => n4595, CK => CLK
                           , Q => n_1701, QN => 
                           DataPath_RF_bus_reg_dataout_1037_port);
   DataPath_RF_BLOCKi_41_Q_reg_13_inst : DFF_X1 port map( D => n4645, CK => CLK
                           , Q => n_1702, QN => 
                           DataPath_RF_bus_reg_dataout_1069_port);
   DataPath_RF_BLOCKi_42_Q_reg_13_inst : DFF_X1 port map( D => n4680, CK => CLK
                           , Q => n_1703, QN => 
                           DataPath_RF_bus_reg_dataout_1101_port);
   DataPath_RF_BLOCKi_43_Q_reg_13_inst : DFF_X1 port map( D => n4715, CK => CLK
                           , Q => n_1704, QN => 
                           DataPath_RF_bus_reg_dataout_1133_port);
   DataPath_RF_BLOCKi_44_Q_reg_13_inst : DFF_X1 port map( D => n4750, CK => CLK
                           , Q => n_1705, QN => 
                           DataPath_RF_bus_reg_dataout_1165_port);
   DataPath_RF_BLOCKi_45_Q_reg_13_inst : DFF_X1 port map( D => n4785, CK => CLK
                           , Q => n_1706, QN => 
                           DataPath_RF_bus_reg_dataout_1197_port);
   DataPath_RF_BLOCKi_46_Q_reg_13_inst : DFF_X1 port map( D => n4820, CK => CLK
                           , Q => n_1707, QN => 
                           DataPath_RF_bus_reg_dataout_1229_port);
   DataPath_RF_BLOCKi_47_Q_reg_13_inst : DFF_X1 port map( D => n4855, CK => CLK
                           , Q => n_1708, QN => 
                           DataPath_RF_bus_reg_dataout_1261_port);
   DataPath_RF_BLOCKi_48_Q_reg_13_inst : DFF_X1 port map( D => n4890, CK => CLK
                           , Q => n_1709, QN => 
                           DataPath_RF_bus_reg_dataout_1293_port);
   DataPath_RF_BLOCKi_49_Q_reg_13_inst : DFF_X1 port map( D => n4925, CK => CLK
                           , Q => n_1710, QN => 
                           DataPath_RF_bus_reg_dataout_1325_port);
   DataPath_RF_BLOCKi_50_Q_reg_13_inst : DFF_X1 port map( D => n4960, CK => CLK
                           , Q => n_1711, QN => 
                           DataPath_RF_bus_reg_dataout_1357_port);
   DataPath_RF_BLOCKi_51_Q_reg_13_inst : DFF_X1 port map( D => n4995, CK => CLK
                           , Q => n_1712, QN => 
                           DataPath_RF_bus_reg_dataout_1389_port);
   DataPath_RF_BLOCKi_52_Q_reg_13_inst : DFF_X1 port map( D => n5030, CK => CLK
                           , Q => n_1713, QN => 
                           DataPath_RF_bus_reg_dataout_1421_port);
   DataPath_RF_BLOCKi_53_Q_reg_13_inst : DFF_X1 port map( D => n5065, CK => CLK
                           , Q => n_1714, QN => 
                           DataPath_RF_bus_reg_dataout_1453_port);
   DataPath_RF_BLOCKi_54_Q_reg_13_inst : DFF_X1 port map( D => n5100, CK => CLK
                           , Q => n_1715, QN => 
                           DataPath_RF_bus_reg_dataout_1485_port);
   DataPath_RF_BLOCKi_55_Q_reg_13_inst : DFF_X1 port map( D => n5135, CK => CLK
                           , Q => n_1716, QN => 
                           DataPath_RF_bus_reg_dataout_1517_port);
   DataPath_RF_BLOCKi_56_Q_reg_13_inst : DFF_X1 port map( D => n5188, CK => CLK
                           , Q => n_1717, QN => 
                           DataPath_RF_bus_reg_dataout_1549_port);
   DataPath_RF_BLOCKi_57_Q_reg_13_inst : DFF_X1 port map( D => n5237, CK => CLK
                           , Q => n_1718, QN => 
                           DataPath_RF_bus_reg_dataout_1581_port);
   DataPath_RF_BLOCKi_58_Q_reg_13_inst : DFF_X1 port map( D => n5273, CK => CLK
                           , Q => n_1719, QN => 
                           DataPath_RF_bus_reg_dataout_1613_port);
   DataPath_RF_BLOCKi_59_Q_reg_13_inst : DFF_X1 port map( D => n5308, CK => CLK
                           , Q => n_1720, QN => 
                           DataPath_RF_bus_reg_dataout_1645_port);
   DataPath_RF_BLOCKi_60_Q_reg_13_inst : DFF_X1 port map( D => n5343, CK => CLK
                           , Q => n_1721, QN => 
                           DataPath_RF_bus_reg_dataout_1677_port);
   DataPath_RF_BLOCKi_61_Q_reg_13_inst : DFF_X1 port map( D => n5378, CK => CLK
                           , Q => n_1722, QN => 
                           DataPath_RF_bus_reg_dataout_1709_port);
   DataPath_RF_BLOCKi_62_Q_reg_13_inst : DFF_X1 port map( D => n5413, CK => CLK
                           , Q => n_1723, QN => 
                           DataPath_RF_bus_reg_dataout_1741_port);
   DataPath_RF_BLOCKi_63_Q_reg_13_inst : DFF_X1 port map( D => n5448, CK => CLK
                           , Q => n_1724, QN => 
                           DataPath_RF_bus_reg_dataout_1773_port);
   DataPath_RF_BLOCKi_64_Q_reg_13_inst : DFF_X1 port map( D => n5483, CK => CLK
                           , Q => n_1725, QN => 
                           DataPath_RF_bus_reg_dataout_1805_port);
   DataPath_RF_BLOCKi_65_Q_reg_13_inst : DFF_X1 port map( D => n5518, CK => CLK
                           , Q => n_1726, QN => 
                           DataPath_RF_bus_reg_dataout_1837_port);
   DataPath_RF_BLOCKi_66_Q_reg_13_inst : DFF_X1 port map( D => n5553, CK => CLK
                           , Q => n_1727, QN => 
                           DataPath_RF_bus_reg_dataout_1869_port);
   DataPath_RF_BLOCKi_67_Q_reg_13_inst : DFF_X1 port map( D => n5588, CK => CLK
                           , Q => n_1728, QN => 
                           DataPath_RF_bus_reg_dataout_1901_port);
   DataPath_RF_BLOCKi_68_Q_reg_13_inst : DFF_X1 port map( D => n5627, CK => CLK
                           , Q => n_1729, QN => 
                           DataPath_RF_bus_reg_dataout_1933_port);
   DataPath_RF_BLOCKi_69_Q_reg_13_inst : DFF_X1 port map( D => n5664, CK => CLK
                           , Q => n_1730, QN => 
                           DataPath_RF_bus_reg_dataout_1965_port);
   DataPath_RF_BLOCKi_70_Q_reg_13_inst : DFF_X1 port map( D => n5701, CK => CLK
                           , Q => n_1731, QN => 
                           DataPath_RF_bus_reg_dataout_1997_port);
   DataPath_RF_BLOCKi_71_Q_reg_13_inst : DFF_X1 port map( D => n5738, CK => CLK
                           , Q => n_1732, QN => 
                           DataPath_RF_bus_reg_dataout_2029_port);
   DataPath_RF_BLOCKi_82_Q_reg_13_inst : DFF_X1 port map( D => n886, CK => CLK,
                           Q => n_1733, QN => 
                           DataPath_RF_bus_reg_dataout_2381_port);
   DataPath_RF_BLOCKi_83_Q_reg_13_inst : DFF_X1 port map( D => n950, CK => CLK,
                           Q => n_1734, QN => 
                           DataPath_RF_bus_reg_dataout_2413_port);
   DataPath_RF_BLOCKi_84_Q_reg_13_inst : DFF_X1 port map( D => n988, CK => CLK,
                           Q => n_1735, QN => 
                           DataPath_RF_bus_reg_dataout_2445_port);
   DataPath_RF_BLOCKi_85_Q_reg_13_inst : DFF_X1 port map( D => n1025, CK => CLK
                           , Q => n_1736, QN => 
                           DataPath_RF_bus_reg_dataout_2477_port);
   DataPath_RF_BLOCKi_86_Q_reg_13_inst : DFF_X1 port map( D => n1062, CK => CLK
                           , Q => n_1737, QN => 
                           DataPath_RF_bus_reg_dataout_2509_port);
   DataPath_RF_BLOCKi_87_Q_reg_13_inst : DFF_X1 port map( D => n1099, CK => CLK
                           , Q => n_1738, QN => 
                           DataPath_RF_bus_reg_dataout_2541_port);
   DataPath_RF_BLOCKi_72_Q_reg_13_inst : DFF_X1 port map( D => n5775, CK => CLK
                           , Q => n_1739, QN => 
                           DataPath_RF_bus_reg_dataout_2061_port);
   DataPath_RF_BLOCKi_73_Q_reg_13_inst : DFF_X1 port map( D => n5814, CK => CLK
                           , Q => n_1740, QN => 
                           DataPath_RF_bus_reg_dataout_2093_port);
   DataPath_RF_BLOCKi_74_Q_reg_13_inst : DFF_X1 port map( D => n5850, CK => CLK
                           , Q => n_1741, QN => 
                           DataPath_RF_bus_reg_dataout_2125_port);
   DataPath_RF_BLOCKi_75_Q_reg_13_inst : DFF_X1 port map( D => n5886, CK => CLK
                           , Q => n_1742, QN => 
                           DataPath_RF_bus_reg_dataout_2157_port);
   DataPath_RF_BLOCKi_76_Q_reg_13_inst : DFF_X1 port map( D => n5922, CK => CLK
                           , Q => n_1743, QN => 
                           DataPath_RF_bus_reg_dataout_2189_port);
   DataPath_RF_BLOCKi_77_Q_reg_13_inst : DFF_X1 port map( D => n5958, CK => CLK
                           , Q => n_1744, QN => 
                           DataPath_RF_bus_reg_dataout_2221_port);
   DataPath_RF_BLOCKi_78_Q_reg_13_inst : DFF_X1 port map( D => n5994, CK => CLK
                           , Q => n_1745, QN => 
                           DataPath_RF_bus_reg_dataout_2253_port);
   DataPath_RF_BLOCKi_79_Q_reg_13_inst : DFF_X1 port map( D => n6030, CK => CLK
                           , Q => n_1746, QN => 
                           DataPath_RF_bus_reg_dataout_2285_port);
   DataPath_RF_BLOCKi_80_Q_reg_13_inst : DFF_X1 port map( D => n6067, CK => CLK
                           , Q => n_1747, QN => 
                           DataPath_RF_bus_reg_dataout_2317_port);
   DataPath_RF_BLOCKi_81_Q_reg_13_inst : DFF_X1 port map( D => n6103, CK => CLK
                           , Q => n_1748, QN => 
                           DataPath_RF_bus_reg_dataout_2349_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_21_inst : DFF_X1 port map( D => n2188, CK 
                           => CLK, Q => n_1749, QN => 
                           DataPath_i_REG_LDSTR_OUT_21_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_29_inst : DFF_X1 port map( D => n2180, CK 
                           => CLK, Q => n_1750, QN => 
                           DataPath_i_REG_LDSTR_OUT_29_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_5_inst : DFF_X1 port map( D => n2204, CK =>
                           CLK, Q => n_1751, QN => 
                           DataPath_i_REG_LDSTR_OUT_5_port);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_5_inst : DFF_X1 port map( D => n6858, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_101_port
                           , QN => n668);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_5_inst : DFF_X1 port map( D => n6890, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_133_port
                           , QN => n700);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_5_inst : DFF_X1 port map( D => n6954, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_197_port
                           , QN => n764);
   DataPath_RF_BLOCKi_8_Q_reg_5_inst : DFF_X1 port map( D => n3362, CK => CLK, 
                           Q => n_1752, QN => 
                           DataPath_RF_bus_reg_dataout_5_port);
   DataPath_RF_BLOCKi_9_Q_reg_5_inst : DFF_X1 port map( D => n3407, CK => CLK, 
                           Q => n_1753, QN => 
                           DataPath_RF_bus_reg_dataout_37_port);
   DataPath_RF_BLOCKi_10_Q_reg_5_inst : DFF_X1 port map( D => n3445, CK => CLK,
                           Q => n_1754, QN => 
                           DataPath_RF_bus_reg_dataout_69_port);
   DataPath_RF_BLOCKi_11_Q_reg_5_inst : DFF_X1 port map( D => n3483, CK => CLK,
                           Q => n_1755, QN => 
                           DataPath_RF_bus_reg_dataout_101_port);
   DataPath_RF_BLOCKi_12_Q_reg_5_inst : DFF_X1 port map( D => n3521, CK => CLK,
                           Q => n_1756, QN => 
                           DataPath_RF_bus_reg_dataout_133_port);
   DataPath_RF_BLOCKi_13_Q_reg_5_inst : DFF_X1 port map( D => n3559, CK => CLK,
                           Q => n_1757, QN => 
                           DataPath_RF_bus_reg_dataout_165_port);
   DataPath_RF_BLOCKi_14_Q_reg_5_inst : DFF_X1 port map( D => n3597, CK => CLK,
                           Q => n_1758, QN => 
                           DataPath_RF_bus_reg_dataout_197_port);
   DataPath_RF_BLOCKi_15_Q_reg_5_inst : DFF_X1 port map( D => n3635, CK => CLK,
                           Q => n_1759, QN => 
                           DataPath_RF_bus_reg_dataout_229_port);
   DataPath_RF_BLOCKi_16_Q_reg_5_inst : DFF_X1 port map( D => n3673, CK => CLK,
                           Q => n_1760, QN => 
                           DataPath_RF_bus_reg_dataout_261_port);
   DataPath_RF_BLOCKi_17_Q_reg_5_inst : DFF_X1 port map( D => n3710, CK => CLK,
                           Q => n_1761, QN => 
                           DataPath_RF_bus_reg_dataout_293_port);
   DataPath_RF_BLOCKi_18_Q_reg_5_inst : DFF_X1 port map( D => n3747, CK => CLK,
                           Q => n_1762, QN => 
                           DataPath_RF_bus_reg_dataout_325_port);
   DataPath_RF_BLOCKi_19_Q_reg_5_inst : DFF_X1 port map( D => n3784, CK => CLK,
                           Q => n_1763, QN => 
                           DataPath_RF_bus_reg_dataout_357_port);
   DataPath_RF_BLOCKi_20_Q_reg_5_inst : DFF_X1 port map( D => n3819, CK => CLK,
                           Q => n_1764, QN => 
                           DataPath_RF_bus_reg_dataout_389_port);
   DataPath_RF_BLOCKi_21_Q_reg_5_inst : DFF_X1 port map( D => n3854, CK => CLK,
                           Q => n_1765, QN => 
                           DataPath_RF_bus_reg_dataout_421_port);
   DataPath_RF_BLOCKi_22_Q_reg_5_inst : DFF_X1 port map( D => n3889, CK => CLK,
                           Q => n_1766, QN => 
                           DataPath_RF_bus_reg_dataout_453_port);
   DataPath_RF_BLOCKi_23_Q_reg_5_inst : DFF_X1 port map( D => n3950, CK => CLK,
                           Q => n_1767, QN => 
                           DataPath_RF_bus_reg_dataout_485_port);
   DataPath_RF_BLOCKi_24_Q_reg_5_inst : DFF_X1 port map( D => n4018, CK => CLK,
                           Q => n_1768, QN => 
                           DataPath_RF_bus_reg_dataout_517_port);
   DataPath_RF_BLOCKi_25_Q_reg_5_inst : DFF_X1 port map( D => n4060, CK => CLK,
                           Q => n_1769, QN => 
                           DataPath_RF_bus_reg_dataout_549_port);
   DataPath_RF_BLOCKi_26_Q_reg_5_inst : DFF_X1 port map( D => n4095, CK => CLK,
                           Q => n_1770, QN => 
                           DataPath_RF_bus_reg_dataout_581_port);
   DataPath_RF_BLOCKi_27_Q_reg_5_inst : DFF_X1 port map( D => n4130, CK => CLK,
                           Q => n_1771, QN => 
                           DataPath_RF_bus_reg_dataout_613_port);
   DataPath_RF_BLOCKi_28_Q_reg_5_inst : DFF_X1 port map( D => n4165, CK => CLK,
                           Q => n_1772, QN => 
                           DataPath_RF_bus_reg_dataout_645_port);
   DataPath_RF_BLOCKi_29_Q_reg_5_inst : DFF_X1 port map( D => n4200, CK => CLK,
                           Q => n_1773, QN => 
                           DataPath_RF_bus_reg_dataout_677_port);
   DataPath_RF_BLOCKi_30_Q_reg_5_inst : DFF_X1 port map( D => n4235, CK => CLK,
                           Q => n_1774, QN => 
                           DataPath_RF_bus_reg_dataout_709_port);
   DataPath_RF_BLOCKi_31_Q_reg_5_inst : DFF_X1 port map( D => n4270, CK => CLK,
                           Q => n_1775, QN => 
                           DataPath_RF_bus_reg_dataout_741_port);
   DataPath_RF_BLOCKi_32_Q_reg_5_inst : DFF_X1 port map( D => n4305, CK => CLK,
                           Q => n_1776, QN => 
                           DataPath_RF_bus_reg_dataout_773_port);
   DataPath_RF_BLOCKi_33_Q_reg_5_inst : DFF_X1 port map( D => n4340, CK => CLK,
                           Q => n_1777, QN => 
                           DataPath_RF_bus_reg_dataout_805_port);
   DataPath_RF_BLOCKi_34_Q_reg_5_inst : DFF_X1 port map( D => n4375, CK => CLK,
                           Q => n_1778, QN => 
                           DataPath_RF_bus_reg_dataout_837_port);
   DataPath_RF_BLOCKi_35_Q_reg_5_inst : DFF_X1 port map( D => n4410, CK => CLK,
                           Q => n_1779, QN => 
                           DataPath_RF_bus_reg_dataout_869_port);
   DataPath_RF_BLOCKi_36_Q_reg_5_inst : DFF_X1 port map( D => n4445, CK => CLK,
                           Q => n_1780, QN => 
                           DataPath_RF_bus_reg_dataout_901_port);
   DataPath_RF_BLOCKi_37_Q_reg_5_inst : DFF_X1 port map( D => n4480, CK => CLK,
                           Q => n_1781, QN => 
                           DataPath_RF_bus_reg_dataout_933_port);
   DataPath_RF_BLOCKi_38_Q_reg_5_inst : DFF_X1 port map( D => n4515, CK => CLK,
                           Q => n_1782, QN => 
                           DataPath_RF_bus_reg_dataout_965_port);
   DataPath_RF_BLOCKi_39_Q_reg_5_inst : DFF_X1 port map( D => n4550, CK => CLK,
                           Q => n_1783, QN => 
                           DataPath_RF_bus_reg_dataout_997_port);
   DataPath_RF_BLOCKi_40_Q_reg_5_inst : DFF_X1 port map( D => n4611, CK => CLK,
                           Q => n_1784, QN => 
                           DataPath_RF_bus_reg_dataout_1029_port);
   DataPath_RF_BLOCKi_41_Q_reg_5_inst : DFF_X1 port map( D => n4653, CK => CLK,
                           Q => n_1785, QN => 
                           DataPath_RF_bus_reg_dataout_1061_port);
   DataPath_RF_BLOCKi_42_Q_reg_5_inst : DFF_X1 port map( D => n4688, CK => CLK,
                           Q => n_1786, QN => 
                           DataPath_RF_bus_reg_dataout_1093_port);
   DataPath_RF_BLOCKi_43_Q_reg_5_inst : DFF_X1 port map( D => n4723, CK => CLK,
                           Q => n_1787, QN => 
                           DataPath_RF_bus_reg_dataout_1125_port);
   DataPath_RF_BLOCKi_44_Q_reg_5_inst : DFF_X1 port map( D => n4758, CK => CLK,
                           Q => n_1788, QN => 
                           DataPath_RF_bus_reg_dataout_1157_port);
   DataPath_RF_BLOCKi_45_Q_reg_5_inst : DFF_X1 port map( D => n4793, CK => CLK,
                           Q => n_1789, QN => 
                           DataPath_RF_bus_reg_dataout_1189_port);
   DataPath_RF_BLOCKi_46_Q_reg_5_inst : DFF_X1 port map( D => n4828, CK => CLK,
                           Q => n_1790, QN => 
                           DataPath_RF_bus_reg_dataout_1221_port);
   DataPath_RF_BLOCKi_47_Q_reg_5_inst : DFF_X1 port map( D => n4863, CK => CLK,
                           Q => n_1791, QN => 
                           DataPath_RF_bus_reg_dataout_1253_port);
   DataPath_RF_BLOCKi_48_Q_reg_5_inst : DFF_X1 port map( D => n4898, CK => CLK,
                           Q => n_1792, QN => 
                           DataPath_RF_bus_reg_dataout_1285_port);
   DataPath_RF_BLOCKi_49_Q_reg_5_inst : DFF_X1 port map( D => n4933, CK => CLK,
                           Q => n_1793, QN => 
                           DataPath_RF_bus_reg_dataout_1317_port);
   DataPath_RF_BLOCKi_50_Q_reg_5_inst : DFF_X1 port map( D => n4968, CK => CLK,
                           Q => n_1794, QN => 
                           DataPath_RF_bus_reg_dataout_1349_port);
   DataPath_RF_BLOCKi_51_Q_reg_5_inst : DFF_X1 port map( D => n5003, CK => CLK,
                           Q => n_1795, QN => 
                           DataPath_RF_bus_reg_dataout_1381_port);
   DataPath_RF_BLOCKi_52_Q_reg_5_inst : DFF_X1 port map( D => n5038, CK => CLK,
                           Q => n_1796, QN => 
                           DataPath_RF_bus_reg_dataout_1413_port);
   DataPath_RF_BLOCKi_53_Q_reg_5_inst : DFF_X1 port map( D => n5073, CK => CLK,
                           Q => n_1797, QN => 
                           DataPath_RF_bus_reg_dataout_1445_port);
   DataPath_RF_BLOCKi_54_Q_reg_5_inst : DFF_X1 port map( D => n5108, CK => CLK,
                           Q => n_1798, QN => 
                           DataPath_RF_bus_reg_dataout_1477_port);
   DataPath_RF_BLOCKi_55_Q_reg_5_inst : DFF_X1 port map( D => n5143, CK => CLK,
                           Q => n_1799, QN => 
                           DataPath_RF_bus_reg_dataout_1509_port);
   DataPath_RF_BLOCKi_56_Q_reg_5_inst : DFF_X1 port map( D => n5204, CK => CLK,
                           Q => n_1800, QN => 
                           DataPath_RF_bus_reg_dataout_1541_port);
   DataPath_RF_BLOCKi_57_Q_reg_5_inst : DFF_X1 port map( D => n5245, CK => CLK,
                           Q => n_1801, QN => 
                           DataPath_RF_bus_reg_dataout_1573_port);
   DataPath_RF_BLOCKi_58_Q_reg_5_inst : DFF_X1 port map( D => n5281, CK => CLK,
                           Q => n_1802, QN => 
                           DataPath_RF_bus_reg_dataout_1605_port);
   DataPath_RF_BLOCKi_59_Q_reg_5_inst : DFF_X1 port map( D => n5316, CK => CLK,
                           Q => n_1803, QN => 
                           DataPath_RF_bus_reg_dataout_1637_port);
   DataPath_RF_BLOCKi_60_Q_reg_5_inst : DFF_X1 port map( D => n5351, CK => CLK,
                           Q => n_1804, QN => 
                           DataPath_RF_bus_reg_dataout_1669_port);
   DataPath_RF_BLOCKi_61_Q_reg_5_inst : DFF_X1 port map( D => n5386, CK => CLK,
                           Q => n_1805, QN => 
                           DataPath_RF_bus_reg_dataout_1701_port);
   DataPath_RF_BLOCKi_62_Q_reg_5_inst : DFF_X1 port map( D => n5421, CK => CLK,
                           Q => n_1806, QN => 
                           DataPath_RF_bus_reg_dataout_1733_port);
   DataPath_RF_BLOCKi_63_Q_reg_5_inst : DFF_X1 port map( D => n5456, CK => CLK,
                           Q => n_1807, QN => 
                           DataPath_RF_bus_reg_dataout_1765_port);
   DataPath_RF_BLOCKi_64_Q_reg_5_inst : DFF_X1 port map( D => n5491, CK => CLK,
                           Q => n_1808, QN => 
                           DataPath_RF_bus_reg_dataout_1797_port);
   DataPath_RF_BLOCKi_65_Q_reg_5_inst : DFF_X1 port map( D => n5526, CK => CLK,
                           Q => n_1809, QN => 
                           DataPath_RF_bus_reg_dataout_1829_port);
   DataPath_RF_BLOCKi_66_Q_reg_5_inst : DFF_X1 port map( D => n5561, CK => CLK,
                           Q => n_1810, QN => 
                           DataPath_RF_bus_reg_dataout_1861_port);
   DataPath_RF_BLOCKi_67_Q_reg_5_inst : DFF_X1 port map( D => n5596, CK => CLK,
                           Q => n_1811, QN => 
                           DataPath_RF_bus_reg_dataout_1893_port);
   DataPath_RF_BLOCKi_68_Q_reg_5_inst : DFF_X1 port map( D => n5635, CK => CLK,
                           Q => n_1812, QN => 
                           DataPath_RF_bus_reg_dataout_1925_port);
   DataPath_RF_BLOCKi_69_Q_reg_5_inst : DFF_X1 port map( D => n5672, CK => CLK,
                           Q => n_1813, QN => 
                           DataPath_RF_bus_reg_dataout_1957_port);
   DataPath_RF_BLOCKi_70_Q_reg_5_inst : DFF_X1 port map( D => n5709, CK => CLK,
                           Q => n_1814, QN => 
                           DataPath_RF_bus_reg_dataout_1989_port);
   DataPath_RF_BLOCKi_71_Q_reg_5_inst : DFF_X1 port map( D => n5746, CK => CLK,
                           Q => n_1815, QN => 
                           DataPath_RF_bus_reg_dataout_2021_port);
   DataPath_RF_BLOCKi_82_Q_reg_5_inst : DFF_X1 port map( D => n902, CK => CLK, 
                           Q => n_1816, QN => 
                           DataPath_RF_bus_reg_dataout_2373_port);
   DataPath_RF_BLOCKi_83_Q_reg_5_inst : DFF_X1 port map( D => n958, CK => CLK, 
                           Q => n_1817, QN => 
                           DataPath_RF_bus_reg_dataout_2405_port);
   DataPath_RF_BLOCKi_84_Q_reg_5_inst : DFF_X1 port map( D => n996, CK => CLK, 
                           Q => n_1818, QN => 
                           DataPath_RF_bus_reg_dataout_2437_port);
   DataPath_RF_BLOCKi_85_Q_reg_5_inst : DFF_X1 port map( D => n1033, CK => CLK,
                           Q => n_1819, QN => 
                           DataPath_RF_bus_reg_dataout_2469_port);
   DataPath_RF_BLOCKi_86_Q_reg_5_inst : DFF_X1 port map( D => n1070, CK => CLK,
                           Q => n_1820, QN => 
                           DataPath_RF_bus_reg_dataout_2501_port);
   DataPath_RF_BLOCKi_87_Q_reg_5_inst : DFF_X1 port map( D => n1107, CK => CLK,
                           Q => n_1821, QN => 
                           DataPath_RF_bus_reg_dataout_2533_port);
   DataPath_RF_BLOCKi_72_Q_reg_5_inst : DFF_X1 port map( D => n5783, CK => CLK,
                           Q => n_1822, QN => 
                           DataPath_RF_bus_reg_dataout_2053_port);
   DataPath_RF_BLOCKi_73_Q_reg_5_inst : DFF_X1 port map( D => n5822, CK => CLK,
                           Q => n_1823, QN => 
                           DataPath_RF_bus_reg_dataout_2085_port);
   DataPath_RF_BLOCKi_74_Q_reg_5_inst : DFF_X1 port map( D => n5858, CK => CLK,
                           Q => n_1824, QN => 
                           DataPath_RF_bus_reg_dataout_2117_port);
   DataPath_RF_BLOCKi_75_Q_reg_5_inst : DFF_X1 port map( D => n5894, CK => CLK,
                           Q => n_1825, QN => 
                           DataPath_RF_bus_reg_dataout_2149_port);
   DataPath_RF_BLOCKi_76_Q_reg_5_inst : DFF_X1 port map( D => n5930, CK => CLK,
                           Q => n_1826, QN => 
                           DataPath_RF_bus_reg_dataout_2181_port);
   DataPath_RF_BLOCKi_77_Q_reg_5_inst : DFF_X1 port map( D => n5966, CK => CLK,
                           Q => n_1827, QN => 
                           DataPath_RF_bus_reg_dataout_2213_port);
   DataPath_RF_BLOCKi_78_Q_reg_5_inst : DFF_X1 port map( D => n6002, CK => CLK,
                           Q => n_1828, QN => 
                           DataPath_RF_bus_reg_dataout_2245_port);
   DataPath_RF_BLOCKi_79_Q_reg_5_inst : DFF_X1 port map( D => n6038, CK => CLK,
                           Q => n_1829, QN => 
                           DataPath_RF_bus_reg_dataout_2277_port);
   DataPath_RF_BLOCKi_80_Q_reg_5_inst : DFF_X1 port map( D => n6075, CK => CLK,
                           Q => n_1830, QN => 
                           DataPath_RF_bus_reg_dataout_2309_port);
   DataPath_RF_BLOCKi_81_Q_reg_5_inst : DFF_X1 port map( D => n6111, CK => CLK,
                           Q => n_1831, QN => 
                           DataPath_RF_bus_reg_dataout_2341_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_12_inst : DFF_X1 port map( D => n2197, CK 
                           => CLK, Q => n_1832, QN => 
                           DataPath_i_REG_LDSTR_OUT_12_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_20_inst : DFF_X1 port map( D => n2189, CK 
                           => CLK, Q => n_1833, QN => 
                           DataPath_i_REG_LDSTR_OUT_20_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_28_inst : DFF_X1 port map( D => n2181, CK 
                           => CLK, Q => n_1834, QN => 
                           DataPath_i_REG_LDSTR_OUT_28_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_4_inst : DFF_X1 port map( D => n2205, CK =>
                           CLK, Q => n_1835, QN => 
                           DataPath_i_REG_LDSTR_OUT_4_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_11_inst : DFF_X1 port map( D => n2198, CK 
                           => CLK, Q => n_1836, QN => 
                           DataPath_i_REG_LDSTR_OUT_11_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_19_inst : DFF_X1 port map( D => n2190, CK 
                           => CLK, Q => n_1837, QN => 
                           DataPath_i_REG_LDSTR_OUT_19_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_27_inst : DFF_X1 port map( D => n2182, CK 
                           => CLK, Q => n_1838, QN => 
                           DataPath_i_REG_LDSTR_OUT_27_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_3_inst : DFF_X1 port map( D => n2206, CK =>
                           CLK, Q => n_1839, QN => 
                           DataPath_i_REG_LDSTR_OUT_3_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_10_inst : DFF_X1 port map( D => n2199, CK 
                           => CLK, Q => n_1840, QN => 
                           DataPath_i_REG_LDSTR_OUT_10_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_18_inst : DFF_X1 port map( D => n2191, CK 
                           => CLK, Q => n_1841, QN => 
                           DataPath_i_REG_LDSTR_OUT_18_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_26_inst : DFF_X1 port map( D => n2183, CK 
                           => CLK, Q => n_1842, QN => 
                           DataPath_i_REG_LDSTR_OUT_26_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_2_inst : DFF_X1 port map( D => n2207, CK =>
                           CLK, Q => n_1843, QN => 
                           DataPath_i_REG_LDSTR_OUT_2_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_16_inst : DFF_X1 port map( D => n2193, CK 
                           => CLK, Q => n_1844, QN => 
                           DataPath_i_REG_LDSTR_OUT_16_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_24_inst : DFF_X1 port map( D => n2185, CK 
                           => CLK, Q => n_1845, QN => 
                           DataPath_i_REG_LDSTR_OUT_24_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_8_inst : DFF_X1 port map( D => n2201, CK =>
                           CLK, Q => n_1846, QN => 
                           DataPath_i_REG_LDSTR_OUT_8_port);
   DataPath_REG_MEM_LDSTR_OUT_Q_reg_0_inst : DFF_X1 port map( D => n2209, CK =>
                           CLK, Q => n_1847, QN => 
                           DataPath_i_REG_LDSTR_OUT_0_port);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_0_inst : DFF_X1 port map( D => n6863, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_96_port,
                           QN => n663);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_0_inst : DFF_X1 port map( D => n6895, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_128_port
                           , QN => n695);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_0_inst : DFF_X1 port map( D => n6959, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_192_port
                           , QN => n759);
   DataPath_RF_BLOCKi_8_Q_reg_0_inst : DFF_X1 port map( D => n3372, CK => CLK, 
                           Q => n_1848, QN => 
                           DataPath_RF_bus_reg_dataout_0_port);
   DataPath_RF_BLOCKi_9_Q_reg_0_inst : DFF_X1 port map( D => n3412, CK => CLK, 
                           Q => n_1849, QN => 
                           DataPath_RF_bus_reg_dataout_32_port);
   DataPath_RF_BLOCKi_10_Q_reg_0_inst : DFF_X1 port map( D => n3450, CK => CLK,
                           Q => n_1850, QN => 
                           DataPath_RF_bus_reg_dataout_64_port);
   DataPath_RF_BLOCKi_11_Q_reg_0_inst : DFF_X1 port map( D => n3488, CK => CLK,
                           Q => n_1851, QN => 
                           DataPath_RF_bus_reg_dataout_96_port);
   DataPath_RF_BLOCKi_12_Q_reg_0_inst : DFF_X1 port map( D => n3526, CK => CLK,
                           Q => n_1852, QN => 
                           DataPath_RF_bus_reg_dataout_128_port);
   DataPath_RF_BLOCKi_13_Q_reg_0_inst : DFF_X1 port map( D => n3564, CK => CLK,
                           Q => n_1853, QN => 
                           DataPath_RF_bus_reg_dataout_160_port);
   DataPath_RF_BLOCKi_14_Q_reg_0_inst : DFF_X1 port map( D => n3602, CK => CLK,
                           Q => n_1854, QN => 
                           DataPath_RF_bus_reg_dataout_192_port);
   DataPath_RF_BLOCKi_15_Q_reg_0_inst : DFF_X1 port map( D => n3640, CK => CLK,
                           Q => n_1855, QN => 
                           DataPath_RF_bus_reg_dataout_224_port);
   DataPath_RF_BLOCKi_16_Q_reg_0_inst : DFF_X1 port map( D => n3678, CK => CLK,
                           Q => n_1856, QN => 
                           DataPath_RF_bus_reg_dataout_256_port);
   DataPath_RF_BLOCKi_17_Q_reg_0_inst : DFF_X1 port map( D => n3715, CK => CLK,
                           Q => n_1857, QN => 
                           DataPath_RF_bus_reg_dataout_288_port);
   DataPath_RF_BLOCKi_18_Q_reg_0_inst : DFF_X1 port map( D => n3752, CK => CLK,
                           Q => n_1858, QN => 
                           DataPath_RF_bus_reg_dataout_320_port);
   DataPath_RF_BLOCKi_19_Q_reg_0_inst : DFF_X1 port map( D => n3789, CK => CLK,
                           Q => n_1859, QN => 
                           DataPath_RF_bus_reg_dataout_352_port);
   DataPath_RF_BLOCKi_20_Q_reg_0_inst : DFF_X1 port map( D => n3824, CK => CLK,
                           Q => n_1860, QN => 
                           DataPath_RF_bus_reg_dataout_384_port);
   DataPath_RF_BLOCKi_21_Q_reg_0_inst : DFF_X1 port map( D => n3859, CK => CLK,
                           Q => n_1861, QN => 
                           DataPath_RF_bus_reg_dataout_416_port);
   DataPath_RF_BLOCKi_22_Q_reg_0_inst : DFF_X1 port map( D => n3894, CK => CLK,
                           Q => n_1862, QN => 
                           DataPath_RF_bus_reg_dataout_448_port);
   DataPath_RF_BLOCKi_23_Q_reg_0_inst : DFF_X1 port map( D => n3960, CK => CLK,
                           Q => n_1863, QN => 
                           DataPath_RF_bus_reg_dataout_480_port);
   DataPath_RF_BLOCKi_24_Q_reg_0_inst : DFF_X1 port map( D => n4028, CK => CLK,
                           Q => n_1864, QN => 
                           DataPath_RF_bus_reg_dataout_512_port);
   DataPath_RF_BLOCKi_25_Q_reg_0_inst : DFF_X1 port map( D => n4065, CK => CLK,
                           Q => n_1865, QN => 
                           DataPath_RF_bus_reg_dataout_544_port);
   DataPath_RF_BLOCKi_26_Q_reg_0_inst : DFF_X1 port map( D => n4100, CK => CLK,
                           Q => n_1866, QN => 
                           DataPath_RF_bus_reg_dataout_576_port);
   DataPath_RF_BLOCKi_27_Q_reg_0_inst : DFF_X1 port map( D => n4135, CK => CLK,
                           Q => n_1867, QN => 
                           DataPath_RF_bus_reg_dataout_608_port);
   DataPath_RF_BLOCKi_28_Q_reg_0_inst : DFF_X1 port map( D => n4170, CK => CLK,
                           Q => n_1868, QN => 
                           DataPath_RF_bus_reg_dataout_640_port);
   DataPath_RF_BLOCKi_29_Q_reg_0_inst : DFF_X1 port map( D => n4205, CK => CLK,
                           Q => n_1869, QN => 
                           DataPath_RF_bus_reg_dataout_672_port);
   DataPath_RF_BLOCKi_30_Q_reg_0_inst : DFF_X1 port map( D => n4240, CK => CLK,
                           Q => n_1870, QN => 
                           DataPath_RF_bus_reg_dataout_704_port);
   DataPath_RF_BLOCKi_31_Q_reg_0_inst : DFF_X1 port map( D => n4275, CK => CLK,
                           Q => n_1871, QN => 
                           DataPath_RF_bus_reg_dataout_736_port);
   DataPath_RF_BLOCKi_32_Q_reg_0_inst : DFF_X1 port map( D => n4310, CK => CLK,
                           Q => n_1872, QN => 
                           DataPath_RF_bus_reg_dataout_768_port);
   DataPath_RF_BLOCKi_33_Q_reg_0_inst : DFF_X1 port map( D => n4345, CK => CLK,
                           Q => n_1873, QN => 
                           DataPath_RF_bus_reg_dataout_800_port);
   DataPath_RF_BLOCKi_34_Q_reg_0_inst : DFF_X1 port map( D => n4380, CK => CLK,
                           Q => n_1874, QN => 
                           DataPath_RF_bus_reg_dataout_832_port);
   DataPath_RF_BLOCKi_35_Q_reg_0_inst : DFF_X1 port map( D => n4415, CK => CLK,
                           Q => n_1875, QN => 
                           DataPath_RF_bus_reg_dataout_864_port);
   DataPath_RF_BLOCKi_36_Q_reg_0_inst : DFF_X1 port map( D => n4450, CK => CLK,
                           Q => n_1876, QN => 
                           DataPath_RF_bus_reg_dataout_896_port);
   DataPath_RF_BLOCKi_37_Q_reg_0_inst : DFF_X1 port map( D => n4485, CK => CLK,
                           Q => n_1877, QN => 
                           DataPath_RF_bus_reg_dataout_928_port);
   DataPath_RF_BLOCKi_38_Q_reg_0_inst : DFF_X1 port map( D => n4520, CK => CLK,
                           Q => n_1878, QN => 
                           DataPath_RF_bus_reg_dataout_960_port);
   DataPath_RF_BLOCKi_39_Q_reg_0_inst : DFF_X1 port map( D => n4555, CK => CLK,
                           Q => n_1879, QN => 
                           DataPath_RF_bus_reg_dataout_992_port);
   DataPath_RF_BLOCKi_40_Q_reg_0_inst : DFF_X1 port map( D => n4621, CK => CLK,
                           Q => n_1880, QN => 
                           DataPath_RF_bus_reg_dataout_1024_port);
   DataPath_RF_BLOCKi_41_Q_reg_0_inst : DFF_X1 port map( D => n4658, CK => CLK,
                           Q => n_1881, QN => 
                           DataPath_RF_bus_reg_dataout_1056_port);
   DataPath_RF_BLOCKi_42_Q_reg_0_inst : DFF_X1 port map( D => n4693, CK => CLK,
                           Q => n_1882, QN => 
                           DataPath_RF_bus_reg_dataout_1088_port);
   DataPath_RF_BLOCKi_43_Q_reg_0_inst : DFF_X1 port map( D => n4728, CK => CLK,
                           Q => n_1883, QN => 
                           DataPath_RF_bus_reg_dataout_1120_port);
   DataPath_RF_BLOCKi_44_Q_reg_0_inst : DFF_X1 port map( D => n4763, CK => CLK,
                           Q => n_1884, QN => 
                           DataPath_RF_bus_reg_dataout_1152_port);
   DataPath_RF_BLOCKi_45_Q_reg_0_inst : DFF_X1 port map( D => n4798, CK => CLK,
                           Q => n_1885, QN => 
                           DataPath_RF_bus_reg_dataout_1184_port);
   DataPath_RF_BLOCKi_46_Q_reg_0_inst : DFF_X1 port map( D => n4833, CK => CLK,
                           Q => n_1886, QN => 
                           DataPath_RF_bus_reg_dataout_1216_port);
   DataPath_RF_BLOCKi_47_Q_reg_0_inst : DFF_X1 port map( D => n4868, CK => CLK,
                           Q => n_1887, QN => 
                           DataPath_RF_bus_reg_dataout_1248_port);
   DataPath_RF_BLOCKi_48_Q_reg_0_inst : DFF_X1 port map( D => n4903, CK => CLK,
                           Q => n_1888, QN => 
                           DataPath_RF_bus_reg_dataout_1280_port);
   DataPath_RF_BLOCKi_49_Q_reg_0_inst : DFF_X1 port map( D => n4938, CK => CLK,
                           Q => n_1889, QN => 
                           DataPath_RF_bus_reg_dataout_1312_port);
   DataPath_RF_BLOCKi_50_Q_reg_0_inst : DFF_X1 port map( D => n4973, CK => CLK,
                           Q => n_1890, QN => 
                           DataPath_RF_bus_reg_dataout_1344_port);
   DataPath_RF_BLOCKi_51_Q_reg_0_inst : DFF_X1 port map( D => n5008, CK => CLK,
                           Q => n_1891, QN => 
                           DataPath_RF_bus_reg_dataout_1376_port);
   DataPath_RF_BLOCKi_52_Q_reg_0_inst : DFF_X1 port map( D => n5043, CK => CLK,
                           Q => n_1892, QN => 
                           DataPath_RF_bus_reg_dataout_1408_port);
   DataPath_RF_BLOCKi_53_Q_reg_0_inst : DFF_X1 port map( D => n5078, CK => CLK,
                           Q => n_1893, QN => 
                           DataPath_RF_bus_reg_dataout_1440_port);
   DataPath_RF_BLOCKi_54_Q_reg_0_inst : DFF_X1 port map( D => n5113, CK => CLK,
                           Q => n_1894, QN => 
                           DataPath_RF_bus_reg_dataout_1472_port);
   DataPath_RF_BLOCKi_55_Q_reg_0_inst : DFF_X1 port map( D => n5148, CK => CLK,
                           Q => n_1895, QN => 
                           DataPath_RF_bus_reg_dataout_1504_port);
   DataPath_RF_BLOCKi_56_Q_reg_0_inst : DFF_X1 port map( D => n5214, CK => CLK,
                           Q => n_1896, QN => 
                           DataPath_RF_bus_reg_dataout_1536_port);
   DataPath_RF_BLOCKi_57_Q_reg_0_inst : DFF_X1 port map( D => n5250, CK => CLK,
                           Q => n_1897, QN => 
                           DataPath_RF_bus_reg_dataout_1568_port);
   DataPath_RF_BLOCKi_58_Q_reg_0_inst : DFF_X1 port map( D => n5286, CK => CLK,
                           Q => n_1898, QN => 
                           DataPath_RF_bus_reg_dataout_1600_port);
   DataPath_RF_BLOCKi_59_Q_reg_0_inst : DFF_X1 port map( D => n5321, CK => CLK,
                           Q => n_1899, QN => 
                           DataPath_RF_bus_reg_dataout_1632_port);
   DataPath_RF_BLOCKi_60_Q_reg_0_inst : DFF_X1 port map( D => n5356, CK => CLK,
                           Q => n_1900, QN => 
                           DataPath_RF_bus_reg_dataout_1664_port);
   DataPath_RF_BLOCKi_61_Q_reg_0_inst : DFF_X1 port map( D => n5391, CK => CLK,
                           Q => n_1901, QN => 
                           DataPath_RF_bus_reg_dataout_1696_port);
   DataPath_RF_BLOCKi_62_Q_reg_0_inst : DFF_X1 port map( D => n5426, CK => CLK,
                           Q => n_1902, QN => 
                           DataPath_RF_bus_reg_dataout_1728_port);
   DataPath_RF_BLOCKi_63_Q_reg_0_inst : DFF_X1 port map( D => n5461, CK => CLK,
                           Q => n_1903, QN => 
                           DataPath_RF_bus_reg_dataout_1760_port);
   DataPath_RF_BLOCKi_64_Q_reg_0_inst : DFF_X1 port map( D => n5496, CK => CLK,
                           Q => n_1904, QN => 
                           DataPath_RF_bus_reg_dataout_1792_port);
   DataPath_RF_BLOCKi_65_Q_reg_0_inst : DFF_X1 port map( D => n5531, CK => CLK,
                           Q => n_1905, QN => 
                           DataPath_RF_bus_reg_dataout_1824_port);
   DataPath_RF_BLOCKi_66_Q_reg_0_inst : DFF_X1 port map( D => n5566, CK => CLK,
                           Q => n_1906, QN => 
                           DataPath_RF_bus_reg_dataout_1856_port);
   DataPath_RF_BLOCKi_67_Q_reg_0_inst : DFF_X1 port map( D => n5601, CK => CLK,
                           Q => n_1907, QN => 
                           DataPath_RF_bus_reg_dataout_1888_port);
   DataPath_RF_BLOCKi_68_Q_reg_0_inst : DFF_X1 port map( D => n5640, CK => CLK,
                           Q => n_1908, QN => 
                           DataPath_RF_bus_reg_dataout_1920_port);
   DataPath_RF_BLOCKi_69_Q_reg_0_inst : DFF_X1 port map( D => n5677, CK => CLK,
                           Q => n_1909, QN => 
                           DataPath_RF_bus_reg_dataout_1952_port);
   DataPath_RF_BLOCKi_70_Q_reg_0_inst : DFF_X1 port map( D => n5714, CK => CLK,
                           Q => n_1910, QN => 
                           DataPath_RF_bus_reg_dataout_1984_port);
   DataPath_RF_BLOCKi_71_Q_reg_0_inst : DFF_X1 port map( D => n5751, CK => CLK,
                           Q => n_1911, QN => 
                           DataPath_RF_bus_reg_dataout_2016_port);
   DataPath_RF_BLOCKi_82_Q_reg_0_inst : DFF_X1 port map( D => n912, CK => CLK, 
                           Q => n_1912, QN => 
                           DataPath_RF_bus_reg_dataout_2368_port);
   DataPath_RF_BLOCKi_83_Q_reg_0_inst : DFF_X1 port map( D => n963, CK => CLK, 
                           Q => n_1913, QN => 
                           DataPath_RF_bus_reg_dataout_2400_port);
   DataPath_RF_BLOCKi_84_Q_reg_0_inst : DFF_X1 port map( D => n1001, CK => CLK,
                           Q => n_1914, QN => 
                           DataPath_RF_bus_reg_dataout_2432_port);
   DataPath_RF_BLOCKi_85_Q_reg_0_inst : DFF_X1 port map( D => n1038, CK => CLK,
                           Q => n_1915, QN => 
                           DataPath_RF_bus_reg_dataout_2464_port);
   DataPath_RF_BLOCKi_86_Q_reg_0_inst : DFF_X1 port map( D => n1075, CK => CLK,
                           Q => n_1916, QN => 
                           DataPath_RF_bus_reg_dataout_2496_port);
   DataPath_RF_BLOCKi_87_Q_reg_0_inst : DFF_X1 port map( D => n1112, CK => CLK,
                           Q => n_1917, QN => 
                           DataPath_RF_bus_reg_dataout_2528_port);
   DataPath_RF_BLOCKi_73_Q_reg_0_inst : DFF_X1 port map( D => n5827, CK => CLK,
                           Q => n_1918, QN => 
                           DataPath_RF_bus_reg_dataout_2080_port);
   DataPath_RF_BLOCKi_74_Q_reg_0_inst : DFF_X1 port map( D => n5863, CK => CLK,
                           Q => n_1919, QN => 
                           DataPath_RF_bus_reg_dataout_2112_port);
   DataPath_RF_BLOCKi_75_Q_reg_0_inst : DFF_X1 port map( D => n5899, CK => CLK,
                           Q => n_1920, QN => 
                           DataPath_RF_bus_reg_dataout_2144_port);
   DataPath_RF_BLOCKi_76_Q_reg_0_inst : DFF_X1 port map( D => n5935, CK => CLK,
                           Q => n_1921, QN => 
                           DataPath_RF_bus_reg_dataout_2176_port);
   DataPath_RF_BLOCKi_77_Q_reg_0_inst : DFF_X1 port map( D => n5971, CK => CLK,
                           Q => n_1922, QN => 
                           DataPath_RF_bus_reg_dataout_2208_port);
   DataPath_RF_BLOCKi_78_Q_reg_0_inst : DFF_X1 port map( D => n6007, CK => CLK,
                           Q => n_1923, QN => 
                           DataPath_RF_bus_reg_dataout_2240_port);
   DataPath_RF_BLOCKi_79_Q_reg_0_inst : DFF_X1 port map( D => n6043, CK => CLK,
                           Q => n_1924, QN => 
                           DataPath_RF_bus_reg_dataout_2272_port);
   DataPath_RF_BLOCKi_80_Q_reg_0_inst : DFF_X1 port map( D => n6080, CK => CLK,
                           Q => n_1925, QN => 
                           DataPath_RF_bus_reg_dataout_2304_port);
   DataPath_RF_BLOCKi_81_Q_reg_0_inst : DFF_X1 port map( D => n6116, CK => CLK,
                           Q => n_1926, QN => 
                           DataPath_RF_bus_reg_dataout_2336_port);
   DataPath_REG_ALU_OUT_Q_reg_21_inst : DFF_X1 port map( D => n7002, CK => CLK,
                           Q => DRAM_ADDRESS_21_port, QN => n8329);
   DataPath_REG_MEM_ALUOUT_Q_reg_21_inst : DFF_X1 port map( D => n1128, CK => 
                           CLK, Q => n_1927, QN => 
                           DataPath_i_REG_MEM_ALUOUT_21_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_21_inst : DFF_X1 port map( D => n6778, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_53_port,
                           QN => n620);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_21_inst : DFF_X1 port map( D => n6810, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_85_port,
                           QN => n652);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_21_inst : DFF_X1 port map( D => n6842, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_117_port
                           , QN => n684);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_21_inst : DFF_X1 port map( D => n6874, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_149_port
                           , QN => n716);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_21_inst : DFF_X1 port map( D => n6906, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_181_port
                           , QN => n748);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_21_inst : DFF_X1 port map( D => n6938, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_213_port
                           , QN => n780);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_21_inst : DFF_X1 port map( D => n6970, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_245_port
                           , QN => n812);
   DataPath_RF_BLOCKi_8_Q_reg_21_inst : DFF_X1 port map( D => n3330, CK => CLK,
                           Q => n_1928, QN => 
                           DataPath_RF_bus_reg_dataout_21_port);
   DataPath_RF_BLOCKi_9_Q_reg_21_inst : DFF_X1 port map( D => n3391, CK => CLK,
                           Q => n_1929, QN => 
                           DataPath_RF_bus_reg_dataout_53_port);
   DataPath_RF_BLOCKi_10_Q_reg_21_inst : DFF_X1 port map( D => n3429, CK => CLK
                           , Q => n_1930, QN => 
                           DataPath_RF_bus_reg_dataout_85_port);
   DataPath_RF_BLOCKi_11_Q_reg_21_inst : DFF_X1 port map( D => n3467, CK => CLK
                           , Q => n_1931, QN => 
                           DataPath_RF_bus_reg_dataout_117_port);
   DataPath_RF_BLOCKi_12_Q_reg_21_inst : DFF_X1 port map( D => n3505, CK => CLK
                           , Q => n_1932, QN => 
                           DataPath_RF_bus_reg_dataout_149_port);
   DataPath_RF_BLOCKi_13_Q_reg_21_inst : DFF_X1 port map( D => n3543, CK => CLK
                           , Q => n_1933, QN => 
                           DataPath_RF_bus_reg_dataout_181_port);
   DataPath_RF_BLOCKi_14_Q_reg_21_inst : DFF_X1 port map( D => n3581, CK => CLK
                           , Q => n_1934, QN => 
                           DataPath_RF_bus_reg_dataout_213_port);
   DataPath_RF_BLOCKi_15_Q_reg_21_inst : DFF_X1 port map( D => n3619, CK => CLK
                           , Q => n_1935, QN => 
                           DataPath_RF_bus_reg_dataout_245_port);
   DataPath_RF_BLOCKi_16_Q_reg_21_inst : DFF_X1 port map( D => n3657, CK => CLK
                           , Q => n_1936, QN => 
                           DataPath_RF_bus_reg_dataout_277_port);
   DataPath_RF_BLOCKi_17_Q_reg_21_inst : DFF_X1 port map( D => n3694, CK => CLK
                           , Q => n_1937, QN => 
                           DataPath_RF_bus_reg_dataout_309_port);
   DataPath_RF_BLOCKi_18_Q_reg_21_inst : DFF_X1 port map( D => n3731, CK => CLK
                           , Q => n_1938, QN => 
                           DataPath_RF_bus_reg_dataout_341_port);
   DataPath_RF_BLOCKi_19_Q_reg_21_inst : DFF_X1 port map( D => n3768, CK => CLK
                           , Q => n_1939, QN => 
                           DataPath_RF_bus_reg_dataout_373_port);
   DataPath_RF_BLOCKi_20_Q_reg_21_inst : DFF_X1 port map( D => n3803, CK => CLK
                           , Q => n_1940, QN => 
                           DataPath_RF_bus_reg_dataout_405_port);
   DataPath_RF_BLOCKi_21_Q_reg_21_inst : DFF_X1 port map( D => n3838, CK => CLK
                           , Q => n_1941, QN => 
                           DataPath_RF_bus_reg_dataout_437_port);
   DataPath_RF_BLOCKi_22_Q_reg_21_inst : DFF_X1 port map( D => n3873, CK => CLK
                           , Q => n_1942, QN => 
                           DataPath_RF_bus_reg_dataout_469_port);
   DataPath_RF_BLOCKi_23_Q_reg_21_inst : DFF_X1 port map( D => n3918, CK => CLK
                           , Q => n_1943, QN => 
                           DataPath_RF_bus_reg_dataout_501_port);
   DataPath_RF_BLOCKi_24_Q_reg_21_inst : DFF_X1 port map( D => n3986, CK => CLK
                           , Q => n_1944, QN => 
                           DataPath_RF_bus_reg_dataout_533_port);
   DataPath_RF_BLOCKi_25_Q_reg_21_inst : DFF_X1 port map( D => n4044, CK => CLK
                           , Q => n_1945, QN => 
                           DataPath_RF_bus_reg_dataout_565_port);
   DataPath_RF_BLOCKi_26_Q_reg_21_inst : DFF_X1 port map( D => n4079, CK => CLK
                           , Q => n_1946, QN => 
                           DataPath_RF_bus_reg_dataout_597_port);
   DataPath_RF_BLOCKi_27_Q_reg_21_inst : DFF_X1 port map( D => n4114, CK => CLK
                           , Q => n_1947, QN => 
                           DataPath_RF_bus_reg_dataout_629_port);
   DataPath_RF_BLOCKi_28_Q_reg_21_inst : DFF_X1 port map( D => n4149, CK => CLK
                           , Q => n_1948, QN => 
                           DataPath_RF_bus_reg_dataout_661_port);
   DataPath_RF_BLOCKi_29_Q_reg_21_inst : DFF_X1 port map( D => n4184, CK => CLK
                           , Q => n_1949, QN => 
                           DataPath_RF_bus_reg_dataout_693_port);
   DataPath_RF_BLOCKi_30_Q_reg_21_inst : DFF_X1 port map( D => n4219, CK => CLK
                           , Q => n_1950, QN => 
                           DataPath_RF_bus_reg_dataout_725_port);
   DataPath_RF_BLOCKi_31_Q_reg_21_inst : DFF_X1 port map( D => n4254, CK => CLK
                           , Q => n_1951, QN => 
                           DataPath_RF_bus_reg_dataout_757_port);
   DataPath_RF_BLOCKi_32_Q_reg_21_inst : DFF_X1 port map( D => n4289, CK => CLK
                           , Q => n_1952, QN => 
                           DataPath_RF_bus_reg_dataout_789_port);
   DataPath_RF_BLOCKi_33_Q_reg_21_inst : DFF_X1 port map( D => n4324, CK => CLK
                           , Q => n_1953, QN => 
                           DataPath_RF_bus_reg_dataout_821_port);
   DataPath_RF_BLOCKi_34_Q_reg_21_inst : DFF_X1 port map( D => n4359, CK => CLK
                           , Q => n_1954, QN => 
                           DataPath_RF_bus_reg_dataout_853_port);
   DataPath_RF_BLOCKi_35_Q_reg_21_inst : DFF_X1 port map( D => n4394, CK => CLK
                           , Q => n_1955, QN => 
                           DataPath_RF_bus_reg_dataout_885_port);
   DataPath_RF_BLOCKi_36_Q_reg_21_inst : DFF_X1 port map( D => n4429, CK => CLK
                           , Q => n_1956, QN => 
                           DataPath_RF_bus_reg_dataout_917_port);
   DataPath_RF_BLOCKi_37_Q_reg_21_inst : DFF_X1 port map( D => n4464, CK => CLK
                           , Q => n_1957, QN => 
                           DataPath_RF_bus_reg_dataout_949_port);
   DataPath_RF_BLOCKi_38_Q_reg_21_inst : DFF_X1 port map( D => n4499, CK => CLK
                           , Q => n_1958, QN => 
                           DataPath_RF_bus_reg_dataout_981_port);
   DataPath_RF_BLOCKi_39_Q_reg_21_inst : DFF_X1 port map( D => n4534, CK => CLK
                           , Q => n_1959, QN => 
                           DataPath_RF_bus_reg_dataout_1013_port);
   DataPath_RF_BLOCKi_40_Q_reg_21_inst : DFF_X1 port map( D => n4579, CK => CLK
                           , Q => n_1960, QN => 
                           DataPath_RF_bus_reg_dataout_1045_port);
   DataPath_RF_BLOCKi_41_Q_reg_21_inst : DFF_X1 port map( D => n4637, CK => CLK
                           , Q => n_1961, QN => 
                           DataPath_RF_bus_reg_dataout_1077_port);
   DataPath_RF_BLOCKi_42_Q_reg_21_inst : DFF_X1 port map( D => n4672, CK => CLK
                           , Q => n_1962, QN => 
                           DataPath_RF_bus_reg_dataout_1109_port);
   DataPath_RF_BLOCKi_43_Q_reg_21_inst : DFF_X1 port map( D => n4707, CK => CLK
                           , Q => n_1963, QN => 
                           DataPath_RF_bus_reg_dataout_1141_port);
   DataPath_RF_BLOCKi_44_Q_reg_21_inst : DFF_X1 port map( D => n4742, CK => CLK
                           , Q => n_1964, QN => 
                           DataPath_RF_bus_reg_dataout_1173_port);
   DataPath_RF_BLOCKi_45_Q_reg_21_inst : DFF_X1 port map( D => n4777, CK => CLK
                           , Q => n_1965, QN => 
                           DataPath_RF_bus_reg_dataout_1205_port);
   DataPath_RF_BLOCKi_46_Q_reg_21_inst : DFF_X1 port map( D => n4812, CK => CLK
                           , Q => n_1966, QN => 
                           DataPath_RF_bus_reg_dataout_1237_port);
   DataPath_RF_BLOCKi_47_Q_reg_21_inst : DFF_X1 port map( D => n4847, CK => CLK
                           , Q => n_1967, QN => 
                           DataPath_RF_bus_reg_dataout_1269_port);
   DataPath_RF_BLOCKi_48_Q_reg_21_inst : DFF_X1 port map( D => n4882, CK => CLK
                           , Q => n_1968, QN => 
                           DataPath_RF_bus_reg_dataout_1301_port);
   DataPath_RF_BLOCKi_49_Q_reg_21_inst : DFF_X1 port map( D => n4917, CK => CLK
                           , Q => n_1969, QN => 
                           DataPath_RF_bus_reg_dataout_1333_port);
   DataPath_RF_BLOCKi_50_Q_reg_21_inst : DFF_X1 port map( D => n4952, CK => CLK
                           , Q => n_1970, QN => 
                           DataPath_RF_bus_reg_dataout_1365_port);
   DataPath_RF_BLOCKi_51_Q_reg_21_inst : DFF_X1 port map( D => n4987, CK => CLK
                           , Q => n_1971, QN => 
                           DataPath_RF_bus_reg_dataout_1397_port);
   DataPath_RF_BLOCKi_52_Q_reg_21_inst : DFF_X1 port map( D => n5022, CK => CLK
                           , Q => n_1972, QN => 
                           DataPath_RF_bus_reg_dataout_1429_port);
   DataPath_RF_BLOCKi_53_Q_reg_21_inst : DFF_X1 port map( D => n5057, CK => CLK
                           , Q => n_1973, QN => 
                           DataPath_RF_bus_reg_dataout_1461_port);
   DataPath_RF_BLOCKi_54_Q_reg_21_inst : DFF_X1 port map( D => n5092, CK => CLK
                           , Q => n_1974, QN => 
                           DataPath_RF_bus_reg_dataout_1493_port);
   DataPath_RF_BLOCKi_55_Q_reg_21_inst : DFF_X1 port map( D => n5127, CK => CLK
                           , Q => n_1975, QN => 
                           DataPath_RF_bus_reg_dataout_1525_port);
   DataPath_RF_BLOCKi_56_Q_reg_21_inst : DFF_X1 port map( D => n5172, CK => CLK
                           , Q => n_1976, QN => 
                           DataPath_RF_bus_reg_dataout_1557_port);
   DataPath_RF_BLOCKi_57_Q_reg_21_inst : DFF_X1 port map( D => n5229, CK => CLK
                           , Q => n_1977, QN => 
                           DataPath_RF_bus_reg_dataout_1589_port);
   DataPath_RF_BLOCKi_58_Q_reg_21_inst : DFF_X1 port map( D => n5265, CK => CLK
                           , Q => n_1978, QN => 
                           DataPath_RF_bus_reg_dataout_1621_port);
   DataPath_RF_BLOCKi_59_Q_reg_21_inst : DFF_X1 port map( D => n5300, CK => CLK
                           , Q => n_1979, QN => 
                           DataPath_RF_bus_reg_dataout_1653_port);
   DataPath_RF_BLOCKi_60_Q_reg_21_inst : DFF_X1 port map( D => n5335, CK => CLK
                           , Q => n_1980, QN => 
                           DataPath_RF_bus_reg_dataout_1685_port);
   DataPath_RF_BLOCKi_61_Q_reg_21_inst : DFF_X1 port map( D => n5370, CK => CLK
                           , Q => n_1981, QN => 
                           DataPath_RF_bus_reg_dataout_1717_port);
   DataPath_RF_BLOCKi_62_Q_reg_21_inst : DFF_X1 port map( D => n5405, CK => CLK
                           , Q => n_1982, QN => 
                           DataPath_RF_bus_reg_dataout_1749_port);
   DataPath_RF_BLOCKi_63_Q_reg_21_inst : DFF_X1 port map( D => n5440, CK => CLK
                           , Q => n_1983, QN => 
                           DataPath_RF_bus_reg_dataout_1781_port);
   DataPath_RF_BLOCKi_64_Q_reg_21_inst : DFF_X1 port map( D => n5475, CK => CLK
                           , Q => n_1984, QN => 
                           DataPath_RF_bus_reg_dataout_1813_port);
   DataPath_RF_BLOCKi_65_Q_reg_21_inst : DFF_X1 port map( D => n5510, CK => CLK
                           , Q => n_1985, QN => 
                           DataPath_RF_bus_reg_dataout_1845_port);
   DataPath_RF_BLOCKi_66_Q_reg_21_inst : DFF_X1 port map( D => n5545, CK => CLK
                           , Q => n_1986, QN => 
                           DataPath_RF_bus_reg_dataout_1877_port);
   DataPath_RF_BLOCKi_67_Q_reg_21_inst : DFF_X1 port map( D => n5580, CK => CLK
                           , Q => n_1987, QN => 
                           DataPath_RF_bus_reg_dataout_1909_port);
   DataPath_RF_BLOCKi_68_Q_reg_21_inst : DFF_X1 port map( D => n5619, CK => CLK
                           , Q => n_1988, QN => 
                           DataPath_RF_bus_reg_dataout_1941_port);
   DataPath_RF_BLOCKi_69_Q_reg_21_inst : DFF_X1 port map( D => n5656, CK => CLK
                           , Q => n_1989, QN => 
                           DataPath_RF_bus_reg_dataout_1973_port);
   DataPath_RF_BLOCKi_70_Q_reg_21_inst : DFF_X1 port map( D => n5693, CK => CLK
                           , Q => n_1990, QN => 
                           DataPath_RF_bus_reg_dataout_2005_port);
   DataPath_RF_BLOCKi_71_Q_reg_21_inst : DFF_X1 port map( D => n5730, CK => CLK
                           , Q => n_1991, QN => 
                           DataPath_RF_bus_reg_dataout_2037_port);
   DataPath_RF_BLOCKi_83_Q_reg_21_inst : DFF_X1 port map( D => n936, CK => CLK,
                           Q => n_1992, QN => 
                           DataPath_RF_bus_reg_dataout_2421_port);
   DataPath_RF_BLOCKi_84_Q_reg_21_inst : DFF_X1 port map( D => n980, CK => CLK,
                           Q => n_1993, QN => 
                           DataPath_RF_bus_reg_dataout_2453_port);
   DataPath_RF_BLOCKi_85_Q_reg_21_inst : DFF_X1 port map( D => n1017, CK => CLK
                           , Q => n_1994, QN => 
                           DataPath_RF_bus_reg_dataout_2485_port);
   DataPath_RF_BLOCKi_86_Q_reg_21_inst : DFF_X1 port map( D => n1054, CK => CLK
                           , Q => n_1995, QN => 
                           DataPath_RF_bus_reg_dataout_2517_port);
   DataPath_RF_BLOCKi_87_Q_reg_21_inst : DFF_X1 port map( D => n1091, CK => CLK
                           , Q => n_1996, QN => 
                           DataPath_RF_bus_reg_dataout_2549_port);
   DataPath_RF_BLOCKi_72_Q_reg_21_inst : DFF_X1 port map( D => n5767, CK => CLK
                           , Q => n_1997, QN => 
                           DataPath_RF_bus_reg_dataout_2069_port);
   DataPath_RF_BLOCKi_73_Q_reg_21_inst : DFF_X1 port map( D => n5806, CK => CLK
                           , Q => n_1998, QN => 
                           DataPath_RF_bus_reg_dataout_2101_port);
   DataPath_RF_BLOCKi_74_Q_reg_21_inst : DFF_X1 port map( D => n5842, CK => CLK
                           , Q => n_1999, QN => 
                           DataPath_RF_bus_reg_dataout_2133_port);
   DataPath_RF_BLOCKi_75_Q_reg_21_inst : DFF_X1 port map( D => n5878, CK => CLK
                           , Q => n_2000, QN => 
                           DataPath_RF_bus_reg_dataout_2165_port);
   DataPath_RF_BLOCKi_76_Q_reg_21_inst : DFF_X1 port map( D => n5914, CK => CLK
                           , Q => n_2001, QN => 
                           DataPath_RF_bus_reg_dataout_2197_port);
   DataPath_RF_BLOCKi_77_Q_reg_21_inst : DFF_X1 port map( D => n5950, CK => CLK
                           , Q => n_2002, QN => 
                           DataPath_RF_bus_reg_dataout_2229_port);
   DataPath_RF_BLOCKi_78_Q_reg_21_inst : DFF_X1 port map( D => n5986, CK => CLK
                           , Q => n_2003, QN => 
                           DataPath_RF_bus_reg_dataout_2261_port);
   DataPath_RF_BLOCKi_79_Q_reg_21_inst : DFF_X1 port map( D => n6022, CK => CLK
                           , Q => n_2004, QN => 
                           DataPath_RF_bus_reg_dataout_2293_port);
   DataPath_RF_BLOCKi_80_Q_reg_21_inst : DFF_X1 port map( D => n6059, CK => CLK
                           , Q => n_2005, QN => 
                           DataPath_RF_bus_reg_dataout_2325_port);
   DataPath_RF_BLOCKi_81_Q_reg_21_inst : DFF_X1 port map( D => n6095, CK => CLK
                           , Q => n_2006, QN => 
                           DataPath_RF_bus_reg_dataout_2357_port);
   DataPath_RF_BLOCKi_82_Q_reg_21_inst : DFF_X1 port map( D => n6129, CK => CLK
                           , Q => n_2007, QN => 
                           DataPath_RF_bus_reg_dataout_2389_port);
   DataPath_REG_ALU_OUT_Q_reg_25_inst : DFF_X1 port map( D => n6998, CK => CLK,
                           Q => DRAM_ADDRESS_25_port, QN => n8328);
   DataPath_REG_MEM_ALUOUT_Q_reg_25_inst : DFF_X1 port map( D => n1124, CK => 
                           CLK, Q => n_2008, QN => 
                           DataPath_i_REG_MEM_ALUOUT_25_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_25_inst : DFF_X1 port map( D => n6774, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_57_port,
                           QN => n624);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_25_inst : DFF_X1 port map( D => n6806, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_89_port,
                           QN => n656);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_25_inst : DFF_X1 port map( D => n6838, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_121_port
                           , QN => n688);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_25_inst : DFF_X1 port map( D => n6870, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_153_port
                           , QN => n720);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_25_inst : DFF_X1 port map( D => n6902, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_185_port
                           , QN => n752);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_25_inst : DFF_X1 port map( D => n6934, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_217_port
                           , QN => n784);
   DataPath_RF_BLOCKi_8_Q_reg_25_inst : DFF_X1 port map( D => n3322, CK => CLK,
                           Q => n_2009, QN => 
                           DataPath_RF_bus_reg_dataout_25_port);
   DataPath_RF_BLOCKi_9_Q_reg_25_inst : DFF_X1 port map( D => n3387, CK => CLK,
                           Q => n_2010, QN => 
                           DataPath_RF_bus_reg_dataout_57_port);
   DataPath_RF_BLOCKi_10_Q_reg_25_inst : DFF_X1 port map( D => n3425, CK => CLK
                           , Q => n_2011, QN => 
                           DataPath_RF_bus_reg_dataout_89_port);
   DataPath_RF_BLOCKi_11_Q_reg_25_inst : DFF_X1 port map( D => n3463, CK => CLK
                           , Q => n_2012, QN => 
                           DataPath_RF_bus_reg_dataout_121_port);
   DataPath_RF_BLOCKi_12_Q_reg_25_inst : DFF_X1 port map( D => n3501, CK => CLK
                           , Q => n_2013, QN => 
                           DataPath_RF_bus_reg_dataout_153_port);
   DataPath_RF_BLOCKi_13_Q_reg_25_inst : DFF_X1 port map( D => n3539, CK => CLK
                           , Q => n_2014, QN => 
                           DataPath_RF_bus_reg_dataout_185_port);
   DataPath_RF_BLOCKi_14_Q_reg_25_inst : DFF_X1 port map( D => n3577, CK => CLK
                           , Q => n_2015, QN => 
                           DataPath_RF_bus_reg_dataout_217_port);
   DataPath_RF_BLOCKi_15_Q_reg_25_inst : DFF_X1 port map( D => n3615, CK => CLK
                           , Q => n_2016, QN => 
                           DataPath_RF_bus_reg_dataout_249_port);
   DataPath_RF_BLOCKi_16_Q_reg_25_inst : DFF_X1 port map( D => n3653, CK => CLK
                           , Q => n_2017, QN => 
                           DataPath_RF_bus_reg_dataout_281_port);
   DataPath_RF_BLOCKi_17_Q_reg_25_inst : DFF_X1 port map( D => n3690, CK => CLK
                           , Q => n_2018, QN => 
                           DataPath_RF_bus_reg_dataout_313_port);
   DataPath_RF_BLOCKi_18_Q_reg_25_inst : DFF_X1 port map( D => n3727, CK => CLK
                           , Q => n_2019, QN => 
                           DataPath_RF_bus_reg_dataout_345_port);
   DataPath_RF_BLOCKi_19_Q_reg_25_inst : DFF_X1 port map( D => n3764, CK => CLK
                           , Q => n_2020, QN => 
                           DataPath_RF_bus_reg_dataout_377_port);
   DataPath_RF_BLOCKi_20_Q_reg_25_inst : DFF_X1 port map( D => n3799, CK => CLK
                           , Q => n_2021, QN => 
                           DataPath_RF_bus_reg_dataout_409_port);
   DataPath_RF_BLOCKi_21_Q_reg_25_inst : DFF_X1 port map( D => n3834, CK => CLK
                           , Q => n_2022, QN => 
                           DataPath_RF_bus_reg_dataout_441_port);
   DataPath_RF_BLOCKi_22_Q_reg_25_inst : DFF_X1 port map( D => n3869, CK => CLK
                           , Q => n_2023, QN => 
                           DataPath_RF_bus_reg_dataout_473_port);
   DataPath_RF_BLOCKi_23_Q_reg_25_inst : DFF_X1 port map( D => n3910, CK => CLK
                           , Q => n_2024, QN => 
                           DataPath_RF_bus_reg_dataout_505_port);
   DataPath_RF_BLOCKi_24_Q_reg_25_inst : DFF_X1 port map( D => n3978, CK => CLK
                           , Q => n_2025, QN => 
                           DataPath_RF_bus_reg_dataout_537_port);
   DataPath_RF_BLOCKi_25_Q_reg_25_inst : DFF_X1 port map( D => n4040, CK => CLK
                           , Q => n_2026, QN => 
                           DataPath_RF_bus_reg_dataout_569_port);
   DataPath_RF_BLOCKi_26_Q_reg_25_inst : DFF_X1 port map( D => n4075, CK => CLK
                           , Q => n_2027, QN => 
                           DataPath_RF_bus_reg_dataout_601_port);
   DataPath_RF_BLOCKi_27_Q_reg_25_inst : DFF_X1 port map( D => n4110, CK => CLK
                           , Q => n_2028, QN => 
                           DataPath_RF_bus_reg_dataout_633_port);
   DataPath_RF_BLOCKi_28_Q_reg_25_inst : DFF_X1 port map( D => n4145, CK => CLK
                           , Q => n_2029, QN => 
                           DataPath_RF_bus_reg_dataout_665_port);
   DataPath_RF_BLOCKi_29_Q_reg_25_inst : DFF_X1 port map( D => n4180, CK => CLK
                           , Q => n_2030, QN => 
                           DataPath_RF_bus_reg_dataout_697_port);
   DataPath_RF_BLOCKi_30_Q_reg_25_inst : DFF_X1 port map( D => n4215, CK => CLK
                           , Q => n_2031, QN => 
                           DataPath_RF_bus_reg_dataout_729_port);
   DataPath_RF_BLOCKi_31_Q_reg_25_inst : DFF_X1 port map( D => n4250, CK => CLK
                           , Q => n_2032, QN => 
                           DataPath_RF_bus_reg_dataout_761_port);
   DataPath_RF_BLOCKi_32_Q_reg_25_inst : DFF_X1 port map( D => n4285, CK => CLK
                           , Q => n_2033, QN => 
                           DataPath_RF_bus_reg_dataout_793_port);
   DataPath_RF_BLOCKi_33_Q_reg_25_inst : DFF_X1 port map( D => n4320, CK => CLK
                           , Q => n_2034, QN => 
                           DataPath_RF_bus_reg_dataout_825_port);
   DataPath_RF_BLOCKi_34_Q_reg_25_inst : DFF_X1 port map( D => n4355, CK => CLK
                           , Q => n_2035, QN => 
                           DataPath_RF_bus_reg_dataout_857_port);
   DataPath_RF_BLOCKi_35_Q_reg_25_inst : DFF_X1 port map( D => n4390, CK => CLK
                           , Q => n_2036, QN => 
                           DataPath_RF_bus_reg_dataout_889_port);
   DataPath_RF_BLOCKi_36_Q_reg_25_inst : DFF_X1 port map( D => n4425, CK => CLK
                           , Q => n_2037, QN => 
                           DataPath_RF_bus_reg_dataout_921_port);
   DataPath_RF_BLOCKi_37_Q_reg_25_inst : DFF_X1 port map( D => n4460, CK => CLK
                           , Q => n_2038, QN => 
                           DataPath_RF_bus_reg_dataout_953_port);
   DataPath_RF_BLOCKi_38_Q_reg_25_inst : DFF_X1 port map( D => n4495, CK => CLK
                           , Q => n_2039, QN => 
                           DataPath_RF_bus_reg_dataout_985_port);
   DataPath_RF_BLOCKi_39_Q_reg_25_inst : DFF_X1 port map( D => n4530, CK => CLK
                           , Q => n_2040, QN => 
                           DataPath_RF_bus_reg_dataout_1017_port);
   DataPath_RF_BLOCKi_40_Q_reg_25_inst : DFF_X1 port map( D => n4571, CK => CLK
                           , Q => n_2041, QN => 
                           DataPath_RF_bus_reg_dataout_1049_port);
   DataPath_RF_BLOCKi_41_Q_reg_25_inst : DFF_X1 port map( D => n4633, CK => CLK
                           , Q => n_2042, QN => 
                           DataPath_RF_bus_reg_dataout_1081_port);
   DataPath_RF_BLOCKi_42_Q_reg_25_inst : DFF_X1 port map( D => n4668, CK => CLK
                           , Q => n_2043, QN => 
                           DataPath_RF_bus_reg_dataout_1113_port);
   DataPath_RF_BLOCKi_43_Q_reg_25_inst : DFF_X1 port map( D => n4703, CK => CLK
                           , Q => n_2044, QN => 
                           DataPath_RF_bus_reg_dataout_1145_port);
   DataPath_RF_BLOCKi_44_Q_reg_25_inst : DFF_X1 port map( D => n4738, CK => CLK
                           , Q => n_2045, QN => 
                           DataPath_RF_bus_reg_dataout_1177_port);
   DataPath_RF_BLOCKi_45_Q_reg_25_inst : DFF_X1 port map( D => n4773, CK => CLK
                           , Q => n_2046, QN => 
                           DataPath_RF_bus_reg_dataout_1209_port);
   DataPath_RF_BLOCKi_46_Q_reg_25_inst : DFF_X1 port map( D => n4808, CK => CLK
                           , Q => n_2047, QN => 
                           DataPath_RF_bus_reg_dataout_1241_port);
   DataPath_RF_BLOCKi_47_Q_reg_25_inst : DFF_X1 port map( D => n4843, CK => CLK
                           , Q => n_2048, QN => 
                           DataPath_RF_bus_reg_dataout_1273_port);
   DataPath_RF_BLOCKi_48_Q_reg_25_inst : DFF_X1 port map( D => n4878, CK => CLK
                           , Q => n_2049, QN => 
                           DataPath_RF_bus_reg_dataout_1305_port);
   DataPath_RF_BLOCKi_49_Q_reg_25_inst : DFF_X1 port map( D => n4913, CK => CLK
                           , Q => n_2050, QN => 
                           DataPath_RF_bus_reg_dataout_1337_port);
   DataPath_RF_BLOCKi_50_Q_reg_25_inst : DFF_X1 port map( D => n4948, CK => CLK
                           , Q => n_2051, QN => 
                           DataPath_RF_bus_reg_dataout_1369_port);
   DataPath_RF_BLOCKi_51_Q_reg_25_inst : DFF_X1 port map( D => n4983, CK => CLK
                           , Q => n_2052, QN => 
                           DataPath_RF_bus_reg_dataout_1401_port);
   DataPath_RF_BLOCKi_52_Q_reg_25_inst : DFF_X1 port map( D => n5018, CK => CLK
                           , Q => n_2053, QN => 
                           DataPath_RF_bus_reg_dataout_1433_port);
   DataPath_RF_BLOCKi_53_Q_reg_25_inst : DFF_X1 port map( D => n5053, CK => CLK
                           , Q => n_2054, QN => 
                           DataPath_RF_bus_reg_dataout_1465_port);
   DataPath_RF_BLOCKi_54_Q_reg_25_inst : DFF_X1 port map( D => n5088, CK => CLK
                           , Q => n_2055, QN => 
                           DataPath_RF_bus_reg_dataout_1497_port);
   DataPath_RF_BLOCKi_55_Q_reg_25_inst : DFF_X1 port map( D => n5123, CK => CLK
                           , Q => n_2056, QN => 
                           DataPath_RF_bus_reg_dataout_1529_port);
   DataPath_RF_BLOCKi_56_Q_reg_25_inst : DFF_X1 port map( D => n5164, CK => CLK
                           , Q => n_2057, QN => 
                           DataPath_RF_bus_reg_dataout_1561_port);
   DataPath_RF_BLOCKi_57_Q_reg_25_inst : DFF_X1 port map( D => n5225, CK => CLK
                           , Q => n_2058, QN => 
                           DataPath_RF_bus_reg_dataout_1593_port);
   DataPath_RF_BLOCKi_58_Q_reg_25_inst : DFF_X1 port map( D => n5261, CK => CLK
                           , Q => n_2059, QN => 
                           DataPath_RF_bus_reg_dataout_1625_port);
   DataPath_RF_BLOCKi_59_Q_reg_25_inst : DFF_X1 port map( D => n5296, CK => CLK
                           , Q => n_2060, QN => 
                           DataPath_RF_bus_reg_dataout_1657_port);
   DataPath_RF_BLOCKi_60_Q_reg_25_inst : DFF_X1 port map( D => n5331, CK => CLK
                           , Q => n_2061, QN => 
                           DataPath_RF_bus_reg_dataout_1689_port);
   DataPath_RF_BLOCKi_61_Q_reg_25_inst : DFF_X1 port map( D => n5366, CK => CLK
                           , Q => n_2062, QN => 
                           DataPath_RF_bus_reg_dataout_1721_port);
   DataPath_RF_BLOCKi_62_Q_reg_25_inst : DFF_X1 port map( D => n5401, CK => CLK
                           , Q => n_2063, QN => 
                           DataPath_RF_bus_reg_dataout_1753_port);
   DataPath_RF_BLOCKi_63_Q_reg_25_inst : DFF_X1 port map( D => n5436, CK => CLK
                           , Q => n_2064, QN => 
                           DataPath_RF_bus_reg_dataout_1785_port);
   DataPath_RF_BLOCKi_64_Q_reg_25_inst : DFF_X1 port map( D => n5471, CK => CLK
                           , Q => n_2065, QN => 
                           DataPath_RF_bus_reg_dataout_1817_port);
   DataPath_RF_BLOCKi_65_Q_reg_25_inst : DFF_X1 port map( D => n5506, CK => CLK
                           , Q => n_2066, QN => 
                           DataPath_RF_bus_reg_dataout_1849_port);
   DataPath_RF_BLOCKi_66_Q_reg_25_inst : DFF_X1 port map( D => n5541, CK => CLK
                           , Q => n_2067, QN => 
                           DataPath_RF_bus_reg_dataout_1881_port);
   DataPath_RF_BLOCKi_67_Q_reg_25_inst : DFF_X1 port map( D => n5576, CK => CLK
                           , Q => n_2068, QN => 
                           DataPath_RF_bus_reg_dataout_1913_port);
   DataPath_RF_BLOCKi_68_Q_reg_25_inst : DFF_X1 port map( D => n5615, CK => CLK
                           , Q => n_2069, QN => 
                           DataPath_RF_bus_reg_dataout_1945_port);
   DataPath_RF_BLOCKi_69_Q_reg_25_inst : DFF_X1 port map( D => n5652, CK => CLK
                           , Q => n_2070, QN => 
                           DataPath_RF_bus_reg_dataout_1977_port);
   DataPath_RF_BLOCKi_70_Q_reg_25_inst : DFF_X1 port map( D => n5689, CK => CLK
                           , Q => n_2071, QN => 
                           DataPath_RF_bus_reg_dataout_2009_port);
   DataPath_RF_BLOCKi_71_Q_reg_25_inst : DFF_X1 port map( D => n5726, CK => CLK
                           , Q => n_2072, QN => 
                           DataPath_RF_bus_reg_dataout_2041_port);
   DataPath_RF_BLOCKi_83_Q_reg_25_inst : DFF_X1 port map( D => n928, CK => CLK,
                           Q => n_2073, QN => 
                           DataPath_RF_bus_reg_dataout_2425_port);
   DataPath_RF_BLOCKi_84_Q_reg_25_inst : DFF_X1 port map( D => n976, CK => CLK,
                           Q => n_2074, QN => 
                           DataPath_RF_bus_reg_dataout_2457_port);
   DataPath_RF_BLOCKi_85_Q_reg_25_inst : DFF_X1 port map( D => n1013, CK => CLK
                           , Q => n_2075, QN => 
                           DataPath_RF_bus_reg_dataout_2489_port);
   DataPath_RF_BLOCKi_86_Q_reg_25_inst : DFF_X1 port map( D => n1050, CK => CLK
                           , Q => n_2076, QN => 
                           DataPath_RF_bus_reg_dataout_2521_port);
   DataPath_RF_BLOCKi_87_Q_reg_25_inst : DFF_X1 port map( D => n1087, CK => CLK
                           , Q => n_2077, QN => 
                           DataPath_RF_bus_reg_dataout_2553_port);
   DataPath_RF_BLOCKi_72_Q_reg_25_inst : DFF_X1 port map( D => n5763, CK => CLK
                           , Q => n_2078, QN => 
                           DataPath_RF_bus_reg_dataout_2073_port);
   DataPath_RF_BLOCKi_73_Q_reg_25_inst : DFF_X1 port map( D => n5802, CK => CLK
                           , Q => n_2079, QN => 
                           DataPath_RF_bus_reg_dataout_2105_port);
   DataPath_RF_BLOCKi_74_Q_reg_25_inst : DFF_X1 port map( D => n5838, CK => CLK
                           , Q => n_2080, QN => 
                           DataPath_RF_bus_reg_dataout_2137_port);
   DataPath_RF_BLOCKi_75_Q_reg_25_inst : DFF_X1 port map( D => n5874, CK => CLK
                           , Q => n_2081, QN => 
                           DataPath_RF_bus_reg_dataout_2169_port);
   DataPath_RF_BLOCKi_76_Q_reg_25_inst : DFF_X1 port map( D => n5910, CK => CLK
                           , Q => n_2082, QN => 
                           DataPath_RF_bus_reg_dataout_2201_port);
   DataPath_RF_BLOCKi_77_Q_reg_25_inst : DFF_X1 port map( D => n5946, CK => CLK
                           , Q => n_2083, QN => 
                           DataPath_RF_bus_reg_dataout_2233_port);
   DataPath_RF_BLOCKi_78_Q_reg_25_inst : DFF_X1 port map( D => n5982, CK => CLK
                           , Q => n_2084, QN => 
                           DataPath_RF_bus_reg_dataout_2265_port);
   DataPath_RF_BLOCKi_79_Q_reg_25_inst : DFF_X1 port map( D => n6018, CK => CLK
                           , Q => n_2085, QN => 
                           DataPath_RF_bus_reg_dataout_2297_port);
   DataPath_RF_BLOCKi_80_Q_reg_25_inst : DFF_X1 port map( D => n6055, CK => CLK
                           , Q => n_2086, QN => 
                           DataPath_RF_bus_reg_dataout_2329_port);
   DataPath_RF_BLOCKi_81_Q_reg_25_inst : DFF_X1 port map( D => n6091, CK => CLK
                           , Q => n_2087, QN => 
                           DataPath_RF_bus_reg_dataout_2361_port);
   DataPath_RF_BLOCKi_82_Q_reg_25_inst : DFF_X1 port map( D => n6125, CK => CLK
                           , Q => n_2088, QN => 
                           DataPath_RF_bus_reg_dataout_2393_port);
   DataPath_REG_ALU_OUT_Q_reg_29_inst : DFF_X1 port map( D => n6994, CK => CLK,
                           Q => DRAM_ADDRESS_29_port, QN => n_2089);
   DataPath_REG_MEM_ALUOUT_Q_reg_29_inst : DFF_X1 port map( D => n1120, CK => 
                           CLK, Q => n_2090, QN => 
                           DataPath_i_REG_MEM_ALUOUT_29_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_29_inst : DFF_X1 port map( D => n6770, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_61_port,
                           QN => n628);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_29_inst : DFF_X1 port map( D => n6802, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_93_port,
                           QN => n660);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_29_inst : DFF_X1 port map( D => n6834, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_125_port
                           , QN => n692);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_29_inst : DFF_X1 port map( D => n6866, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_157_port
                           , QN => n724);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_29_inst : DFF_X1 port map( D => n6898, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_189_port
                           , QN => n756);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_29_inst : DFF_X1 port map( D => n6930, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_221_port
                           , QN => n788);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_29_inst : DFF_X1 port map( D => n6962, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_253_port
                           , QN => n820);
   DataPath_RF_BLOCKi_8_Q_reg_29_inst : DFF_X1 port map( D => n3314, CK => CLK,
                           Q => n_2091, QN => 
                           DataPath_RF_bus_reg_dataout_29_port);
   DataPath_RF_BLOCKi_9_Q_reg_29_inst : DFF_X1 port map( D => n3383, CK => CLK,
                           Q => n_2092, QN => 
                           DataPath_RF_bus_reg_dataout_61_port);
   DataPath_RF_BLOCKi_10_Q_reg_29_inst : DFF_X1 port map( D => n3421, CK => CLK
                           , Q => n_2093, QN => 
                           DataPath_RF_bus_reg_dataout_93_port);
   DataPath_RF_BLOCKi_11_Q_reg_29_inst : DFF_X1 port map( D => n3459, CK => CLK
                           , Q => n_2094, QN => 
                           DataPath_RF_bus_reg_dataout_125_port);
   DataPath_RF_BLOCKi_12_Q_reg_29_inst : DFF_X1 port map( D => n3497, CK => CLK
                           , Q => n_2095, QN => 
                           DataPath_RF_bus_reg_dataout_157_port);
   DataPath_RF_BLOCKi_13_Q_reg_29_inst : DFF_X1 port map( D => n3535, CK => CLK
                           , Q => n_2096, QN => 
                           DataPath_RF_bus_reg_dataout_189_port);
   DataPath_RF_BLOCKi_14_Q_reg_29_inst : DFF_X1 port map( D => n3573, CK => CLK
                           , Q => n_2097, QN => 
                           DataPath_RF_bus_reg_dataout_221_port);
   DataPath_RF_BLOCKi_15_Q_reg_29_inst : DFF_X1 port map( D => n3611, CK => CLK
                           , Q => n_2098, QN => 
                           DataPath_RF_bus_reg_dataout_253_port);
   DataPath_RF_BLOCKi_16_Q_reg_29_inst : DFF_X1 port map( D => n3649, CK => CLK
                           , Q => n_2099, QN => 
                           DataPath_RF_bus_reg_dataout_285_port);
   DataPath_RF_BLOCKi_17_Q_reg_29_inst : DFF_X1 port map( D => n3686, CK => CLK
                           , Q => n_2100, QN => 
                           DataPath_RF_bus_reg_dataout_317_port);
   DataPath_RF_BLOCKi_18_Q_reg_29_inst : DFF_X1 port map( D => n3723, CK => CLK
                           , Q => n_2101, QN => 
                           DataPath_RF_bus_reg_dataout_349_port);
   DataPath_RF_BLOCKi_19_Q_reg_29_inst : DFF_X1 port map( D => n3760, CK => CLK
                           , Q => n_2102, QN => 
                           DataPath_RF_bus_reg_dataout_381_port);
   DataPath_RF_BLOCKi_20_Q_reg_29_inst : DFF_X1 port map( D => n3795, CK => CLK
                           , Q => n_2103, QN => 
                           DataPath_RF_bus_reg_dataout_413_port);
   DataPath_RF_BLOCKi_21_Q_reg_29_inst : DFF_X1 port map( D => n3830, CK => CLK
                           , Q => n_2104, QN => 
                           DataPath_RF_bus_reg_dataout_445_port);
   DataPath_RF_BLOCKi_22_Q_reg_29_inst : DFF_X1 port map( D => n3865, CK => CLK
                           , Q => n_2105, QN => 
                           DataPath_RF_bus_reg_dataout_477_port);
   DataPath_RF_BLOCKi_23_Q_reg_29_inst : DFF_X1 port map( D => n3902, CK => CLK
                           , Q => n_2106, QN => 
                           DataPath_RF_bus_reg_dataout_509_port);
   DataPath_RF_BLOCKi_24_Q_reg_29_inst : DFF_X1 port map( D => n3970, CK => CLK
                           , Q => n_2107, QN => 
                           DataPath_RF_bus_reg_dataout_541_port);
   DataPath_RF_BLOCKi_25_Q_reg_29_inst : DFF_X1 port map( D => n4036, CK => CLK
                           , Q => n_2108, QN => 
                           DataPath_RF_bus_reg_dataout_573_port);
   DataPath_RF_BLOCKi_26_Q_reg_29_inst : DFF_X1 port map( D => n4071, CK => CLK
                           , Q => n_2109, QN => 
                           DataPath_RF_bus_reg_dataout_605_port);
   DataPath_RF_BLOCKi_27_Q_reg_29_inst : DFF_X1 port map( D => n4106, CK => CLK
                           , Q => n_2110, QN => 
                           DataPath_RF_bus_reg_dataout_637_port);
   DataPath_RF_BLOCKi_28_Q_reg_29_inst : DFF_X1 port map( D => n4141, CK => CLK
                           , Q => n_2111, QN => 
                           DataPath_RF_bus_reg_dataout_669_port);
   DataPath_RF_BLOCKi_29_Q_reg_29_inst : DFF_X1 port map( D => n4176, CK => CLK
                           , Q => n_2112, QN => 
                           DataPath_RF_bus_reg_dataout_701_port);
   DataPath_RF_BLOCKi_30_Q_reg_29_inst : DFF_X1 port map( D => n4211, CK => CLK
                           , Q => n_2113, QN => 
                           DataPath_RF_bus_reg_dataout_733_port);
   DataPath_RF_BLOCKi_31_Q_reg_29_inst : DFF_X1 port map( D => n4246, CK => CLK
                           , Q => n_2114, QN => 
                           DataPath_RF_bus_reg_dataout_765_port);
   DataPath_RF_BLOCKi_32_Q_reg_29_inst : DFF_X1 port map( D => n4281, CK => CLK
                           , Q => n_2115, QN => 
                           DataPath_RF_bus_reg_dataout_797_port);
   DataPath_RF_BLOCKi_33_Q_reg_29_inst : DFF_X1 port map( D => n4316, CK => CLK
                           , Q => n_2116, QN => 
                           DataPath_RF_bus_reg_dataout_829_port);
   DataPath_RF_BLOCKi_34_Q_reg_29_inst : DFF_X1 port map( D => n4351, CK => CLK
                           , Q => n_2117, QN => 
                           DataPath_RF_bus_reg_dataout_861_port);
   DataPath_RF_BLOCKi_35_Q_reg_29_inst : DFF_X1 port map( D => n4386, CK => CLK
                           , Q => n_2118, QN => 
                           DataPath_RF_bus_reg_dataout_893_port);
   DataPath_RF_BLOCKi_36_Q_reg_29_inst : DFF_X1 port map( D => n4421, CK => CLK
                           , Q => n_2119, QN => 
                           DataPath_RF_bus_reg_dataout_925_port);
   DataPath_RF_BLOCKi_37_Q_reg_29_inst : DFF_X1 port map( D => n4456, CK => CLK
                           , Q => n_2120, QN => 
                           DataPath_RF_bus_reg_dataout_957_port);
   DataPath_RF_BLOCKi_38_Q_reg_29_inst : DFF_X1 port map( D => n4491, CK => CLK
                           , Q => n_2121, QN => 
                           DataPath_RF_bus_reg_dataout_989_port);
   DataPath_RF_BLOCKi_39_Q_reg_29_inst : DFF_X1 port map( D => n4526, CK => CLK
                           , Q => n_2122, QN => 
                           DataPath_RF_bus_reg_dataout_1021_port);
   DataPath_RF_BLOCKi_40_Q_reg_29_inst : DFF_X1 port map( D => n4563, CK => CLK
                           , Q => n_2123, QN => 
                           DataPath_RF_bus_reg_dataout_1053_port);
   DataPath_RF_BLOCKi_41_Q_reg_29_inst : DFF_X1 port map( D => n4629, CK => CLK
                           , Q => n_2124, QN => 
                           DataPath_RF_bus_reg_dataout_1085_port);
   DataPath_RF_BLOCKi_42_Q_reg_29_inst : DFF_X1 port map( D => n4664, CK => CLK
                           , Q => n_2125, QN => 
                           DataPath_RF_bus_reg_dataout_1117_port);
   DataPath_RF_BLOCKi_43_Q_reg_29_inst : DFF_X1 port map( D => n4699, CK => CLK
                           , Q => n_2126, QN => 
                           DataPath_RF_bus_reg_dataout_1149_port);
   DataPath_RF_BLOCKi_44_Q_reg_29_inst : DFF_X1 port map( D => n4734, CK => CLK
                           , Q => n_2127, QN => 
                           DataPath_RF_bus_reg_dataout_1181_port);
   DataPath_RF_BLOCKi_45_Q_reg_29_inst : DFF_X1 port map( D => n4769, CK => CLK
                           , Q => n_2128, QN => 
                           DataPath_RF_bus_reg_dataout_1213_port);
   DataPath_RF_BLOCKi_46_Q_reg_29_inst : DFF_X1 port map( D => n4804, CK => CLK
                           , Q => n_2129, QN => 
                           DataPath_RF_bus_reg_dataout_1245_port);
   DataPath_RF_BLOCKi_47_Q_reg_29_inst : DFF_X1 port map( D => n4839, CK => CLK
                           , Q => n_2130, QN => 
                           DataPath_RF_bus_reg_dataout_1277_port);
   DataPath_RF_BLOCKi_48_Q_reg_29_inst : DFF_X1 port map( D => n4874, CK => CLK
                           , Q => n_2131, QN => 
                           DataPath_RF_bus_reg_dataout_1309_port);
   DataPath_RF_BLOCKi_49_Q_reg_29_inst : DFF_X1 port map( D => n4909, CK => CLK
                           , Q => n_2132, QN => 
                           DataPath_RF_bus_reg_dataout_1341_port);
   DataPath_RF_BLOCKi_50_Q_reg_29_inst : DFF_X1 port map( D => n4944, CK => CLK
                           , Q => n_2133, QN => 
                           DataPath_RF_bus_reg_dataout_1373_port);
   DataPath_RF_BLOCKi_51_Q_reg_29_inst : DFF_X1 port map( D => n4979, CK => CLK
                           , Q => n_2134, QN => 
                           DataPath_RF_bus_reg_dataout_1405_port);
   DataPath_RF_BLOCKi_52_Q_reg_29_inst : DFF_X1 port map( D => n5014, CK => CLK
                           , Q => n_2135, QN => 
                           DataPath_RF_bus_reg_dataout_1437_port);
   DataPath_RF_BLOCKi_53_Q_reg_29_inst : DFF_X1 port map( D => n5049, CK => CLK
                           , Q => n_2136, QN => 
                           DataPath_RF_bus_reg_dataout_1469_port);
   DataPath_RF_BLOCKi_54_Q_reg_29_inst : DFF_X1 port map( D => n5084, CK => CLK
                           , Q => n_2137, QN => 
                           DataPath_RF_bus_reg_dataout_1501_port);
   DataPath_RF_BLOCKi_55_Q_reg_29_inst : DFF_X1 port map( D => n5119, CK => CLK
                           , Q => n_2138, QN => 
                           DataPath_RF_bus_reg_dataout_1533_port);
   DataPath_RF_BLOCKi_56_Q_reg_29_inst : DFF_X1 port map( D => n5156, CK => CLK
                           , Q => n_2139, QN => 
                           DataPath_RF_bus_reg_dataout_1565_port);
   DataPath_RF_BLOCKi_57_Q_reg_29_inst : DFF_X1 port map( D => n5221, CK => CLK
                           , Q => n_2140, QN => 
                           DataPath_RF_bus_reg_dataout_1597_port);
   DataPath_RF_BLOCKi_58_Q_reg_29_inst : DFF_X1 port map( D => n5257, CK => CLK
                           , Q => n_2141, QN => 
                           DataPath_RF_bus_reg_dataout_1629_port);
   DataPath_RF_BLOCKi_59_Q_reg_29_inst : DFF_X1 port map( D => n5292, CK => CLK
                           , Q => n_2142, QN => 
                           DataPath_RF_bus_reg_dataout_1661_port);
   DataPath_RF_BLOCKi_60_Q_reg_29_inst : DFF_X1 port map( D => n5327, CK => CLK
                           , Q => n_2143, QN => 
                           DataPath_RF_bus_reg_dataout_1693_port);
   DataPath_RF_BLOCKi_61_Q_reg_29_inst : DFF_X1 port map( D => n5362, CK => CLK
                           , Q => n_2144, QN => 
                           DataPath_RF_bus_reg_dataout_1725_port);
   DataPath_RF_BLOCKi_62_Q_reg_29_inst : DFF_X1 port map( D => n5397, CK => CLK
                           , Q => n_2145, QN => 
                           DataPath_RF_bus_reg_dataout_1757_port);
   DataPath_RF_BLOCKi_63_Q_reg_29_inst : DFF_X1 port map( D => n5432, CK => CLK
                           , Q => n_2146, QN => 
                           DataPath_RF_bus_reg_dataout_1789_port);
   DataPath_RF_BLOCKi_64_Q_reg_29_inst : DFF_X1 port map( D => n5467, CK => CLK
                           , Q => n_2147, QN => 
                           DataPath_RF_bus_reg_dataout_1821_port);
   DataPath_RF_BLOCKi_65_Q_reg_29_inst : DFF_X1 port map( D => n5502, CK => CLK
                           , Q => n_2148, QN => 
                           DataPath_RF_bus_reg_dataout_1853_port);
   DataPath_RF_BLOCKi_66_Q_reg_29_inst : DFF_X1 port map( D => n5537, CK => CLK
                           , Q => n_2149, QN => 
                           DataPath_RF_bus_reg_dataout_1885_port);
   DataPath_RF_BLOCKi_67_Q_reg_29_inst : DFF_X1 port map( D => n5572, CK => CLK
                           , Q => n_2150, QN => 
                           DataPath_RF_bus_reg_dataout_1917_port);
   DataPath_RF_BLOCKi_68_Q_reg_29_inst : DFF_X1 port map( D => n5611, CK => CLK
                           , Q => n_2151, QN => 
                           DataPath_RF_bus_reg_dataout_1949_port);
   DataPath_RF_BLOCKi_69_Q_reg_29_inst : DFF_X1 port map( D => n5648, CK => CLK
                           , Q => n_2152, QN => 
                           DataPath_RF_bus_reg_dataout_1981_port);
   DataPath_RF_BLOCKi_70_Q_reg_29_inst : DFF_X1 port map( D => n5685, CK => CLK
                           , Q => n_2153, QN => 
                           DataPath_RF_bus_reg_dataout_2013_port);
   DataPath_RF_BLOCKi_71_Q_reg_29_inst : DFF_X1 port map( D => n5722, CK => CLK
                           , Q => n_2154, QN => 
                           DataPath_RF_bus_reg_dataout_2045_port);
   DataPath_RF_BLOCKi_83_Q_reg_29_inst : DFF_X1 port map( D => n920, CK => CLK,
                           Q => n_2155, QN => 
                           DataPath_RF_bus_reg_dataout_2429_port);
   DataPath_RF_BLOCKi_84_Q_reg_29_inst : DFF_X1 port map( D => n972, CK => CLK,
                           Q => n_2156, QN => 
                           DataPath_RF_bus_reg_dataout_2461_port);
   DataPath_RF_BLOCKi_85_Q_reg_29_inst : DFF_X1 port map( D => n1009, CK => CLK
                           , Q => n_2157, QN => 
                           DataPath_RF_bus_reg_dataout_2493_port);
   DataPath_RF_BLOCKi_86_Q_reg_29_inst : DFF_X1 port map( D => n1046, CK => CLK
                           , Q => n_2158, QN => 
                           DataPath_RF_bus_reg_dataout_2525_port);
   DataPath_RF_BLOCKi_87_Q_reg_29_inst : DFF_X1 port map( D => n1083, CK => CLK
                           , Q => n_2159, QN => 
                           DataPath_RF_bus_reg_dataout_2557_port);
   DataPath_RF_BLOCKi_72_Q_reg_29_inst : DFF_X1 port map( D => n5759, CK => CLK
                           , Q => n_2160, QN => 
                           DataPath_RF_bus_reg_dataout_2077_port);
   DataPath_RF_BLOCKi_73_Q_reg_29_inst : DFF_X1 port map( D => n5798, CK => CLK
                           , Q => n_2161, QN => 
                           DataPath_RF_bus_reg_dataout_2109_port);
   DataPath_RF_BLOCKi_74_Q_reg_29_inst : DFF_X1 port map( D => n5834, CK => CLK
                           , Q => n_2162, QN => 
                           DataPath_RF_bus_reg_dataout_2141_port);
   DataPath_RF_BLOCKi_75_Q_reg_29_inst : DFF_X1 port map( D => n5870, CK => CLK
                           , Q => n_2163, QN => 
                           DataPath_RF_bus_reg_dataout_2173_port);
   DataPath_RF_BLOCKi_76_Q_reg_29_inst : DFF_X1 port map( D => n5906, CK => CLK
                           , Q => n_2164, QN => 
                           DataPath_RF_bus_reg_dataout_2205_port);
   DataPath_RF_BLOCKi_77_Q_reg_29_inst : DFF_X1 port map( D => n5942, CK => CLK
                           , Q => n_2165, QN => 
                           DataPath_RF_bus_reg_dataout_2237_port);
   DataPath_RF_BLOCKi_78_Q_reg_29_inst : DFF_X1 port map( D => n5978, CK => CLK
                           , Q => n_2166, QN => 
                           DataPath_RF_bus_reg_dataout_2269_port);
   DataPath_RF_BLOCKi_79_Q_reg_29_inst : DFF_X1 port map( D => n6014, CK => CLK
                           , Q => n_2167, QN => 
                           DataPath_RF_bus_reg_dataout_2301_port);
   DataPath_RF_BLOCKi_80_Q_reg_29_inst : DFF_X1 port map( D => n6051, CK => CLK
                           , Q => n_2168, QN => 
                           DataPath_RF_bus_reg_dataout_2333_port);
   DataPath_RF_BLOCKi_81_Q_reg_29_inst : DFF_X1 port map( D => n6087, CK => CLK
                           , Q => n_2169, QN => 
                           DataPath_RF_bus_reg_dataout_2365_port);
   DataPath_RF_BLOCKi_82_Q_reg_29_inst : DFF_X1 port map( D => n6121, CK => CLK
                           , Q => n_2170, QN => 
                           DataPath_RF_bus_reg_dataout_2397_port);
   DataPath_REG_ALU_OUT_Q_reg_2_inst : DFF_X1 port map( D => n2151, CK => CLK, 
                           Q => n_2171, QN => DRAM_ADDRESS_2_port);
   DataPath_REG_MEM_ALUOUT_Q_reg_2_inst : DFF_X1 port map( D => n1147, CK => 
                           CLK, Q => n_2172, QN => 
                           DataPath_i_REG_MEM_ALUOUT_2_port);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_2_inst : DFF_X1 port map( D => n6861, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_98_port,
                           QN => n665);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_2_inst : DFF_X1 port map( D => n6893, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_130_port
                           , QN => n697);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_2_inst : DFF_X1 port map( D => n6957, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_194_port
                           , QN => n761);
   DataPath_RF_BLOCKi_8_Q_reg_2_inst : DFF_X1 port map( D => n3368, CK => CLK, 
                           Q => n_2173, QN => 
                           DataPath_RF_bus_reg_dataout_2_port);
   DataPath_RF_BLOCKi_9_Q_reg_2_inst : DFF_X1 port map( D => n3410, CK => CLK, 
                           Q => n_2174, QN => 
                           DataPath_RF_bus_reg_dataout_34_port);
   DataPath_RF_BLOCKi_10_Q_reg_2_inst : DFF_X1 port map( D => n3448, CK => CLK,
                           Q => n_2175, QN => 
                           DataPath_RF_bus_reg_dataout_66_port);
   DataPath_RF_BLOCKi_11_Q_reg_2_inst : DFF_X1 port map( D => n3486, CK => CLK,
                           Q => n_2176, QN => 
                           DataPath_RF_bus_reg_dataout_98_port);
   DataPath_RF_BLOCKi_12_Q_reg_2_inst : DFF_X1 port map( D => n3524, CK => CLK,
                           Q => n_2177, QN => 
                           DataPath_RF_bus_reg_dataout_130_port);
   DataPath_RF_BLOCKi_13_Q_reg_2_inst : DFF_X1 port map( D => n3562, CK => CLK,
                           Q => n_2178, QN => 
                           DataPath_RF_bus_reg_dataout_162_port);
   DataPath_RF_BLOCKi_14_Q_reg_2_inst : DFF_X1 port map( D => n3600, CK => CLK,
                           Q => n_2179, QN => 
                           DataPath_RF_bus_reg_dataout_194_port);
   DataPath_RF_BLOCKi_15_Q_reg_2_inst : DFF_X1 port map( D => n3638, CK => CLK,
                           Q => n_2180, QN => 
                           DataPath_RF_bus_reg_dataout_226_port);
   DataPath_RF_BLOCKi_16_Q_reg_2_inst : DFF_X1 port map( D => n3676, CK => CLK,
                           Q => n_2181, QN => 
                           DataPath_RF_bus_reg_dataout_258_port);
   DataPath_RF_BLOCKi_17_Q_reg_2_inst : DFF_X1 port map( D => n3713, CK => CLK,
                           Q => n_2182, QN => 
                           DataPath_RF_bus_reg_dataout_290_port);
   DataPath_RF_BLOCKi_18_Q_reg_2_inst : DFF_X1 port map( D => n3750, CK => CLK,
                           Q => n_2183, QN => 
                           DataPath_RF_bus_reg_dataout_322_port);
   DataPath_RF_BLOCKi_19_Q_reg_2_inst : DFF_X1 port map( D => n3787, CK => CLK,
                           Q => n_2184, QN => 
                           DataPath_RF_bus_reg_dataout_354_port);
   DataPath_RF_BLOCKi_20_Q_reg_2_inst : DFF_X1 port map( D => n3822, CK => CLK,
                           Q => n_2185, QN => 
                           DataPath_RF_bus_reg_dataout_386_port);
   DataPath_RF_BLOCKi_21_Q_reg_2_inst : DFF_X1 port map( D => n3857, CK => CLK,
                           Q => n_2186, QN => 
                           DataPath_RF_bus_reg_dataout_418_port);
   DataPath_RF_BLOCKi_22_Q_reg_2_inst : DFF_X1 port map( D => n3892, CK => CLK,
                           Q => n_2187, QN => 
                           DataPath_RF_bus_reg_dataout_450_port);
   DataPath_RF_BLOCKi_23_Q_reg_2_inst : DFF_X1 port map( D => n3956, CK => CLK,
                           Q => n_2188, QN => 
                           DataPath_RF_bus_reg_dataout_482_port);
   DataPath_RF_BLOCKi_24_Q_reg_2_inst : DFF_X1 port map( D => n4024, CK => CLK,
                           Q => n_2189, QN => 
                           DataPath_RF_bus_reg_dataout_514_port);
   DataPath_RF_BLOCKi_25_Q_reg_2_inst : DFF_X1 port map( D => n4063, CK => CLK,
                           Q => n_2190, QN => 
                           DataPath_RF_bus_reg_dataout_546_port);
   DataPath_RF_BLOCKi_26_Q_reg_2_inst : DFF_X1 port map( D => n4098, CK => CLK,
                           Q => n_2191, QN => 
                           DataPath_RF_bus_reg_dataout_578_port);
   DataPath_RF_BLOCKi_27_Q_reg_2_inst : DFF_X1 port map( D => n4133, CK => CLK,
                           Q => n_2192, QN => 
                           DataPath_RF_bus_reg_dataout_610_port);
   DataPath_RF_BLOCKi_28_Q_reg_2_inst : DFF_X1 port map( D => n4168, CK => CLK,
                           Q => n_2193, QN => 
                           DataPath_RF_bus_reg_dataout_642_port);
   DataPath_RF_BLOCKi_29_Q_reg_2_inst : DFF_X1 port map( D => n4203, CK => CLK,
                           Q => n_2194, QN => 
                           DataPath_RF_bus_reg_dataout_674_port);
   DataPath_RF_BLOCKi_30_Q_reg_2_inst : DFF_X1 port map( D => n4238, CK => CLK,
                           Q => n_2195, QN => 
                           DataPath_RF_bus_reg_dataout_706_port);
   DataPath_RF_BLOCKi_31_Q_reg_2_inst : DFF_X1 port map( D => n4273, CK => CLK,
                           Q => n_2196, QN => 
                           DataPath_RF_bus_reg_dataout_738_port);
   DataPath_RF_BLOCKi_32_Q_reg_2_inst : DFF_X1 port map( D => n4308, CK => CLK,
                           Q => n_2197, QN => 
                           DataPath_RF_bus_reg_dataout_770_port);
   DataPath_RF_BLOCKi_33_Q_reg_2_inst : DFF_X1 port map( D => n4343, CK => CLK,
                           Q => n_2198, QN => 
                           DataPath_RF_bus_reg_dataout_802_port);
   DataPath_RF_BLOCKi_34_Q_reg_2_inst : DFF_X1 port map( D => n4378, CK => CLK,
                           Q => n_2199, QN => 
                           DataPath_RF_bus_reg_dataout_834_port);
   DataPath_RF_BLOCKi_35_Q_reg_2_inst : DFF_X1 port map( D => n4413, CK => CLK,
                           Q => n_2200, QN => 
                           DataPath_RF_bus_reg_dataout_866_port);
   DataPath_RF_BLOCKi_36_Q_reg_2_inst : DFF_X1 port map( D => n4448, CK => CLK,
                           Q => n_2201, QN => 
                           DataPath_RF_bus_reg_dataout_898_port);
   DataPath_RF_BLOCKi_37_Q_reg_2_inst : DFF_X1 port map( D => n4483, CK => CLK,
                           Q => n_2202, QN => 
                           DataPath_RF_bus_reg_dataout_930_port);
   DataPath_RF_BLOCKi_38_Q_reg_2_inst : DFF_X1 port map( D => n4518, CK => CLK,
                           Q => n_2203, QN => 
                           DataPath_RF_bus_reg_dataout_962_port);
   DataPath_RF_BLOCKi_39_Q_reg_2_inst : DFF_X1 port map( D => n4553, CK => CLK,
                           Q => n_2204, QN => 
                           DataPath_RF_bus_reg_dataout_994_port);
   DataPath_RF_BLOCKi_40_Q_reg_2_inst : DFF_X1 port map( D => n4617, CK => CLK,
                           Q => n_2205, QN => 
                           DataPath_RF_bus_reg_dataout_1026_port);
   DataPath_RF_BLOCKi_41_Q_reg_2_inst : DFF_X1 port map( D => n4656, CK => CLK,
                           Q => n_2206, QN => 
                           DataPath_RF_bus_reg_dataout_1058_port);
   DataPath_RF_BLOCKi_42_Q_reg_2_inst : DFF_X1 port map( D => n4691, CK => CLK,
                           Q => n_2207, QN => 
                           DataPath_RF_bus_reg_dataout_1090_port);
   DataPath_RF_BLOCKi_43_Q_reg_2_inst : DFF_X1 port map( D => n4726, CK => CLK,
                           Q => n_2208, QN => 
                           DataPath_RF_bus_reg_dataout_1122_port);
   DataPath_RF_BLOCKi_44_Q_reg_2_inst : DFF_X1 port map( D => n4761, CK => CLK,
                           Q => n_2209, QN => 
                           DataPath_RF_bus_reg_dataout_1154_port);
   DataPath_RF_BLOCKi_45_Q_reg_2_inst : DFF_X1 port map( D => n4796, CK => CLK,
                           Q => n_2210, QN => 
                           DataPath_RF_bus_reg_dataout_1186_port);
   DataPath_RF_BLOCKi_46_Q_reg_2_inst : DFF_X1 port map( D => n4831, CK => CLK,
                           Q => n_2211, QN => 
                           DataPath_RF_bus_reg_dataout_1218_port);
   DataPath_RF_BLOCKi_47_Q_reg_2_inst : DFF_X1 port map( D => n4866, CK => CLK,
                           Q => n_2212, QN => 
                           DataPath_RF_bus_reg_dataout_1250_port);
   DataPath_RF_BLOCKi_48_Q_reg_2_inst : DFF_X1 port map( D => n4901, CK => CLK,
                           Q => n_2213, QN => 
                           DataPath_RF_bus_reg_dataout_1282_port);
   DataPath_RF_BLOCKi_49_Q_reg_2_inst : DFF_X1 port map( D => n4936, CK => CLK,
                           Q => n_2214, QN => 
                           DataPath_RF_bus_reg_dataout_1314_port);
   DataPath_RF_BLOCKi_50_Q_reg_2_inst : DFF_X1 port map( D => n4971, CK => CLK,
                           Q => n_2215, QN => 
                           DataPath_RF_bus_reg_dataout_1346_port);
   DataPath_RF_BLOCKi_51_Q_reg_2_inst : DFF_X1 port map( D => n5006, CK => CLK,
                           Q => n_2216, QN => 
                           DataPath_RF_bus_reg_dataout_1378_port);
   DataPath_RF_BLOCKi_52_Q_reg_2_inst : DFF_X1 port map( D => n5041, CK => CLK,
                           Q => n_2217, QN => 
                           DataPath_RF_bus_reg_dataout_1410_port);
   DataPath_RF_BLOCKi_53_Q_reg_2_inst : DFF_X1 port map( D => n5076, CK => CLK,
                           Q => n_2218, QN => 
                           DataPath_RF_bus_reg_dataout_1442_port);
   DataPath_RF_BLOCKi_54_Q_reg_2_inst : DFF_X1 port map( D => n5111, CK => CLK,
                           Q => n_2219, QN => 
                           DataPath_RF_bus_reg_dataout_1474_port);
   DataPath_RF_BLOCKi_55_Q_reg_2_inst : DFF_X1 port map( D => n5146, CK => CLK,
                           Q => n_2220, QN => 
                           DataPath_RF_bus_reg_dataout_1506_port);
   DataPath_RF_BLOCKi_56_Q_reg_2_inst : DFF_X1 port map( D => n5210, CK => CLK,
                           Q => n_2221, QN => 
                           DataPath_RF_bus_reg_dataout_1538_port);
   DataPath_RF_BLOCKi_57_Q_reg_2_inst : DFF_X1 port map( D => n5248, CK => CLK,
                           Q => n_2222, QN => 
                           DataPath_RF_bus_reg_dataout_1570_port);
   DataPath_RF_BLOCKi_58_Q_reg_2_inst : DFF_X1 port map( D => n5284, CK => CLK,
                           Q => n_2223, QN => 
                           DataPath_RF_bus_reg_dataout_1602_port);
   DataPath_RF_BLOCKi_59_Q_reg_2_inst : DFF_X1 port map( D => n5319, CK => CLK,
                           Q => n_2224, QN => 
                           DataPath_RF_bus_reg_dataout_1634_port);
   DataPath_RF_BLOCKi_60_Q_reg_2_inst : DFF_X1 port map( D => n5354, CK => CLK,
                           Q => n_2225, QN => 
                           DataPath_RF_bus_reg_dataout_1666_port);
   DataPath_RF_BLOCKi_61_Q_reg_2_inst : DFF_X1 port map( D => n5389, CK => CLK,
                           Q => n_2226, QN => 
                           DataPath_RF_bus_reg_dataout_1698_port);
   DataPath_RF_BLOCKi_62_Q_reg_2_inst : DFF_X1 port map( D => n5424, CK => CLK,
                           Q => n_2227, QN => 
                           DataPath_RF_bus_reg_dataout_1730_port);
   DataPath_RF_BLOCKi_63_Q_reg_2_inst : DFF_X1 port map( D => n5459, CK => CLK,
                           Q => n_2228, QN => 
                           DataPath_RF_bus_reg_dataout_1762_port);
   DataPath_RF_BLOCKi_64_Q_reg_2_inst : DFF_X1 port map( D => n5494, CK => CLK,
                           Q => n_2229, QN => 
                           DataPath_RF_bus_reg_dataout_1794_port);
   DataPath_RF_BLOCKi_65_Q_reg_2_inst : DFF_X1 port map( D => n5529, CK => CLK,
                           Q => n_2230, QN => 
                           DataPath_RF_bus_reg_dataout_1826_port);
   DataPath_RF_BLOCKi_66_Q_reg_2_inst : DFF_X1 port map( D => n5564, CK => CLK,
                           Q => n_2231, QN => 
                           DataPath_RF_bus_reg_dataout_1858_port);
   DataPath_RF_BLOCKi_67_Q_reg_2_inst : DFF_X1 port map( D => n5599, CK => CLK,
                           Q => n_2232, QN => 
                           DataPath_RF_bus_reg_dataout_1890_port);
   DataPath_RF_BLOCKi_68_Q_reg_2_inst : DFF_X1 port map( D => n5638, CK => CLK,
                           Q => n_2233, QN => 
                           DataPath_RF_bus_reg_dataout_1922_port);
   DataPath_RF_BLOCKi_69_Q_reg_2_inst : DFF_X1 port map( D => n5675, CK => CLK,
                           Q => n_2234, QN => 
                           DataPath_RF_bus_reg_dataout_1954_port);
   DataPath_RF_BLOCKi_70_Q_reg_2_inst : DFF_X1 port map( D => n5712, CK => CLK,
                           Q => n_2235, QN => 
                           DataPath_RF_bus_reg_dataout_1986_port);
   DataPath_RF_BLOCKi_71_Q_reg_2_inst : DFF_X1 port map( D => n5749, CK => CLK,
                           Q => n_2236, QN => 
                           DataPath_RF_bus_reg_dataout_2018_port);
   DataPath_RF_BLOCKi_82_Q_reg_2_inst : DFF_X1 port map( D => n908, CK => CLK, 
                           Q => n_2237, QN => 
                           DataPath_RF_bus_reg_dataout_2370_port);
   DataPath_RF_BLOCKi_83_Q_reg_2_inst : DFF_X1 port map( D => n961, CK => CLK, 
                           Q => n_2238, QN => 
                           DataPath_RF_bus_reg_dataout_2402_port);
   DataPath_RF_BLOCKi_84_Q_reg_2_inst : DFF_X1 port map( D => n999, CK => CLK, 
                           Q => n_2239, QN => 
                           DataPath_RF_bus_reg_dataout_2434_port);
   DataPath_RF_BLOCKi_85_Q_reg_2_inst : DFF_X1 port map( D => n1036, CK => CLK,
                           Q => n_2240, QN => 
                           DataPath_RF_bus_reg_dataout_2466_port);
   DataPath_RF_BLOCKi_86_Q_reg_2_inst : DFF_X1 port map( D => n1073, CK => CLK,
                           Q => n_2241, QN => 
                           DataPath_RF_bus_reg_dataout_2498_port);
   DataPath_RF_BLOCKi_87_Q_reg_2_inst : DFF_X1 port map( D => n1110, CK => CLK,
                           Q => n_2242, QN => 
                           DataPath_RF_bus_reg_dataout_2530_port);
   DataPath_RF_BLOCKi_72_Q_reg_2_inst : DFF_X1 port map( D => n5786, CK => CLK,
                           Q => n_2243, QN => 
                           DataPath_RF_bus_reg_dataout_2050_port);
   DataPath_RF_BLOCKi_73_Q_reg_2_inst : DFF_X1 port map( D => n5825, CK => CLK,
                           Q => n_2244, QN => 
                           DataPath_RF_bus_reg_dataout_2082_port);
   DataPath_RF_BLOCKi_74_Q_reg_2_inst : DFF_X1 port map( D => n5861, CK => CLK,
                           Q => n_2245, QN => 
                           DataPath_RF_bus_reg_dataout_2114_port);
   DataPath_RF_BLOCKi_75_Q_reg_2_inst : DFF_X1 port map( D => n5897, CK => CLK,
                           Q => n_2246, QN => 
                           DataPath_RF_bus_reg_dataout_2146_port);
   DataPath_RF_BLOCKi_76_Q_reg_2_inst : DFF_X1 port map( D => n5933, CK => CLK,
                           Q => n_2247, QN => 
                           DataPath_RF_bus_reg_dataout_2178_port);
   DataPath_RF_BLOCKi_77_Q_reg_2_inst : DFF_X1 port map( D => n5969, CK => CLK,
                           Q => n_2248, QN => 
                           DataPath_RF_bus_reg_dataout_2210_port);
   DataPath_RF_BLOCKi_78_Q_reg_2_inst : DFF_X1 port map( D => n6005, CK => CLK,
                           Q => n_2249, QN => 
                           DataPath_RF_bus_reg_dataout_2242_port);
   DataPath_RF_BLOCKi_79_Q_reg_2_inst : DFF_X1 port map( D => n6041, CK => CLK,
                           Q => n_2250, QN => 
                           DataPath_RF_bus_reg_dataout_2274_port);
   DataPath_RF_BLOCKi_80_Q_reg_2_inst : DFF_X1 port map( D => n6078, CK => CLK,
                           Q => n_2251, QN => 
                           DataPath_RF_bus_reg_dataout_2306_port);
   DataPath_RF_BLOCKi_81_Q_reg_2_inst : DFF_X1 port map( D => n6114, CK => CLK,
                           Q => n_2252, QN => 
                           DataPath_RF_bus_reg_dataout_2338_port);
   DataPath_REG_ALU_OUT_Q_reg_3_inst : DFF_X1 port map( D => n2119, CK => CLK, 
                           Q => n_2253, QN => DRAM_ADDRESS_3_port);
   DataPath_REG_MEM_ALUOUT_Q_reg_3_inst : DFF_X1 port map( D => n1146, CK => 
                           CLK, Q => n_2254, QN => 
                           DataPath_i_REG_MEM_ALUOUT_3_port);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_3_inst : DFF_X1 port map( D => n6860, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_99_port,
                           QN => n666);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_3_inst : DFF_X1 port map( D => n6892, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_131_port
                           , QN => n698);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_3_inst : DFF_X1 port map( D => n6956, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_195_port
                           , QN => n762);
   DataPath_RF_BLOCKi_8_Q_reg_3_inst : DFF_X1 port map( D => n3366, CK => CLK, 
                           Q => n_2255, QN => 
                           DataPath_RF_bus_reg_dataout_3_port);
   DataPath_RF_BLOCKi_9_Q_reg_3_inst : DFF_X1 port map( D => n3409, CK => CLK, 
                           Q => n_2256, QN => 
                           DataPath_RF_bus_reg_dataout_35_port);
   DataPath_RF_BLOCKi_10_Q_reg_3_inst : DFF_X1 port map( D => n3447, CK => CLK,
                           Q => n_2257, QN => 
                           DataPath_RF_bus_reg_dataout_67_port);
   DataPath_RF_BLOCKi_11_Q_reg_3_inst : DFF_X1 port map( D => n3485, CK => CLK,
                           Q => n_2258, QN => 
                           DataPath_RF_bus_reg_dataout_99_port);
   DataPath_RF_BLOCKi_12_Q_reg_3_inst : DFF_X1 port map( D => n3523, CK => CLK,
                           Q => n_2259, QN => 
                           DataPath_RF_bus_reg_dataout_131_port);
   DataPath_RF_BLOCKi_13_Q_reg_3_inst : DFF_X1 port map( D => n3561, CK => CLK,
                           Q => n_2260, QN => 
                           DataPath_RF_bus_reg_dataout_163_port);
   DataPath_RF_BLOCKi_14_Q_reg_3_inst : DFF_X1 port map( D => n3599, CK => CLK,
                           Q => n_2261, QN => 
                           DataPath_RF_bus_reg_dataout_195_port);
   DataPath_RF_BLOCKi_15_Q_reg_3_inst : DFF_X1 port map( D => n3637, CK => CLK,
                           Q => n_2262, QN => 
                           DataPath_RF_bus_reg_dataout_227_port);
   DataPath_RF_BLOCKi_16_Q_reg_3_inst : DFF_X1 port map( D => n3675, CK => CLK,
                           Q => n_2263, QN => 
                           DataPath_RF_bus_reg_dataout_259_port);
   DataPath_RF_BLOCKi_17_Q_reg_3_inst : DFF_X1 port map( D => n3712, CK => CLK,
                           Q => n_2264, QN => 
                           DataPath_RF_bus_reg_dataout_291_port);
   DataPath_RF_BLOCKi_18_Q_reg_3_inst : DFF_X1 port map( D => n3749, CK => CLK,
                           Q => n_2265, QN => 
                           DataPath_RF_bus_reg_dataout_323_port);
   DataPath_RF_BLOCKi_19_Q_reg_3_inst : DFF_X1 port map( D => n3786, CK => CLK,
                           Q => n_2266, QN => 
                           DataPath_RF_bus_reg_dataout_355_port);
   DataPath_RF_BLOCKi_20_Q_reg_3_inst : DFF_X1 port map( D => n3821, CK => CLK,
                           Q => n_2267, QN => 
                           DataPath_RF_bus_reg_dataout_387_port);
   DataPath_RF_BLOCKi_21_Q_reg_3_inst : DFF_X1 port map( D => n3856, CK => CLK,
                           Q => n_2268, QN => 
                           DataPath_RF_bus_reg_dataout_419_port);
   DataPath_RF_BLOCKi_22_Q_reg_3_inst : DFF_X1 port map( D => n3891, CK => CLK,
                           Q => n_2269, QN => 
                           DataPath_RF_bus_reg_dataout_451_port);
   DataPath_RF_BLOCKi_23_Q_reg_3_inst : DFF_X1 port map( D => n3954, CK => CLK,
                           Q => n_2270, QN => 
                           DataPath_RF_bus_reg_dataout_483_port);
   DataPath_RF_BLOCKi_24_Q_reg_3_inst : DFF_X1 port map( D => n4022, CK => CLK,
                           Q => n_2271, QN => 
                           DataPath_RF_bus_reg_dataout_515_port);
   DataPath_RF_BLOCKi_25_Q_reg_3_inst : DFF_X1 port map( D => n4062, CK => CLK,
                           Q => n_2272, QN => 
                           DataPath_RF_bus_reg_dataout_547_port);
   DataPath_RF_BLOCKi_26_Q_reg_3_inst : DFF_X1 port map( D => n4097, CK => CLK,
                           Q => n_2273, QN => 
                           DataPath_RF_bus_reg_dataout_579_port);
   DataPath_RF_BLOCKi_27_Q_reg_3_inst : DFF_X1 port map( D => n4132, CK => CLK,
                           Q => n_2274, QN => 
                           DataPath_RF_bus_reg_dataout_611_port);
   DataPath_RF_BLOCKi_28_Q_reg_3_inst : DFF_X1 port map( D => n4167, CK => CLK,
                           Q => n_2275, QN => 
                           DataPath_RF_bus_reg_dataout_643_port);
   DataPath_RF_BLOCKi_29_Q_reg_3_inst : DFF_X1 port map( D => n4202, CK => CLK,
                           Q => n_2276, QN => 
                           DataPath_RF_bus_reg_dataout_675_port);
   DataPath_RF_BLOCKi_30_Q_reg_3_inst : DFF_X1 port map( D => n4237, CK => CLK,
                           Q => n_2277, QN => 
                           DataPath_RF_bus_reg_dataout_707_port);
   DataPath_RF_BLOCKi_31_Q_reg_3_inst : DFF_X1 port map( D => n4272, CK => CLK,
                           Q => n_2278, QN => 
                           DataPath_RF_bus_reg_dataout_739_port);
   DataPath_RF_BLOCKi_32_Q_reg_3_inst : DFF_X1 port map( D => n4307, CK => CLK,
                           Q => n_2279, QN => 
                           DataPath_RF_bus_reg_dataout_771_port);
   DataPath_RF_BLOCKi_33_Q_reg_3_inst : DFF_X1 port map( D => n4342, CK => CLK,
                           Q => n_2280, QN => 
                           DataPath_RF_bus_reg_dataout_803_port);
   DataPath_RF_BLOCKi_34_Q_reg_3_inst : DFF_X1 port map( D => n4377, CK => CLK,
                           Q => n_2281, QN => 
                           DataPath_RF_bus_reg_dataout_835_port);
   DataPath_RF_BLOCKi_35_Q_reg_3_inst : DFF_X1 port map( D => n4412, CK => CLK,
                           Q => n_2282, QN => 
                           DataPath_RF_bus_reg_dataout_867_port);
   DataPath_RF_BLOCKi_36_Q_reg_3_inst : DFF_X1 port map( D => n4447, CK => CLK,
                           Q => n_2283, QN => 
                           DataPath_RF_bus_reg_dataout_899_port);
   DataPath_RF_BLOCKi_37_Q_reg_3_inst : DFF_X1 port map( D => n4482, CK => CLK,
                           Q => n_2284, QN => 
                           DataPath_RF_bus_reg_dataout_931_port);
   DataPath_RF_BLOCKi_38_Q_reg_3_inst : DFF_X1 port map( D => n4517, CK => CLK,
                           Q => n_2285, QN => 
                           DataPath_RF_bus_reg_dataout_963_port);
   DataPath_RF_BLOCKi_39_Q_reg_3_inst : DFF_X1 port map( D => n4552, CK => CLK,
                           Q => n_2286, QN => 
                           DataPath_RF_bus_reg_dataout_995_port);
   DataPath_RF_BLOCKi_40_Q_reg_3_inst : DFF_X1 port map( D => n4615, CK => CLK,
                           Q => n_2287, QN => 
                           DataPath_RF_bus_reg_dataout_1027_port);
   DataPath_RF_BLOCKi_41_Q_reg_3_inst : DFF_X1 port map( D => n4655, CK => CLK,
                           Q => n_2288, QN => 
                           DataPath_RF_bus_reg_dataout_1059_port);
   DataPath_RF_BLOCKi_42_Q_reg_3_inst : DFF_X1 port map( D => n4690, CK => CLK,
                           Q => n_2289, QN => 
                           DataPath_RF_bus_reg_dataout_1091_port);
   DataPath_RF_BLOCKi_43_Q_reg_3_inst : DFF_X1 port map( D => n4725, CK => CLK,
                           Q => n_2290, QN => 
                           DataPath_RF_bus_reg_dataout_1123_port);
   DataPath_RF_BLOCKi_44_Q_reg_3_inst : DFF_X1 port map( D => n4760, CK => CLK,
                           Q => n_2291, QN => 
                           DataPath_RF_bus_reg_dataout_1155_port);
   DataPath_RF_BLOCKi_45_Q_reg_3_inst : DFF_X1 port map( D => n4795, CK => CLK,
                           Q => n_2292, QN => 
                           DataPath_RF_bus_reg_dataout_1187_port);
   DataPath_RF_BLOCKi_46_Q_reg_3_inst : DFF_X1 port map( D => n4830, CK => CLK,
                           Q => n_2293, QN => 
                           DataPath_RF_bus_reg_dataout_1219_port);
   DataPath_RF_BLOCKi_47_Q_reg_3_inst : DFF_X1 port map( D => n4865, CK => CLK,
                           Q => n_2294, QN => 
                           DataPath_RF_bus_reg_dataout_1251_port);
   DataPath_RF_BLOCKi_48_Q_reg_3_inst : DFF_X1 port map( D => n4900, CK => CLK,
                           Q => n_2295, QN => 
                           DataPath_RF_bus_reg_dataout_1283_port);
   DataPath_RF_BLOCKi_49_Q_reg_3_inst : DFF_X1 port map( D => n4935, CK => CLK,
                           Q => n_2296, QN => 
                           DataPath_RF_bus_reg_dataout_1315_port);
   DataPath_RF_BLOCKi_50_Q_reg_3_inst : DFF_X1 port map( D => n4970, CK => CLK,
                           Q => n_2297, QN => 
                           DataPath_RF_bus_reg_dataout_1347_port);
   DataPath_RF_BLOCKi_51_Q_reg_3_inst : DFF_X1 port map( D => n5005, CK => CLK,
                           Q => n_2298, QN => 
                           DataPath_RF_bus_reg_dataout_1379_port);
   DataPath_RF_BLOCKi_52_Q_reg_3_inst : DFF_X1 port map( D => n5040, CK => CLK,
                           Q => n_2299, QN => 
                           DataPath_RF_bus_reg_dataout_1411_port);
   DataPath_RF_BLOCKi_53_Q_reg_3_inst : DFF_X1 port map( D => n5075, CK => CLK,
                           Q => n_2300, QN => 
                           DataPath_RF_bus_reg_dataout_1443_port);
   DataPath_RF_BLOCKi_54_Q_reg_3_inst : DFF_X1 port map( D => n5110, CK => CLK,
                           Q => n_2301, QN => 
                           DataPath_RF_bus_reg_dataout_1475_port);
   DataPath_RF_BLOCKi_55_Q_reg_3_inst : DFF_X1 port map( D => n5145, CK => CLK,
                           Q => n_2302, QN => 
                           DataPath_RF_bus_reg_dataout_1507_port);
   DataPath_RF_BLOCKi_56_Q_reg_3_inst : DFF_X1 port map( D => n5208, CK => CLK,
                           Q => n_2303, QN => 
                           DataPath_RF_bus_reg_dataout_1539_port);
   DataPath_RF_BLOCKi_57_Q_reg_3_inst : DFF_X1 port map( D => n5247, CK => CLK,
                           Q => n_2304, QN => 
                           DataPath_RF_bus_reg_dataout_1571_port);
   DataPath_RF_BLOCKi_58_Q_reg_3_inst : DFF_X1 port map( D => n5283, CK => CLK,
                           Q => n_2305, QN => 
                           DataPath_RF_bus_reg_dataout_1603_port);
   DataPath_RF_BLOCKi_59_Q_reg_3_inst : DFF_X1 port map( D => n5318, CK => CLK,
                           Q => n_2306, QN => 
                           DataPath_RF_bus_reg_dataout_1635_port);
   DataPath_RF_BLOCKi_60_Q_reg_3_inst : DFF_X1 port map( D => n5353, CK => CLK,
                           Q => n_2307, QN => 
                           DataPath_RF_bus_reg_dataout_1667_port);
   DataPath_RF_BLOCKi_61_Q_reg_3_inst : DFF_X1 port map( D => n5388, CK => CLK,
                           Q => n_2308, QN => 
                           DataPath_RF_bus_reg_dataout_1699_port);
   DataPath_RF_BLOCKi_62_Q_reg_3_inst : DFF_X1 port map( D => n5423, CK => CLK,
                           Q => n_2309, QN => 
                           DataPath_RF_bus_reg_dataout_1731_port);
   DataPath_RF_BLOCKi_63_Q_reg_3_inst : DFF_X1 port map( D => n5458, CK => CLK,
                           Q => n_2310, QN => 
                           DataPath_RF_bus_reg_dataout_1763_port);
   DataPath_RF_BLOCKi_64_Q_reg_3_inst : DFF_X1 port map( D => n5493, CK => CLK,
                           Q => n_2311, QN => 
                           DataPath_RF_bus_reg_dataout_1795_port);
   DataPath_RF_BLOCKi_65_Q_reg_3_inst : DFF_X1 port map( D => n5528, CK => CLK,
                           Q => n_2312, QN => 
                           DataPath_RF_bus_reg_dataout_1827_port);
   DataPath_RF_BLOCKi_66_Q_reg_3_inst : DFF_X1 port map( D => n5563, CK => CLK,
                           Q => n_2313, QN => 
                           DataPath_RF_bus_reg_dataout_1859_port);
   DataPath_RF_BLOCKi_67_Q_reg_3_inst : DFF_X1 port map( D => n5598, CK => CLK,
                           Q => n_2314, QN => 
                           DataPath_RF_bus_reg_dataout_1891_port);
   DataPath_RF_BLOCKi_68_Q_reg_3_inst : DFF_X1 port map( D => n5637, CK => CLK,
                           Q => n_2315, QN => 
                           DataPath_RF_bus_reg_dataout_1923_port);
   DataPath_RF_BLOCKi_69_Q_reg_3_inst : DFF_X1 port map( D => n5674, CK => CLK,
                           Q => n_2316, QN => 
                           DataPath_RF_bus_reg_dataout_1955_port);
   DataPath_RF_BLOCKi_70_Q_reg_3_inst : DFF_X1 port map( D => n5711, CK => CLK,
                           Q => n_2317, QN => 
                           DataPath_RF_bus_reg_dataout_1987_port);
   DataPath_RF_BLOCKi_71_Q_reg_3_inst : DFF_X1 port map( D => n5748, CK => CLK,
                           Q => n_2318, QN => 
                           DataPath_RF_bus_reg_dataout_2019_port);
   DataPath_RF_BLOCKi_82_Q_reg_3_inst : DFF_X1 port map( D => n906, CK => CLK, 
                           Q => n_2319, QN => 
                           DataPath_RF_bus_reg_dataout_2371_port);
   DataPath_RF_BLOCKi_83_Q_reg_3_inst : DFF_X1 port map( D => n960, CK => CLK, 
                           Q => n_2320, QN => 
                           DataPath_RF_bus_reg_dataout_2403_port);
   DataPath_RF_BLOCKi_84_Q_reg_3_inst : DFF_X1 port map( D => n998, CK => CLK, 
                           Q => n_2321, QN => 
                           DataPath_RF_bus_reg_dataout_2435_port);
   DataPath_RF_BLOCKi_85_Q_reg_3_inst : DFF_X1 port map( D => n1035, CK => CLK,
                           Q => n_2322, QN => 
                           DataPath_RF_bus_reg_dataout_2467_port);
   DataPath_RF_BLOCKi_86_Q_reg_3_inst : DFF_X1 port map( D => n1072, CK => CLK,
                           Q => n_2323, QN => 
                           DataPath_RF_bus_reg_dataout_2499_port);
   DataPath_RF_BLOCKi_87_Q_reg_3_inst : DFF_X1 port map( D => n1109, CK => CLK,
                           Q => n_2324, QN => 
                           DataPath_RF_bus_reg_dataout_2531_port);
   DataPath_RF_BLOCKi_72_Q_reg_3_inst : DFF_X1 port map( D => n5785, CK => CLK,
                           Q => n_2325, QN => 
                           DataPath_RF_bus_reg_dataout_2051_port);
   DataPath_RF_BLOCKi_73_Q_reg_3_inst : DFF_X1 port map( D => n5824, CK => CLK,
                           Q => n_2326, QN => 
                           DataPath_RF_bus_reg_dataout_2083_port);
   DataPath_RF_BLOCKi_74_Q_reg_3_inst : DFF_X1 port map( D => n5860, CK => CLK,
                           Q => n_2327, QN => 
                           DataPath_RF_bus_reg_dataout_2115_port);
   DataPath_RF_BLOCKi_75_Q_reg_3_inst : DFF_X1 port map( D => n5896, CK => CLK,
                           Q => n_2328, QN => 
                           DataPath_RF_bus_reg_dataout_2147_port);
   DataPath_RF_BLOCKi_76_Q_reg_3_inst : DFF_X1 port map( D => n5932, CK => CLK,
                           Q => n_2329, QN => 
                           DataPath_RF_bus_reg_dataout_2179_port);
   DataPath_RF_BLOCKi_77_Q_reg_3_inst : DFF_X1 port map( D => n5968, CK => CLK,
                           Q => n_2330, QN => 
                           DataPath_RF_bus_reg_dataout_2211_port);
   DataPath_RF_BLOCKi_78_Q_reg_3_inst : DFF_X1 port map( D => n6004, CK => CLK,
                           Q => n_2331, QN => 
                           DataPath_RF_bus_reg_dataout_2243_port);
   DataPath_RF_BLOCKi_79_Q_reg_3_inst : DFF_X1 port map( D => n6040, CK => CLK,
                           Q => n_2332, QN => 
                           DataPath_RF_bus_reg_dataout_2275_port);
   DataPath_RF_BLOCKi_80_Q_reg_3_inst : DFF_X1 port map( D => n6077, CK => CLK,
                           Q => n_2333, QN => 
                           DataPath_RF_bus_reg_dataout_2307_port);
   DataPath_RF_BLOCKi_81_Q_reg_3_inst : DFF_X1 port map( D => n6113, CK => CLK,
                           Q => n_2334, QN => 
                           DataPath_RF_bus_reg_dataout_2339_port);
   DataPath_REG_ALU_OUT_Q_reg_4_inst : DFF_X1 port map( D => n7018, CK => CLK, 
                           Q => DRAM_ADDRESS_4_port, QN => n496);
   DataPath_REG_MEM_ALUOUT_Q_reg_4_inst : DFF_X1 port map( D => n1145, CK => 
                           CLK, Q => n_2335, QN => 
                           DataPath_i_REG_MEM_ALUOUT_4_port);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_4_inst : DFF_X1 port map( D => n6859, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_100_port
                           , QN => n667);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_4_inst : DFF_X1 port map( D => n6891, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_132_port
                           , QN => n699);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_4_inst : DFF_X1 port map( D => n6955, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_196_port
                           , QN => n763);
   DataPath_RF_BLOCKi_8_Q_reg_4_inst : DFF_X1 port map( D => n3364, CK => CLK, 
                           Q => n_2336, QN => 
                           DataPath_RF_bus_reg_dataout_4_port);
   DataPath_RF_BLOCKi_9_Q_reg_4_inst : DFF_X1 port map( D => n3408, CK => CLK, 
                           Q => n_2337, QN => 
                           DataPath_RF_bus_reg_dataout_36_port);
   DataPath_RF_BLOCKi_10_Q_reg_4_inst : DFF_X1 port map( D => n3446, CK => CLK,
                           Q => n_2338, QN => 
                           DataPath_RF_bus_reg_dataout_68_port);
   DataPath_RF_BLOCKi_11_Q_reg_4_inst : DFF_X1 port map( D => n3484, CK => CLK,
                           Q => n_2339, QN => 
                           DataPath_RF_bus_reg_dataout_100_port);
   DataPath_RF_BLOCKi_12_Q_reg_4_inst : DFF_X1 port map( D => n3522, CK => CLK,
                           Q => n_2340, QN => 
                           DataPath_RF_bus_reg_dataout_132_port);
   DataPath_RF_BLOCKi_13_Q_reg_4_inst : DFF_X1 port map( D => n3560, CK => CLK,
                           Q => n_2341, QN => 
                           DataPath_RF_bus_reg_dataout_164_port);
   DataPath_RF_BLOCKi_14_Q_reg_4_inst : DFF_X1 port map( D => n3598, CK => CLK,
                           Q => n_2342, QN => 
                           DataPath_RF_bus_reg_dataout_196_port);
   DataPath_RF_BLOCKi_15_Q_reg_4_inst : DFF_X1 port map( D => n3636, CK => CLK,
                           Q => n_2343, QN => 
                           DataPath_RF_bus_reg_dataout_228_port);
   DataPath_RF_BLOCKi_16_Q_reg_4_inst : DFF_X1 port map( D => n3674, CK => CLK,
                           Q => n_2344, QN => 
                           DataPath_RF_bus_reg_dataout_260_port);
   DataPath_RF_BLOCKi_17_Q_reg_4_inst : DFF_X1 port map( D => n3711, CK => CLK,
                           Q => n_2345, QN => 
                           DataPath_RF_bus_reg_dataout_292_port);
   DataPath_RF_BLOCKi_18_Q_reg_4_inst : DFF_X1 port map( D => n3748, CK => CLK,
                           Q => n_2346, QN => 
                           DataPath_RF_bus_reg_dataout_324_port);
   DataPath_RF_BLOCKi_19_Q_reg_4_inst : DFF_X1 port map( D => n3785, CK => CLK,
                           Q => n_2347, QN => 
                           DataPath_RF_bus_reg_dataout_356_port);
   DataPath_RF_BLOCKi_20_Q_reg_4_inst : DFF_X1 port map( D => n3820, CK => CLK,
                           Q => n_2348, QN => 
                           DataPath_RF_bus_reg_dataout_388_port);
   DataPath_RF_BLOCKi_21_Q_reg_4_inst : DFF_X1 port map( D => n3855, CK => CLK,
                           Q => n_2349, QN => 
                           DataPath_RF_bus_reg_dataout_420_port);
   DataPath_RF_BLOCKi_22_Q_reg_4_inst : DFF_X1 port map( D => n3890, CK => CLK,
                           Q => n_2350, QN => 
                           DataPath_RF_bus_reg_dataout_452_port);
   DataPath_RF_BLOCKi_23_Q_reg_4_inst : DFF_X1 port map( D => n3952, CK => CLK,
                           Q => n_2351, QN => 
                           DataPath_RF_bus_reg_dataout_484_port);
   DataPath_RF_BLOCKi_24_Q_reg_4_inst : DFF_X1 port map( D => n4020, CK => CLK,
                           Q => n_2352, QN => 
                           DataPath_RF_bus_reg_dataout_516_port);
   DataPath_RF_BLOCKi_25_Q_reg_4_inst : DFF_X1 port map( D => n4061, CK => CLK,
                           Q => n_2353, QN => 
                           DataPath_RF_bus_reg_dataout_548_port);
   DataPath_RF_BLOCKi_26_Q_reg_4_inst : DFF_X1 port map( D => n4096, CK => CLK,
                           Q => n_2354, QN => 
                           DataPath_RF_bus_reg_dataout_580_port);
   DataPath_RF_BLOCKi_27_Q_reg_4_inst : DFF_X1 port map( D => n4131, CK => CLK,
                           Q => n_2355, QN => 
                           DataPath_RF_bus_reg_dataout_612_port);
   DataPath_RF_BLOCKi_28_Q_reg_4_inst : DFF_X1 port map( D => n4166, CK => CLK,
                           Q => n_2356, QN => 
                           DataPath_RF_bus_reg_dataout_644_port);
   DataPath_RF_BLOCKi_29_Q_reg_4_inst : DFF_X1 port map( D => n4201, CK => CLK,
                           Q => n_2357, QN => 
                           DataPath_RF_bus_reg_dataout_676_port);
   DataPath_RF_BLOCKi_30_Q_reg_4_inst : DFF_X1 port map( D => n4236, CK => CLK,
                           Q => n_2358, QN => 
                           DataPath_RF_bus_reg_dataout_708_port);
   DataPath_RF_BLOCKi_31_Q_reg_4_inst : DFF_X1 port map( D => n4271, CK => CLK,
                           Q => n_2359, QN => 
                           DataPath_RF_bus_reg_dataout_740_port);
   DataPath_RF_BLOCKi_32_Q_reg_4_inst : DFF_X1 port map( D => n4306, CK => CLK,
                           Q => n_2360, QN => 
                           DataPath_RF_bus_reg_dataout_772_port);
   DataPath_RF_BLOCKi_33_Q_reg_4_inst : DFF_X1 port map( D => n4341, CK => CLK,
                           Q => n_2361, QN => 
                           DataPath_RF_bus_reg_dataout_804_port);
   DataPath_RF_BLOCKi_34_Q_reg_4_inst : DFF_X1 port map( D => n4376, CK => CLK,
                           Q => n_2362, QN => 
                           DataPath_RF_bus_reg_dataout_836_port);
   DataPath_RF_BLOCKi_35_Q_reg_4_inst : DFF_X1 port map( D => n4411, CK => CLK,
                           Q => n_2363, QN => 
                           DataPath_RF_bus_reg_dataout_868_port);
   DataPath_RF_BLOCKi_36_Q_reg_4_inst : DFF_X1 port map( D => n4446, CK => CLK,
                           Q => n_2364, QN => 
                           DataPath_RF_bus_reg_dataout_900_port);
   DataPath_RF_BLOCKi_37_Q_reg_4_inst : DFF_X1 port map( D => n4481, CK => CLK,
                           Q => n_2365, QN => 
                           DataPath_RF_bus_reg_dataout_932_port);
   DataPath_RF_BLOCKi_38_Q_reg_4_inst : DFF_X1 port map( D => n4516, CK => CLK,
                           Q => n_2366, QN => 
                           DataPath_RF_bus_reg_dataout_964_port);
   DataPath_RF_BLOCKi_39_Q_reg_4_inst : DFF_X1 port map( D => n4551, CK => CLK,
                           Q => n_2367, QN => 
                           DataPath_RF_bus_reg_dataout_996_port);
   DataPath_RF_BLOCKi_40_Q_reg_4_inst : DFF_X1 port map( D => n4613, CK => CLK,
                           Q => n_2368, QN => 
                           DataPath_RF_bus_reg_dataout_1028_port);
   DataPath_RF_BLOCKi_41_Q_reg_4_inst : DFF_X1 port map( D => n4654, CK => CLK,
                           Q => n_2369, QN => 
                           DataPath_RF_bus_reg_dataout_1060_port);
   DataPath_RF_BLOCKi_42_Q_reg_4_inst : DFF_X1 port map( D => n4689, CK => CLK,
                           Q => n_2370, QN => 
                           DataPath_RF_bus_reg_dataout_1092_port);
   DataPath_RF_BLOCKi_43_Q_reg_4_inst : DFF_X1 port map( D => n4724, CK => CLK,
                           Q => n_2371, QN => 
                           DataPath_RF_bus_reg_dataout_1124_port);
   DataPath_RF_BLOCKi_44_Q_reg_4_inst : DFF_X1 port map( D => n4759, CK => CLK,
                           Q => n_2372, QN => 
                           DataPath_RF_bus_reg_dataout_1156_port);
   DataPath_RF_BLOCKi_45_Q_reg_4_inst : DFF_X1 port map( D => n4794, CK => CLK,
                           Q => n_2373, QN => 
                           DataPath_RF_bus_reg_dataout_1188_port);
   DataPath_RF_BLOCKi_46_Q_reg_4_inst : DFF_X1 port map( D => n4829, CK => CLK,
                           Q => n_2374, QN => 
                           DataPath_RF_bus_reg_dataout_1220_port);
   DataPath_RF_BLOCKi_47_Q_reg_4_inst : DFF_X1 port map( D => n4864, CK => CLK,
                           Q => n_2375, QN => 
                           DataPath_RF_bus_reg_dataout_1252_port);
   DataPath_RF_BLOCKi_48_Q_reg_4_inst : DFF_X1 port map( D => n4899, CK => CLK,
                           Q => n_2376, QN => 
                           DataPath_RF_bus_reg_dataout_1284_port);
   DataPath_RF_BLOCKi_49_Q_reg_4_inst : DFF_X1 port map( D => n4934, CK => CLK,
                           Q => n_2377, QN => 
                           DataPath_RF_bus_reg_dataout_1316_port);
   DataPath_RF_BLOCKi_50_Q_reg_4_inst : DFF_X1 port map( D => n4969, CK => CLK,
                           Q => n_2378, QN => 
                           DataPath_RF_bus_reg_dataout_1348_port);
   DataPath_RF_BLOCKi_51_Q_reg_4_inst : DFF_X1 port map( D => n5004, CK => CLK,
                           Q => n_2379, QN => 
                           DataPath_RF_bus_reg_dataout_1380_port);
   DataPath_RF_BLOCKi_52_Q_reg_4_inst : DFF_X1 port map( D => n5039, CK => CLK,
                           Q => n_2380, QN => 
                           DataPath_RF_bus_reg_dataout_1412_port);
   DataPath_RF_BLOCKi_53_Q_reg_4_inst : DFF_X1 port map( D => n5074, CK => CLK,
                           Q => n_2381, QN => 
                           DataPath_RF_bus_reg_dataout_1444_port);
   DataPath_RF_BLOCKi_54_Q_reg_4_inst : DFF_X1 port map( D => n5109, CK => CLK,
                           Q => n_2382, QN => 
                           DataPath_RF_bus_reg_dataout_1476_port);
   DataPath_RF_BLOCKi_55_Q_reg_4_inst : DFF_X1 port map( D => n5144, CK => CLK,
                           Q => n_2383, QN => 
                           DataPath_RF_bus_reg_dataout_1508_port);
   DataPath_RF_BLOCKi_56_Q_reg_4_inst : DFF_X1 port map( D => n5206, CK => CLK,
                           Q => n_2384, QN => 
                           DataPath_RF_bus_reg_dataout_1540_port);
   DataPath_RF_BLOCKi_57_Q_reg_4_inst : DFF_X1 port map( D => n5246, CK => CLK,
                           Q => n_2385, QN => 
                           DataPath_RF_bus_reg_dataout_1572_port);
   DataPath_RF_BLOCKi_58_Q_reg_4_inst : DFF_X1 port map( D => n5282, CK => CLK,
                           Q => n_2386, QN => 
                           DataPath_RF_bus_reg_dataout_1604_port);
   DataPath_RF_BLOCKi_59_Q_reg_4_inst : DFF_X1 port map( D => n5317, CK => CLK,
                           Q => n_2387, QN => 
                           DataPath_RF_bus_reg_dataout_1636_port);
   DataPath_RF_BLOCKi_60_Q_reg_4_inst : DFF_X1 port map( D => n5352, CK => CLK,
                           Q => n_2388, QN => 
                           DataPath_RF_bus_reg_dataout_1668_port);
   DataPath_RF_BLOCKi_61_Q_reg_4_inst : DFF_X1 port map( D => n5387, CK => CLK,
                           Q => n_2389, QN => 
                           DataPath_RF_bus_reg_dataout_1700_port);
   DataPath_RF_BLOCKi_62_Q_reg_4_inst : DFF_X1 port map( D => n5422, CK => CLK,
                           Q => n_2390, QN => 
                           DataPath_RF_bus_reg_dataout_1732_port);
   DataPath_RF_BLOCKi_63_Q_reg_4_inst : DFF_X1 port map( D => n5457, CK => CLK,
                           Q => n_2391, QN => 
                           DataPath_RF_bus_reg_dataout_1764_port);
   DataPath_RF_BLOCKi_64_Q_reg_4_inst : DFF_X1 port map( D => n5492, CK => CLK,
                           Q => n_2392, QN => 
                           DataPath_RF_bus_reg_dataout_1796_port);
   DataPath_RF_BLOCKi_65_Q_reg_4_inst : DFF_X1 port map( D => n5527, CK => CLK,
                           Q => n_2393, QN => 
                           DataPath_RF_bus_reg_dataout_1828_port);
   DataPath_RF_BLOCKi_66_Q_reg_4_inst : DFF_X1 port map( D => n5562, CK => CLK,
                           Q => n_2394, QN => 
                           DataPath_RF_bus_reg_dataout_1860_port);
   DataPath_RF_BLOCKi_67_Q_reg_4_inst : DFF_X1 port map( D => n5597, CK => CLK,
                           Q => n_2395, QN => 
                           DataPath_RF_bus_reg_dataout_1892_port);
   DataPath_RF_BLOCKi_68_Q_reg_4_inst : DFF_X1 port map( D => n5636, CK => CLK,
                           Q => n_2396, QN => 
                           DataPath_RF_bus_reg_dataout_1924_port);
   DataPath_RF_BLOCKi_69_Q_reg_4_inst : DFF_X1 port map( D => n5673, CK => CLK,
                           Q => n_2397, QN => 
                           DataPath_RF_bus_reg_dataout_1956_port);
   DataPath_RF_BLOCKi_70_Q_reg_4_inst : DFF_X1 port map( D => n5710, CK => CLK,
                           Q => n_2398, QN => 
                           DataPath_RF_bus_reg_dataout_1988_port);
   DataPath_RF_BLOCKi_71_Q_reg_4_inst : DFF_X1 port map( D => n5747, CK => CLK,
                           Q => n_2399, QN => 
                           DataPath_RF_bus_reg_dataout_2020_port);
   DataPath_RF_BLOCKi_82_Q_reg_4_inst : DFF_X1 port map( D => n904, CK => CLK, 
                           Q => n_2400, QN => 
                           DataPath_RF_bus_reg_dataout_2372_port);
   DataPath_RF_BLOCKi_83_Q_reg_4_inst : DFF_X1 port map( D => n959, CK => CLK, 
                           Q => n_2401, QN => 
                           DataPath_RF_bus_reg_dataout_2404_port);
   DataPath_RF_BLOCKi_84_Q_reg_4_inst : DFF_X1 port map( D => n997, CK => CLK, 
                           Q => n_2402, QN => 
                           DataPath_RF_bus_reg_dataout_2436_port);
   DataPath_RF_BLOCKi_85_Q_reg_4_inst : DFF_X1 port map( D => n1034, CK => CLK,
                           Q => n_2403, QN => 
                           DataPath_RF_bus_reg_dataout_2468_port);
   DataPath_RF_BLOCKi_86_Q_reg_4_inst : DFF_X1 port map( D => n1071, CK => CLK,
                           Q => n_2404, QN => 
                           DataPath_RF_bus_reg_dataout_2500_port);
   DataPath_RF_BLOCKi_87_Q_reg_4_inst : DFF_X1 port map( D => n1108, CK => CLK,
                           Q => n_2405, QN => 
                           DataPath_RF_bus_reg_dataout_2532_port);
   DataPath_RF_BLOCKi_72_Q_reg_4_inst : DFF_X1 port map( D => n5784, CK => CLK,
                           Q => n_2406, QN => 
                           DataPath_RF_bus_reg_dataout_2052_port);
   DataPath_RF_BLOCKi_73_Q_reg_4_inst : DFF_X1 port map( D => n5823, CK => CLK,
                           Q => n_2407, QN => 
                           DataPath_RF_bus_reg_dataout_2084_port);
   DataPath_RF_BLOCKi_74_Q_reg_4_inst : DFF_X1 port map( D => n5859, CK => CLK,
                           Q => n_2408, QN => 
                           DataPath_RF_bus_reg_dataout_2116_port);
   DataPath_RF_BLOCKi_75_Q_reg_4_inst : DFF_X1 port map( D => n5895, CK => CLK,
                           Q => n_2409, QN => 
                           DataPath_RF_bus_reg_dataout_2148_port);
   DataPath_RF_BLOCKi_76_Q_reg_4_inst : DFF_X1 port map( D => n5931, CK => CLK,
                           Q => n_2410, QN => 
                           DataPath_RF_bus_reg_dataout_2180_port);
   DataPath_RF_BLOCKi_77_Q_reg_4_inst : DFF_X1 port map( D => n5967, CK => CLK,
                           Q => n_2411, QN => 
                           DataPath_RF_bus_reg_dataout_2212_port);
   DataPath_RF_BLOCKi_78_Q_reg_4_inst : DFF_X1 port map( D => n6003, CK => CLK,
                           Q => n_2412, QN => 
                           DataPath_RF_bus_reg_dataout_2244_port);
   DataPath_RF_BLOCKi_79_Q_reg_4_inst : DFF_X1 port map( D => n6039, CK => CLK,
                           Q => n_2413, QN => 
                           DataPath_RF_bus_reg_dataout_2276_port);
   DataPath_RF_BLOCKi_80_Q_reg_4_inst : DFF_X1 port map( D => n6076, CK => CLK,
                           Q => n_2414, QN => 
                           DataPath_RF_bus_reg_dataout_2308_port);
   DataPath_RF_BLOCKi_81_Q_reg_4_inst : DFF_X1 port map( D => n6112, CK => CLK,
                           Q => n_2415, QN => 
                           DataPath_RF_bus_reg_dataout_2340_port);
   DataPath_REG_ALU_OUT_Q_reg_8_inst : DFF_X1 port map( D => n7015, CK => CLK, 
                           Q => DRAM_ADDRESS_8_port, QN => n498);
   DataPath_REG_MEM_ALUOUT_Q_reg_8_inst : DFF_X1 port map( D => n1141, CK => 
                           CLK, Q => n_2416, QN => 
                           DataPath_i_REG_MEM_ALUOUT_8_port);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_8_inst : DFF_X1 port map( D => n6855, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_104_port
                           , QN => n671);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_8_inst : DFF_X1 port map( D => n6887, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_136_port
                           , QN => n703);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_8_inst : DFF_X1 port map( D => n6951, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_200_port
                           , QN => n767);
   DataPath_RF_BLOCKi_8_Q_reg_8_inst : DFF_X1 port map( D => n3356, CK => CLK, 
                           Q => n_2417, QN => 
                           DataPath_RF_bus_reg_dataout_8_port);
   DataPath_RF_BLOCKi_9_Q_reg_8_inst : DFF_X1 port map( D => n3404, CK => CLK, 
                           Q => n_2418, QN => 
                           DataPath_RF_bus_reg_dataout_40_port);
   DataPath_RF_BLOCKi_10_Q_reg_8_inst : DFF_X1 port map( D => n3442, CK => CLK,
                           Q => n_2419, QN => 
                           DataPath_RF_bus_reg_dataout_72_port);
   DataPath_RF_BLOCKi_11_Q_reg_8_inst : DFF_X1 port map( D => n3480, CK => CLK,
                           Q => n_2420, QN => 
                           DataPath_RF_bus_reg_dataout_104_port);
   DataPath_RF_BLOCKi_12_Q_reg_8_inst : DFF_X1 port map( D => n3518, CK => CLK,
                           Q => n_2421, QN => 
                           DataPath_RF_bus_reg_dataout_136_port);
   DataPath_RF_BLOCKi_13_Q_reg_8_inst : DFF_X1 port map( D => n3556, CK => CLK,
                           Q => n_2422, QN => 
                           DataPath_RF_bus_reg_dataout_168_port);
   DataPath_RF_BLOCKi_14_Q_reg_8_inst : DFF_X1 port map( D => n3594, CK => CLK,
                           Q => n_2423, QN => 
                           DataPath_RF_bus_reg_dataout_200_port);
   DataPath_RF_BLOCKi_15_Q_reg_8_inst : DFF_X1 port map( D => n3632, CK => CLK,
                           Q => n_2424, QN => 
                           DataPath_RF_bus_reg_dataout_232_port);
   DataPath_RF_BLOCKi_16_Q_reg_8_inst : DFF_X1 port map( D => n3670, CK => CLK,
                           Q => n_2425, QN => 
                           DataPath_RF_bus_reg_dataout_264_port);
   DataPath_RF_BLOCKi_17_Q_reg_8_inst : DFF_X1 port map( D => n3707, CK => CLK,
                           Q => n_2426, QN => 
                           DataPath_RF_bus_reg_dataout_296_port);
   DataPath_RF_BLOCKi_18_Q_reg_8_inst : DFF_X1 port map( D => n3744, CK => CLK,
                           Q => n_2427, QN => 
                           DataPath_RF_bus_reg_dataout_328_port);
   DataPath_RF_BLOCKi_19_Q_reg_8_inst : DFF_X1 port map( D => n3781, CK => CLK,
                           Q => n_2428, QN => 
                           DataPath_RF_bus_reg_dataout_360_port);
   DataPath_RF_BLOCKi_20_Q_reg_8_inst : DFF_X1 port map( D => n3816, CK => CLK,
                           Q => n_2429, QN => 
                           DataPath_RF_bus_reg_dataout_392_port);
   DataPath_RF_BLOCKi_21_Q_reg_8_inst : DFF_X1 port map( D => n3851, CK => CLK,
                           Q => n_2430, QN => 
                           DataPath_RF_bus_reg_dataout_424_port);
   DataPath_RF_BLOCKi_22_Q_reg_8_inst : DFF_X1 port map( D => n3886, CK => CLK,
                           Q => n_2431, QN => 
                           DataPath_RF_bus_reg_dataout_456_port);
   DataPath_RF_BLOCKi_23_Q_reg_8_inst : DFF_X1 port map( D => n3944, CK => CLK,
                           Q => n_2432, QN => 
                           DataPath_RF_bus_reg_dataout_488_port);
   DataPath_RF_BLOCKi_24_Q_reg_8_inst : DFF_X1 port map( D => n4012, CK => CLK,
                           Q => n_2433, QN => 
                           DataPath_RF_bus_reg_dataout_520_port);
   DataPath_RF_BLOCKi_25_Q_reg_8_inst : DFF_X1 port map( D => n4057, CK => CLK,
                           Q => n_2434, QN => 
                           DataPath_RF_bus_reg_dataout_552_port);
   DataPath_RF_BLOCKi_26_Q_reg_8_inst : DFF_X1 port map( D => n4092, CK => CLK,
                           Q => n_2435, QN => 
                           DataPath_RF_bus_reg_dataout_584_port);
   DataPath_RF_BLOCKi_27_Q_reg_8_inst : DFF_X1 port map( D => n4127, CK => CLK,
                           Q => n_2436, QN => 
                           DataPath_RF_bus_reg_dataout_616_port);
   DataPath_RF_BLOCKi_28_Q_reg_8_inst : DFF_X1 port map( D => n4162, CK => CLK,
                           Q => n_2437, QN => 
                           DataPath_RF_bus_reg_dataout_648_port);
   DataPath_RF_BLOCKi_29_Q_reg_8_inst : DFF_X1 port map( D => n4197, CK => CLK,
                           Q => n_2438, QN => 
                           DataPath_RF_bus_reg_dataout_680_port);
   DataPath_RF_BLOCKi_30_Q_reg_8_inst : DFF_X1 port map( D => n4232, CK => CLK,
                           Q => n_2439, QN => 
                           DataPath_RF_bus_reg_dataout_712_port);
   DataPath_RF_BLOCKi_31_Q_reg_8_inst : DFF_X1 port map( D => n4267, CK => CLK,
                           Q => n_2440, QN => 
                           DataPath_RF_bus_reg_dataout_744_port);
   DataPath_RF_BLOCKi_32_Q_reg_8_inst : DFF_X1 port map( D => n4302, CK => CLK,
                           Q => n_2441, QN => 
                           DataPath_RF_bus_reg_dataout_776_port);
   DataPath_RF_BLOCKi_33_Q_reg_8_inst : DFF_X1 port map( D => n4337, CK => CLK,
                           Q => n_2442, QN => 
                           DataPath_RF_bus_reg_dataout_808_port);
   DataPath_RF_BLOCKi_34_Q_reg_8_inst : DFF_X1 port map( D => n4372, CK => CLK,
                           Q => n_2443, QN => 
                           DataPath_RF_bus_reg_dataout_840_port);
   DataPath_RF_BLOCKi_35_Q_reg_8_inst : DFF_X1 port map( D => n4407, CK => CLK,
                           Q => n_2444, QN => 
                           DataPath_RF_bus_reg_dataout_872_port);
   DataPath_RF_BLOCKi_36_Q_reg_8_inst : DFF_X1 port map( D => n4442, CK => CLK,
                           Q => n_2445, QN => 
                           DataPath_RF_bus_reg_dataout_904_port);
   DataPath_RF_BLOCKi_37_Q_reg_8_inst : DFF_X1 port map( D => n4477, CK => CLK,
                           Q => n_2446, QN => 
                           DataPath_RF_bus_reg_dataout_936_port);
   DataPath_RF_BLOCKi_38_Q_reg_8_inst : DFF_X1 port map( D => n4512, CK => CLK,
                           Q => n_2447, QN => 
                           DataPath_RF_bus_reg_dataout_968_port);
   DataPath_RF_BLOCKi_39_Q_reg_8_inst : DFF_X1 port map( D => n4547, CK => CLK,
                           Q => n_2448, QN => 
                           DataPath_RF_bus_reg_dataout_1000_port);
   DataPath_RF_BLOCKi_40_Q_reg_8_inst : DFF_X1 port map( D => n4605, CK => CLK,
                           Q => n_2449, QN => 
                           DataPath_RF_bus_reg_dataout_1032_port);
   DataPath_RF_BLOCKi_41_Q_reg_8_inst : DFF_X1 port map( D => n4650, CK => CLK,
                           Q => n_2450, QN => 
                           DataPath_RF_bus_reg_dataout_1064_port);
   DataPath_RF_BLOCKi_42_Q_reg_8_inst : DFF_X1 port map( D => n4685, CK => CLK,
                           Q => n_2451, QN => 
                           DataPath_RF_bus_reg_dataout_1096_port);
   DataPath_RF_BLOCKi_43_Q_reg_8_inst : DFF_X1 port map( D => n4720, CK => CLK,
                           Q => n_2452, QN => 
                           DataPath_RF_bus_reg_dataout_1128_port);
   DataPath_RF_BLOCKi_44_Q_reg_8_inst : DFF_X1 port map( D => n4755, CK => CLK,
                           Q => n_2453, QN => 
                           DataPath_RF_bus_reg_dataout_1160_port);
   DataPath_RF_BLOCKi_45_Q_reg_8_inst : DFF_X1 port map( D => n4790, CK => CLK,
                           Q => n_2454, QN => 
                           DataPath_RF_bus_reg_dataout_1192_port);
   DataPath_RF_BLOCKi_46_Q_reg_8_inst : DFF_X1 port map( D => n4825, CK => CLK,
                           Q => n_2455, QN => 
                           DataPath_RF_bus_reg_dataout_1224_port);
   DataPath_RF_BLOCKi_47_Q_reg_8_inst : DFF_X1 port map( D => n4860, CK => CLK,
                           Q => n_2456, QN => 
                           DataPath_RF_bus_reg_dataout_1256_port);
   DataPath_RF_BLOCKi_48_Q_reg_8_inst : DFF_X1 port map( D => n4895, CK => CLK,
                           Q => n_2457, QN => 
                           DataPath_RF_bus_reg_dataout_1288_port);
   DataPath_RF_BLOCKi_49_Q_reg_8_inst : DFF_X1 port map( D => n4930, CK => CLK,
                           Q => n_2458, QN => 
                           DataPath_RF_bus_reg_dataout_1320_port);
   DataPath_RF_BLOCKi_50_Q_reg_8_inst : DFF_X1 port map( D => n4965, CK => CLK,
                           Q => n_2459, QN => 
                           DataPath_RF_bus_reg_dataout_1352_port);
   DataPath_RF_BLOCKi_51_Q_reg_8_inst : DFF_X1 port map( D => n5000, CK => CLK,
                           Q => n_2460, QN => 
                           DataPath_RF_bus_reg_dataout_1384_port);
   DataPath_RF_BLOCKi_52_Q_reg_8_inst : DFF_X1 port map( D => n5035, CK => CLK,
                           Q => n_2461, QN => 
                           DataPath_RF_bus_reg_dataout_1416_port);
   DataPath_RF_BLOCKi_53_Q_reg_8_inst : DFF_X1 port map( D => n5070, CK => CLK,
                           Q => n_2462, QN => 
                           DataPath_RF_bus_reg_dataout_1448_port);
   DataPath_RF_BLOCKi_54_Q_reg_8_inst : DFF_X1 port map( D => n5105, CK => CLK,
                           Q => n_2463, QN => 
                           DataPath_RF_bus_reg_dataout_1480_port);
   DataPath_RF_BLOCKi_55_Q_reg_8_inst : DFF_X1 port map( D => n5140, CK => CLK,
                           Q => n_2464, QN => 
                           DataPath_RF_bus_reg_dataout_1512_port);
   DataPath_RF_BLOCKi_56_Q_reg_8_inst : DFF_X1 port map( D => n5198, CK => CLK,
                           Q => n_2465, QN => 
                           DataPath_RF_bus_reg_dataout_1544_port);
   DataPath_RF_BLOCKi_57_Q_reg_8_inst : DFF_X1 port map( D => n5242, CK => CLK,
                           Q => n_2466, QN => 
                           DataPath_RF_bus_reg_dataout_1576_port);
   DataPath_RF_BLOCKi_58_Q_reg_8_inst : DFF_X1 port map( D => n5278, CK => CLK,
                           Q => n_2467, QN => 
                           DataPath_RF_bus_reg_dataout_1608_port);
   DataPath_RF_BLOCKi_59_Q_reg_8_inst : DFF_X1 port map( D => n5313, CK => CLK,
                           Q => n_2468, QN => 
                           DataPath_RF_bus_reg_dataout_1640_port);
   DataPath_RF_BLOCKi_60_Q_reg_8_inst : DFF_X1 port map( D => n5348, CK => CLK,
                           Q => n_2469, QN => 
                           DataPath_RF_bus_reg_dataout_1672_port);
   DataPath_RF_BLOCKi_61_Q_reg_8_inst : DFF_X1 port map( D => n5383, CK => CLK,
                           Q => n_2470, QN => 
                           DataPath_RF_bus_reg_dataout_1704_port);
   DataPath_RF_BLOCKi_62_Q_reg_8_inst : DFF_X1 port map( D => n5418, CK => CLK,
                           Q => n_2471, QN => 
                           DataPath_RF_bus_reg_dataout_1736_port);
   DataPath_RF_BLOCKi_63_Q_reg_8_inst : DFF_X1 port map( D => n5453, CK => CLK,
                           Q => n_2472, QN => 
                           DataPath_RF_bus_reg_dataout_1768_port);
   DataPath_RF_BLOCKi_64_Q_reg_8_inst : DFF_X1 port map( D => n5488, CK => CLK,
                           Q => n_2473, QN => 
                           DataPath_RF_bus_reg_dataout_1800_port);
   DataPath_RF_BLOCKi_65_Q_reg_8_inst : DFF_X1 port map( D => n5523, CK => CLK,
                           Q => n_2474, QN => 
                           DataPath_RF_bus_reg_dataout_1832_port);
   DataPath_RF_BLOCKi_66_Q_reg_8_inst : DFF_X1 port map( D => n5558, CK => CLK,
                           Q => n_2475, QN => 
                           DataPath_RF_bus_reg_dataout_1864_port);
   DataPath_RF_BLOCKi_67_Q_reg_8_inst : DFF_X1 port map( D => n5593, CK => CLK,
                           Q => n_2476, QN => 
                           DataPath_RF_bus_reg_dataout_1896_port);
   DataPath_RF_BLOCKi_68_Q_reg_8_inst : DFF_X1 port map( D => n5632, CK => CLK,
                           Q => n_2477, QN => 
                           DataPath_RF_bus_reg_dataout_1928_port);
   DataPath_RF_BLOCKi_69_Q_reg_8_inst : DFF_X1 port map( D => n5669, CK => CLK,
                           Q => n_2478, QN => 
                           DataPath_RF_bus_reg_dataout_1960_port);
   DataPath_RF_BLOCKi_70_Q_reg_8_inst : DFF_X1 port map( D => n5706, CK => CLK,
                           Q => n_2479, QN => 
                           DataPath_RF_bus_reg_dataout_1992_port);
   DataPath_RF_BLOCKi_71_Q_reg_8_inst : DFF_X1 port map( D => n5743, CK => CLK,
                           Q => n_2480, QN => 
                           DataPath_RF_bus_reg_dataout_2024_port);
   DataPath_RF_BLOCKi_82_Q_reg_8_inst : DFF_X1 port map( D => n896, CK => CLK, 
                           Q => n_2481, QN => 
                           DataPath_RF_bus_reg_dataout_2376_port);
   DataPath_RF_BLOCKi_83_Q_reg_8_inst : DFF_X1 port map( D => n955, CK => CLK, 
                           Q => n_2482, QN => 
                           DataPath_RF_bus_reg_dataout_2408_port);
   DataPath_RF_BLOCKi_84_Q_reg_8_inst : DFF_X1 port map( D => n993, CK => CLK, 
                           Q => n_2483, QN => 
                           DataPath_RF_bus_reg_dataout_2440_port);
   DataPath_RF_BLOCKi_85_Q_reg_8_inst : DFF_X1 port map( D => n1030, CK => CLK,
                           Q => n_2484, QN => 
                           DataPath_RF_bus_reg_dataout_2472_port);
   DataPath_RF_BLOCKi_86_Q_reg_8_inst : DFF_X1 port map( D => n1067, CK => CLK,
                           Q => n_2485, QN => 
                           DataPath_RF_bus_reg_dataout_2504_port);
   DataPath_RF_BLOCKi_87_Q_reg_8_inst : DFF_X1 port map( D => n1104, CK => CLK,
                           Q => n_2486, QN => 
                           DataPath_RF_bus_reg_dataout_2536_port);
   DataPath_RF_BLOCKi_72_Q_reg_8_inst : DFF_X1 port map( D => n5780, CK => CLK,
                           Q => n_2487, QN => 
                           DataPath_RF_bus_reg_dataout_2056_port);
   DataPath_RF_BLOCKi_73_Q_reg_8_inst : DFF_X1 port map( D => n5819, CK => CLK,
                           Q => n_2488, QN => 
                           DataPath_RF_bus_reg_dataout_2088_port);
   DataPath_RF_BLOCKi_74_Q_reg_8_inst : DFF_X1 port map( D => n5855, CK => CLK,
                           Q => n_2489, QN => 
                           DataPath_RF_bus_reg_dataout_2120_port);
   DataPath_RF_BLOCKi_75_Q_reg_8_inst : DFF_X1 port map( D => n5891, CK => CLK,
                           Q => n_2490, QN => 
                           DataPath_RF_bus_reg_dataout_2152_port);
   DataPath_RF_BLOCKi_76_Q_reg_8_inst : DFF_X1 port map( D => n5927, CK => CLK,
                           Q => n_2491, QN => 
                           DataPath_RF_bus_reg_dataout_2184_port);
   DataPath_RF_BLOCKi_77_Q_reg_8_inst : DFF_X1 port map( D => n5963, CK => CLK,
                           Q => n_2492, QN => 
                           DataPath_RF_bus_reg_dataout_2216_port);
   DataPath_RF_BLOCKi_78_Q_reg_8_inst : DFF_X1 port map( D => n5999, CK => CLK,
                           Q => n_2493, QN => 
                           DataPath_RF_bus_reg_dataout_2248_port);
   DataPath_RF_BLOCKi_79_Q_reg_8_inst : DFF_X1 port map( D => n6035, CK => CLK,
                           Q => n_2494, QN => 
                           DataPath_RF_bus_reg_dataout_2280_port);
   DataPath_RF_BLOCKi_80_Q_reg_8_inst : DFF_X1 port map( D => n6072, CK => CLK,
                           Q => n_2495, QN => 
                           DataPath_RF_bus_reg_dataout_2312_port);
   DataPath_RF_BLOCKi_81_Q_reg_8_inst : DFF_X1 port map( D => n6108, CK => CLK,
                           Q => n_2496, QN => 
                           DataPath_RF_bus_reg_dataout_2344_port);
   DataPath_REG_ALU_OUT_Q_reg_10_inst : DFF_X1 port map( D => n7013, CK => CLK,
                           Q => DRAM_ADDRESS_10_port, QN => n499);
   DataPath_REG_MEM_ALUOUT_Q_reg_10_inst : DFF_X1 port map( D => n1139, CK => 
                           CLK, Q => n_2497, QN => 
                           DataPath_i_REG_MEM_ALUOUT_10_port);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_10_inst : DFF_X1 port map( D => n6821, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_74_port,
                           QN => n641);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_10_inst : DFF_X1 port map( D => n6853, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_106_port
                           , QN => n673);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_10_inst : DFF_X1 port map( D => n6885, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_138_port
                           , QN => n705);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_10_inst : DFF_X1 port map( D => n6949, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_202_port
                           , QN => n769);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_10_inst : DFF_X1 port map( D => n6981, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_234_port
                           , QN => n801);
   DataPath_RF_BLOCKi_8_Q_reg_10_inst : DFF_X1 port map( D => n3352, CK => CLK,
                           Q => n_2498, QN => 
                           DataPath_RF_bus_reg_dataout_10_port);
   DataPath_RF_BLOCKi_9_Q_reg_10_inst : DFF_X1 port map( D => n3402, CK => CLK,
                           Q => n_2499, QN => 
                           DataPath_RF_bus_reg_dataout_42_port);
   DataPath_RF_BLOCKi_10_Q_reg_10_inst : DFF_X1 port map( D => n3440, CK => CLK
                           , Q => n_2500, QN => 
                           DataPath_RF_bus_reg_dataout_74_port);
   DataPath_RF_BLOCKi_11_Q_reg_10_inst : DFF_X1 port map( D => n3478, CK => CLK
                           , Q => n_2501, QN => 
                           DataPath_RF_bus_reg_dataout_106_port);
   DataPath_RF_BLOCKi_12_Q_reg_10_inst : DFF_X1 port map( D => n3516, CK => CLK
                           , Q => n_2502, QN => 
                           DataPath_RF_bus_reg_dataout_138_port);
   DataPath_RF_BLOCKi_13_Q_reg_10_inst : DFF_X1 port map( D => n3554, CK => CLK
                           , Q => n_2503, QN => 
                           DataPath_RF_bus_reg_dataout_170_port);
   DataPath_RF_BLOCKi_14_Q_reg_10_inst : DFF_X1 port map( D => n3592, CK => CLK
                           , Q => n_2504, QN => 
                           DataPath_RF_bus_reg_dataout_202_port);
   DataPath_RF_BLOCKi_15_Q_reg_10_inst : DFF_X1 port map( D => n3630, CK => CLK
                           , Q => n_2505, QN => 
                           DataPath_RF_bus_reg_dataout_234_port);
   DataPath_RF_BLOCKi_16_Q_reg_10_inst : DFF_X1 port map( D => n3668, CK => CLK
                           , Q => n_2506, QN => 
                           DataPath_RF_bus_reg_dataout_266_port);
   DataPath_RF_BLOCKi_17_Q_reg_10_inst : DFF_X1 port map( D => n3705, CK => CLK
                           , Q => n_2507, QN => 
                           DataPath_RF_bus_reg_dataout_298_port);
   DataPath_RF_BLOCKi_18_Q_reg_10_inst : DFF_X1 port map( D => n3742, CK => CLK
                           , Q => n_2508, QN => 
                           DataPath_RF_bus_reg_dataout_330_port);
   DataPath_RF_BLOCKi_19_Q_reg_10_inst : DFF_X1 port map( D => n3779, CK => CLK
                           , Q => n_2509, QN => 
                           DataPath_RF_bus_reg_dataout_362_port);
   DataPath_RF_BLOCKi_20_Q_reg_10_inst : DFF_X1 port map( D => n3814, CK => CLK
                           , Q => n_2510, QN => 
                           DataPath_RF_bus_reg_dataout_394_port);
   DataPath_RF_BLOCKi_21_Q_reg_10_inst : DFF_X1 port map( D => n3849, CK => CLK
                           , Q => n_2511, QN => 
                           DataPath_RF_bus_reg_dataout_426_port);
   DataPath_RF_BLOCKi_22_Q_reg_10_inst : DFF_X1 port map( D => n3884, CK => CLK
                           , Q => n_2512, QN => 
                           DataPath_RF_bus_reg_dataout_458_port);
   DataPath_RF_BLOCKi_23_Q_reg_10_inst : DFF_X1 port map( D => n3940, CK => CLK
                           , Q => n_2513, QN => 
                           DataPath_RF_bus_reg_dataout_490_port);
   DataPath_RF_BLOCKi_24_Q_reg_10_inst : DFF_X1 port map( D => n4008, CK => CLK
                           , Q => n_2514, QN => 
                           DataPath_RF_bus_reg_dataout_522_port);
   DataPath_RF_BLOCKi_25_Q_reg_10_inst : DFF_X1 port map( D => n4055, CK => CLK
                           , Q => n_2515, QN => 
                           DataPath_RF_bus_reg_dataout_554_port);
   DataPath_RF_BLOCKi_26_Q_reg_10_inst : DFF_X1 port map( D => n4090, CK => CLK
                           , Q => n_2516, QN => 
                           DataPath_RF_bus_reg_dataout_586_port);
   DataPath_RF_BLOCKi_27_Q_reg_10_inst : DFF_X1 port map( D => n4125, CK => CLK
                           , Q => n_2517, QN => 
                           DataPath_RF_bus_reg_dataout_618_port);
   DataPath_RF_BLOCKi_28_Q_reg_10_inst : DFF_X1 port map( D => n4160, CK => CLK
                           , Q => n_2518, QN => 
                           DataPath_RF_bus_reg_dataout_650_port);
   DataPath_RF_BLOCKi_29_Q_reg_10_inst : DFF_X1 port map( D => n4195, CK => CLK
                           , Q => n_2519, QN => 
                           DataPath_RF_bus_reg_dataout_682_port);
   DataPath_RF_BLOCKi_30_Q_reg_10_inst : DFF_X1 port map( D => n4230, CK => CLK
                           , Q => n_2520, QN => 
                           DataPath_RF_bus_reg_dataout_714_port);
   DataPath_RF_BLOCKi_31_Q_reg_10_inst : DFF_X1 port map( D => n4265, CK => CLK
                           , Q => n_2521, QN => 
                           DataPath_RF_bus_reg_dataout_746_port);
   DataPath_RF_BLOCKi_32_Q_reg_10_inst : DFF_X1 port map( D => n4300, CK => CLK
                           , Q => n_2522, QN => 
                           DataPath_RF_bus_reg_dataout_778_port);
   DataPath_RF_BLOCKi_33_Q_reg_10_inst : DFF_X1 port map( D => n4335, CK => CLK
                           , Q => n_2523, QN => 
                           DataPath_RF_bus_reg_dataout_810_port);
   DataPath_RF_BLOCKi_34_Q_reg_10_inst : DFF_X1 port map( D => n4370, CK => CLK
                           , Q => n_2524, QN => 
                           DataPath_RF_bus_reg_dataout_842_port);
   DataPath_RF_BLOCKi_35_Q_reg_10_inst : DFF_X1 port map( D => n4405, CK => CLK
                           , Q => n_2525, QN => 
                           DataPath_RF_bus_reg_dataout_874_port);
   DataPath_RF_BLOCKi_36_Q_reg_10_inst : DFF_X1 port map( D => n4440, CK => CLK
                           , Q => n_2526, QN => 
                           DataPath_RF_bus_reg_dataout_906_port);
   DataPath_RF_BLOCKi_37_Q_reg_10_inst : DFF_X1 port map( D => n4475, CK => CLK
                           , Q => n_2527, QN => 
                           DataPath_RF_bus_reg_dataout_938_port);
   DataPath_RF_BLOCKi_38_Q_reg_10_inst : DFF_X1 port map( D => n4510, CK => CLK
                           , Q => n_2528, QN => 
                           DataPath_RF_bus_reg_dataout_970_port);
   DataPath_RF_BLOCKi_39_Q_reg_10_inst : DFF_X1 port map( D => n4545, CK => CLK
                           , Q => n_2529, QN => 
                           DataPath_RF_bus_reg_dataout_1002_port);
   DataPath_RF_BLOCKi_40_Q_reg_10_inst : DFF_X1 port map( D => n4601, CK => CLK
                           , Q => n_2530, QN => 
                           DataPath_RF_bus_reg_dataout_1034_port);
   DataPath_RF_BLOCKi_41_Q_reg_10_inst : DFF_X1 port map( D => n4648, CK => CLK
                           , Q => n_2531, QN => 
                           DataPath_RF_bus_reg_dataout_1066_port);
   DataPath_RF_BLOCKi_42_Q_reg_10_inst : DFF_X1 port map( D => n4683, CK => CLK
                           , Q => n_2532, QN => 
                           DataPath_RF_bus_reg_dataout_1098_port);
   DataPath_RF_BLOCKi_43_Q_reg_10_inst : DFF_X1 port map( D => n4718, CK => CLK
                           , Q => n_2533, QN => 
                           DataPath_RF_bus_reg_dataout_1130_port);
   DataPath_RF_BLOCKi_44_Q_reg_10_inst : DFF_X1 port map( D => n4753, CK => CLK
                           , Q => n_2534, QN => 
                           DataPath_RF_bus_reg_dataout_1162_port);
   DataPath_RF_BLOCKi_45_Q_reg_10_inst : DFF_X1 port map( D => n4788, CK => CLK
                           , Q => n_2535, QN => 
                           DataPath_RF_bus_reg_dataout_1194_port);
   DataPath_RF_BLOCKi_46_Q_reg_10_inst : DFF_X1 port map( D => n4823, CK => CLK
                           , Q => n_2536, QN => 
                           DataPath_RF_bus_reg_dataout_1226_port);
   DataPath_RF_BLOCKi_47_Q_reg_10_inst : DFF_X1 port map( D => n4858, CK => CLK
                           , Q => n_2537, QN => 
                           DataPath_RF_bus_reg_dataout_1258_port);
   DataPath_RF_BLOCKi_48_Q_reg_10_inst : DFF_X1 port map( D => n4893, CK => CLK
                           , Q => n_2538, QN => 
                           DataPath_RF_bus_reg_dataout_1290_port);
   DataPath_RF_BLOCKi_49_Q_reg_10_inst : DFF_X1 port map( D => n4928, CK => CLK
                           , Q => n_2539, QN => 
                           DataPath_RF_bus_reg_dataout_1322_port);
   DataPath_RF_BLOCKi_50_Q_reg_10_inst : DFF_X1 port map( D => n4963, CK => CLK
                           , Q => n_2540, QN => 
                           DataPath_RF_bus_reg_dataout_1354_port);
   DataPath_RF_BLOCKi_51_Q_reg_10_inst : DFF_X1 port map( D => n4998, CK => CLK
                           , Q => n_2541, QN => 
                           DataPath_RF_bus_reg_dataout_1386_port);
   DataPath_RF_BLOCKi_52_Q_reg_10_inst : DFF_X1 port map( D => n5033, CK => CLK
                           , Q => n_2542, QN => 
                           DataPath_RF_bus_reg_dataout_1418_port);
   DataPath_RF_BLOCKi_53_Q_reg_10_inst : DFF_X1 port map( D => n5068, CK => CLK
                           , Q => n_2543, QN => 
                           DataPath_RF_bus_reg_dataout_1450_port);
   DataPath_RF_BLOCKi_54_Q_reg_10_inst : DFF_X1 port map( D => n5103, CK => CLK
                           , Q => n_2544, QN => 
                           DataPath_RF_bus_reg_dataout_1482_port);
   DataPath_RF_BLOCKi_55_Q_reg_10_inst : DFF_X1 port map( D => n5138, CK => CLK
                           , Q => n_2545, QN => 
                           DataPath_RF_bus_reg_dataout_1514_port);
   DataPath_RF_BLOCKi_56_Q_reg_10_inst : DFF_X1 port map( D => n5194, CK => CLK
                           , Q => n_2546, QN => 
                           DataPath_RF_bus_reg_dataout_1546_port);
   DataPath_RF_BLOCKi_57_Q_reg_10_inst : DFF_X1 port map( D => n5240, CK => CLK
                           , Q => n_2547, QN => 
                           DataPath_RF_bus_reg_dataout_1578_port);
   DataPath_RF_BLOCKi_58_Q_reg_10_inst : DFF_X1 port map( D => n5276, CK => CLK
                           , Q => n_2548, QN => 
                           DataPath_RF_bus_reg_dataout_1610_port);
   DataPath_RF_BLOCKi_59_Q_reg_10_inst : DFF_X1 port map( D => n5311, CK => CLK
                           , Q => n_2549, QN => 
                           DataPath_RF_bus_reg_dataout_1642_port);
   DataPath_RF_BLOCKi_60_Q_reg_10_inst : DFF_X1 port map( D => n5346, CK => CLK
                           , Q => n_2550, QN => 
                           DataPath_RF_bus_reg_dataout_1674_port);
   DataPath_RF_BLOCKi_61_Q_reg_10_inst : DFF_X1 port map( D => n5381, CK => CLK
                           , Q => n_2551, QN => 
                           DataPath_RF_bus_reg_dataout_1706_port);
   DataPath_RF_BLOCKi_62_Q_reg_10_inst : DFF_X1 port map( D => n5416, CK => CLK
                           , Q => n_2552, QN => 
                           DataPath_RF_bus_reg_dataout_1738_port);
   DataPath_RF_BLOCKi_63_Q_reg_10_inst : DFF_X1 port map( D => n5451, CK => CLK
                           , Q => n_2553, QN => 
                           DataPath_RF_bus_reg_dataout_1770_port);
   DataPath_RF_BLOCKi_64_Q_reg_10_inst : DFF_X1 port map( D => n5486, CK => CLK
                           , Q => n_2554, QN => 
                           DataPath_RF_bus_reg_dataout_1802_port);
   DataPath_RF_BLOCKi_65_Q_reg_10_inst : DFF_X1 port map( D => n5521, CK => CLK
                           , Q => n_2555, QN => 
                           DataPath_RF_bus_reg_dataout_1834_port);
   DataPath_RF_BLOCKi_66_Q_reg_10_inst : DFF_X1 port map( D => n5556, CK => CLK
                           , Q => n_2556, QN => 
                           DataPath_RF_bus_reg_dataout_1866_port);
   DataPath_RF_BLOCKi_67_Q_reg_10_inst : DFF_X1 port map( D => n5591, CK => CLK
                           , Q => n_2557, QN => 
                           DataPath_RF_bus_reg_dataout_1898_port);
   DataPath_RF_BLOCKi_68_Q_reg_10_inst : DFF_X1 port map( D => n5630, CK => CLK
                           , Q => n_2558, QN => 
                           DataPath_RF_bus_reg_dataout_1930_port);
   DataPath_RF_BLOCKi_69_Q_reg_10_inst : DFF_X1 port map( D => n5667, CK => CLK
                           , Q => n_2559, QN => 
                           DataPath_RF_bus_reg_dataout_1962_port);
   DataPath_RF_BLOCKi_70_Q_reg_10_inst : DFF_X1 port map( D => n5704, CK => CLK
                           , Q => n_2560, QN => 
                           DataPath_RF_bus_reg_dataout_1994_port);
   DataPath_RF_BLOCKi_71_Q_reg_10_inst : DFF_X1 port map( D => n5741, CK => CLK
                           , Q => n_2561, QN => 
                           DataPath_RF_bus_reg_dataout_2026_port);
   DataPath_RF_BLOCKi_82_Q_reg_10_inst : DFF_X1 port map( D => n892, CK => CLK,
                           Q => n_2562, QN => 
                           DataPath_RF_bus_reg_dataout_2378_port);
   DataPath_RF_BLOCKi_83_Q_reg_10_inst : DFF_X1 port map( D => n953, CK => CLK,
                           Q => n_2563, QN => 
                           DataPath_RF_bus_reg_dataout_2410_port);
   DataPath_RF_BLOCKi_84_Q_reg_10_inst : DFF_X1 port map( D => n991, CK => CLK,
                           Q => n_2564, QN => 
                           DataPath_RF_bus_reg_dataout_2442_port);
   DataPath_RF_BLOCKi_85_Q_reg_10_inst : DFF_X1 port map( D => n1028, CK => CLK
                           , Q => n_2565, QN => 
                           DataPath_RF_bus_reg_dataout_2474_port);
   DataPath_RF_BLOCKi_86_Q_reg_10_inst : DFF_X1 port map( D => n1065, CK => CLK
                           , Q => n_2566, QN => 
                           DataPath_RF_bus_reg_dataout_2506_port);
   DataPath_RF_BLOCKi_87_Q_reg_10_inst : DFF_X1 port map( D => n1102, CK => CLK
                           , Q => n_2567, QN => 
                           DataPath_RF_bus_reg_dataout_2538_port);
   DataPath_RF_BLOCKi_72_Q_reg_10_inst : DFF_X1 port map( D => n5778, CK => CLK
                           , Q => n_2568, QN => 
                           DataPath_RF_bus_reg_dataout_2058_port);
   DataPath_RF_BLOCKi_73_Q_reg_10_inst : DFF_X1 port map( D => n5817, CK => CLK
                           , Q => n_2569, QN => 
                           DataPath_RF_bus_reg_dataout_2090_port);
   DataPath_RF_BLOCKi_74_Q_reg_10_inst : DFF_X1 port map( D => n5853, CK => CLK
                           , Q => n_2570, QN => 
                           DataPath_RF_bus_reg_dataout_2122_port);
   DataPath_RF_BLOCKi_75_Q_reg_10_inst : DFF_X1 port map( D => n5889, CK => CLK
                           , Q => n_2571, QN => 
                           DataPath_RF_bus_reg_dataout_2154_port);
   DataPath_RF_BLOCKi_76_Q_reg_10_inst : DFF_X1 port map( D => n5925, CK => CLK
                           , Q => n_2572, QN => 
                           DataPath_RF_bus_reg_dataout_2186_port);
   DataPath_RF_BLOCKi_77_Q_reg_10_inst : DFF_X1 port map( D => n5961, CK => CLK
                           , Q => n_2573, QN => 
                           DataPath_RF_bus_reg_dataout_2218_port);
   DataPath_RF_BLOCKi_78_Q_reg_10_inst : DFF_X1 port map( D => n5997, CK => CLK
                           , Q => n_2574, QN => 
                           DataPath_RF_bus_reg_dataout_2250_port);
   DataPath_RF_BLOCKi_79_Q_reg_10_inst : DFF_X1 port map( D => n6033, CK => CLK
                           , Q => n_2575, QN => 
                           DataPath_RF_bus_reg_dataout_2282_port);
   DataPath_RF_BLOCKi_80_Q_reg_10_inst : DFF_X1 port map( D => n6070, CK => CLK
                           , Q => n_2576, QN => 
                           DataPath_RF_bus_reg_dataout_2314_port);
   DataPath_RF_BLOCKi_81_Q_reg_10_inst : DFF_X1 port map( D => n6106, CK => CLK
                           , Q => n_2577, QN => 
                           DataPath_RF_bus_reg_dataout_2346_port);
   DataPath_REG_ALU_OUT_Q_reg_11_inst : DFF_X1 port map( D => n7012, CK => CLK,
                           Q => DRAM_ADDRESS_11_port, QN => n500);
   DataPath_REG_MEM_ALUOUT_Q_reg_11_inst : DFF_X1 port map( D => n1138, CK => 
                           CLK, Q => n_2578, QN => 
                           DataPath_i_REG_MEM_ALUOUT_11_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_11_inst : DFF_X1 port map( D => n6788, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_43_port,
                           QN => n610);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_11_inst : DFF_X1 port map( D => n6820, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_75_port,
                           QN => n642);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_11_inst : DFF_X1 port map( D => n6852, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_107_port
                           , QN => n674);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_11_inst : DFF_X1 port map( D => n6884, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_139_port
                           , QN => n706);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_11_inst : DFF_X1 port map( D => n6916, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_171_port
                           , QN => n738);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_11_inst : DFF_X1 port map( D => n6948, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_203_port
                           , QN => n770);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_11_inst : DFF_X1 port map( D => n6980, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_235_port
                           , QN => n802);
   DataPath_RF_BLOCKi_8_Q_reg_11_inst : DFF_X1 port map( D => n3350, CK => CLK,
                           Q => n_2579, QN => 
                           DataPath_RF_bus_reg_dataout_11_port);
   DataPath_RF_BLOCKi_9_Q_reg_11_inst : DFF_X1 port map( D => n3401, CK => CLK,
                           Q => n_2580, QN => 
                           DataPath_RF_bus_reg_dataout_43_port);
   DataPath_RF_BLOCKi_10_Q_reg_11_inst : DFF_X1 port map( D => n3439, CK => CLK
                           , Q => n_2581, QN => 
                           DataPath_RF_bus_reg_dataout_75_port);
   DataPath_RF_BLOCKi_11_Q_reg_11_inst : DFF_X1 port map( D => n3477, CK => CLK
                           , Q => n_2582, QN => 
                           DataPath_RF_bus_reg_dataout_107_port);
   DataPath_RF_BLOCKi_12_Q_reg_11_inst : DFF_X1 port map( D => n3515, CK => CLK
                           , Q => n_2583, QN => 
                           DataPath_RF_bus_reg_dataout_139_port);
   DataPath_RF_BLOCKi_13_Q_reg_11_inst : DFF_X1 port map( D => n3553, CK => CLK
                           , Q => n_2584, QN => 
                           DataPath_RF_bus_reg_dataout_171_port);
   DataPath_RF_BLOCKi_14_Q_reg_11_inst : DFF_X1 port map( D => n3591, CK => CLK
                           , Q => n_2585, QN => 
                           DataPath_RF_bus_reg_dataout_203_port);
   DataPath_RF_BLOCKi_15_Q_reg_11_inst : DFF_X1 port map( D => n3629, CK => CLK
                           , Q => n_2586, QN => 
                           DataPath_RF_bus_reg_dataout_235_port);
   DataPath_RF_BLOCKi_16_Q_reg_11_inst : DFF_X1 port map( D => n3667, CK => CLK
                           , Q => n_2587, QN => 
                           DataPath_RF_bus_reg_dataout_267_port);
   DataPath_RF_BLOCKi_17_Q_reg_11_inst : DFF_X1 port map( D => n3704, CK => CLK
                           , Q => n_2588, QN => 
                           DataPath_RF_bus_reg_dataout_299_port);
   DataPath_RF_BLOCKi_18_Q_reg_11_inst : DFF_X1 port map( D => n3741, CK => CLK
                           , Q => n_2589, QN => 
                           DataPath_RF_bus_reg_dataout_331_port);
   DataPath_RF_BLOCKi_19_Q_reg_11_inst : DFF_X1 port map( D => n3778, CK => CLK
                           , Q => n_2590, QN => 
                           DataPath_RF_bus_reg_dataout_363_port);
   DataPath_RF_BLOCKi_20_Q_reg_11_inst : DFF_X1 port map( D => n3813, CK => CLK
                           , Q => n_2591, QN => 
                           DataPath_RF_bus_reg_dataout_395_port);
   DataPath_RF_BLOCKi_21_Q_reg_11_inst : DFF_X1 port map( D => n3848, CK => CLK
                           , Q => n_2592, QN => 
                           DataPath_RF_bus_reg_dataout_427_port);
   DataPath_RF_BLOCKi_22_Q_reg_11_inst : DFF_X1 port map( D => n3883, CK => CLK
                           , Q => n_2593, QN => 
                           DataPath_RF_bus_reg_dataout_459_port);
   DataPath_RF_BLOCKi_23_Q_reg_11_inst : DFF_X1 port map( D => n3938, CK => CLK
                           , Q => n_2594, QN => 
                           DataPath_RF_bus_reg_dataout_491_port);
   DataPath_RF_BLOCKi_24_Q_reg_11_inst : DFF_X1 port map( D => n4006, CK => CLK
                           , Q => n_2595, QN => 
                           DataPath_RF_bus_reg_dataout_523_port);
   DataPath_RF_BLOCKi_25_Q_reg_11_inst : DFF_X1 port map( D => n4054, CK => CLK
                           , Q => n_2596, QN => 
                           DataPath_RF_bus_reg_dataout_555_port);
   DataPath_RF_BLOCKi_26_Q_reg_11_inst : DFF_X1 port map( D => n4089, CK => CLK
                           , Q => n_2597, QN => 
                           DataPath_RF_bus_reg_dataout_587_port);
   DataPath_RF_BLOCKi_27_Q_reg_11_inst : DFF_X1 port map( D => n4124, CK => CLK
                           , Q => n_2598, QN => 
                           DataPath_RF_bus_reg_dataout_619_port);
   DataPath_RF_BLOCKi_28_Q_reg_11_inst : DFF_X1 port map( D => n4159, CK => CLK
                           , Q => n_2599, QN => 
                           DataPath_RF_bus_reg_dataout_651_port);
   DataPath_RF_BLOCKi_29_Q_reg_11_inst : DFF_X1 port map( D => n4194, CK => CLK
                           , Q => n_2600, QN => 
                           DataPath_RF_bus_reg_dataout_683_port);
   DataPath_RF_BLOCKi_30_Q_reg_11_inst : DFF_X1 port map( D => n4229, CK => CLK
                           , Q => n_2601, QN => 
                           DataPath_RF_bus_reg_dataout_715_port);
   DataPath_RF_BLOCKi_31_Q_reg_11_inst : DFF_X1 port map( D => n4264, CK => CLK
                           , Q => n_2602, QN => 
                           DataPath_RF_bus_reg_dataout_747_port);
   DataPath_RF_BLOCKi_32_Q_reg_11_inst : DFF_X1 port map( D => n4299, CK => CLK
                           , Q => n_2603, QN => 
                           DataPath_RF_bus_reg_dataout_779_port);
   DataPath_RF_BLOCKi_33_Q_reg_11_inst : DFF_X1 port map( D => n4334, CK => CLK
                           , Q => n_2604, QN => 
                           DataPath_RF_bus_reg_dataout_811_port);
   DataPath_RF_BLOCKi_34_Q_reg_11_inst : DFF_X1 port map( D => n4369, CK => CLK
                           , Q => n_2605, QN => 
                           DataPath_RF_bus_reg_dataout_843_port);
   DataPath_RF_BLOCKi_35_Q_reg_11_inst : DFF_X1 port map( D => n4404, CK => CLK
                           , Q => n_2606, QN => 
                           DataPath_RF_bus_reg_dataout_875_port);
   DataPath_RF_BLOCKi_36_Q_reg_11_inst : DFF_X1 port map( D => n4439, CK => CLK
                           , Q => n_2607, QN => 
                           DataPath_RF_bus_reg_dataout_907_port);
   DataPath_RF_BLOCKi_37_Q_reg_11_inst : DFF_X1 port map( D => n4474, CK => CLK
                           , Q => n_2608, QN => 
                           DataPath_RF_bus_reg_dataout_939_port);
   DataPath_RF_BLOCKi_38_Q_reg_11_inst : DFF_X1 port map( D => n4509, CK => CLK
                           , Q => n_2609, QN => 
                           DataPath_RF_bus_reg_dataout_971_port);
   DataPath_RF_BLOCKi_39_Q_reg_11_inst : DFF_X1 port map( D => n4544, CK => CLK
                           , Q => n_2610, QN => 
                           DataPath_RF_bus_reg_dataout_1003_port);
   DataPath_RF_BLOCKi_40_Q_reg_11_inst : DFF_X1 port map( D => n4599, CK => CLK
                           , Q => n_2611, QN => 
                           DataPath_RF_bus_reg_dataout_1035_port);
   DataPath_RF_BLOCKi_41_Q_reg_11_inst : DFF_X1 port map( D => n4647, CK => CLK
                           , Q => n_2612, QN => 
                           DataPath_RF_bus_reg_dataout_1067_port);
   DataPath_RF_BLOCKi_42_Q_reg_11_inst : DFF_X1 port map( D => n4682, CK => CLK
                           , Q => n_2613, QN => 
                           DataPath_RF_bus_reg_dataout_1099_port);
   DataPath_RF_BLOCKi_43_Q_reg_11_inst : DFF_X1 port map( D => n4717, CK => CLK
                           , Q => n_2614, QN => 
                           DataPath_RF_bus_reg_dataout_1131_port);
   DataPath_RF_BLOCKi_44_Q_reg_11_inst : DFF_X1 port map( D => n4752, CK => CLK
                           , Q => n_2615, QN => 
                           DataPath_RF_bus_reg_dataout_1163_port);
   DataPath_RF_BLOCKi_45_Q_reg_11_inst : DFF_X1 port map( D => n4787, CK => CLK
                           , Q => n_2616, QN => 
                           DataPath_RF_bus_reg_dataout_1195_port);
   DataPath_RF_BLOCKi_46_Q_reg_11_inst : DFF_X1 port map( D => n4822, CK => CLK
                           , Q => n_2617, QN => 
                           DataPath_RF_bus_reg_dataout_1227_port);
   DataPath_RF_BLOCKi_47_Q_reg_11_inst : DFF_X1 port map( D => n4857, CK => CLK
                           , Q => n_2618, QN => 
                           DataPath_RF_bus_reg_dataout_1259_port);
   DataPath_RF_BLOCKi_48_Q_reg_11_inst : DFF_X1 port map( D => n4892, CK => CLK
                           , Q => n_2619, QN => 
                           DataPath_RF_bus_reg_dataout_1291_port);
   DataPath_RF_BLOCKi_49_Q_reg_11_inst : DFF_X1 port map( D => n4927, CK => CLK
                           , Q => n_2620, QN => 
                           DataPath_RF_bus_reg_dataout_1323_port);
   DataPath_RF_BLOCKi_50_Q_reg_11_inst : DFF_X1 port map( D => n4962, CK => CLK
                           , Q => n_2621, QN => 
                           DataPath_RF_bus_reg_dataout_1355_port);
   DataPath_RF_BLOCKi_51_Q_reg_11_inst : DFF_X1 port map( D => n4997, CK => CLK
                           , Q => n_2622, QN => 
                           DataPath_RF_bus_reg_dataout_1387_port);
   DataPath_RF_BLOCKi_52_Q_reg_11_inst : DFF_X1 port map( D => n5032, CK => CLK
                           , Q => n_2623, QN => 
                           DataPath_RF_bus_reg_dataout_1419_port);
   DataPath_RF_BLOCKi_53_Q_reg_11_inst : DFF_X1 port map( D => n5067, CK => CLK
                           , Q => n_2624, QN => 
                           DataPath_RF_bus_reg_dataout_1451_port);
   DataPath_RF_BLOCKi_54_Q_reg_11_inst : DFF_X1 port map( D => n5102, CK => CLK
                           , Q => n_2625, QN => 
                           DataPath_RF_bus_reg_dataout_1483_port);
   DataPath_RF_BLOCKi_55_Q_reg_11_inst : DFF_X1 port map( D => n5137, CK => CLK
                           , Q => n_2626, QN => 
                           DataPath_RF_bus_reg_dataout_1515_port);
   DataPath_RF_BLOCKi_56_Q_reg_11_inst : DFF_X1 port map( D => n5192, CK => CLK
                           , Q => n_2627, QN => 
                           DataPath_RF_bus_reg_dataout_1547_port);
   DataPath_RF_BLOCKi_57_Q_reg_11_inst : DFF_X1 port map( D => n5239, CK => CLK
                           , Q => n_2628, QN => 
                           DataPath_RF_bus_reg_dataout_1579_port);
   DataPath_RF_BLOCKi_58_Q_reg_11_inst : DFF_X1 port map( D => n5275, CK => CLK
                           , Q => n_2629, QN => 
                           DataPath_RF_bus_reg_dataout_1611_port);
   DataPath_RF_BLOCKi_59_Q_reg_11_inst : DFF_X1 port map( D => n5310, CK => CLK
                           , Q => n_2630, QN => 
                           DataPath_RF_bus_reg_dataout_1643_port);
   DataPath_RF_BLOCKi_60_Q_reg_11_inst : DFF_X1 port map( D => n5345, CK => CLK
                           , Q => n_2631, QN => 
                           DataPath_RF_bus_reg_dataout_1675_port);
   DataPath_RF_BLOCKi_61_Q_reg_11_inst : DFF_X1 port map( D => n5380, CK => CLK
                           , Q => n_2632, QN => 
                           DataPath_RF_bus_reg_dataout_1707_port);
   DataPath_RF_BLOCKi_62_Q_reg_11_inst : DFF_X1 port map( D => n5415, CK => CLK
                           , Q => n_2633, QN => 
                           DataPath_RF_bus_reg_dataout_1739_port);
   DataPath_RF_BLOCKi_63_Q_reg_11_inst : DFF_X1 port map( D => n5450, CK => CLK
                           , Q => n_2634, QN => 
                           DataPath_RF_bus_reg_dataout_1771_port);
   DataPath_RF_BLOCKi_64_Q_reg_11_inst : DFF_X1 port map( D => n5485, CK => CLK
                           , Q => n_2635, QN => 
                           DataPath_RF_bus_reg_dataout_1803_port);
   DataPath_RF_BLOCKi_65_Q_reg_11_inst : DFF_X1 port map( D => n5520, CK => CLK
                           , Q => n_2636, QN => 
                           DataPath_RF_bus_reg_dataout_1835_port);
   DataPath_RF_BLOCKi_66_Q_reg_11_inst : DFF_X1 port map( D => n5555, CK => CLK
                           , Q => n_2637, QN => 
                           DataPath_RF_bus_reg_dataout_1867_port);
   DataPath_RF_BLOCKi_67_Q_reg_11_inst : DFF_X1 port map( D => n5590, CK => CLK
                           , Q => n_2638, QN => 
                           DataPath_RF_bus_reg_dataout_1899_port);
   DataPath_RF_BLOCKi_68_Q_reg_11_inst : DFF_X1 port map( D => n5629, CK => CLK
                           , Q => n_2639, QN => 
                           DataPath_RF_bus_reg_dataout_1931_port);
   DataPath_RF_BLOCKi_69_Q_reg_11_inst : DFF_X1 port map( D => n5666, CK => CLK
                           , Q => n_2640, QN => 
                           DataPath_RF_bus_reg_dataout_1963_port);
   DataPath_RF_BLOCKi_70_Q_reg_11_inst : DFF_X1 port map( D => n5703, CK => CLK
                           , Q => n_2641, QN => 
                           DataPath_RF_bus_reg_dataout_1995_port);
   DataPath_RF_BLOCKi_71_Q_reg_11_inst : DFF_X1 port map( D => n5740, CK => CLK
                           , Q => n_2642, QN => 
                           DataPath_RF_bus_reg_dataout_2027_port);
   DataPath_RF_BLOCKi_82_Q_reg_11_inst : DFF_X1 port map( D => n890, CK => CLK,
                           Q => n_2643, QN => 
                           DataPath_RF_bus_reg_dataout_2379_port);
   DataPath_RF_BLOCKi_83_Q_reg_11_inst : DFF_X1 port map( D => n952, CK => CLK,
                           Q => n_2644, QN => 
                           DataPath_RF_bus_reg_dataout_2411_port);
   DataPath_RF_BLOCKi_84_Q_reg_11_inst : DFF_X1 port map( D => n990, CK => CLK,
                           Q => n_2645, QN => 
                           DataPath_RF_bus_reg_dataout_2443_port);
   DataPath_RF_BLOCKi_85_Q_reg_11_inst : DFF_X1 port map( D => n1027, CK => CLK
                           , Q => n_2646, QN => 
                           DataPath_RF_bus_reg_dataout_2475_port);
   DataPath_RF_BLOCKi_86_Q_reg_11_inst : DFF_X1 port map( D => n1064, CK => CLK
                           , Q => n_2647, QN => 
                           DataPath_RF_bus_reg_dataout_2507_port);
   DataPath_RF_BLOCKi_87_Q_reg_11_inst : DFF_X1 port map( D => n1101, CK => CLK
                           , Q => n_2648, QN => 
                           DataPath_RF_bus_reg_dataout_2539_port);
   DataPath_RF_BLOCKi_72_Q_reg_11_inst : DFF_X1 port map( D => n5777, CK => CLK
                           , Q => n_2649, QN => 
                           DataPath_RF_bus_reg_dataout_2059_port);
   DataPath_RF_BLOCKi_73_Q_reg_11_inst : DFF_X1 port map( D => n5816, CK => CLK
                           , Q => n_2650, QN => 
                           DataPath_RF_bus_reg_dataout_2091_port);
   DataPath_RF_BLOCKi_74_Q_reg_11_inst : DFF_X1 port map( D => n5852, CK => CLK
                           , Q => n_2651, QN => 
                           DataPath_RF_bus_reg_dataout_2123_port);
   DataPath_RF_BLOCKi_75_Q_reg_11_inst : DFF_X1 port map( D => n5888, CK => CLK
                           , Q => n_2652, QN => 
                           DataPath_RF_bus_reg_dataout_2155_port);
   DataPath_RF_BLOCKi_76_Q_reg_11_inst : DFF_X1 port map( D => n5924, CK => CLK
                           , Q => n_2653, QN => 
                           DataPath_RF_bus_reg_dataout_2187_port);
   DataPath_RF_BLOCKi_77_Q_reg_11_inst : DFF_X1 port map( D => n5960, CK => CLK
                           , Q => n_2654, QN => 
                           DataPath_RF_bus_reg_dataout_2219_port);
   DataPath_RF_BLOCKi_78_Q_reg_11_inst : DFF_X1 port map( D => n5996, CK => CLK
                           , Q => n_2655, QN => 
                           DataPath_RF_bus_reg_dataout_2251_port);
   DataPath_RF_BLOCKi_79_Q_reg_11_inst : DFF_X1 port map( D => n6032, CK => CLK
                           , Q => n_2656, QN => 
                           DataPath_RF_bus_reg_dataout_2283_port);
   DataPath_RF_BLOCKi_80_Q_reg_11_inst : DFF_X1 port map( D => n6069, CK => CLK
                           , Q => n_2657, QN => 
                           DataPath_RF_bus_reg_dataout_2315_port);
   DataPath_RF_BLOCKi_81_Q_reg_11_inst : DFF_X1 port map( D => n6105, CK => CLK
                           , Q => n_2658, QN => 
                           DataPath_RF_bus_reg_dataout_2347_port);
   DataPath_REG_ALU_OUT_Q_reg_12_inst : DFF_X1 port map( D => n7011, CK => CLK,
                           Q => DRAM_ADDRESS_12_port, QN => n501);
   DataPath_REG_MEM_ALUOUT_Q_reg_12_inst : DFF_X1 port map( D => n1137, CK => 
                           CLK, Q => n_2659, QN => 
                           DataPath_i_REG_MEM_ALUOUT_12_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_12_inst : DFF_X1 port map( D => n6787, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_44_port,
                           QN => n611);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_12_inst : DFF_X1 port map( D => n6819, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_76_port,
                           QN => n643);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_12_inst : DFF_X1 port map( D => n6851, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_108_port
                           , QN => n675);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_12_inst : DFF_X1 port map( D => n6883, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_140_port
                           , QN => n707);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_12_inst : DFF_X1 port map( D => n6915, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_172_port
                           , QN => n739);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_12_inst : DFF_X1 port map( D => n6947, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_204_port
                           , QN => n771);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_12_inst : DFF_X1 port map( D => n6979, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_236_port
                           , QN => n803);
   DataPath_RF_BLOCKi_8_Q_reg_12_inst : DFF_X1 port map( D => n3348, CK => CLK,
                           Q => n_2660, QN => 
                           DataPath_RF_bus_reg_dataout_12_port);
   DataPath_RF_BLOCKi_9_Q_reg_12_inst : DFF_X1 port map( D => n3400, CK => CLK,
                           Q => n_2661, QN => 
                           DataPath_RF_bus_reg_dataout_44_port);
   DataPath_RF_BLOCKi_10_Q_reg_12_inst : DFF_X1 port map( D => n3438, CK => CLK
                           , Q => n_2662, QN => 
                           DataPath_RF_bus_reg_dataout_76_port);
   DataPath_RF_BLOCKi_11_Q_reg_12_inst : DFF_X1 port map( D => n3476, CK => CLK
                           , Q => n_2663, QN => 
                           DataPath_RF_bus_reg_dataout_108_port);
   DataPath_RF_BLOCKi_12_Q_reg_12_inst : DFF_X1 port map( D => n3514, CK => CLK
                           , Q => n_2664, QN => 
                           DataPath_RF_bus_reg_dataout_140_port);
   DataPath_RF_BLOCKi_13_Q_reg_12_inst : DFF_X1 port map( D => n3552, CK => CLK
                           , Q => n_2665, QN => 
                           DataPath_RF_bus_reg_dataout_172_port);
   DataPath_RF_BLOCKi_14_Q_reg_12_inst : DFF_X1 port map( D => n3590, CK => CLK
                           , Q => n_2666, QN => 
                           DataPath_RF_bus_reg_dataout_204_port);
   DataPath_RF_BLOCKi_15_Q_reg_12_inst : DFF_X1 port map( D => n3628, CK => CLK
                           , Q => n_2667, QN => 
                           DataPath_RF_bus_reg_dataout_236_port);
   DataPath_RF_BLOCKi_16_Q_reg_12_inst : DFF_X1 port map( D => n3666, CK => CLK
                           , Q => n_2668, QN => 
                           DataPath_RF_bus_reg_dataout_268_port);
   DataPath_RF_BLOCKi_17_Q_reg_12_inst : DFF_X1 port map( D => n3703, CK => CLK
                           , Q => n_2669, QN => 
                           DataPath_RF_bus_reg_dataout_300_port);
   DataPath_RF_BLOCKi_18_Q_reg_12_inst : DFF_X1 port map( D => n3740, CK => CLK
                           , Q => n_2670, QN => 
                           DataPath_RF_bus_reg_dataout_332_port);
   DataPath_RF_BLOCKi_19_Q_reg_12_inst : DFF_X1 port map( D => n3777, CK => CLK
                           , Q => n_2671, QN => 
                           DataPath_RF_bus_reg_dataout_364_port);
   DataPath_RF_BLOCKi_20_Q_reg_12_inst : DFF_X1 port map( D => n3812, CK => CLK
                           , Q => n_2672, QN => 
                           DataPath_RF_bus_reg_dataout_396_port);
   DataPath_RF_BLOCKi_21_Q_reg_12_inst : DFF_X1 port map( D => n3847, CK => CLK
                           , Q => n_2673, QN => 
                           DataPath_RF_bus_reg_dataout_428_port);
   DataPath_RF_BLOCKi_22_Q_reg_12_inst : DFF_X1 port map( D => n3882, CK => CLK
                           , Q => n_2674, QN => 
                           DataPath_RF_bus_reg_dataout_460_port);
   DataPath_RF_BLOCKi_23_Q_reg_12_inst : DFF_X1 port map( D => n3936, CK => CLK
                           , Q => n_2675, QN => 
                           DataPath_RF_bus_reg_dataout_492_port);
   DataPath_RF_BLOCKi_24_Q_reg_12_inst : DFF_X1 port map( D => n4004, CK => CLK
                           , Q => n_2676, QN => 
                           DataPath_RF_bus_reg_dataout_524_port);
   DataPath_RF_BLOCKi_25_Q_reg_12_inst : DFF_X1 port map( D => n4053, CK => CLK
                           , Q => n_2677, QN => 
                           DataPath_RF_bus_reg_dataout_556_port);
   DataPath_RF_BLOCKi_26_Q_reg_12_inst : DFF_X1 port map( D => n4088, CK => CLK
                           , Q => n_2678, QN => 
                           DataPath_RF_bus_reg_dataout_588_port);
   DataPath_RF_BLOCKi_27_Q_reg_12_inst : DFF_X1 port map( D => n4123, CK => CLK
                           , Q => n_2679, QN => 
                           DataPath_RF_bus_reg_dataout_620_port);
   DataPath_RF_BLOCKi_28_Q_reg_12_inst : DFF_X1 port map( D => n4158, CK => CLK
                           , Q => n_2680, QN => 
                           DataPath_RF_bus_reg_dataout_652_port);
   DataPath_RF_BLOCKi_29_Q_reg_12_inst : DFF_X1 port map( D => n4193, CK => CLK
                           , Q => n_2681, QN => 
                           DataPath_RF_bus_reg_dataout_684_port);
   DataPath_RF_BLOCKi_30_Q_reg_12_inst : DFF_X1 port map( D => n4228, CK => CLK
                           , Q => n_2682, QN => 
                           DataPath_RF_bus_reg_dataout_716_port);
   DataPath_RF_BLOCKi_31_Q_reg_12_inst : DFF_X1 port map( D => n4263, CK => CLK
                           , Q => n_2683, QN => 
                           DataPath_RF_bus_reg_dataout_748_port);
   DataPath_RF_BLOCKi_32_Q_reg_12_inst : DFF_X1 port map( D => n4298, CK => CLK
                           , Q => n_2684, QN => 
                           DataPath_RF_bus_reg_dataout_780_port);
   DataPath_RF_BLOCKi_33_Q_reg_12_inst : DFF_X1 port map( D => n4333, CK => CLK
                           , Q => n_2685, QN => 
                           DataPath_RF_bus_reg_dataout_812_port);
   DataPath_RF_BLOCKi_34_Q_reg_12_inst : DFF_X1 port map( D => n4368, CK => CLK
                           , Q => n_2686, QN => 
                           DataPath_RF_bus_reg_dataout_844_port);
   DataPath_RF_BLOCKi_35_Q_reg_12_inst : DFF_X1 port map( D => n4403, CK => CLK
                           , Q => n_2687, QN => 
                           DataPath_RF_bus_reg_dataout_876_port);
   DataPath_RF_BLOCKi_36_Q_reg_12_inst : DFF_X1 port map( D => n4438, CK => CLK
                           , Q => n_2688, QN => 
                           DataPath_RF_bus_reg_dataout_908_port);
   DataPath_RF_BLOCKi_37_Q_reg_12_inst : DFF_X1 port map( D => n4473, CK => CLK
                           , Q => n_2689, QN => 
                           DataPath_RF_bus_reg_dataout_940_port);
   DataPath_RF_BLOCKi_38_Q_reg_12_inst : DFF_X1 port map( D => n4508, CK => CLK
                           , Q => n_2690, QN => 
                           DataPath_RF_bus_reg_dataout_972_port);
   DataPath_RF_BLOCKi_39_Q_reg_12_inst : DFF_X1 port map( D => n4543, CK => CLK
                           , Q => n_2691, QN => 
                           DataPath_RF_bus_reg_dataout_1004_port);
   DataPath_RF_BLOCKi_40_Q_reg_12_inst : DFF_X1 port map( D => n4597, CK => CLK
                           , Q => n_2692, QN => 
                           DataPath_RF_bus_reg_dataout_1036_port);
   DataPath_RF_BLOCKi_41_Q_reg_12_inst : DFF_X1 port map( D => n4646, CK => CLK
                           , Q => n_2693, QN => 
                           DataPath_RF_bus_reg_dataout_1068_port);
   DataPath_RF_BLOCKi_42_Q_reg_12_inst : DFF_X1 port map( D => n4681, CK => CLK
                           , Q => n_2694, QN => 
                           DataPath_RF_bus_reg_dataout_1100_port);
   DataPath_RF_BLOCKi_43_Q_reg_12_inst : DFF_X1 port map( D => n4716, CK => CLK
                           , Q => n_2695, QN => 
                           DataPath_RF_bus_reg_dataout_1132_port);
   DataPath_RF_BLOCKi_44_Q_reg_12_inst : DFF_X1 port map( D => n4751, CK => CLK
                           , Q => n_2696, QN => 
                           DataPath_RF_bus_reg_dataout_1164_port);
   DataPath_RF_BLOCKi_45_Q_reg_12_inst : DFF_X1 port map( D => n4786, CK => CLK
                           , Q => n_2697, QN => 
                           DataPath_RF_bus_reg_dataout_1196_port);
   DataPath_RF_BLOCKi_46_Q_reg_12_inst : DFF_X1 port map( D => n4821, CK => CLK
                           , Q => n_2698, QN => 
                           DataPath_RF_bus_reg_dataout_1228_port);
   DataPath_RF_BLOCKi_47_Q_reg_12_inst : DFF_X1 port map( D => n4856, CK => CLK
                           , Q => n_2699, QN => 
                           DataPath_RF_bus_reg_dataout_1260_port);
   DataPath_RF_BLOCKi_48_Q_reg_12_inst : DFF_X1 port map( D => n4891, CK => CLK
                           , Q => n_2700, QN => 
                           DataPath_RF_bus_reg_dataout_1292_port);
   DataPath_RF_BLOCKi_49_Q_reg_12_inst : DFF_X1 port map( D => n4926, CK => CLK
                           , Q => n_2701, QN => 
                           DataPath_RF_bus_reg_dataout_1324_port);
   DataPath_RF_BLOCKi_50_Q_reg_12_inst : DFF_X1 port map( D => n4961, CK => CLK
                           , Q => n_2702, QN => 
                           DataPath_RF_bus_reg_dataout_1356_port);
   DataPath_RF_BLOCKi_51_Q_reg_12_inst : DFF_X1 port map( D => n4996, CK => CLK
                           , Q => n_2703, QN => 
                           DataPath_RF_bus_reg_dataout_1388_port);
   DataPath_RF_BLOCKi_52_Q_reg_12_inst : DFF_X1 port map( D => n5031, CK => CLK
                           , Q => n_2704, QN => 
                           DataPath_RF_bus_reg_dataout_1420_port);
   DataPath_RF_BLOCKi_53_Q_reg_12_inst : DFF_X1 port map( D => n5066, CK => CLK
                           , Q => n_2705, QN => 
                           DataPath_RF_bus_reg_dataout_1452_port);
   DataPath_RF_BLOCKi_54_Q_reg_12_inst : DFF_X1 port map( D => n5101, CK => CLK
                           , Q => n_2706, QN => 
                           DataPath_RF_bus_reg_dataout_1484_port);
   DataPath_RF_BLOCKi_55_Q_reg_12_inst : DFF_X1 port map( D => n5136, CK => CLK
                           , Q => n_2707, QN => 
                           DataPath_RF_bus_reg_dataout_1516_port);
   DataPath_RF_BLOCKi_56_Q_reg_12_inst : DFF_X1 port map( D => n5190, CK => CLK
                           , Q => n_2708, QN => 
                           DataPath_RF_bus_reg_dataout_1548_port);
   DataPath_RF_BLOCKi_57_Q_reg_12_inst : DFF_X1 port map( D => n5238, CK => CLK
                           , Q => n_2709, QN => 
                           DataPath_RF_bus_reg_dataout_1580_port);
   DataPath_RF_BLOCKi_58_Q_reg_12_inst : DFF_X1 port map( D => n5274, CK => CLK
                           , Q => n_2710, QN => 
                           DataPath_RF_bus_reg_dataout_1612_port);
   DataPath_RF_BLOCKi_59_Q_reg_12_inst : DFF_X1 port map( D => n5309, CK => CLK
                           , Q => n_2711, QN => 
                           DataPath_RF_bus_reg_dataout_1644_port);
   DataPath_RF_BLOCKi_60_Q_reg_12_inst : DFF_X1 port map( D => n5344, CK => CLK
                           , Q => n_2712, QN => 
                           DataPath_RF_bus_reg_dataout_1676_port);
   DataPath_RF_BLOCKi_61_Q_reg_12_inst : DFF_X1 port map( D => n5379, CK => CLK
                           , Q => n_2713, QN => 
                           DataPath_RF_bus_reg_dataout_1708_port);
   DataPath_RF_BLOCKi_62_Q_reg_12_inst : DFF_X1 port map( D => n5414, CK => CLK
                           , Q => n_2714, QN => 
                           DataPath_RF_bus_reg_dataout_1740_port);
   DataPath_RF_BLOCKi_63_Q_reg_12_inst : DFF_X1 port map( D => n5449, CK => CLK
                           , Q => n_2715, QN => 
                           DataPath_RF_bus_reg_dataout_1772_port);
   DataPath_RF_BLOCKi_64_Q_reg_12_inst : DFF_X1 port map( D => n5484, CK => CLK
                           , Q => n_2716, QN => 
                           DataPath_RF_bus_reg_dataout_1804_port);
   DataPath_RF_BLOCKi_65_Q_reg_12_inst : DFF_X1 port map( D => n5519, CK => CLK
                           , Q => n_2717, QN => 
                           DataPath_RF_bus_reg_dataout_1836_port);
   DataPath_RF_BLOCKi_66_Q_reg_12_inst : DFF_X1 port map( D => n5554, CK => CLK
                           , Q => n_2718, QN => 
                           DataPath_RF_bus_reg_dataout_1868_port);
   DataPath_RF_BLOCKi_67_Q_reg_12_inst : DFF_X1 port map( D => n5589, CK => CLK
                           , Q => n_2719, QN => 
                           DataPath_RF_bus_reg_dataout_1900_port);
   DataPath_RF_BLOCKi_68_Q_reg_12_inst : DFF_X1 port map( D => n5628, CK => CLK
                           , Q => n_2720, QN => 
                           DataPath_RF_bus_reg_dataout_1932_port);
   DataPath_RF_BLOCKi_69_Q_reg_12_inst : DFF_X1 port map( D => n5665, CK => CLK
                           , Q => n_2721, QN => 
                           DataPath_RF_bus_reg_dataout_1964_port);
   DataPath_RF_BLOCKi_70_Q_reg_12_inst : DFF_X1 port map( D => n5702, CK => CLK
                           , Q => n_2722, QN => 
                           DataPath_RF_bus_reg_dataout_1996_port);
   DataPath_RF_BLOCKi_71_Q_reg_12_inst : DFF_X1 port map( D => n5739, CK => CLK
                           , Q => n_2723, QN => 
                           DataPath_RF_bus_reg_dataout_2028_port);
   DataPath_RF_BLOCKi_82_Q_reg_12_inst : DFF_X1 port map( D => n888, CK => CLK,
                           Q => n_2724, QN => 
                           DataPath_RF_bus_reg_dataout_2380_port);
   DataPath_RF_BLOCKi_83_Q_reg_12_inst : DFF_X1 port map( D => n951, CK => CLK,
                           Q => n_2725, QN => 
                           DataPath_RF_bus_reg_dataout_2412_port);
   DataPath_RF_BLOCKi_84_Q_reg_12_inst : DFF_X1 port map( D => n989, CK => CLK,
                           Q => n_2726, QN => 
                           DataPath_RF_bus_reg_dataout_2444_port);
   DataPath_RF_BLOCKi_85_Q_reg_12_inst : DFF_X1 port map( D => n1026, CK => CLK
                           , Q => n_2727, QN => 
                           DataPath_RF_bus_reg_dataout_2476_port);
   DataPath_RF_BLOCKi_86_Q_reg_12_inst : DFF_X1 port map( D => n1063, CK => CLK
                           , Q => n_2728, QN => 
                           DataPath_RF_bus_reg_dataout_2508_port);
   DataPath_RF_BLOCKi_87_Q_reg_12_inst : DFF_X1 port map( D => n1100, CK => CLK
                           , Q => n_2729, QN => 
                           DataPath_RF_bus_reg_dataout_2540_port);
   DataPath_RF_BLOCKi_72_Q_reg_12_inst : DFF_X1 port map( D => n5776, CK => CLK
                           , Q => n_2730, QN => 
                           DataPath_RF_bus_reg_dataout_2060_port);
   DataPath_RF_BLOCKi_73_Q_reg_12_inst : DFF_X1 port map( D => n5815, CK => CLK
                           , Q => n_2731, QN => 
                           DataPath_RF_bus_reg_dataout_2092_port);
   DataPath_RF_BLOCKi_74_Q_reg_12_inst : DFF_X1 port map( D => n5851, CK => CLK
                           , Q => n_2732, QN => 
                           DataPath_RF_bus_reg_dataout_2124_port);
   DataPath_RF_BLOCKi_75_Q_reg_12_inst : DFF_X1 port map( D => n5887, CK => CLK
                           , Q => n_2733, QN => 
                           DataPath_RF_bus_reg_dataout_2156_port);
   DataPath_RF_BLOCKi_76_Q_reg_12_inst : DFF_X1 port map( D => n5923, CK => CLK
                           , Q => n_2734, QN => 
                           DataPath_RF_bus_reg_dataout_2188_port);
   DataPath_RF_BLOCKi_77_Q_reg_12_inst : DFF_X1 port map( D => n5959, CK => CLK
                           , Q => n_2735, QN => 
                           DataPath_RF_bus_reg_dataout_2220_port);
   DataPath_RF_BLOCKi_78_Q_reg_12_inst : DFF_X1 port map( D => n5995, CK => CLK
                           , Q => n_2736, QN => 
                           DataPath_RF_bus_reg_dataout_2252_port);
   DataPath_RF_BLOCKi_79_Q_reg_12_inst : DFF_X1 port map( D => n6031, CK => CLK
                           , Q => n_2737, QN => 
                           DataPath_RF_bus_reg_dataout_2284_port);
   DataPath_RF_BLOCKi_80_Q_reg_12_inst : DFF_X1 port map( D => n6068, CK => CLK
                           , Q => n_2738, QN => 
                           DataPath_RF_bus_reg_dataout_2316_port);
   DataPath_RF_BLOCKi_81_Q_reg_12_inst : DFF_X1 port map( D => n6104, CK => CLK
                           , Q => n_2739, QN => 
                           DataPath_RF_bus_reg_dataout_2348_port);
   DataPath_REG_ALU_OUT_Q_reg_14_inst : DFF_X1 port map( D => n7009, CK => CLK,
                           Q => DRAM_ADDRESS_14_port, QN => n502);
   DataPath_REG_MEM_ALUOUT_Q_reg_14_inst : DFF_X1 port map( D => n1135, CK => 
                           CLK, Q => n_2740, QN => 
                           DataPath_i_REG_MEM_ALUOUT_14_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_14_inst : DFF_X1 port map( D => n6785, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_46_port,
                           QN => n613);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_14_inst : DFF_X1 port map( D => n6817, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_78_port,
                           QN => n645);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_14_inst : DFF_X1 port map( D => n6849, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_110_port
                           , QN => n677);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_14_inst : DFF_X1 port map( D => n6881, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_142_port
                           , QN => n709);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_14_inst : DFF_X1 port map( D => n6913, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_174_port
                           , QN => n741);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_14_inst : DFF_X1 port map( D => n6945, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_206_port
                           , QN => n773);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_14_inst : DFF_X1 port map( D => n6977, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_238_port
                           , QN => n805);
   DataPath_RF_BLOCKi_8_Q_reg_14_inst : DFF_X1 port map( D => n3344, CK => CLK,
                           Q => n_2741, QN => 
                           DataPath_RF_bus_reg_dataout_14_port);
   DataPath_RF_BLOCKi_9_Q_reg_14_inst : DFF_X1 port map( D => n3398, CK => CLK,
                           Q => n_2742, QN => 
                           DataPath_RF_bus_reg_dataout_46_port);
   DataPath_RF_BLOCKi_10_Q_reg_14_inst : DFF_X1 port map( D => n3436, CK => CLK
                           , Q => n_2743, QN => 
                           DataPath_RF_bus_reg_dataout_78_port);
   DataPath_RF_BLOCKi_11_Q_reg_14_inst : DFF_X1 port map( D => n3474, CK => CLK
                           , Q => n_2744, QN => 
                           DataPath_RF_bus_reg_dataout_110_port);
   DataPath_RF_BLOCKi_12_Q_reg_14_inst : DFF_X1 port map( D => n3512, CK => CLK
                           , Q => n_2745, QN => 
                           DataPath_RF_bus_reg_dataout_142_port);
   DataPath_RF_BLOCKi_13_Q_reg_14_inst : DFF_X1 port map( D => n3550, CK => CLK
                           , Q => n_2746, QN => 
                           DataPath_RF_bus_reg_dataout_174_port);
   DataPath_RF_BLOCKi_14_Q_reg_14_inst : DFF_X1 port map( D => n3588, CK => CLK
                           , Q => n_2747, QN => 
                           DataPath_RF_bus_reg_dataout_206_port);
   DataPath_RF_BLOCKi_15_Q_reg_14_inst : DFF_X1 port map( D => n3626, CK => CLK
                           , Q => n_2748, QN => 
                           DataPath_RF_bus_reg_dataout_238_port);
   DataPath_RF_BLOCKi_16_Q_reg_14_inst : DFF_X1 port map( D => n3664, CK => CLK
                           , Q => n_2749, QN => 
                           DataPath_RF_bus_reg_dataout_270_port);
   DataPath_RF_BLOCKi_17_Q_reg_14_inst : DFF_X1 port map( D => n3701, CK => CLK
                           , Q => n_2750, QN => 
                           DataPath_RF_bus_reg_dataout_302_port);
   DataPath_RF_BLOCKi_18_Q_reg_14_inst : DFF_X1 port map( D => n3738, CK => CLK
                           , Q => n_2751, QN => 
                           DataPath_RF_bus_reg_dataout_334_port);
   DataPath_RF_BLOCKi_19_Q_reg_14_inst : DFF_X1 port map( D => n3775, CK => CLK
                           , Q => n_2752, QN => 
                           DataPath_RF_bus_reg_dataout_366_port);
   DataPath_RF_BLOCKi_20_Q_reg_14_inst : DFF_X1 port map( D => n3810, CK => CLK
                           , Q => n_2753, QN => 
                           DataPath_RF_bus_reg_dataout_398_port);
   DataPath_RF_BLOCKi_21_Q_reg_14_inst : DFF_X1 port map( D => n3845, CK => CLK
                           , Q => n_2754, QN => 
                           DataPath_RF_bus_reg_dataout_430_port);
   DataPath_RF_BLOCKi_22_Q_reg_14_inst : DFF_X1 port map( D => n3880, CK => CLK
                           , Q => n_2755, QN => 
                           DataPath_RF_bus_reg_dataout_462_port);
   DataPath_RF_BLOCKi_23_Q_reg_14_inst : DFF_X1 port map( D => n3932, CK => CLK
                           , Q => n_2756, QN => 
                           DataPath_RF_bus_reg_dataout_494_port);
   DataPath_RF_BLOCKi_24_Q_reg_14_inst : DFF_X1 port map( D => n4000, CK => CLK
                           , Q => n_2757, QN => 
                           DataPath_RF_bus_reg_dataout_526_port);
   DataPath_RF_BLOCKi_25_Q_reg_14_inst : DFF_X1 port map( D => n4051, CK => CLK
                           , Q => n_2758, QN => 
                           DataPath_RF_bus_reg_dataout_558_port);
   DataPath_RF_BLOCKi_26_Q_reg_14_inst : DFF_X1 port map( D => n4086, CK => CLK
                           , Q => n_2759, QN => 
                           DataPath_RF_bus_reg_dataout_590_port);
   DataPath_RF_BLOCKi_27_Q_reg_14_inst : DFF_X1 port map( D => n4121, CK => CLK
                           , Q => n_2760, QN => 
                           DataPath_RF_bus_reg_dataout_622_port);
   DataPath_RF_BLOCKi_28_Q_reg_14_inst : DFF_X1 port map( D => n4156, CK => CLK
                           , Q => n_2761, QN => 
                           DataPath_RF_bus_reg_dataout_654_port);
   DataPath_RF_BLOCKi_29_Q_reg_14_inst : DFF_X1 port map( D => n4191, CK => CLK
                           , Q => n_2762, QN => 
                           DataPath_RF_bus_reg_dataout_686_port);
   DataPath_RF_BLOCKi_30_Q_reg_14_inst : DFF_X1 port map( D => n4226, CK => CLK
                           , Q => n_2763, QN => 
                           DataPath_RF_bus_reg_dataout_718_port);
   DataPath_RF_BLOCKi_31_Q_reg_14_inst : DFF_X1 port map( D => n4261, CK => CLK
                           , Q => n_2764, QN => 
                           DataPath_RF_bus_reg_dataout_750_port);
   DataPath_RF_BLOCKi_32_Q_reg_14_inst : DFF_X1 port map( D => n4296, CK => CLK
                           , Q => n_2765, QN => 
                           DataPath_RF_bus_reg_dataout_782_port);
   DataPath_RF_BLOCKi_33_Q_reg_14_inst : DFF_X1 port map( D => n4331, CK => CLK
                           , Q => n_2766, QN => 
                           DataPath_RF_bus_reg_dataout_814_port);
   DataPath_RF_BLOCKi_34_Q_reg_14_inst : DFF_X1 port map( D => n4366, CK => CLK
                           , Q => n_2767, QN => 
                           DataPath_RF_bus_reg_dataout_846_port);
   DataPath_RF_BLOCKi_35_Q_reg_14_inst : DFF_X1 port map( D => n4401, CK => CLK
                           , Q => n_2768, QN => 
                           DataPath_RF_bus_reg_dataout_878_port);
   DataPath_RF_BLOCKi_36_Q_reg_14_inst : DFF_X1 port map( D => n4436, CK => CLK
                           , Q => n_2769, QN => 
                           DataPath_RF_bus_reg_dataout_910_port);
   DataPath_RF_BLOCKi_37_Q_reg_14_inst : DFF_X1 port map( D => n4471, CK => CLK
                           , Q => n_2770, QN => 
                           DataPath_RF_bus_reg_dataout_942_port);
   DataPath_RF_BLOCKi_38_Q_reg_14_inst : DFF_X1 port map( D => n4506, CK => CLK
                           , Q => n_2771, QN => 
                           DataPath_RF_bus_reg_dataout_974_port);
   DataPath_RF_BLOCKi_39_Q_reg_14_inst : DFF_X1 port map( D => n4541, CK => CLK
                           , Q => n_2772, QN => 
                           DataPath_RF_bus_reg_dataout_1006_port);
   DataPath_RF_BLOCKi_40_Q_reg_14_inst : DFF_X1 port map( D => n4593, CK => CLK
                           , Q => n_2773, QN => 
                           DataPath_RF_bus_reg_dataout_1038_port);
   DataPath_RF_BLOCKi_41_Q_reg_14_inst : DFF_X1 port map( D => n4644, CK => CLK
                           , Q => n_2774, QN => 
                           DataPath_RF_bus_reg_dataout_1070_port);
   DataPath_RF_BLOCKi_42_Q_reg_14_inst : DFF_X1 port map( D => n4679, CK => CLK
                           , Q => n_2775, QN => 
                           DataPath_RF_bus_reg_dataout_1102_port);
   DataPath_RF_BLOCKi_43_Q_reg_14_inst : DFF_X1 port map( D => n4714, CK => CLK
                           , Q => n_2776, QN => 
                           DataPath_RF_bus_reg_dataout_1134_port);
   DataPath_RF_BLOCKi_44_Q_reg_14_inst : DFF_X1 port map( D => n4749, CK => CLK
                           , Q => n_2777, QN => 
                           DataPath_RF_bus_reg_dataout_1166_port);
   DataPath_RF_BLOCKi_45_Q_reg_14_inst : DFF_X1 port map( D => n4784, CK => CLK
                           , Q => n_2778, QN => 
                           DataPath_RF_bus_reg_dataout_1198_port);
   DataPath_RF_BLOCKi_46_Q_reg_14_inst : DFF_X1 port map( D => n4819, CK => CLK
                           , Q => n_2779, QN => 
                           DataPath_RF_bus_reg_dataout_1230_port);
   DataPath_RF_BLOCKi_47_Q_reg_14_inst : DFF_X1 port map( D => n4854, CK => CLK
                           , Q => n_2780, QN => 
                           DataPath_RF_bus_reg_dataout_1262_port);
   DataPath_RF_BLOCKi_48_Q_reg_14_inst : DFF_X1 port map( D => n4889, CK => CLK
                           , Q => n_2781, QN => 
                           DataPath_RF_bus_reg_dataout_1294_port);
   DataPath_RF_BLOCKi_49_Q_reg_14_inst : DFF_X1 port map( D => n4924, CK => CLK
                           , Q => n_2782, QN => 
                           DataPath_RF_bus_reg_dataout_1326_port);
   DataPath_RF_BLOCKi_50_Q_reg_14_inst : DFF_X1 port map( D => n4959, CK => CLK
                           , Q => n_2783, QN => 
                           DataPath_RF_bus_reg_dataout_1358_port);
   DataPath_RF_BLOCKi_51_Q_reg_14_inst : DFF_X1 port map( D => n4994, CK => CLK
                           , Q => n_2784, QN => 
                           DataPath_RF_bus_reg_dataout_1390_port);
   DataPath_RF_BLOCKi_52_Q_reg_14_inst : DFF_X1 port map( D => n5029, CK => CLK
                           , Q => n_2785, QN => 
                           DataPath_RF_bus_reg_dataout_1422_port);
   DataPath_RF_BLOCKi_53_Q_reg_14_inst : DFF_X1 port map( D => n5064, CK => CLK
                           , Q => n_2786, QN => 
                           DataPath_RF_bus_reg_dataout_1454_port);
   DataPath_RF_BLOCKi_54_Q_reg_14_inst : DFF_X1 port map( D => n5099, CK => CLK
                           , Q => n_2787, QN => 
                           DataPath_RF_bus_reg_dataout_1486_port);
   DataPath_RF_BLOCKi_55_Q_reg_14_inst : DFF_X1 port map( D => n5134, CK => CLK
                           , Q => n_2788, QN => 
                           DataPath_RF_bus_reg_dataout_1518_port);
   DataPath_RF_BLOCKi_56_Q_reg_14_inst : DFF_X1 port map( D => n5186, CK => CLK
                           , Q => n_2789, QN => 
                           DataPath_RF_bus_reg_dataout_1550_port);
   DataPath_RF_BLOCKi_57_Q_reg_14_inst : DFF_X1 port map( D => n5236, CK => CLK
                           , Q => n_2790, QN => 
                           DataPath_RF_bus_reg_dataout_1582_port);
   DataPath_RF_BLOCKi_58_Q_reg_14_inst : DFF_X1 port map( D => n5272, CK => CLK
                           , Q => n_2791, QN => 
                           DataPath_RF_bus_reg_dataout_1614_port);
   DataPath_RF_BLOCKi_59_Q_reg_14_inst : DFF_X1 port map( D => n5307, CK => CLK
                           , Q => n_2792, QN => 
                           DataPath_RF_bus_reg_dataout_1646_port);
   DataPath_RF_BLOCKi_60_Q_reg_14_inst : DFF_X1 port map( D => n5342, CK => CLK
                           , Q => n_2793, QN => 
                           DataPath_RF_bus_reg_dataout_1678_port);
   DataPath_RF_BLOCKi_61_Q_reg_14_inst : DFF_X1 port map( D => n5377, CK => CLK
                           , Q => n_2794, QN => 
                           DataPath_RF_bus_reg_dataout_1710_port);
   DataPath_RF_BLOCKi_62_Q_reg_14_inst : DFF_X1 port map( D => n5412, CK => CLK
                           , Q => n_2795, QN => 
                           DataPath_RF_bus_reg_dataout_1742_port);
   DataPath_RF_BLOCKi_63_Q_reg_14_inst : DFF_X1 port map( D => n5447, CK => CLK
                           , Q => n_2796, QN => 
                           DataPath_RF_bus_reg_dataout_1774_port);
   DataPath_RF_BLOCKi_64_Q_reg_14_inst : DFF_X1 port map( D => n5482, CK => CLK
                           , Q => n_2797, QN => 
                           DataPath_RF_bus_reg_dataout_1806_port);
   DataPath_RF_BLOCKi_65_Q_reg_14_inst : DFF_X1 port map( D => n5517, CK => CLK
                           , Q => n_2798, QN => 
                           DataPath_RF_bus_reg_dataout_1838_port);
   DataPath_RF_BLOCKi_66_Q_reg_14_inst : DFF_X1 port map( D => n5552, CK => CLK
                           , Q => n_2799, QN => 
                           DataPath_RF_bus_reg_dataout_1870_port);
   DataPath_RF_BLOCKi_67_Q_reg_14_inst : DFF_X1 port map( D => n5587, CK => CLK
                           , Q => n_2800, QN => 
                           DataPath_RF_bus_reg_dataout_1902_port);
   DataPath_RF_BLOCKi_68_Q_reg_14_inst : DFF_X1 port map( D => n5626, CK => CLK
                           , Q => n_2801, QN => 
                           DataPath_RF_bus_reg_dataout_1934_port);
   DataPath_RF_BLOCKi_69_Q_reg_14_inst : DFF_X1 port map( D => n5663, CK => CLK
                           , Q => n_2802, QN => 
                           DataPath_RF_bus_reg_dataout_1966_port);
   DataPath_RF_BLOCKi_70_Q_reg_14_inst : DFF_X1 port map( D => n5700, CK => CLK
                           , Q => n_2803, QN => 
                           DataPath_RF_bus_reg_dataout_1998_port);
   DataPath_RF_BLOCKi_71_Q_reg_14_inst : DFF_X1 port map( D => n5737, CK => CLK
                           , Q => n_2804, QN => 
                           DataPath_RF_bus_reg_dataout_2030_port);
   DataPath_RF_BLOCKi_82_Q_reg_14_inst : DFF_X1 port map( D => n884, CK => CLK,
                           Q => n_2805, QN => 
                           DataPath_RF_bus_reg_dataout_2382_port);
   DataPath_RF_BLOCKi_83_Q_reg_14_inst : DFF_X1 port map( D => n949, CK => CLK,
                           Q => n_2806, QN => 
                           DataPath_RF_bus_reg_dataout_2414_port);
   DataPath_RF_BLOCKi_84_Q_reg_14_inst : DFF_X1 port map( D => n987, CK => CLK,
                           Q => n_2807, QN => 
                           DataPath_RF_bus_reg_dataout_2446_port);
   DataPath_RF_BLOCKi_85_Q_reg_14_inst : DFF_X1 port map( D => n1024, CK => CLK
                           , Q => n_2808, QN => 
                           DataPath_RF_bus_reg_dataout_2478_port);
   DataPath_RF_BLOCKi_86_Q_reg_14_inst : DFF_X1 port map( D => n1061, CK => CLK
                           , Q => n_2809, QN => 
                           DataPath_RF_bus_reg_dataout_2510_port);
   DataPath_RF_BLOCKi_87_Q_reg_14_inst : DFF_X1 port map( D => n1098, CK => CLK
                           , Q => n_2810, QN => 
                           DataPath_RF_bus_reg_dataout_2542_port);
   DataPath_RF_BLOCKi_72_Q_reg_14_inst : DFF_X1 port map( D => n5774, CK => CLK
                           , Q => n_2811, QN => 
                           DataPath_RF_bus_reg_dataout_2062_port);
   DataPath_RF_BLOCKi_73_Q_reg_14_inst : DFF_X1 port map( D => n5813, CK => CLK
                           , Q => n_2812, QN => 
                           DataPath_RF_bus_reg_dataout_2094_port);
   DataPath_RF_BLOCKi_74_Q_reg_14_inst : DFF_X1 port map( D => n5849, CK => CLK
                           , Q => n_2813, QN => 
                           DataPath_RF_bus_reg_dataout_2126_port);
   DataPath_RF_BLOCKi_75_Q_reg_14_inst : DFF_X1 port map( D => n5885, CK => CLK
                           , Q => n_2814, QN => 
                           DataPath_RF_bus_reg_dataout_2158_port);
   DataPath_RF_BLOCKi_76_Q_reg_14_inst : DFF_X1 port map( D => n5921, CK => CLK
                           , Q => n_2815, QN => 
                           DataPath_RF_bus_reg_dataout_2190_port);
   DataPath_RF_BLOCKi_77_Q_reg_14_inst : DFF_X1 port map( D => n5957, CK => CLK
                           , Q => n_2816, QN => 
                           DataPath_RF_bus_reg_dataout_2222_port);
   DataPath_RF_BLOCKi_78_Q_reg_14_inst : DFF_X1 port map( D => n5993, CK => CLK
                           , Q => n_2817, QN => 
                           DataPath_RF_bus_reg_dataout_2254_port);
   DataPath_RF_BLOCKi_79_Q_reg_14_inst : DFF_X1 port map( D => n6029, CK => CLK
                           , Q => n_2818, QN => 
                           DataPath_RF_bus_reg_dataout_2286_port);
   DataPath_RF_BLOCKi_80_Q_reg_14_inst : DFF_X1 port map( D => n6066, CK => CLK
                           , Q => n_2819, QN => 
                           DataPath_RF_bus_reg_dataout_2318_port);
   DataPath_RF_BLOCKi_81_Q_reg_14_inst : DFF_X1 port map( D => n6102, CK => CLK
                           , Q => n_2820, QN => 
                           DataPath_RF_bus_reg_dataout_2350_port);
   DataPath_REG_ALU_OUT_Q_reg_15_inst : DFF_X1 port map( D => n7008, CK => CLK,
                           Q => DRAM_ADDRESS_15_port, QN => n503);
   DataPath_REG_MEM_ALUOUT_Q_reg_15_inst : DFF_X1 port map( D => n1134, CK => 
                           CLK, Q => n_2821, QN => 
                           DataPath_i_REG_MEM_ALUOUT_15_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_15_inst : DFF_X1 port map( D => n6784, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_47_port,
                           QN => n614);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_15_inst : DFF_X1 port map( D => n6816, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_79_port,
                           QN => n646);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_15_inst : DFF_X1 port map( D => n6848, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_111_port
                           , QN => n678);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_15_inst : DFF_X1 port map( D => n6880, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_143_port
                           , QN => n710);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_15_inst : DFF_X1 port map( D => n6912, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_175_port
                           , QN => n742);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_15_inst : DFF_X1 port map( D => n6944, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_207_port
                           , QN => n774);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_15_inst : DFF_X1 port map( D => n6976, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_239_port
                           , QN => n806);
   DataPath_RF_BLOCKi_8_Q_reg_15_inst : DFF_X1 port map( D => n3342, CK => CLK,
                           Q => n_2822, QN => 
                           DataPath_RF_bus_reg_dataout_15_port);
   DataPath_RF_BLOCKi_9_Q_reg_15_inst : DFF_X1 port map( D => n3397, CK => CLK,
                           Q => n_2823, QN => 
                           DataPath_RF_bus_reg_dataout_47_port);
   DataPath_RF_BLOCKi_10_Q_reg_15_inst : DFF_X1 port map( D => n3435, CK => CLK
                           , Q => n_2824, QN => 
                           DataPath_RF_bus_reg_dataout_79_port);
   DataPath_RF_BLOCKi_11_Q_reg_15_inst : DFF_X1 port map( D => n3473, CK => CLK
                           , Q => n_2825, QN => 
                           DataPath_RF_bus_reg_dataout_111_port);
   DataPath_RF_BLOCKi_12_Q_reg_15_inst : DFF_X1 port map( D => n3511, CK => CLK
                           , Q => n_2826, QN => 
                           DataPath_RF_bus_reg_dataout_143_port);
   DataPath_RF_BLOCKi_13_Q_reg_15_inst : DFF_X1 port map( D => n3549, CK => CLK
                           , Q => n_2827, QN => 
                           DataPath_RF_bus_reg_dataout_175_port);
   DataPath_RF_BLOCKi_14_Q_reg_15_inst : DFF_X1 port map( D => n3587, CK => CLK
                           , Q => n_2828, QN => 
                           DataPath_RF_bus_reg_dataout_207_port);
   DataPath_RF_BLOCKi_15_Q_reg_15_inst : DFF_X1 port map( D => n3625, CK => CLK
                           , Q => n_2829, QN => 
                           DataPath_RF_bus_reg_dataout_239_port);
   DataPath_RF_BLOCKi_16_Q_reg_15_inst : DFF_X1 port map( D => n3663, CK => CLK
                           , Q => n_2830, QN => 
                           DataPath_RF_bus_reg_dataout_271_port);
   DataPath_RF_BLOCKi_17_Q_reg_15_inst : DFF_X1 port map( D => n3700, CK => CLK
                           , Q => n_2831, QN => 
                           DataPath_RF_bus_reg_dataout_303_port);
   DataPath_RF_BLOCKi_18_Q_reg_15_inst : DFF_X1 port map( D => n3737, CK => CLK
                           , Q => n_2832, QN => 
                           DataPath_RF_bus_reg_dataout_335_port);
   DataPath_RF_BLOCKi_19_Q_reg_15_inst : DFF_X1 port map( D => n3774, CK => CLK
                           , Q => n_2833, QN => 
                           DataPath_RF_bus_reg_dataout_367_port);
   DataPath_RF_BLOCKi_20_Q_reg_15_inst : DFF_X1 port map( D => n3809, CK => CLK
                           , Q => n_2834, QN => 
                           DataPath_RF_bus_reg_dataout_399_port);
   DataPath_RF_BLOCKi_21_Q_reg_15_inst : DFF_X1 port map( D => n3844, CK => CLK
                           , Q => n_2835, QN => 
                           DataPath_RF_bus_reg_dataout_431_port);
   DataPath_RF_BLOCKi_22_Q_reg_15_inst : DFF_X1 port map( D => n3879, CK => CLK
                           , Q => n_2836, QN => 
                           DataPath_RF_bus_reg_dataout_463_port);
   DataPath_RF_BLOCKi_23_Q_reg_15_inst : DFF_X1 port map( D => n3930, CK => CLK
                           , Q => n_2837, QN => 
                           DataPath_RF_bus_reg_dataout_495_port);
   DataPath_RF_BLOCKi_24_Q_reg_15_inst : DFF_X1 port map( D => n3998, CK => CLK
                           , Q => n_2838, QN => 
                           DataPath_RF_bus_reg_dataout_527_port);
   DataPath_RF_BLOCKi_25_Q_reg_15_inst : DFF_X1 port map( D => n4050, CK => CLK
                           , Q => n_2839, QN => 
                           DataPath_RF_bus_reg_dataout_559_port);
   DataPath_RF_BLOCKi_26_Q_reg_15_inst : DFF_X1 port map( D => n4085, CK => CLK
                           , Q => n_2840, QN => 
                           DataPath_RF_bus_reg_dataout_591_port);
   DataPath_RF_BLOCKi_27_Q_reg_15_inst : DFF_X1 port map( D => n4120, CK => CLK
                           , Q => n_2841, QN => 
                           DataPath_RF_bus_reg_dataout_623_port);
   DataPath_RF_BLOCKi_28_Q_reg_15_inst : DFF_X1 port map( D => n4155, CK => CLK
                           , Q => n_2842, QN => 
                           DataPath_RF_bus_reg_dataout_655_port);
   DataPath_RF_BLOCKi_29_Q_reg_15_inst : DFF_X1 port map( D => n4190, CK => CLK
                           , Q => n_2843, QN => 
                           DataPath_RF_bus_reg_dataout_687_port);
   DataPath_RF_BLOCKi_30_Q_reg_15_inst : DFF_X1 port map( D => n4225, CK => CLK
                           , Q => n_2844, QN => 
                           DataPath_RF_bus_reg_dataout_719_port);
   DataPath_RF_BLOCKi_31_Q_reg_15_inst : DFF_X1 port map( D => n4260, CK => CLK
                           , Q => n_2845, QN => 
                           DataPath_RF_bus_reg_dataout_751_port);
   DataPath_RF_BLOCKi_32_Q_reg_15_inst : DFF_X1 port map( D => n4295, CK => CLK
                           , Q => n_2846, QN => 
                           DataPath_RF_bus_reg_dataout_783_port);
   DataPath_RF_BLOCKi_33_Q_reg_15_inst : DFF_X1 port map( D => n4330, CK => CLK
                           , Q => n_2847, QN => 
                           DataPath_RF_bus_reg_dataout_815_port);
   DataPath_RF_BLOCKi_34_Q_reg_15_inst : DFF_X1 port map( D => n4365, CK => CLK
                           , Q => n_2848, QN => 
                           DataPath_RF_bus_reg_dataout_847_port);
   DataPath_RF_BLOCKi_35_Q_reg_15_inst : DFF_X1 port map( D => n4400, CK => CLK
                           , Q => n_2849, QN => 
                           DataPath_RF_bus_reg_dataout_879_port);
   DataPath_RF_BLOCKi_36_Q_reg_15_inst : DFF_X1 port map( D => n4435, CK => CLK
                           , Q => n_2850, QN => 
                           DataPath_RF_bus_reg_dataout_911_port);
   DataPath_RF_BLOCKi_37_Q_reg_15_inst : DFF_X1 port map( D => n4470, CK => CLK
                           , Q => n_2851, QN => 
                           DataPath_RF_bus_reg_dataout_943_port);
   DataPath_RF_BLOCKi_38_Q_reg_15_inst : DFF_X1 port map( D => n4505, CK => CLK
                           , Q => n_2852, QN => 
                           DataPath_RF_bus_reg_dataout_975_port);
   DataPath_RF_BLOCKi_39_Q_reg_15_inst : DFF_X1 port map( D => n4540, CK => CLK
                           , Q => n_2853, QN => 
                           DataPath_RF_bus_reg_dataout_1007_port);
   DataPath_RF_BLOCKi_40_Q_reg_15_inst : DFF_X1 port map( D => n4591, CK => CLK
                           , Q => n_2854, QN => 
                           DataPath_RF_bus_reg_dataout_1039_port);
   DataPath_RF_BLOCKi_41_Q_reg_15_inst : DFF_X1 port map( D => n4643, CK => CLK
                           , Q => n_2855, QN => 
                           DataPath_RF_bus_reg_dataout_1071_port);
   DataPath_RF_BLOCKi_42_Q_reg_15_inst : DFF_X1 port map( D => n4678, CK => CLK
                           , Q => n_2856, QN => 
                           DataPath_RF_bus_reg_dataout_1103_port);
   DataPath_RF_BLOCKi_43_Q_reg_15_inst : DFF_X1 port map( D => n4713, CK => CLK
                           , Q => n_2857, QN => 
                           DataPath_RF_bus_reg_dataout_1135_port);
   DataPath_RF_BLOCKi_44_Q_reg_15_inst : DFF_X1 port map( D => n4748, CK => CLK
                           , Q => n_2858, QN => 
                           DataPath_RF_bus_reg_dataout_1167_port);
   DataPath_RF_BLOCKi_45_Q_reg_15_inst : DFF_X1 port map( D => n4783, CK => CLK
                           , Q => n_2859, QN => 
                           DataPath_RF_bus_reg_dataout_1199_port);
   DataPath_RF_BLOCKi_46_Q_reg_15_inst : DFF_X1 port map( D => n4818, CK => CLK
                           , Q => n_2860, QN => 
                           DataPath_RF_bus_reg_dataout_1231_port);
   DataPath_RF_BLOCKi_47_Q_reg_15_inst : DFF_X1 port map( D => n4853, CK => CLK
                           , Q => n_2861, QN => 
                           DataPath_RF_bus_reg_dataout_1263_port);
   DataPath_RF_BLOCKi_48_Q_reg_15_inst : DFF_X1 port map( D => n4888, CK => CLK
                           , Q => n_2862, QN => 
                           DataPath_RF_bus_reg_dataout_1295_port);
   DataPath_RF_BLOCKi_49_Q_reg_15_inst : DFF_X1 port map( D => n4923, CK => CLK
                           , Q => n_2863, QN => 
                           DataPath_RF_bus_reg_dataout_1327_port);
   DataPath_RF_BLOCKi_50_Q_reg_15_inst : DFF_X1 port map( D => n4958, CK => CLK
                           , Q => n_2864, QN => 
                           DataPath_RF_bus_reg_dataout_1359_port);
   DataPath_RF_BLOCKi_51_Q_reg_15_inst : DFF_X1 port map( D => n4993, CK => CLK
                           , Q => n_2865, QN => 
                           DataPath_RF_bus_reg_dataout_1391_port);
   DataPath_RF_BLOCKi_52_Q_reg_15_inst : DFF_X1 port map( D => n5028, CK => CLK
                           , Q => n_2866, QN => 
                           DataPath_RF_bus_reg_dataout_1423_port);
   DataPath_RF_BLOCKi_53_Q_reg_15_inst : DFF_X1 port map( D => n5063, CK => CLK
                           , Q => n_2867, QN => 
                           DataPath_RF_bus_reg_dataout_1455_port);
   DataPath_RF_BLOCKi_54_Q_reg_15_inst : DFF_X1 port map( D => n5098, CK => CLK
                           , Q => n_2868, QN => 
                           DataPath_RF_bus_reg_dataout_1487_port);
   DataPath_RF_BLOCKi_55_Q_reg_15_inst : DFF_X1 port map( D => n5133, CK => CLK
                           , Q => n_2869, QN => 
                           DataPath_RF_bus_reg_dataout_1519_port);
   DataPath_RF_BLOCKi_56_Q_reg_15_inst : DFF_X1 port map( D => n5184, CK => CLK
                           , Q => n_2870, QN => 
                           DataPath_RF_bus_reg_dataout_1551_port);
   DataPath_RF_BLOCKi_57_Q_reg_15_inst : DFF_X1 port map( D => n5235, CK => CLK
                           , Q => n_2871, QN => 
                           DataPath_RF_bus_reg_dataout_1583_port);
   DataPath_RF_BLOCKi_58_Q_reg_15_inst : DFF_X1 port map( D => n5271, CK => CLK
                           , Q => n_2872, QN => 
                           DataPath_RF_bus_reg_dataout_1615_port);
   DataPath_RF_BLOCKi_59_Q_reg_15_inst : DFF_X1 port map( D => n5306, CK => CLK
                           , Q => n_2873, QN => 
                           DataPath_RF_bus_reg_dataout_1647_port);
   DataPath_RF_BLOCKi_60_Q_reg_15_inst : DFF_X1 port map( D => n5341, CK => CLK
                           , Q => n_2874, QN => 
                           DataPath_RF_bus_reg_dataout_1679_port);
   DataPath_RF_BLOCKi_61_Q_reg_15_inst : DFF_X1 port map( D => n5376, CK => CLK
                           , Q => n_2875, QN => 
                           DataPath_RF_bus_reg_dataout_1711_port);
   DataPath_RF_BLOCKi_62_Q_reg_15_inst : DFF_X1 port map( D => n5411, CK => CLK
                           , Q => n_2876, QN => 
                           DataPath_RF_bus_reg_dataout_1743_port);
   DataPath_RF_BLOCKi_63_Q_reg_15_inst : DFF_X1 port map( D => n5446, CK => CLK
                           , Q => n_2877, QN => 
                           DataPath_RF_bus_reg_dataout_1775_port);
   DataPath_RF_BLOCKi_64_Q_reg_15_inst : DFF_X1 port map( D => n5481, CK => CLK
                           , Q => n_2878, QN => 
                           DataPath_RF_bus_reg_dataout_1807_port);
   DataPath_RF_BLOCKi_65_Q_reg_15_inst : DFF_X1 port map( D => n5516, CK => CLK
                           , Q => n_2879, QN => 
                           DataPath_RF_bus_reg_dataout_1839_port);
   DataPath_RF_BLOCKi_66_Q_reg_15_inst : DFF_X1 port map( D => n5551, CK => CLK
                           , Q => n_2880, QN => 
                           DataPath_RF_bus_reg_dataout_1871_port);
   DataPath_RF_BLOCKi_67_Q_reg_15_inst : DFF_X1 port map( D => n5586, CK => CLK
                           , Q => n_2881, QN => 
                           DataPath_RF_bus_reg_dataout_1903_port);
   DataPath_RF_BLOCKi_68_Q_reg_15_inst : DFF_X1 port map( D => n5625, CK => CLK
                           , Q => n_2882, QN => 
                           DataPath_RF_bus_reg_dataout_1935_port);
   DataPath_RF_BLOCKi_69_Q_reg_15_inst : DFF_X1 port map( D => n5662, CK => CLK
                           , Q => n_2883, QN => 
                           DataPath_RF_bus_reg_dataout_1967_port);
   DataPath_RF_BLOCKi_70_Q_reg_15_inst : DFF_X1 port map( D => n5699, CK => CLK
                           , Q => n_2884, QN => 
                           DataPath_RF_bus_reg_dataout_1999_port);
   DataPath_RF_BLOCKi_71_Q_reg_15_inst : DFF_X1 port map( D => n5736, CK => CLK
                           , Q => n_2885, QN => 
                           DataPath_RF_bus_reg_dataout_2031_port);
   DataPath_RF_BLOCKi_82_Q_reg_15_inst : DFF_X1 port map( D => n880, CK => CLK,
                           Q => n_2886, QN => 
                           DataPath_RF_bus_reg_dataout_2383_port);
   DataPath_RF_BLOCKi_83_Q_reg_15_inst : DFF_X1 port map( D => n948, CK => CLK,
                           Q => n_2887, QN => 
                           DataPath_RF_bus_reg_dataout_2415_port);
   DataPath_RF_BLOCKi_84_Q_reg_15_inst : DFF_X1 port map( D => n986, CK => CLK,
                           Q => n_2888, QN => 
                           DataPath_RF_bus_reg_dataout_2447_port);
   DataPath_RF_BLOCKi_85_Q_reg_15_inst : DFF_X1 port map( D => n1023, CK => CLK
                           , Q => n_2889, QN => 
                           DataPath_RF_bus_reg_dataout_2479_port);
   DataPath_RF_BLOCKi_86_Q_reg_15_inst : DFF_X1 port map( D => n1060, CK => CLK
                           , Q => n_2890, QN => 
                           DataPath_RF_bus_reg_dataout_2511_port);
   DataPath_RF_BLOCKi_87_Q_reg_15_inst : DFF_X1 port map( D => n1097, CK => CLK
                           , Q => n_2891, QN => 
                           DataPath_RF_bus_reg_dataout_2543_port);
   DataPath_RF_BLOCKi_72_Q_reg_15_inst : DFF_X1 port map( D => n5773, CK => CLK
                           , Q => n_2892, QN => 
                           DataPath_RF_bus_reg_dataout_2063_port);
   DataPath_RF_BLOCKi_73_Q_reg_15_inst : DFF_X1 port map( D => n5812, CK => CLK
                           , Q => n_2893, QN => 
                           DataPath_RF_bus_reg_dataout_2095_port);
   DataPath_RF_BLOCKi_74_Q_reg_15_inst : DFF_X1 port map( D => n5848, CK => CLK
                           , Q => n_2894, QN => 
                           DataPath_RF_bus_reg_dataout_2127_port);
   DataPath_RF_BLOCKi_75_Q_reg_15_inst : DFF_X1 port map( D => n5884, CK => CLK
                           , Q => n_2895, QN => 
                           DataPath_RF_bus_reg_dataout_2159_port);
   DataPath_RF_BLOCKi_76_Q_reg_15_inst : DFF_X1 port map( D => n5920, CK => CLK
                           , Q => n_2896, QN => 
                           DataPath_RF_bus_reg_dataout_2191_port);
   DataPath_RF_BLOCKi_77_Q_reg_15_inst : DFF_X1 port map( D => n5956, CK => CLK
                           , Q => n_2897, QN => 
                           DataPath_RF_bus_reg_dataout_2223_port);
   DataPath_RF_BLOCKi_78_Q_reg_15_inst : DFF_X1 port map( D => n5992, CK => CLK
                           , Q => n_2898, QN => 
                           DataPath_RF_bus_reg_dataout_2255_port);
   DataPath_RF_BLOCKi_79_Q_reg_15_inst : DFF_X1 port map( D => n6028, CK => CLK
                           , Q => n_2899, QN => 
                           DataPath_RF_bus_reg_dataout_2287_port);
   DataPath_RF_BLOCKi_80_Q_reg_15_inst : DFF_X1 port map( D => n6065, CK => CLK
                           , Q => n_2900, QN => 
                           DataPath_RF_bus_reg_dataout_2319_port);
   DataPath_RF_BLOCKi_81_Q_reg_15_inst : DFF_X1 port map( D => n6101, CK => CLK
                           , Q => n_2901, QN => 
                           DataPath_RF_bus_reg_dataout_2351_port);
   DataPath_REG_ALU_OUT_Q_reg_16_inst : DFF_X1 port map( D => n7007, CK => CLK,
                           Q => DRAM_ADDRESS_16_port, QN => n504);
   DataPath_REG_MEM_ALUOUT_Q_reg_16_inst : DFF_X1 port map( D => n1133, CK => 
                           CLK, Q => n_2902, QN => 
                           DataPath_i_REG_MEM_ALUOUT_16_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_16_inst : DFF_X1 port map( D => n6783, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_48_port,
                           QN => n615);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_16_inst : DFF_X1 port map( D => n6815, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_80_port,
                           QN => n647);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_16_inst : DFF_X1 port map( D => n6847, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_112_port
                           , QN => n679);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_16_inst : DFF_X1 port map( D => n6879, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_144_port
                           , QN => n711);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_16_inst : DFF_X1 port map( D => n6911, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_176_port
                           , QN => n743);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_16_inst : DFF_X1 port map( D => n6943, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_208_port
                           , QN => n775);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_16_inst : DFF_X1 port map( D => n6975, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_240_port
                           , QN => n807);
   DataPath_RF_BLOCKi_8_Q_reg_16_inst : DFF_X1 port map( D => n3340, CK => CLK,
                           Q => n_2903, QN => 
                           DataPath_RF_bus_reg_dataout_16_port);
   DataPath_RF_BLOCKi_9_Q_reg_16_inst : DFF_X1 port map( D => n3396, CK => CLK,
                           Q => n_2904, QN => 
                           DataPath_RF_bus_reg_dataout_48_port);
   DataPath_RF_BLOCKi_10_Q_reg_16_inst : DFF_X1 port map( D => n3434, CK => CLK
                           , Q => n_2905, QN => 
                           DataPath_RF_bus_reg_dataout_80_port);
   DataPath_RF_BLOCKi_11_Q_reg_16_inst : DFF_X1 port map( D => n3472, CK => CLK
                           , Q => n_2906, QN => 
                           DataPath_RF_bus_reg_dataout_112_port);
   DataPath_RF_BLOCKi_12_Q_reg_16_inst : DFF_X1 port map( D => n3510, CK => CLK
                           , Q => n_2907, QN => 
                           DataPath_RF_bus_reg_dataout_144_port);
   DataPath_RF_BLOCKi_13_Q_reg_16_inst : DFF_X1 port map( D => n3548, CK => CLK
                           , Q => n_2908, QN => 
                           DataPath_RF_bus_reg_dataout_176_port);
   DataPath_RF_BLOCKi_14_Q_reg_16_inst : DFF_X1 port map( D => n3586, CK => CLK
                           , Q => n_2909, QN => 
                           DataPath_RF_bus_reg_dataout_208_port);
   DataPath_RF_BLOCKi_15_Q_reg_16_inst : DFF_X1 port map( D => n3624, CK => CLK
                           , Q => n_2910, QN => 
                           DataPath_RF_bus_reg_dataout_240_port);
   DataPath_RF_BLOCKi_16_Q_reg_16_inst : DFF_X1 port map( D => n3662, CK => CLK
                           , Q => n_2911, QN => 
                           DataPath_RF_bus_reg_dataout_272_port);
   DataPath_RF_BLOCKi_17_Q_reg_16_inst : DFF_X1 port map( D => n3699, CK => CLK
                           , Q => n_2912, QN => 
                           DataPath_RF_bus_reg_dataout_304_port);
   DataPath_RF_BLOCKi_18_Q_reg_16_inst : DFF_X1 port map( D => n3736, CK => CLK
                           , Q => n_2913, QN => 
                           DataPath_RF_bus_reg_dataout_336_port);
   DataPath_RF_BLOCKi_19_Q_reg_16_inst : DFF_X1 port map( D => n3773, CK => CLK
                           , Q => n_2914, QN => 
                           DataPath_RF_bus_reg_dataout_368_port);
   DataPath_RF_BLOCKi_20_Q_reg_16_inst : DFF_X1 port map( D => n3808, CK => CLK
                           , Q => n_2915, QN => 
                           DataPath_RF_bus_reg_dataout_400_port);
   DataPath_RF_BLOCKi_21_Q_reg_16_inst : DFF_X1 port map( D => n3843, CK => CLK
                           , Q => n_2916, QN => 
                           DataPath_RF_bus_reg_dataout_432_port);
   DataPath_RF_BLOCKi_22_Q_reg_16_inst : DFF_X1 port map( D => n3878, CK => CLK
                           , Q => n_2917, QN => 
                           DataPath_RF_bus_reg_dataout_464_port);
   DataPath_RF_BLOCKi_23_Q_reg_16_inst : DFF_X1 port map( D => n3928, CK => CLK
                           , Q => n_2918, QN => 
                           DataPath_RF_bus_reg_dataout_496_port);
   DataPath_RF_BLOCKi_24_Q_reg_16_inst : DFF_X1 port map( D => n3996, CK => CLK
                           , Q => n_2919, QN => 
                           DataPath_RF_bus_reg_dataout_528_port);
   DataPath_RF_BLOCKi_25_Q_reg_16_inst : DFF_X1 port map( D => n4049, CK => CLK
                           , Q => n_2920, QN => 
                           DataPath_RF_bus_reg_dataout_560_port);
   DataPath_RF_BLOCKi_26_Q_reg_16_inst : DFF_X1 port map( D => n4084, CK => CLK
                           , Q => n_2921, QN => 
                           DataPath_RF_bus_reg_dataout_592_port);
   DataPath_RF_BLOCKi_27_Q_reg_16_inst : DFF_X1 port map( D => n4119, CK => CLK
                           , Q => n_2922, QN => 
                           DataPath_RF_bus_reg_dataout_624_port);
   DataPath_RF_BLOCKi_28_Q_reg_16_inst : DFF_X1 port map( D => n4154, CK => CLK
                           , Q => n_2923, QN => 
                           DataPath_RF_bus_reg_dataout_656_port);
   DataPath_RF_BLOCKi_29_Q_reg_16_inst : DFF_X1 port map( D => n4189, CK => CLK
                           , Q => n_2924, QN => 
                           DataPath_RF_bus_reg_dataout_688_port);
   DataPath_RF_BLOCKi_30_Q_reg_16_inst : DFF_X1 port map( D => n4224, CK => CLK
                           , Q => n_2925, QN => 
                           DataPath_RF_bus_reg_dataout_720_port);
   DataPath_RF_BLOCKi_31_Q_reg_16_inst : DFF_X1 port map( D => n4259, CK => CLK
                           , Q => n_2926, QN => 
                           DataPath_RF_bus_reg_dataout_752_port);
   DataPath_RF_BLOCKi_32_Q_reg_16_inst : DFF_X1 port map( D => n4294, CK => CLK
                           , Q => n_2927, QN => 
                           DataPath_RF_bus_reg_dataout_784_port);
   DataPath_RF_BLOCKi_33_Q_reg_16_inst : DFF_X1 port map( D => n4329, CK => CLK
                           , Q => n_2928, QN => 
                           DataPath_RF_bus_reg_dataout_816_port);
   DataPath_RF_BLOCKi_34_Q_reg_16_inst : DFF_X1 port map( D => n4364, CK => CLK
                           , Q => n_2929, QN => 
                           DataPath_RF_bus_reg_dataout_848_port);
   DataPath_RF_BLOCKi_35_Q_reg_16_inst : DFF_X1 port map( D => n4399, CK => CLK
                           , Q => n_2930, QN => 
                           DataPath_RF_bus_reg_dataout_880_port);
   DataPath_RF_BLOCKi_36_Q_reg_16_inst : DFF_X1 port map( D => n4434, CK => CLK
                           , Q => n_2931, QN => 
                           DataPath_RF_bus_reg_dataout_912_port);
   DataPath_RF_BLOCKi_37_Q_reg_16_inst : DFF_X1 port map( D => n4469, CK => CLK
                           , Q => n_2932, QN => 
                           DataPath_RF_bus_reg_dataout_944_port);
   DataPath_RF_BLOCKi_38_Q_reg_16_inst : DFF_X1 port map( D => n4504, CK => CLK
                           , Q => n_2933, QN => 
                           DataPath_RF_bus_reg_dataout_976_port);
   DataPath_RF_BLOCKi_39_Q_reg_16_inst : DFF_X1 port map( D => n4539, CK => CLK
                           , Q => n_2934, QN => 
                           DataPath_RF_bus_reg_dataout_1008_port);
   DataPath_RF_BLOCKi_40_Q_reg_16_inst : DFF_X1 port map( D => n4589, CK => CLK
                           , Q => n_2935, QN => 
                           DataPath_RF_bus_reg_dataout_1040_port);
   DataPath_RF_BLOCKi_41_Q_reg_16_inst : DFF_X1 port map( D => n4642, CK => CLK
                           , Q => n_2936, QN => 
                           DataPath_RF_bus_reg_dataout_1072_port);
   DataPath_RF_BLOCKi_42_Q_reg_16_inst : DFF_X1 port map( D => n4677, CK => CLK
                           , Q => n_2937, QN => 
                           DataPath_RF_bus_reg_dataout_1104_port);
   DataPath_RF_BLOCKi_43_Q_reg_16_inst : DFF_X1 port map( D => n4712, CK => CLK
                           , Q => n_2938, QN => 
                           DataPath_RF_bus_reg_dataout_1136_port);
   DataPath_RF_BLOCKi_44_Q_reg_16_inst : DFF_X1 port map( D => n4747, CK => CLK
                           , Q => n_2939, QN => 
                           DataPath_RF_bus_reg_dataout_1168_port);
   DataPath_RF_BLOCKi_45_Q_reg_16_inst : DFF_X1 port map( D => n4782, CK => CLK
                           , Q => n_2940, QN => 
                           DataPath_RF_bus_reg_dataout_1200_port);
   DataPath_RF_BLOCKi_46_Q_reg_16_inst : DFF_X1 port map( D => n4817, CK => CLK
                           , Q => n_2941, QN => 
                           DataPath_RF_bus_reg_dataout_1232_port);
   DataPath_RF_BLOCKi_47_Q_reg_16_inst : DFF_X1 port map( D => n4852, CK => CLK
                           , Q => n_2942, QN => 
                           DataPath_RF_bus_reg_dataout_1264_port);
   DataPath_RF_BLOCKi_48_Q_reg_16_inst : DFF_X1 port map( D => n4887, CK => CLK
                           , Q => n_2943, QN => 
                           DataPath_RF_bus_reg_dataout_1296_port);
   DataPath_RF_BLOCKi_49_Q_reg_16_inst : DFF_X1 port map( D => n4922, CK => CLK
                           , Q => n_2944, QN => 
                           DataPath_RF_bus_reg_dataout_1328_port);
   DataPath_RF_BLOCKi_50_Q_reg_16_inst : DFF_X1 port map( D => n4957, CK => CLK
                           , Q => n_2945, QN => 
                           DataPath_RF_bus_reg_dataout_1360_port);
   DataPath_RF_BLOCKi_51_Q_reg_16_inst : DFF_X1 port map( D => n4992, CK => CLK
                           , Q => n_2946, QN => 
                           DataPath_RF_bus_reg_dataout_1392_port);
   DataPath_RF_BLOCKi_52_Q_reg_16_inst : DFF_X1 port map( D => n5027, CK => CLK
                           , Q => n_2947, QN => 
                           DataPath_RF_bus_reg_dataout_1424_port);
   DataPath_RF_BLOCKi_53_Q_reg_16_inst : DFF_X1 port map( D => n5062, CK => CLK
                           , Q => n_2948, QN => 
                           DataPath_RF_bus_reg_dataout_1456_port);
   DataPath_RF_BLOCKi_54_Q_reg_16_inst : DFF_X1 port map( D => n5097, CK => CLK
                           , Q => n_2949, QN => 
                           DataPath_RF_bus_reg_dataout_1488_port);
   DataPath_RF_BLOCKi_55_Q_reg_16_inst : DFF_X1 port map( D => n5132, CK => CLK
                           , Q => n_2950, QN => 
                           DataPath_RF_bus_reg_dataout_1520_port);
   DataPath_RF_BLOCKi_56_Q_reg_16_inst : DFF_X1 port map( D => n5182, CK => CLK
                           , Q => n_2951, QN => 
                           DataPath_RF_bus_reg_dataout_1552_port);
   DataPath_RF_BLOCKi_57_Q_reg_16_inst : DFF_X1 port map( D => n5234, CK => CLK
                           , Q => n_2952, QN => 
                           DataPath_RF_bus_reg_dataout_1584_port);
   DataPath_RF_BLOCKi_58_Q_reg_16_inst : DFF_X1 port map( D => n5270, CK => CLK
                           , Q => n_2953, QN => 
                           DataPath_RF_bus_reg_dataout_1616_port);
   DataPath_RF_BLOCKi_59_Q_reg_16_inst : DFF_X1 port map( D => n5305, CK => CLK
                           , Q => n_2954, QN => 
                           DataPath_RF_bus_reg_dataout_1648_port);
   DataPath_RF_BLOCKi_60_Q_reg_16_inst : DFF_X1 port map( D => n5340, CK => CLK
                           , Q => n_2955, QN => 
                           DataPath_RF_bus_reg_dataout_1680_port);
   DataPath_RF_BLOCKi_61_Q_reg_16_inst : DFF_X1 port map( D => n5375, CK => CLK
                           , Q => n_2956, QN => 
                           DataPath_RF_bus_reg_dataout_1712_port);
   DataPath_RF_BLOCKi_62_Q_reg_16_inst : DFF_X1 port map( D => n5410, CK => CLK
                           , Q => n_2957, QN => 
                           DataPath_RF_bus_reg_dataout_1744_port);
   DataPath_RF_BLOCKi_63_Q_reg_16_inst : DFF_X1 port map( D => n5445, CK => CLK
                           , Q => n_2958, QN => 
                           DataPath_RF_bus_reg_dataout_1776_port);
   DataPath_RF_BLOCKi_64_Q_reg_16_inst : DFF_X1 port map( D => n5480, CK => CLK
                           , Q => n_2959, QN => 
                           DataPath_RF_bus_reg_dataout_1808_port);
   DataPath_RF_BLOCKi_65_Q_reg_16_inst : DFF_X1 port map( D => n5515, CK => CLK
                           , Q => n_2960, QN => 
                           DataPath_RF_bus_reg_dataout_1840_port);
   DataPath_RF_BLOCKi_66_Q_reg_16_inst : DFF_X1 port map( D => n5550, CK => CLK
                           , Q => n_2961, QN => 
                           DataPath_RF_bus_reg_dataout_1872_port);
   DataPath_RF_BLOCKi_67_Q_reg_16_inst : DFF_X1 port map( D => n5585, CK => CLK
                           , Q => n_2962, QN => 
                           DataPath_RF_bus_reg_dataout_1904_port);
   DataPath_RF_BLOCKi_68_Q_reg_16_inst : DFF_X1 port map( D => n5624, CK => CLK
                           , Q => n_2963, QN => 
                           DataPath_RF_bus_reg_dataout_1936_port);
   DataPath_RF_BLOCKi_69_Q_reg_16_inst : DFF_X1 port map( D => n5661, CK => CLK
                           , Q => n_2964, QN => 
                           DataPath_RF_bus_reg_dataout_1968_port);
   DataPath_RF_BLOCKi_70_Q_reg_16_inst : DFF_X1 port map( D => n5698, CK => CLK
                           , Q => n_2965, QN => 
                           DataPath_RF_bus_reg_dataout_2000_port);
   DataPath_RF_BLOCKi_71_Q_reg_16_inst : DFF_X1 port map( D => n5735, CK => CLK
                           , Q => n_2966, QN => 
                           DataPath_RF_bus_reg_dataout_2032_port);
   DataPath_RF_BLOCKi_83_Q_reg_16_inst : DFF_X1 port map( D => n946, CK => CLK,
                           Q => n_2967, QN => 
                           DataPath_RF_bus_reg_dataout_2416_port);
   DataPath_RF_BLOCKi_84_Q_reg_16_inst : DFF_X1 port map( D => n985, CK => CLK,
                           Q => n_2968, QN => 
                           DataPath_RF_bus_reg_dataout_2448_port);
   DataPath_RF_BLOCKi_85_Q_reg_16_inst : DFF_X1 port map( D => n1022, CK => CLK
                           , Q => n_2969, QN => 
                           DataPath_RF_bus_reg_dataout_2480_port);
   DataPath_RF_BLOCKi_86_Q_reg_16_inst : DFF_X1 port map( D => n1059, CK => CLK
                           , Q => n_2970, QN => 
                           DataPath_RF_bus_reg_dataout_2512_port);
   DataPath_RF_BLOCKi_87_Q_reg_16_inst : DFF_X1 port map( D => n1096, CK => CLK
                           , Q => n_2971, QN => 
                           DataPath_RF_bus_reg_dataout_2544_port);
   DataPath_RF_BLOCKi_72_Q_reg_16_inst : DFF_X1 port map( D => n5772, CK => CLK
                           , Q => n_2972, QN => 
                           DataPath_RF_bus_reg_dataout_2064_port);
   DataPath_RF_BLOCKi_73_Q_reg_16_inst : DFF_X1 port map( D => n5811, CK => CLK
                           , Q => n_2973, QN => 
                           DataPath_RF_bus_reg_dataout_2096_port);
   DataPath_RF_BLOCKi_74_Q_reg_16_inst : DFF_X1 port map( D => n5847, CK => CLK
                           , Q => n_2974, QN => 
                           DataPath_RF_bus_reg_dataout_2128_port);
   DataPath_RF_BLOCKi_75_Q_reg_16_inst : DFF_X1 port map( D => n5883, CK => CLK
                           , Q => n_2975, QN => 
                           DataPath_RF_bus_reg_dataout_2160_port);
   DataPath_RF_BLOCKi_76_Q_reg_16_inst : DFF_X1 port map( D => n5919, CK => CLK
                           , Q => n_2976, QN => 
                           DataPath_RF_bus_reg_dataout_2192_port);
   DataPath_RF_BLOCKi_77_Q_reg_16_inst : DFF_X1 port map( D => n5955, CK => CLK
                           , Q => n_2977, QN => 
                           DataPath_RF_bus_reg_dataout_2224_port);
   DataPath_RF_BLOCKi_78_Q_reg_16_inst : DFF_X1 port map( D => n5991, CK => CLK
                           , Q => n_2978, QN => 
                           DataPath_RF_bus_reg_dataout_2256_port);
   DataPath_RF_BLOCKi_79_Q_reg_16_inst : DFF_X1 port map( D => n6027, CK => CLK
                           , Q => n_2979, QN => 
                           DataPath_RF_bus_reg_dataout_2288_port);
   DataPath_RF_BLOCKi_80_Q_reg_16_inst : DFF_X1 port map( D => n6064, CK => CLK
                           , Q => n_2980, QN => 
                           DataPath_RF_bus_reg_dataout_2320_port);
   DataPath_RF_BLOCKi_81_Q_reg_16_inst : DFF_X1 port map( D => n6100, CK => CLK
                           , Q => n_2981, QN => 
                           DataPath_RF_bus_reg_dataout_2352_port);
   DataPath_RF_BLOCKi_82_Q_reg_16_inst : DFF_X1 port map( D => n6134, CK => CLK
                           , Q => n_2982, QN => 
                           DataPath_RF_bus_reg_dataout_2384_port);
   DataPath_REG_ALU_OUT_Q_reg_18_inst : DFF_X1 port map( D => n7005, CK => CLK,
                           Q => DRAM_ADDRESS_18_port, QN => n505);
   DataPath_REG_MEM_ALUOUT_Q_reg_18_inst : DFF_X1 port map( D => n1131, CK => 
                           CLK, Q => n_2983, QN => 
                           DataPath_i_REG_MEM_ALUOUT_18_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_18_inst : DFF_X1 port map( D => n6781, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_50_port,
                           QN => n617);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_18_inst : DFF_X1 port map( D => n6813, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_82_port,
                           QN => n649);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_18_inst : DFF_X1 port map( D => n6845, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_114_port
                           , QN => n681);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_18_inst : DFF_X1 port map( D => n6877, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_146_port
                           , QN => n713);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_18_inst : DFF_X1 port map( D => n6909, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_178_port
                           , QN => n745);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_18_inst : DFF_X1 port map( D => n6941, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_210_port
                           , QN => n777);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_18_inst : DFF_X1 port map( D => n6973, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_242_port
                           , QN => n809);
   DataPath_RF_BLOCKi_8_Q_reg_18_inst : DFF_X1 port map( D => n3336, CK => CLK,
                           Q => n_2984, QN => 
                           DataPath_RF_bus_reg_dataout_18_port);
   DataPath_RF_BLOCKi_9_Q_reg_18_inst : DFF_X1 port map( D => n3394, CK => CLK,
                           Q => n_2985, QN => 
                           DataPath_RF_bus_reg_dataout_50_port);
   DataPath_RF_BLOCKi_10_Q_reg_18_inst : DFF_X1 port map( D => n3432, CK => CLK
                           , Q => n_2986, QN => 
                           DataPath_RF_bus_reg_dataout_82_port);
   DataPath_RF_BLOCKi_11_Q_reg_18_inst : DFF_X1 port map( D => n3470, CK => CLK
                           , Q => n_2987, QN => 
                           DataPath_RF_bus_reg_dataout_114_port);
   DataPath_RF_BLOCKi_12_Q_reg_18_inst : DFF_X1 port map( D => n3508, CK => CLK
                           , Q => n_2988, QN => 
                           DataPath_RF_bus_reg_dataout_146_port);
   DataPath_RF_BLOCKi_13_Q_reg_18_inst : DFF_X1 port map( D => n3546, CK => CLK
                           , Q => n_2989, QN => 
                           DataPath_RF_bus_reg_dataout_178_port);
   DataPath_RF_BLOCKi_14_Q_reg_18_inst : DFF_X1 port map( D => n3584, CK => CLK
                           , Q => n_2990, QN => 
                           DataPath_RF_bus_reg_dataout_210_port);
   DataPath_RF_BLOCKi_15_Q_reg_18_inst : DFF_X1 port map( D => n3622, CK => CLK
                           , Q => n_2991, QN => 
                           DataPath_RF_bus_reg_dataout_242_port);
   DataPath_RF_BLOCKi_16_Q_reg_18_inst : DFF_X1 port map( D => n3660, CK => CLK
                           , Q => n_2992, QN => 
                           DataPath_RF_bus_reg_dataout_274_port);
   DataPath_RF_BLOCKi_17_Q_reg_18_inst : DFF_X1 port map( D => n3697, CK => CLK
                           , Q => n_2993, QN => 
                           DataPath_RF_bus_reg_dataout_306_port);
   DataPath_RF_BLOCKi_18_Q_reg_18_inst : DFF_X1 port map( D => n3734, CK => CLK
                           , Q => n_2994, QN => 
                           DataPath_RF_bus_reg_dataout_338_port);
   DataPath_RF_BLOCKi_19_Q_reg_18_inst : DFF_X1 port map( D => n3771, CK => CLK
                           , Q => n_2995, QN => 
                           DataPath_RF_bus_reg_dataout_370_port);
   DataPath_RF_BLOCKi_20_Q_reg_18_inst : DFF_X1 port map( D => n3806, CK => CLK
                           , Q => n_2996, QN => 
                           DataPath_RF_bus_reg_dataout_402_port);
   DataPath_RF_BLOCKi_21_Q_reg_18_inst : DFF_X1 port map( D => n3841, CK => CLK
                           , Q => n_2997, QN => 
                           DataPath_RF_bus_reg_dataout_434_port);
   DataPath_RF_BLOCKi_22_Q_reg_18_inst : DFF_X1 port map( D => n3876, CK => CLK
                           , Q => n_2998, QN => 
                           DataPath_RF_bus_reg_dataout_466_port);
   DataPath_RF_BLOCKi_23_Q_reg_18_inst : DFF_X1 port map( D => n3924, CK => CLK
                           , Q => n_2999, QN => 
                           DataPath_RF_bus_reg_dataout_498_port);
   DataPath_RF_BLOCKi_24_Q_reg_18_inst : DFF_X1 port map( D => n3992, CK => CLK
                           , Q => n_3000, QN => 
                           DataPath_RF_bus_reg_dataout_530_port);
   DataPath_RF_BLOCKi_25_Q_reg_18_inst : DFF_X1 port map( D => n4047, CK => CLK
                           , Q => n_3001, QN => 
                           DataPath_RF_bus_reg_dataout_562_port);
   DataPath_RF_BLOCKi_26_Q_reg_18_inst : DFF_X1 port map( D => n4082, CK => CLK
                           , Q => n_3002, QN => 
                           DataPath_RF_bus_reg_dataout_594_port);
   DataPath_RF_BLOCKi_27_Q_reg_18_inst : DFF_X1 port map( D => n4117, CK => CLK
                           , Q => n_3003, QN => 
                           DataPath_RF_bus_reg_dataout_626_port);
   DataPath_RF_BLOCKi_28_Q_reg_18_inst : DFF_X1 port map( D => n4152, CK => CLK
                           , Q => n_3004, QN => 
                           DataPath_RF_bus_reg_dataout_658_port);
   DataPath_RF_BLOCKi_29_Q_reg_18_inst : DFF_X1 port map( D => n4187, CK => CLK
                           , Q => n_3005, QN => 
                           DataPath_RF_bus_reg_dataout_690_port);
   DataPath_RF_BLOCKi_30_Q_reg_18_inst : DFF_X1 port map( D => n4222, CK => CLK
                           , Q => n_3006, QN => 
                           DataPath_RF_bus_reg_dataout_722_port);
   DataPath_RF_BLOCKi_31_Q_reg_18_inst : DFF_X1 port map( D => n4257, CK => CLK
                           , Q => n_3007, QN => 
                           DataPath_RF_bus_reg_dataout_754_port);
   DataPath_RF_BLOCKi_32_Q_reg_18_inst : DFF_X1 port map( D => n4292, CK => CLK
                           , Q => n_3008, QN => 
                           DataPath_RF_bus_reg_dataout_786_port);
   DataPath_RF_BLOCKi_33_Q_reg_18_inst : DFF_X1 port map( D => n4327, CK => CLK
                           , Q => n_3009, QN => 
                           DataPath_RF_bus_reg_dataout_818_port);
   DataPath_RF_BLOCKi_34_Q_reg_18_inst : DFF_X1 port map( D => n4362, CK => CLK
                           , Q => n_3010, QN => 
                           DataPath_RF_bus_reg_dataout_850_port);
   DataPath_RF_BLOCKi_35_Q_reg_18_inst : DFF_X1 port map( D => n4397, CK => CLK
                           , Q => n_3011, QN => 
                           DataPath_RF_bus_reg_dataout_882_port);
   DataPath_RF_BLOCKi_36_Q_reg_18_inst : DFF_X1 port map( D => n4432, CK => CLK
                           , Q => n_3012, QN => 
                           DataPath_RF_bus_reg_dataout_914_port);
   DataPath_RF_BLOCKi_37_Q_reg_18_inst : DFF_X1 port map( D => n4467, CK => CLK
                           , Q => n_3013, QN => 
                           DataPath_RF_bus_reg_dataout_946_port);
   DataPath_RF_BLOCKi_38_Q_reg_18_inst : DFF_X1 port map( D => n4502, CK => CLK
                           , Q => n_3014, QN => 
                           DataPath_RF_bus_reg_dataout_978_port);
   DataPath_RF_BLOCKi_39_Q_reg_18_inst : DFF_X1 port map( D => n4537, CK => CLK
                           , Q => n_3015, QN => 
                           DataPath_RF_bus_reg_dataout_1010_port);
   DataPath_RF_BLOCKi_40_Q_reg_18_inst : DFF_X1 port map( D => n4585, CK => CLK
                           , Q => n_3016, QN => 
                           DataPath_RF_bus_reg_dataout_1042_port);
   DataPath_RF_BLOCKi_41_Q_reg_18_inst : DFF_X1 port map( D => n4640, CK => CLK
                           , Q => n_3017, QN => 
                           DataPath_RF_bus_reg_dataout_1074_port);
   DataPath_RF_BLOCKi_42_Q_reg_18_inst : DFF_X1 port map( D => n4675, CK => CLK
                           , Q => n_3018, QN => 
                           DataPath_RF_bus_reg_dataout_1106_port);
   DataPath_RF_BLOCKi_43_Q_reg_18_inst : DFF_X1 port map( D => n4710, CK => CLK
                           , Q => n_3019, QN => 
                           DataPath_RF_bus_reg_dataout_1138_port);
   DataPath_RF_BLOCKi_44_Q_reg_18_inst : DFF_X1 port map( D => n4745, CK => CLK
                           , Q => n_3020, QN => 
                           DataPath_RF_bus_reg_dataout_1170_port);
   DataPath_RF_BLOCKi_45_Q_reg_18_inst : DFF_X1 port map( D => n4780, CK => CLK
                           , Q => n_3021, QN => 
                           DataPath_RF_bus_reg_dataout_1202_port);
   DataPath_RF_BLOCKi_46_Q_reg_18_inst : DFF_X1 port map( D => n4815, CK => CLK
                           , Q => n_3022, QN => 
                           DataPath_RF_bus_reg_dataout_1234_port);
   DataPath_RF_BLOCKi_47_Q_reg_18_inst : DFF_X1 port map( D => n4850, CK => CLK
                           , Q => n_3023, QN => 
                           DataPath_RF_bus_reg_dataout_1266_port);
   DataPath_RF_BLOCKi_48_Q_reg_18_inst : DFF_X1 port map( D => n4885, CK => CLK
                           , Q => n_3024, QN => 
                           DataPath_RF_bus_reg_dataout_1298_port);
   DataPath_RF_BLOCKi_49_Q_reg_18_inst : DFF_X1 port map( D => n4920, CK => CLK
                           , Q => n_3025, QN => 
                           DataPath_RF_bus_reg_dataout_1330_port);
   DataPath_RF_BLOCKi_50_Q_reg_18_inst : DFF_X1 port map( D => n4955, CK => CLK
                           , Q => n_3026, QN => 
                           DataPath_RF_bus_reg_dataout_1362_port);
   DataPath_RF_BLOCKi_51_Q_reg_18_inst : DFF_X1 port map( D => n4990, CK => CLK
                           , Q => n_3027, QN => 
                           DataPath_RF_bus_reg_dataout_1394_port);
   DataPath_RF_BLOCKi_52_Q_reg_18_inst : DFF_X1 port map( D => n5025, CK => CLK
                           , Q => n_3028, QN => 
                           DataPath_RF_bus_reg_dataout_1426_port);
   DataPath_RF_BLOCKi_53_Q_reg_18_inst : DFF_X1 port map( D => n5060, CK => CLK
                           , Q => n_3029, QN => 
                           DataPath_RF_bus_reg_dataout_1458_port);
   DataPath_RF_BLOCKi_54_Q_reg_18_inst : DFF_X1 port map( D => n5095, CK => CLK
                           , Q => n_3030, QN => 
                           DataPath_RF_bus_reg_dataout_1490_port);
   DataPath_RF_BLOCKi_55_Q_reg_18_inst : DFF_X1 port map( D => n5130, CK => CLK
                           , Q => n_3031, QN => 
                           DataPath_RF_bus_reg_dataout_1522_port);
   DataPath_RF_BLOCKi_56_Q_reg_18_inst : DFF_X1 port map( D => n5178, CK => CLK
                           , Q => n_3032, QN => 
                           DataPath_RF_bus_reg_dataout_1554_port);
   DataPath_RF_BLOCKi_57_Q_reg_18_inst : DFF_X1 port map( D => n5232, CK => CLK
                           , Q => n_3033, QN => 
                           DataPath_RF_bus_reg_dataout_1586_port);
   DataPath_RF_BLOCKi_58_Q_reg_18_inst : DFF_X1 port map( D => n5268, CK => CLK
                           , Q => n_3034, QN => 
                           DataPath_RF_bus_reg_dataout_1618_port);
   DataPath_RF_BLOCKi_59_Q_reg_18_inst : DFF_X1 port map( D => n5303, CK => CLK
                           , Q => n_3035, QN => 
                           DataPath_RF_bus_reg_dataout_1650_port);
   DataPath_RF_BLOCKi_60_Q_reg_18_inst : DFF_X1 port map( D => n5338, CK => CLK
                           , Q => n_3036, QN => 
                           DataPath_RF_bus_reg_dataout_1682_port);
   DataPath_RF_BLOCKi_61_Q_reg_18_inst : DFF_X1 port map( D => n5373, CK => CLK
                           , Q => n_3037, QN => 
                           DataPath_RF_bus_reg_dataout_1714_port);
   DataPath_RF_BLOCKi_62_Q_reg_18_inst : DFF_X1 port map( D => n5408, CK => CLK
                           , Q => n_3038, QN => 
                           DataPath_RF_bus_reg_dataout_1746_port);
   DataPath_RF_BLOCKi_63_Q_reg_18_inst : DFF_X1 port map( D => n5443, CK => CLK
                           , Q => n_3039, QN => 
                           DataPath_RF_bus_reg_dataout_1778_port);
   DataPath_RF_BLOCKi_64_Q_reg_18_inst : DFF_X1 port map( D => n5478, CK => CLK
                           , Q => n_3040, QN => 
                           DataPath_RF_bus_reg_dataout_1810_port);
   DataPath_RF_BLOCKi_65_Q_reg_18_inst : DFF_X1 port map( D => n5513, CK => CLK
                           , Q => n_3041, QN => 
                           DataPath_RF_bus_reg_dataout_1842_port);
   DataPath_RF_BLOCKi_66_Q_reg_18_inst : DFF_X1 port map( D => n5548, CK => CLK
                           , Q => n_3042, QN => 
                           DataPath_RF_bus_reg_dataout_1874_port);
   DataPath_RF_BLOCKi_67_Q_reg_18_inst : DFF_X1 port map( D => n5583, CK => CLK
                           , Q => n_3043, QN => 
                           DataPath_RF_bus_reg_dataout_1906_port);
   DataPath_RF_BLOCKi_68_Q_reg_18_inst : DFF_X1 port map( D => n5622, CK => CLK
                           , Q => n_3044, QN => 
                           DataPath_RF_bus_reg_dataout_1938_port);
   DataPath_RF_BLOCKi_69_Q_reg_18_inst : DFF_X1 port map( D => n5659, CK => CLK
                           , Q => n_3045, QN => 
                           DataPath_RF_bus_reg_dataout_1970_port);
   DataPath_RF_BLOCKi_70_Q_reg_18_inst : DFF_X1 port map( D => n5696, CK => CLK
                           , Q => n_3046, QN => 
                           DataPath_RF_bus_reg_dataout_2002_port);
   DataPath_RF_BLOCKi_71_Q_reg_18_inst : DFF_X1 port map( D => n5733, CK => CLK
                           , Q => n_3047, QN => 
                           DataPath_RF_bus_reg_dataout_2034_port);
   DataPath_RF_BLOCKi_83_Q_reg_18_inst : DFF_X1 port map( D => n942, CK => CLK,
                           Q => n_3048, QN => 
                           DataPath_RF_bus_reg_dataout_2418_port);
   DataPath_RF_BLOCKi_84_Q_reg_18_inst : DFF_X1 port map( D => n983, CK => CLK,
                           Q => n_3049, QN => 
                           DataPath_RF_bus_reg_dataout_2450_port);
   DataPath_RF_BLOCKi_85_Q_reg_18_inst : DFF_X1 port map( D => n1020, CK => CLK
                           , Q => n_3050, QN => 
                           DataPath_RF_bus_reg_dataout_2482_port);
   DataPath_RF_BLOCKi_86_Q_reg_18_inst : DFF_X1 port map( D => n1057, CK => CLK
                           , Q => n_3051, QN => 
                           DataPath_RF_bus_reg_dataout_2514_port);
   DataPath_RF_BLOCKi_87_Q_reg_18_inst : DFF_X1 port map( D => n1094, CK => CLK
                           , Q => n_3052, QN => 
                           DataPath_RF_bus_reg_dataout_2546_port);
   DataPath_RF_BLOCKi_72_Q_reg_18_inst : DFF_X1 port map( D => n5770, CK => CLK
                           , Q => n_3053, QN => 
                           DataPath_RF_bus_reg_dataout_2066_port);
   DataPath_RF_BLOCKi_73_Q_reg_18_inst : DFF_X1 port map( D => n5809, CK => CLK
                           , Q => n_3054, QN => 
                           DataPath_RF_bus_reg_dataout_2098_port);
   DataPath_RF_BLOCKi_74_Q_reg_18_inst : DFF_X1 port map( D => n5845, CK => CLK
                           , Q => n_3055, QN => 
                           DataPath_RF_bus_reg_dataout_2130_port);
   DataPath_RF_BLOCKi_75_Q_reg_18_inst : DFF_X1 port map( D => n5881, CK => CLK
                           , Q => n_3056, QN => 
                           DataPath_RF_bus_reg_dataout_2162_port);
   DataPath_RF_BLOCKi_76_Q_reg_18_inst : DFF_X1 port map( D => n5917, CK => CLK
                           , Q => n_3057, QN => 
                           DataPath_RF_bus_reg_dataout_2194_port);
   DataPath_RF_BLOCKi_77_Q_reg_18_inst : DFF_X1 port map( D => n5953, CK => CLK
                           , Q => n_3058, QN => 
                           DataPath_RF_bus_reg_dataout_2226_port);
   DataPath_RF_BLOCKi_78_Q_reg_18_inst : DFF_X1 port map( D => n5989, CK => CLK
                           , Q => n_3059, QN => 
                           DataPath_RF_bus_reg_dataout_2258_port);
   DataPath_RF_BLOCKi_79_Q_reg_18_inst : DFF_X1 port map( D => n6025, CK => CLK
                           , Q => n_3060, QN => 
                           DataPath_RF_bus_reg_dataout_2290_port);
   DataPath_RF_BLOCKi_80_Q_reg_18_inst : DFF_X1 port map( D => n6062, CK => CLK
                           , Q => n_3061, QN => 
                           DataPath_RF_bus_reg_dataout_2322_port);
   DataPath_RF_BLOCKi_81_Q_reg_18_inst : DFF_X1 port map( D => n6098, CK => CLK
                           , Q => n_3062, QN => 
                           DataPath_RF_bus_reg_dataout_2354_port);
   DataPath_RF_BLOCKi_82_Q_reg_18_inst : DFF_X1 port map( D => n6132, CK => CLK
                           , Q => n_3063, QN => 
                           DataPath_RF_bus_reg_dataout_2386_port);
   DataPath_REG_ALU_OUT_Q_reg_19_inst : DFF_X1 port map( D => n7004, CK => CLK,
                           Q => DRAM_ADDRESS_19_port, QN => n506);
   DataPath_REG_MEM_ALUOUT_Q_reg_19_inst : DFF_X1 port map( D => n1130, CK => 
                           CLK, Q => n_3064, QN => 
                           DataPath_i_REG_MEM_ALUOUT_19_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_19_inst : DFF_X1 port map( D => n6780, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_51_port,
                           QN => n618);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_19_inst : DFF_X1 port map( D => n6812, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_83_port,
                           QN => n650);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_19_inst : DFF_X1 port map( D => n6844, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_115_port
                           , QN => n682);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_19_inst : DFF_X1 port map( D => n6876, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_147_port
                           , QN => n714);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_19_inst : DFF_X1 port map( D => n6908, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_179_port
                           , QN => n746);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_19_inst : DFF_X1 port map( D => n6940, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_211_port
                           , QN => n778);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_19_inst : DFF_X1 port map( D => n6972, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_243_port
                           , QN => n810);
   DataPath_RF_BLOCKi_8_Q_reg_19_inst : DFF_X1 port map( D => n3334, CK => CLK,
                           Q => n_3065, QN => 
                           DataPath_RF_bus_reg_dataout_19_port);
   DataPath_RF_BLOCKi_9_Q_reg_19_inst : DFF_X1 port map( D => n3393, CK => CLK,
                           Q => n_3066, QN => 
                           DataPath_RF_bus_reg_dataout_51_port);
   DataPath_RF_BLOCKi_10_Q_reg_19_inst : DFF_X1 port map( D => n3431, CK => CLK
                           , Q => n_3067, QN => 
                           DataPath_RF_bus_reg_dataout_83_port);
   DataPath_RF_BLOCKi_11_Q_reg_19_inst : DFF_X1 port map( D => n3469, CK => CLK
                           , Q => n_3068, QN => 
                           DataPath_RF_bus_reg_dataout_115_port);
   DataPath_RF_BLOCKi_12_Q_reg_19_inst : DFF_X1 port map( D => n3507, CK => CLK
                           , Q => n_3069, QN => 
                           DataPath_RF_bus_reg_dataout_147_port);
   DataPath_RF_BLOCKi_13_Q_reg_19_inst : DFF_X1 port map( D => n3545, CK => CLK
                           , Q => n_3070, QN => 
                           DataPath_RF_bus_reg_dataout_179_port);
   DataPath_RF_BLOCKi_14_Q_reg_19_inst : DFF_X1 port map( D => n3583, CK => CLK
                           , Q => n_3071, QN => 
                           DataPath_RF_bus_reg_dataout_211_port);
   DataPath_RF_BLOCKi_15_Q_reg_19_inst : DFF_X1 port map( D => n3621, CK => CLK
                           , Q => n_3072, QN => 
                           DataPath_RF_bus_reg_dataout_243_port);
   DataPath_RF_BLOCKi_16_Q_reg_19_inst : DFF_X1 port map( D => n3659, CK => CLK
                           , Q => n_3073, QN => 
                           DataPath_RF_bus_reg_dataout_275_port);
   DataPath_RF_BLOCKi_17_Q_reg_19_inst : DFF_X1 port map( D => n3696, CK => CLK
                           , Q => n_3074, QN => 
                           DataPath_RF_bus_reg_dataout_307_port);
   DataPath_RF_BLOCKi_18_Q_reg_19_inst : DFF_X1 port map( D => n3733, CK => CLK
                           , Q => n_3075, QN => 
                           DataPath_RF_bus_reg_dataout_339_port);
   DataPath_RF_BLOCKi_19_Q_reg_19_inst : DFF_X1 port map( D => n3770, CK => CLK
                           , Q => n_3076, QN => 
                           DataPath_RF_bus_reg_dataout_371_port);
   DataPath_RF_BLOCKi_20_Q_reg_19_inst : DFF_X1 port map( D => n3805, CK => CLK
                           , Q => n_3077, QN => 
                           DataPath_RF_bus_reg_dataout_403_port);
   DataPath_RF_BLOCKi_21_Q_reg_19_inst : DFF_X1 port map( D => n3840, CK => CLK
                           , Q => n_3078, QN => 
                           DataPath_RF_bus_reg_dataout_435_port);
   DataPath_RF_BLOCKi_22_Q_reg_19_inst : DFF_X1 port map( D => n3875, CK => CLK
                           , Q => n_3079, QN => 
                           DataPath_RF_bus_reg_dataout_467_port);
   DataPath_RF_BLOCKi_23_Q_reg_19_inst : DFF_X1 port map( D => n3922, CK => CLK
                           , Q => n_3080, QN => 
                           DataPath_RF_bus_reg_dataout_499_port);
   DataPath_RF_BLOCKi_24_Q_reg_19_inst : DFF_X1 port map( D => n3990, CK => CLK
                           , Q => n_3081, QN => 
                           DataPath_RF_bus_reg_dataout_531_port);
   DataPath_RF_BLOCKi_25_Q_reg_19_inst : DFF_X1 port map( D => n4046, CK => CLK
                           , Q => n_3082, QN => 
                           DataPath_RF_bus_reg_dataout_563_port);
   DataPath_RF_BLOCKi_26_Q_reg_19_inst : DFF_X1 port map( D => n4081, CK => CLK
                           , Q => n_3083, QN => 
                           DataPath_RF_bus_reg_dataout_595_port);
   DataPath_RF_BLOCKi_27_Q_reg_19_inst : DFF_X1 port map( D => n4116, CK => CLK
                           , Q => n_3084, QN => 
                           DataPath_RF_bus_reg_dataout_627_port);
   DataPath_RF_BLOCKi_28_Q_reg_19_inst : DFF_X1 port map( D => n4151, CK => CLK
                           , Q => n_3085, QN => 
                           DataPath_RF_bus_reg_dataout_659_port);
   DataPath_RF_BLOCKi_29_Q_reg_19_inst : DFF_X1 port map( D => n4186, CK => CLK
                           , Q => n_3086, QN => 
                           DataPath_RF_bus_reg_dataout_691_port);
   DataPath_RF_BLOCKi_30_Q_reg_19_inst : DFF_X1 port map( D => n4221, CK => CLK
                           , Q => n_3087, QN => 
                           DataPath_RF_bus_reg_dataout_723_port);
   DataPath_RF_BLOCKi_31_Q_reg_19_inst : DFF_X1 port map( D => n4256, CK => CLK
                           , Q => n_3088, QN => 
                           DataPath_RF_bus_reg_dataout_755_port);
   DataPath_RF_BLOCKi_32_Q_reg_19_inst : DFF_X1 port map( D => n4291, CK => CLK
                           , Q => n_3089, QN => 
                           DataPath_RF_bus_reg_dataout_787_port);
   DataPath_RF_BLOCKi_33_Q_reg_19_inst : DFF_X1 port map( D => n4326, CK => CLK
                           , Q => n_3090, QN => 
                           DataPath_RF_bus_reg_dataout_819_port);
   DataPath_RF_BLOCKi_34_Q_reg_19_inst : DFF_X1 port map( D => n4361, CK => CLK
                           , Q => n_3091, QN => 
                           DataPath_RF_bus_reg_dataout_851_port);
   DataPath_RF_BLOCKi_35_Q_reg_19_inst : DFF_X1 port map( D => n4396, CK => CLK
                           , Q => n_3092, QN => 
                           DataPath_RF_bus_reg_dataout_883_port);
   DataPath_RF_BLOCKi_36_Q_reg_19_inst : DFF_X1 port map( D => n4431, CK => CLK
                           , Q => n_3093, QN => 
                           DataPath_RF_bus_reg_dataout_915_port);
   DataPath_RF_BLOCKi_37_Q_reg_19_inst : DFF_X1 port map( D => n4466, CK => CLK
                           , Q => n_3094, QN => 
                           DataPath_RF_bus_reg_dataout_947_port);
   DataPath_RF_BLOCKi_38_Q_reg_19_inst : DFF_X1 port map( D => n4501, CK => CLK
                           , Q => n_3095, QN => 
                           DataPath_RF_bus_reg_dataout_979_port);
   DataPath_RF_BLOCKi_39_Q_reg_19_inst : DFF_X1 port map( D => n4536, CK => CLK
                           , Q => n_3096, QN => 
                           DataPath_RF_bus_reg_dataout_1011_port);
   DataPath_RF_BLOCKi_40_Q_reg_19_inst : DFF_X1 port map( D => n4583, CK => CLK
                           , Q => n_3097, QN => 
                           DataPath_RF_bus_reg_dataout_1043_port);
   DataPath_RF_BLOCKi_41_Q_reg_19_inst : DFF_X1 port map( D => n4639, CK => CLK
                           , Q => n_3098, QN => 
                           DataPath_RF_bus_reg_dataout_1075_port);
   DataPath_RF_BLOCKi_42_Q_reg_19_inst : DFF_X1 port map( D => n4674, CK => CLK
                           , Q => n_3099, QN => 
                           DataPath_RF_bus_reg_dataout_1107_port);
   DataPath_RF_BLOCKi_43_Q_reg_19_inst : DFF_X1 port map( D => n4709, CK => CLK
                           , Q => n_3100, QN => 
                           DataPath_RF_bus_reg_dataout_1139_port);
   DataPath_RF_BLOCKi_44_Q_reg_19_inst : DFF_X1 port map( D => n4744, CK => CLK
                           , Q => n_3101, QN => 
                           DataPath_RF_bus_reg_dataout_1171_port);
   DataPath_RF_BLOCKi_45_Q_reg_19_inst : DFF_X1 port map( D => n4779, CK => CLK
                           , Q => n_3102, QN => 
                           DataPath_RF_bus_reg_dataout_1203_port);
   DataPath_RF_BLOCKi_46_Q_reg_19_inst : DFF_X1 port map( D => n4814, CK => CLK
                           , Q => n_3103, QN => 
                           DataPath_RF_bus_reg_dataout_1235_port);
   DataPath_RF_BLOCKi_47_Q_reg_19_inst : DFF_X1 port map( D => n4849, CK => CLK
                           , Q => n_3104, QN => 
                           DataPath_RF_bus_reg_dataout_1267_port);
   DataPath_RF_BLOCKi_48_Q_reg_19_inst : DFF_X1 port map( D => n4884, CK => CLK
                           , Q => n_3105, QN => 
                           DataPath_RF_bus_reg_dataout_1299_port);
   DataPath_RF_BLOCKi_49_Q_reg_19_inst : DFF_X1 port map( D => n4919, CK => CLK
                           , Q => n_3106, QN => 
                           DataPath_RF_bus_reg_dataout_1331_port);
   DataPath_RF_BLOCKi_50_Q_reg_19_inst : DFF_X1 port map( D => n4954, CK => CLK
                           , Q => n_3107, QN => 
                           DataPath_RF_bus_reg_dataout_1363_port);
   DataPath_RF_BLOCKi_51_Q_reg_19_inst : DFF_X1 port map( D => n4989, CK => CLK
                           , Q => n_3108, QN => 
                           DataPath_RF_bus_reg_dataout_1395_port);
   DataPath_RF_BLOCKi_52_Q_reg_19_inst : DFF_X1 port map( D => n5024, CK => CLK
                           , Q => n_3109, QN => 
                           DataPath_RF_bus_reg_dataout_1427_port);
   DataPath_RF_BLOCKi_53_Q_reg_19_inst : DFF_X1 port map( D => n5059, CK => CLK
                           , Q => n_3110, QN => 
                           DataPath_RF_bus_reg_dataout_1459_port);
   DataPath_RF_BLOCKi_54_Q_reg_19_inst : DFF_X1 port map( D => n5094, CK => CLK
                           , Q => n_3111, QN => 
                           DataPath_RF_bus_reg_dataout_1491_port);
   DataPath_RF_BLOCKi_55_Q_reg_19_inst : DFF_X1 port map( D => n5129, CK => CLK
                           , Q => n_3112, QN => 
                           DataPath_RF_bus_reg_dataout_1523_port);
   DataPath_RF_BLOCKi_56_Q_reg_19_inst : DFF_X1 port map( D => n5176, CK => CLK
                           , Q => n_3113, QN => 
                           DataPath_RF_bus_reg_dataout_1555_port);
   DataPath_RF_BLOCKi_57_Q_reg_19_inst : DFF_X1 port map( D => n5231, CK => CLK
                           , Q => n_3114, QN => 
                           DataPath_RF_bus_reg_dataout_1587_port);
   DataPath_RF_BLOCKi_58_Q_reg_19_inst : DFF_X1 port map( D => n5267, CK => CLK
                           , Q => n_3115, QN => 
                           DataPath_RF_bus_reg_dataout_1619_port);
   DataPath_RF_BLOCKi_59_Q_reg_19_inst : DFF_X1 port map( D => n5302, CK => CLK
                           , Q => n_3116, QN => 
                           DataPath_RF_bus_reg_dataout_1651_port);
   DataPath_RF_BLOCKi_60_Q_reg_19_inst : DFF_X1 port map( D => n5337, CK => CLK
                           , Q => n_3117, QN => 
                           DataPath_RF_bus_reg_dataout_1683_port);
   DataPath_RF_BLOCKi_61_Q_reg_19_inst : DFF_X1 port map( D => n5372, CK => CLK
                           , Q => n_3118, QN => 
                           DataPath_RF_bus_reg_dataout_1715_port);
   DataPath_RF_BLOCKi_62_Q_reg_19_inst : DFF_X1 port map( D => n5407, CK => CLK
                           , Q => n_3119, QN => 
                           DataPath_RF_bus_reg_dataout_1747_port);
   DataPath_RF_BLOCKi_63_Q_reg_19_inst : DFF_X1 port map( D => n5442, CK => CLK
                           , Q => n_3120, QN => 
                           DataPath_RF_bus_reg_dataout_1779_port);
   DataPath_RF_BLOCKi_64_Q_reg_19_inst : DFF_X1 port map( D => n5477, CK => CLK
                           , Q => n_3121, QN => 
                           DataPath_RF_bus_reg_dataout_1811_port);
   DataPath_RF_BLOCKi_65_Q_reg_19_inst : DFF_X1 port map( D => n5512, CK => CLK
                           , Q => n_3122, QN => 
                           DataPath_RF_bus_reg_dataout_1843_port);
   DataPath_RF_BLOCKi_66_Q_reg_19_inst : DFF_X1 port map( D => n5547, CK => CLK
                           , Q => n_3123, QN => 
                           DataPath_RF_bus_reg_dataout_1875_port);
   DataPath_RF_BLOCKi_67_Q_reg_19_inst : DFF_X1 port map( D => n5582, CK => CLK
                           , Q => n_3124, QN => 
                           DataPath_RF_bus_reg_dataout_1907_port);
   DataPath_RF_BLOCKi_68_Q_reg_19_inst : DFF_X1 port map( D => n5621, CK => CLK
                           , Q => n_3125, QN => 
                           DataPath_RF_bus_reg_dataout_1939_port);
   DataPath_RF_BLOCKi_69_Q_reg_19_inst : DFF_X1 port map( D => n5658, CK => CLK
                           , Q => n_3126, QN => 
                           DataPath_RF_bus_reg_dataout_1971_port);
   DataPath_RF_BLOCKi_70_Q_reg_19_inst : DFF_X1 port map( D => n5695, CK => CLK
                           , Q => n_3127, QN => 
                           DataPath_RF_bus_reg_dataout_2003_port);
   DataPath_RF_BLOCKi_71_Q_reg_19_inst : DFF_X1 port map( D => n5732, CK => CLK
                           , Q => n_3128, QN => 
                           DataPath_RF_bus_reg_dataout_2035_port);
   DataPath_RF_BLOCKi_83_Q_reg_19_inst : DFF_X1 port map( D => n940, CK => CLK,
                           Q => n_3129, QN => 
                           DataPath_RF_bus_reg_dataout_2419_port);
   DataPath_RF_BLOCKi_84_Q_reg_19_inst : DFF_X1 port map( D => n982, CK => CLK,
                           Q => n_3130, QN => 
                           DataPath_RF_bus_reg_dataout_2451_port);
   DataPath_RF_BLOCKi_85_Q_reg_19_inst : DFF_X1 port map( D => n1019, CK => CLK
                           , Q => n_3131, QN => 
                           DataPath_RF_bus_reg_dataout_2483_port);
   DataPath_RF_BLOCKi_86_Q_reg_19_inst : DFF_X1 port map( D => n1056, CK => CLK
                           , Q => n_3132, QN => 
                           DataPath_RF_bus_reg_dataout_2515_port);
   DataPath_RF_BLOCKi_87_Q_reg_19_inst : DFF_X1 port map( D => n1093, CK => CLK
                           , Q => n_3133, QN => 
                           DataPath_RF_bus_reg_dataout_2547_port);
   DataPath_RF_BLOCKi_72_Q_reg_19_inst : DFF_X1 port map( D => n5769, CK => CLK
                           , Q => n_3134, QN => 
                           DataPath_RF_bus_reg_dataout_2067_port);
   DataPath_RF_BLOCKi_73_Q_reg_19_inst : DFF_X1 port map( D => n5808, CK => CLK
                           , Q => n_3135, QN => 
                           DataPath_RF_bus_reg_dataout_2099_port);
   DataPath_RF_BLOCKi_74_Q_reg_19_inst : DFF_X1 port map( D => n5844, CK => CLK
                           , Q => n_3136, QN => 
                           DataPath_RF_bus_reg_dataout_2131_port);
   DataPath_RF_BLOCKi_75_Q_reg_19_inst : DFF_X1 port map( D => n5880, CK => CLK
                           , Q => n_3137, QN => 
                           DataPath_RF_bus_reg_dataout_2163_port);
   DataPath_RF_BLOCKi_76_Q_reg_19_inst : DFF_X1 port map( D => n5916, CK => CLK
                           , Q => n_3138, QN => 
                           DataPath_RF_bus_reg_dataout_2195_port);
   DataPath_RF_BLOCKi_77_Q_reg_19_inst : DFF_X1 port map( D => n5952, CK => CLK
                           , Q => n_3139, QN => 
                           DataPath_RF_bus_reg_dataout_2227_port);
   DataPath_RF_BLOCKi_78_Q_reg_19_inst : DFF_X1 port map( D => n5988, CK => CLK
                           , Q => n_3140, QN => 
                           DataPath_RF_bus_reg_dataout_2259_port);
   DataPath_RF_BLOCKi_79_Q_reg_19_inst : DFF_X1 port map( D => n6024, CK => CLK
                           , Q => n_3141, QN => 
                           DataPath_RF_bus_reg_dataout_2291_port);
   DataPath_RF_BLOCKi_80_Q_reg_19_inst : DFF_X1 port map( D => n6061, CK => CLK
                           , Q => n_3142, QN => 
                           DataPath_RF_bus_reg_dataout_2323_port);
   DataPath_RF_BLOCKi_81_Q_reg_19_inst : DFF_X1 port map( D => n6097, CK => CLK
                           , Q => n_3143, QN => 
                           DataPath_RF_bus_reg_dataout_2355_port);
   DataPath_RF_BLOCKi_82_Q_reg_19_inst : DFF_X1 port map( D => n6131, CK => CLK
                           , Q => n_3144, QN => 
                           DataPath_RF_bus_reg_dataout_2387_port);
   DataPath_REG_ALU_OUT_Q_reg_20_inst : DFF_X1 port map( D => n7003, CK => CLK,
                           Q => DRAM_ADDRESS_20_port, QN => n507);
   DataPath_REG_MEM_ALUOUT_Q_reg_20_inst : DFF_X1 port map( D => n1129, CK => 
                           CLK, Q => n_3145, QN => 
                           DataPath_i_REG_MEM_ALUOUT_20_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_20_inst : DFF_X1 port map( D => n6779, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_52_port,
                           QN => n619);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_20_inst : DFF_X1 port map( D => n6811, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_84_port,
                           QN => n651);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_20_inst : DFF_X1 port map( D => n6843, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_116_port
                           , QN => n683);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_20_inst : DFF_X1 port map( D => n6875, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_148_port
                           , QN => n715);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_20_inst : DFF_X1 port map( D => n6907, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_180_port
                           , QN => n747);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_20_inst : DFF_X1 port map( D => n6939, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_212_port
                           , QN => n779);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_20_inst : DFF_X1 port map( D => n6971, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_244_port
                           , QN => n811);
   DataPath_RF_BLOCKi_8_Q_reg_20_inst : DFF_X1 port map( D => n3332, CK => CLK,
                           Q => n_3146, QN => 
                           DataPath_RF_bus_reg_dataout_20_port);
   DataPath_RF_BLOCKi_9_Q_reg_20_inst : DFF_X1 port map( D => n3392, CK => CLK,
                           Q => n_3147, QN => 
                           DataPath_RF_bus_reg_dataout_52_port);
   DataPath_RF_BLOCKi_10_Q_reg_20_inst : DFF_X1 port map( D => n3430, CK => CLK
                           , Q => n_3148, QN => 
                           DataPath_RF_bus_reg_dataout_84_port);
   DataPath_RF_BLOCKi_11_Q_reg_20_inst : DFF_X1 port map( D => n3468, CK => CLK
                           , Q => n_3149, QN => 
                           DataPath_RF_bus_reg_dataout_116_port);
   DataPath_RF_BLOCKi_12_Q_reg_20_inst : DFF_X1 port map( D => n3506, CK => CLK
                           , Q => n_3150, QN => 
                           DataPath_RF_bus_reg_dataout_148_port);
   DataPath_RF_BLOCKi_13_Q_reg_20_inst : DFF_X1 port map( D => n3544, CK => CLK
                           , Q => n_3151, QN => 
                           DataPath_RF_bus_reg_dataout_180_port);
   DataPath_RF_BLOCKi_14_Q_reg_20_inst : DFF_X1 port map( D => n3582, CK => CLK
                           , Q => n_3152, QN => 
                           DataPath_RF_bus_reg_dataout_212_port);
   DataPath_RF_BLOCKi_15_Q_reg_20_inst : DFF_X1 port map( D => n3620, CK => CLK
                           , Q => n_3153, QN => 
                           DataPath_RF_bus_reg_dataout_244_port);
   DataPath_RF_BLOCKi_16_Q_reg_20_inst : DFF_X1 port map( D => n3658, CK => CLK
                           , Q => n_3154, QN => 
                           DataPath_RF_bus_reg_dataout_276_port);
   DataPath_RF_BLOCKi_17_Q_reg_20_inst : DFF_X1 port map( D => n3695, CK => CLK
                           , Q => n_3155, QN => 
                           DataPath_RF_bus_reg_dataout_308_port);
   DataPath_RF_BLOCKi_18_Q_reg_20_inst : DFF_X1 port map( D => n3732, CK => CLK
                           , Q => n_3156, QN => 
                           DataPath_RF_bus_reg_dataout_340_port);
   DataPath_RF_BLOCKi_19_Q_reg_20_inst : DFF_X1 port map( D => n3769, CK => CLK
                           , Q => n_3157, QN => 
                           DataPath_RF_bus_reg_dataout_372_port);
   DataPath_RF_BLOCKi_20_Q_reg_20_inst : DFF_X1 port map( D => n3804, CK => CLK
                           , Q => n_3158, QN => 
                           DataPath_RF_bus_reg_dataout_404_port);
   DataPath_RF_BLOCKi_21_Q_reg_20_inst : DFF_X1 port map( D => n3839, CK => CLK
                           , Q => n_3159, QN => 
                           DataPath_RF_bus_reg_dataout_436_port);
   DataPath_RF_BLOCKi_22_Q_reg_20_inst : DFF_X1 port map( D => n3874, CK => CLK
                           , Q => n_3160, QN => 
                           DataPath_RF_bus_reg_dataout_468_port);
   DataPath_RF_BLOCKi_23_Q_reg_20_inst : DFF_X1 port map( D => n3920, CK => CLK
                           , Q => n_3161, QN => 
                           DataPath_RF_bus_reg_dataout_500_port);
   DataPath_RF_BLOCKi_24_Q_reg_20_inst : DFF_X1 port map( D => n3988, CK => CLK
                           , Q => n_3162, QN => 
                           DataPath_RF_bus_reg_dataout_532_port);
   DataPath_RF_BLOCKi_25_Q_reg_20_inst : DFF_X1 port map( D => n4045, CK => CLK
                           , Q => n_3163, QN => 
                           DataPath_RF_bus_reg_dataout_564_port);
   DataPath_RF_BLOCKi_26_Q_reg_20_inst : DFF_X1 port map( D => n4080, CK => CLK
                           , Q => n_3164, QN => 
                           DataPath_RF_bus_reg_dataout_596_port);
   DataPath_RF_BLOCKi_27_Q_reg_20_inst : DFF_X1 port map( D => n4115, CK => CLK
                           , Q => n_3165, QN => 
                           DataPath_RF_bus_reg_dataout_628_port);
   DataPath_RF_BLOCKi_28_Q_reg_20_inst : DFF_X1 port map( D => n4150, CK => CLK
                           , Q => n_3166, QN => 
                           DataPath_RF_bus_reg_dataout_660_port);
   DataPath_RF_BLOCKi_29_Q_reg_20_inst : DFF_X1 port map( D => n4185, CK => CLK
                           , Q => n_3167, QN => 
                           DataPath_RF_bus_reg_dataout_692_port);
   DataPath_RF_BLOCKi_30_Q_reg_20_inst : DFF_X1 port map( D => n4220, CK => CLK
                           , Q => n_3168, QN => 
                           DataPath_RF_bus_reg_dataout_724_port);
   DataPath_RF_BLOCKi_31_Q_reg_20_inst : DFF_X1 port map( D => n4255, CK => CLK
                           , Q => n_3169, QN => 
                           DataPath_RF_bus_reg_dataout_756_port);
   DataPath_RF_BLOCKi_32_Q_reg_20_inst : DFF_X1 port map( D => n4290, CK => CLK
                           , Q => n_3170, QN => 
                           DataPath_RF_bus_reg_dataout_788_port);
   DataPath_RF_BLOCKi_33_Q_reg_20_inst : DFF_X1 port map( D => n4325, CK => CLK
                           , Q => n_3171, QN => 
                           DataPath_RF_bus_reg_dataout_820_port);
   DataPath_RF_BLOCKi_34_Q_reg_20_inst : DFF_X1 port map( D => n4360, CK => CLK
                           , Q => n_3172, QN => 
                           DataPath_RF_bus_reg_dataout_852_port);
   DataPath_RF_BLOCKi_35_Q_reg_20_inst : DFF_X1 port map( D => n4395, CK => CLK
                           , Q => n_3173, QN => 
                           DataPath_RF_bus_reg_dataout_884_port);
   DataPath_RF_BLOCKi_36_Q_reg_20_inst : DFF_X1 port map( D => n4430, CK => CLK
                           , Q => n_3174, QN => 
                           DataPath_RF_bus_reg_dataout_916_port);
   DataPath_RF_BLOCKi_37_Q_reg_20_inst : DFF_X1 port map( D => n4465, CK => CLK
                           , Q => n_3175, QN => 
                           DataPath_RF_bus_reg_dataout_948_port);
   DataPath_RF_BLOCKi_38_Q_reg_20_inst : DFF_X1 port map( D => n4500, CK => CLK
                           , Q => n_3176, QN => 
                           DataPath_RF_bus_reg_dataout_980_port);
   DataPath_RF_BLOCKi_39_Q_reg_20_inst : DFF_X1 port map( D => n4535, CK => CLK
                           , Q => n_3177, QN => 
                           DataPath_RF_bus_reg_dataout_1012_port);
   DataPath_RF_BLOCKi_40_Q_reg_20_inst : DFF_X1 port map( D => n4581, CK => CLK
                           , Q => n_3178, QN => 
                           DataPath_RF_bus_reg_dataout_1044_port);
   DataPath_RF_BLOCKi_41_Q_reg_20_inst : DFF_X1 port map( D => n4638, CK => CLK
                           , Q => n_3179, QN => 
                           DataPath_RF_bus_reg_dataout_1076_port);
   DataPath_RF_BLOCKi_42_Q_reg_20_inst : DFF_X1 port map( D => n4673, CK => CLK
                           , Q => n_3180, QN => 
                           DataPath_RF_bus_reg_dataout_1108_port);
   DataPath_RF_BLOCKi_43_Q_reg_20_inst : DFF_X1 port map( D => n4708, CK => CLK
                           , Q => n_3181, QN => 
                           DataPath_RF_bus_reg_dataout_1140_port);
   DataPath_RF_BLOCKi_44_Q_reg_20_inst : DFF_X1 port map( D => n4743, CK => CLK
                           , Q => n_3182, QN => 
                           DataPath_RF_bus_reg_dataout_1172_port);
   DataPath_RF_BLOCKi_45_Q_reg_20_inst : DFF_X1 port map( D => n4778, CK => CLK
                           , Q => n_3183, QN => 
                           DataPath_RF_bus_reg_dataout_1204_port);
   DataPath_RF_BLOCKi_46_Q_reg_20_inst : DFF_X1 port map( D => n4813, CK => CLK
                           , Q => n_3184, QN => 
                           DataPath_RF_bus_reg_dataout_1236_port);
   DataPath_RF_BLOCKi_47_Q_reg_20_inst : DFF_X1 port map( D => n4848, CK => CLK
                           , Q => n_3185, QN => 
                           DataPath_RF_bus_reg_dataout_1268_port);
   DataPath_RF_BLOCKi_48_Q_reg_20_inst : DFF_X1 port map( D => n4883, CK => CLK
                           , Q => n_3186, QN => 
                           DataPath_RF_bus_reg_dataout_1300_port);
   DataPath_RF_BLOCKi_49_Q_reg_20_inst : DFF_X1 port map( D => n4918, CK => CLK
                           , Q => n_3187, QN => 
                           DataPath_RF_bus_reg_dataout_1332_port);
   DataPath_RF_BLOCKi_50_Q_reg_20_inst : DFF_X1 port map( D => n4953, CK => CLK
                           , Q => n_3188, QN => 
                           DataPath_RF_bus_reg_dataout_1364_port);
   DataPath_RF_BLOCKi_51_Q_reg_20_inst : DFF_X1 port map( D => n4988, CK => CLK
                           , Q => n_3189, QN => 
                           DataPath_RF_bus_reg_dataout_1396_port);
   DataPath_RF_BLOCKi_52_Q_reg_20_inst : DFF_X1 port map( D => n5023, CK => CLK
                           , Q => n_3190, QN => 
                           DataPath_RF_bus_reg_dataout_1428_port);
   DataPath_RF_BLOCKi_53_Q_reg_20_inst : DFF_X1 port map( D => n5058, CK => CLK
                           , Q => n_3191, QN => 
                           DataPath_RF_bus_reg_dataout_1460_port);
   DataPath_RF_BLOCKi_54_Q_reg_20_inst : DFF_X1 port map( D => n5093, CK => CLK
                           , Q => n_3192, QN => 
                           DataPath_RF_bus_reg_dataout_1492_port);
   DataPath_RF_BLOCKi_55_Q_reg_20_inst : DFF_X1 port map( D => n5128, CK => CLK
                           , Q => n_3193, QN => 
                           DataPath_RF_bus_reg_dataout_1524_port);
   DataPath_RF_BLOCKi_56_Q_reg_20_inst : DFF_X1 port map( D => n5174, CK => CLK
                           , Q => n_3194, QN => 
                           DataPath_RF_bus_reg_dataout_1556_port);
   DataPath_RF_BLOCKi_57_Q_reg_20_inst : DFF_X1 port map( D => n5230, CK => CLK
                           , Q => n_3195, QN => 
                           DataPath_RF_bus_reg_dataout_1588_port);
   DataPath_RF_BLOCKi_58_Q_reg_20_inst : DFF_X1 port map( D => n5266, CK => CLK
                           , Q => n_3196, QN => 
                           DataPath_RF_bus_reg_dataout_1620_port);
   DataPath_RF_BLOCKi_59_Q_reg_20_inst : DFF_X1 port map( D => n5301, CK => CLK
                           , Q => n_3197, QN => 
                           DataPath_RF_bus_reg_dataout_1652_port);
   DataPath_RF_BLOCKi_60_Q_reg_20_inst : DFF_X1 port map( D => n5336, CK => CLK
                           , Q => n_3198, QN => 
                           DataPath_RF_bus_reg_dataout_1684_port);
   DataPath_RF_BLOCKi_61_Q_reg_20_inst : DFF_X1 port map( D => n5371, CK => CLK
                           , Q => n_3199, QN => 
                           DataPath_RF_bus_reg_dataout_1716_port);
   DataPath_RF_BLOCKi_62_Q_reg_20_inst : DFF_X1 port map( D => n5406, CK => CLK
                           , Q => n_3200, QN => 
                           DataPath_RF_bus_reg_dataout_1748_port);
   DataPath_RF_BLOCKi_63_Q_reg_20_inst : DFF_X1 port map( D => n5441, CK => CLK
                           , Q => n_3201, QN => 
                           DataPath_RF_bus_reg_dataout_1780_port);
   DataPath_RF_BLOCKi_64_Q_reg_20_inst : DFF_X1 port map( D => n5476, CK => CLK
                           , Q => n_3202, QN => 
                           DataPath_RF_bus_reg_dataout_1812_port);
   DataPath_RF_BLOCKi_65_Q_reg_20_inst : DFF_X1 port map( D => n5511, CK => CLK
                           , Q => n_3203, QN => 
                           DataPath_RF_bus_reg_dataout_1844_port);
   DataPath_RF_BLOCKi_66_Q_reg_20_inst : DFF_X1 port map( D => n5546, CK => CLK
                           , Q => n_3204, QN => 
                           DataPath_RF_bus_reg_dataout_1876_port);
   DataPath_RF_BLOCKi_67_Q_reg_20_inst : DFF_X1 port map( D => n5581, CK => CLK
                           , Q => n_3205, QN => 
                           DataPath_RF_bus_reg_dataout_1908_port);
   DataPath_RF_BLOCKi_68_Q_reg_20_inst : DFF_X1 port map( D => n5620, CK => CLK
                           , Q => n_3206, QN => 
                           DataPath_RF_bus_reg_dataout_1940_port);
   DataPath_RF_BLOCKi_69_Q_reg_20_inst : DFF_X1 port map( D => n5657, CK => CLK
                           , Q => n_3207, QN => 
                           DataPath_RF_bus_reg_dataout_1972_port);
   DataPath_RF_BLOCKi_70_Q_reg_20_inst : DFF_X1 port map( D => n5694, CK => CLK
                           , Q => n_3208, QN => 
                           DataPath_RF_bus_reg_dataout_2004_port);
   DataPath_RF_BLOCKi_71_Q_reg_20_inst : DFF_X1 port map( D => n5731, CK => CLK
                           , Q => n_3209, QN => 
                           DataPath_RF_bus_reg_dataout_2036_port);
   DataPath_RF_BLOCKi_83_Q_reg_20_inst : DFF_X1 port map( D => n938, CK => CLK,
                           Q => n_3210, QN => 
                           DataPath_RF_bus_reg_dataout_2420_port);
   DataPath_RF_BLOCKi_84_Q_reg_20_inst : DFF_X1 port map( D => n981, CK => CLK,
                           Q => n_3211, QN => 
                           DataPath_RF_bus_reg_dataout_2452_port);
   DataPath_RF_BLOCKi_85_Q_reg_20_inst : DFF_X1 port map( D => n1018, CK => CLK
                           , Q => n_3212, QN => 
                           DataPath_RF_bus_reg_dataout_2484_port);
   DataPath_RF_BLOCKi_86_Q_reg_20_inst : DFF_X1 port map( D => n1055, CK => CLK
                           , Q => n_3213, QN => 
                           DataPath_RF_bus_reg_dataout_2516_port);
   DataPath_RF_BLOCKi_87_Q_reg_20_inst : DFF_X1 port map( D => n1092, CK => CLK
                           , Q => n_3214, QN => 
                           DataPath_RF_bus_reg_dataout_2548_port);
   DataPath_RF_BLOCKi_72_Q_reg_20_inst : DFF_X1 port map( D => n5768, CK => CLK
                           , Q => n_3215, QN => 
                           DataPath_RF_bus_reg_dataout_2068_port);
   DataPath_RF_BLOCKi_73_Q_reg_20_inst : DFF_X1 port map( D => n5807, CK => CLK
                           , Q => n_3216, QN => 
                           DataPath_RF_bus_reg_dataout_2100_port);
   DataPath_RF_BLOCKi_74_Q_reg_20_inst : DFF_X1 port map( D => n5843, CK => CLK
                           , Q => n_3217, QN => 
                           DataPath_RF_bus_reg_dataout_2132_port);
   DataPath_RF_BLOCKi_75_Q_reg_20_inst : DFF_X1 port map( D => n5879, CK => CLK
                           , Q => n_3218, QN => 
                           DataPath_RF_bus_reg_dataout_2164_port);
   DataPath_RF_BLOCKi_76_Q_reg_20_inst : DFF_X1 port map( D => n5915, CK => CLK
                           , Q => n_3219, QN => 
                           DataPath_RF_bus_reg_dataout_2196_port);
   DataPath_RF_BLOCKi_77_Q_reg_20_inst : DFF_X1 port map( D => n5951, CK => CLK
                           , Q => n_3220, QN => 
                           DataPath_RF_bus_reg_dataout_2228_port);
   DataPath_RF_BLOCKi_78_Q_reg_20_inst : DFF_X1 port map( D => n5987, CK => CLK
                           , Q => n_3221, QN => 
                           DataPath_RF_bus_reg_dataout_2260_port);
   DataPath_RF_BLOCKi_79_Q_reg_20_inst : DFF_X1 port map( D => n6023, CK => CLK
                           , Q => n_3222, QN => 
                           DataPath_RF_bus_reg_dataout_2292_port);
   DataPath_RF_BLOCKi_80_Q_reg_20_inst : DFF_X1 port map( D => n6060, CK => CLK
                           , Q => n_3223, QN => 
                           DataPath_RF_bus_reg_dataout_2324_port);
   DataPath_RF_BLOCKi_81_Q_reg_20_inst : DFF_X1 port map( D => n6096, CK => CLK
                           , Q => n_3224, QN => 
                           DataPath_RF_bus_reg_dataout_2356_port);
   DataPath_RF_BLOCKi_82_Q_reg_20_inst : DFF_X1 port map( D => n6130, CK => CLK
                           , Q => n_3225, QN => 
                           DataPath_RF_bus_reg_dataout_2388_port);
   DataPath_REG_ALU_OUT_Q_reg_22_inst : DFF_X1 port map( D => n7001, CK => CLK,
                           Q => DRAM_ADDRESS_22_port, QN => n508);
   DataPath_REG_MEM_ALUOUT_Q_reg_22_inst : DFF_X1 port map( D => n1127, CK => 
                           CLK, Q => n_3226, QN => 
                           DataPath_i_REG_MEM_ALUOUT_22_port);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_22_inst : DFF_X1 port map( D => n6841, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_118_port
                           , QN => n685);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_22_inst : DFF_X1 port map( D => n6873, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_150_port
                           , QN => n717);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_22_inst : DFF_X1 port map( D => n6937, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_214_port
                           , QN => n781);
   DataPath_RF_BLOCKi_8_Q_reg_22_inst : DFF_X1 port map( D => n3328, CK => CLK,
                           Q => n_3227, QN => 
                           DataPath_RF_bus_reg_dataout_22_port);
   DataPath_RF_BLOCKi_9_Q_reg_22_inst : DFF_X1 port map( D => n3390, CK => CLK,
                           Q => n_3228, QN => 
                           DataPath_RF_bus_reg_dataout_54_port);
   DataPath_RF_BLOCKi_10_Q_reg_22_inst : DFF_X1 port map( D => n3428, CK => CLK
                           , Q => n_3229, QN => 
                           DataPath_RF_bus_reg_dataout_86_port);
   DataPath_RF_BLOCKi_11_Q_reg_22_inst : DFF_X1 port map( D => n3466, CK => CLK
                           , Q => n_3230, QN => 
                           DataPath_RF_bus_reg_dataout_118_port);
   DataPath_RF_BLOCKi_12_Q_reg_22_inst : DFF_X1 port map( D => n3504, CK => CLK
                           , Q => n_3231, QN => 
                           DataPath_RF_bus_reg_dataout_150_port);
   DataPath_RF_BLOCKi_13_Q_reg_22_inst : DFF_X1 port map( D => n3542, CK => CLK
                           , Q => n_3232, QN => 
                           DataPath_RF_bus_reg_dataout_182_port);
   DataPath_RF_BLOCKi_14_Q_reg_22_inst : DFF_X1 port map( D => n3580, CK => CLK
                           , Q => n_3233, QN => 
                           DataPath_RF_bus_reg_dataout_214_port);
   DataPath_RF_BLOCKi_15_Q_reg_22_inst : DFF_X1 port map( D => n3618, CK => CLK
                           , Q => n_3234, QN => 
                           DataPath_RF_bus_reg_dataout_246_port);
   DataPath_RF_BLOCKi_16_Q_reg_22_inst : DFF_X1 port map( D => n3656, CK => CLK
                           , Q => n_3235, QN => 
                           DataPath_RF_bus_reg_dataout_278_port);
   DataPath_RF_BLOCKi_17_Q_reg_22_inst : DFF_X1 port map( D => n3693, CK => CLK
                           , Q => n_3236, QN => 
                           DataPath_RF_bus_reg_dataout_310_port);
   DataPath_RF_BLOCKi_18_Q_reg_22_inst : DFF_X1 port map( D => n3730, CK => CLK
                           , Q => n_3237, QN => 
                           DataPath_RF_bus_reg_dataout_342_port);
   DataPath_RF_BLOCKi_19_Q_reg_22_inst : DFF_X1 port map( D => n3767, CK => CLK
                           , Q => n_3238, QN => 
                           DataPath_RF_bus_reg_dataout_374_port);
   DataPath_RF_BLOCKi_20_Q_reg_22_inst : DFF_X1 port map( D => n3802, CK => CLK
                           , Q => n_3239, QN => 
                           DataPath_RF_bus_reg_dataout_406_port);
   DataPath_RF_BLOCKi_21_Q_reg_22_inst : DFF_X1 port map( D => n3837, CK => CLK
                           , Q => n_3240, QN => 
                           DataPath_RF_bus_reg_dataout_438_port);
   DataPath_RF_BLOCKi_22_Q_reg_22_inst : DFF_X1 port map( D => n3872, CK => CLK
                           , Q => n_3241, QN => 
                           DataPath_RF_bus_reg_dataout_470_port);
   DataPath_RF_BLOCKi_23_Q_reg_22_inst : DFF_X1 port map( D => n3916, CK => CLK
                           , Q => n_3242, QN => 
                           DataPath_RF_bus_reg_dataout_502_port);
   DataPath_RF_BLOCKi_24_Q_reg_22_inst : DFF_X1 port map( D => n3984, CK => CLK
                           , Q => n_3243, QN => 
                           DataPath_RF_bus_reg_dataout_534_port);
   DataPath_RF_BLOCKi_25_Q_reg_22_inst : DFF_X1 port map( D => n4043, CK => CLK
                           , Q => n_3244, QN => 
                           DataPath_RF_bus_reg_dataout_566_port);
   DataPath_RF_BLOCKi_26_Q_reg_22_inst : DFF_X1 port map( D => n4078, CK => CLK
                           , Q => n_3245, QN => 
                           DataPath_RF_bus_reg_dataout_598_port);
   DataPath_RF_BLOCKi_27_Q_reg_22_inst : DFF_X1 port map( D => n4113, CK => CLK
                           , Q => n_3246, QN => 
                           DataPath_RF_bus_reg_dataout_630_port);
   DataPath_RF_BLOCKi_28_Q_reg_22_inst : DFF_X1 port map( D => n4148, CK => CLK
                           , Q => n_3247, QN => 
                           DataPath_RF_bus_reg_dataout_662_port);
   DataPath_RF_BLOCKi_29_Q_reg_22_inst : DFF_X1 port map( D => n4183, CK => CLK
                           , Q => n_3248, QN => 
                           DataPath_RF_bus_reg_dataout_694_port);
   DataPath_RF_BLOCKi_30_Q_reg_22_inst : DFF_X1 port map( D => n4218, CK => CLK
                           , Q => n_3249, QN => 
                           DataPath_RF_bus_reg_dataout_726_port);
   DataPath_RF_BLOCKi_31_Q_reg_22_inst : DFF_X1 port map( D => n4253, CK => CLK
                           , Q => n_3250, QN => 
                           DataPath_RF_bus_reg_dataout_758_port);
   DataPath_RF_BLOCKi_32_Q_reg_22_inst : DFF_X1 port map( D => n4288, CK => CLK
                           , Q => n_3251, QN => 
                           DataPath_RF_bus_reg_dataout_790_port);
   DataPath_RF_BLOCKi_33_Q_reg_22_inst : DFF_X1 port map( D => n4323, CK => CLK
                           , Q => n_3252, QN => 
                           DataPath_RF_bus_reg_dataout_822_port);
   DataPath_RF_BLOCKi_34_Q_reg_22_inst : DFF_X1 port map( D => n4358, CK => CLK
                           , Q => n_3253, QN => 
                           DataPath_RF_bus_reg_dataout_854_port);
   DataPath_RF_BLOCKi_35_Q_reg_22_inst : DFF_X1 port map( D => n4393, CK => CLK
                           , Q => n_3254, QN => 
                           DataPath_RF_bus_reg_dataout_886_port);
   DataPath_RF_BLOCKi_36_Q_reg_22_inst : DFF_X1 port map( D => n4428, CK => CLK
                           , Q => n_3255, QN => 
                           DataPath_RF_bus_reg_dataout_918_port);
   DataPath_RF_BLOCKi_37_Q_reg_22_inst : DFF_X1 port map( D => n4463, CK => CLK
                           , Q => n_3256, QN => 
                           DataPath_RF_bus_reg_dataout_950_port);
   DataPath_RF_BLOCKi_38_Q_reg_22_inst : DFF_X1 port map( D => n4498, CK => CLK
                           , Q => n_3257, QN => 
                           DataPath_RF_bus_reg_dataout_982_port);
   DataPath_RF_BLOCKi_39_Q_reg_22_inst : DFF_X1 port map( D => n4533, CK => CLK
                           , Q => n_3258, QN => 
                           DataPath_RF_bus_reg_dataout_1014_port);
   DataPath_RF_BLOCKi_40_Q_reg_22_inst : DFF_X1 port map( D => n4577, CK => CLK
                           , Q => n_3259, QN => 
                           DataPath_RF_bus_reg_dataout_1046_port);
   DataPath_RF_BLOCKi_41_Q_reg_22_inst : DFF_X1 port map( D => n4636, CK => CLK
                           , Q => n_3260, QN => 
                           DataPath_RF_bus_reg_dataout_1078_port);
   DataPath_RF_BLOCKi_42_Q_reg_22_inst : DFF_X1 port map( D => n4671, CK => CLK
                           , Q => n_3261, QN => 
                           DataPath_RF_bus_reg_dataout_1110_port);
   DataPath_RF_BLOCKi_43_Q_reg_22_inst : DFF_X1 port map( D => n4706, CK => CLK
                           , Q => n_3262, QN => 
                           DataPath_RF_bus_reg_dataout_1142_port);
   DataPath_RF_BLOCKi_44_Q_reg_22_inst : DFF_X1 port map( D => n4741, CK => CLK
                           , Q => n_3263, QN => 
                           DataPath_RF_bus_reg_dataout_1174_port);
   DataPath_RF_BLOCKi_45_Q_reg_22_inst : DFF_X1 port map( D => n4776, CK => CLK
                           , Q => n_3264, QN => 
                           DataPath_RF_bus_reg_dataout_1206_port);
   DataPath_RF_BLOCKi_46_Q_reg_22_inst : DFF_X1 port map( D => n4811, CK => CLK
                           , Q => n_3265, QN => 
                           DataPath_RF_bus_reg_dataout_1238_port);
   DataPath_RF_BLOCKi_47_Q_reg_22_inst : DFF_X1 port map( D => n4846, CK => CLK
                           , Q => n_3266, QN => 
                           DataPath_RF_bus_reg_dataout_1270_port);
   DataPath_RF_BLOCKi_48_Q_reg_22_inst : DFF_X1 port map( D => n4881, CK => CLK
                           , Q => n_3267, QN => 
                           DataPath_RF_bus_reg_dataout_1302_port);
   DataPath_RF_BLOCKi_49_Q_reg_22_inst : DFF_X1 port map( D => n4916, CK => CLK
                           , Q => n_3268, QN => 
                           DataPath_RF_bus_reg_dataout_1334_port);
   DataPath_RF_BLOCKi_50_Q_reg_22_inst : DFF_X1 port map( D => n4951, CK => CLK
                           , Q => n_3269, QN => 
                           DataPath_RF_bus_reg_dataout_1366_port);
   DataPath_RF_BLOCKi_51_Q_reg_22_inst : DFF_X1 port map( D => n4986, CK => CLK
                           , Q => n_3270, QN => 
                           DataPath_RF_bus_reg_dataout_1398_port);
   DataPath_RF_BLOCKi_52_Q_reg_22_inst : DFF_X1 port map( D => n5021, CK => CLK
                           , Q => n_3271, QN => 
                           DataPath_RF_bus_reg_dataout_1430_port);
   DataPath_RF_BLOCKi_53_Q_reg_22_inst : DFF_X1 port map( D => n5056, CK => CLK
                           , Q => n_3272, QN => 
                           DataPath_RF_bus_reg_dataout_1462_port);
   DataPath_RF_BLOCKi_54_Q_reg_22_inst : DFF_X1 port map( D => n5091, CK => CLK
                           , Q => n_3273, QN => 
                           DataPath_RF_bus_reg_dataout_1494_port);
   DataPath_RF_BLOCKi_55_Q_reg_22_inst : DFF_X1 port map( D => n5126, CK => CLK
                           , Q => n_3274, QN => 
                           DataPath_RF_bus_reg_dataout_1526_port);
   DataPath_RF_BLOCKi_56_Q_reg_22_inst : DFF_X1 port map( D => n5170, CK => CLK
                           , Q => n_3275, QN => 
                           DataPath_RF_bus_reg_dataout_1558_port);
   DataPath_RF_BLOCKi_57_Q_reg_22_inst : DFF_X1 port map( D => n5228, CK => CLK
                           , Q => n_3276, QN => 
                           DataPath_RF_bus_reg_dataout_1590_port);
   DataPath_RF_BLOCKi_58_Q_reg_22_inst : DFF_X1 port map( D => n5264, CK => CLK
                           , Q => n_3277, QN => 
                           DataPath_RF_bus_reg_dataout_1622_port);
   DataPath_RF_BLOCKi_59_Q_reg_22_inst : DFF_X1 port map( D => n5299, CK => CLK
                           , Q => n_3278, QN => 
                           DataPath_RF_bus_reg_dataout_1654_port);
   DataPath_RF_BLOCKi_60_Q_reg_22_inst : DFF_X1 port map( D => n5334, CK => CLK
                           , Q => n_3279, QN => 
                           DataPath_RF_bus_reg_dataout_1686_port);
   DataPath_RF_BLOCKi_61_Q_reg_22_inst : DFF_X1 port map( D => n5369, CK => CLK
                           , Q => n_3280, QN => 
                           DataPath_RF_bus_reg_dataout_1718_port);
   DataPath_RF_BLOCKi_62_Q_reg_22_inst : DFF_X1 port map( D => n5404, CK => CLK
                           , Q => n_3281, QN => 
                           DataPath_RF_bus_reg_dataout_1750_port);
   DataPath_RF_BLOCKi_63_Q_reg_22_inst : DFF_X1 port map( D => n5439, CK => CLK
                           , Q => n_3282, QN => 
                           DataPath_RF_bus_reg_dataout_1782_port);
   DataPath_RF_BLOCKi_64_Q_reg_22_inst : DFF_X1 port map( D => n5474, CK => CLK
                           , Q => n_3283, QN => 
                           DataPath_RF_bus_reg_dataout_1814_port);
   DataPath_RF_BLOCKi_65_Q_reg_22_inst : DFF_X1 port map( D => n5509, CK => CLK
                           , Q => n_3284, QN => 
                           DataPath_RF_bus_reg_dataout_1846_port);
   DataPath_RF_BLOCKi_66_Q_reg_22_inst : DFF_X1 port map( D => n5544, CK => CLK
                           , Q => n_3285, QN => 
                           DataPath_RF_bus_reg_dataout_1878_port);
   DataPath_RF_BLOCKi_67_Q_reg_22_inst : DFF_X1 port map( D => n5579, CK => CLK
                           , Q => n_3286, QN => 
                           DataPath_RF_bus_reg_dataout_1910_port);
   DataPath_RF_BLOCKi_68_Q_reg_22_inst : DFF_X1 port map( D => n5618, CK => CLK
                           , Q => n_3287, QN => 
                           DataPath_RF_bus_reg_dataout_1942_port);
   DataPath_RF_BLOCKi_69_Q_reg_22_inst : DFF_X1 port map( D => n5655, CK => CLK
                           , Q => n_3288, QN => 
                           DataPath_RF_bus_reg_dataout_1974_port);
   DataPath_RF_BLOCKi_70_Q_reg_22_inst : DFF_X1 port map( D => n5692, CK => CLK
                           , Q => n_3289, QN => 
                           DataPath_RF_bus_reg_dataout_2006_port);
   DataPath_RF_BLOCKi_71_Q_reg_22_inst : DFF_X1 port map( D => n5729, CK => CLK
                           , Q => n_3290, QN => 
                           DataPath_RF_bus_reg_dataout_2038_port);
   DataPath_RF_BLOCKi_83_Q_reg_22_inst : DFF_X1 port map( D => n934, CK => CLK,
                           Q => n_3291, QN => 
                           DataPath_RF_bus_reg_dataout_2422_port);
   DataPath_RF_BLOCKi_84_Q_reg_22_inst : DFF_X1 port map( D => n979, CK => CLK,
                           Q => n_3292, QN => 
                           DataPath_RF_bus_reg_dataout_2454_port);
   DataPath_RF_BLOCKi_85_Q_reg_22_inst : DFF_X1 port map( D => n1016, CK => CLK
                           , Q => n_3293, QN => 
                           DataPath_RF_bus_reg_dataout_2486_port);
   DataPath_RF_BLOCKi_86_Q_reg_22_inst : DFF_X1 port map( D => n1053, CK => CLK
                           , Q => n_3294, QN => 
                           DataPath_RF_bus_reg_dataout_2518_port);
   DataPath_RF_BLOCKi_87_Q_reg_22_inst : DFF_X1 port map( D => n1090, CK => CLK
                           , Q => n_3295, QN => 
                           DataPath_RF_bus_reg_dataout_2550_port);
   DataPath_RF_BLOCKi_72_Q_reg_22_inst : DFF_X1 port map( D => n5766, CK => CLK
                           , Q => n_3296, QN => 
                           DataPath_RF_bus_reg_dataout_2070_port);
   DataPath_RF_BLOCKi_73_Q_reg_22_inst : DFF_X1 port map( D => n5805, CK => CLK
                           , Q => n_3297, QN => 
                           DataPath_RF_bus_reg_dataout_2102_port);
   DataPath_RF_BLOCKi_74_Q_reg_22_inst : DFF_X1 port map( D => n5841, CK => CLK
                           , Q => n_3298, QN => 
                           DataPath_RF_bus_reg_dataout_2134_port);
   DataPath_RF_BLOCKi_75_Q_reg_22_inst : DFF_X1 port map( D => n5877, CK => CLK
                           , Q => n_3299, QN => 
                           DataPath_RF_bus_reg_dataout_2166_port);
   DataPath_RF_BLOCKi_76_Q_reg_22_inst : DFF_X1 port map( D => n5913, CK => CLK
                           , Q => n_3300, QN => 
                           DataPath_RF_bus_reg_dataout_2198_port);
   DataPath_RF_BLOCKi_77_Q_reg_22_inst : DFF_X1 port map( D => n5949, CK => CLK
                           , Q => n_3301, QN => 
                           DataPath_RF_bus_reg_dataout_2230_port);
   DataPath_RF_BLOCKi_78_Q_reg_22_inst : DFF_X1 port map( D => n5985, CK => CLK
                           , Q => n_3302, QN => 
                           DataPath_RF_bus_reg_dataout_2262_port);
   DataPath_RF_BLOCKi_79_Q_reg_22_inst : DFF_X1 port map( D => n6021, CK => CLK
                           , Q => n_3303, QN => 
                           DataPath_RF_bus_reg_dataout_2294_port);
   DataPath_RF_BLOCKi_80_Q_reg_22_inst : DFF_X1 port map( D => n6058, CK => CLK
                           , Q => n_3304, QN => 
                           DataPath_RF_bus_reg_dataout_2326_port);
   DataPath_RF_BLOCKi_81_Q_reg_22_inst : DFF_X1 port map( D => n6094, CK => CLK
                           , Q => n_3305, QN => 
                           DataPath_RF_bus_reg_dataout_2358_port);
   DataPath_RF_BLOCKi_82_Q_reg_22_inst : DFF_X1 port map( D => n6128, CK => CLK
                           , Q => n_3306, QN => 
                           DataPath_RF_bus_reg_dataout_2390_port);
   DataPath_REG_ALU_OUT_Q_reg_23_inst : DFF_X1 port map( D => n7000, CK => CLK,
                           Q => DRAM_ADDRESS_23_port, QN => n509);
   DataPath_REG_MEM_ALUOUT_Q_reg_23_inst : DFF_X1 port map( D => n1126, CK => 
                           CLK, Q => n_3307, QN => 
                           DataPath_i_REG_MEM_ALUOUT_23_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_23_inst : DFF_X1 port map( D => n6776, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_55_port,
                           QN => n622);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_23_inst : DFF_X1 port map( D => n6808, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_87_port,
                           QN => n654);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_23_inst : DFF_X1 port map( D => n6840, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_119_port
                           , QN => n686);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_23_inst : DFF_X1 port map( D => n6872, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_151_port
                           , QN => n718);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_23_inst : DFF_X1 port map( D => n6904, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_183_port
                           , QN => n750);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_23_inst : DFF_X1 port map( D => n6936, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_215_port
                           , QN => n782);
   DataPath_RF_BLOCKi_8_Q_reg_23_inst : DFF_X1 port map( D => n3326, CK => CLK,
                           Q => n_3308, QN => 
                           DataPath_RF_bus_reg_dataout_23_port);
   DataPath_RF_BLOCKi_9_Q_reg_23_inst : DFF_X1 port map( D => n3389, CK => CLK,
                           Q => n_3309, QN => 
                           DataPath_RF_bus_reg_dataout_55_port);
   DataPath_RF_BLOCKi_10_Q_reg_23_inst : DFF_X1 port map( D => n3427, CK => CLK
                           , Q => n_3310, QN => 
                           DataPath_RF_bus_reg_dataout_87_port);
   DataPath_RF_BLOCKi_11_Q_reg_23_inst : DFF_X1 port map( D => n3465, CK => CLK
                           , Q => n_3311, QN => 
                           DataPath_RF_bus_reg_dataout_119_port);
   DataPath_RF_BLOCKi_12_Q_reg_23_inst : DFF_X1 port map( D => n3503, CK => CLK
                           , Q => n_3312, QN => 
                           DataPath_RF_bus_reg_dataout_151_port);
   DataPath_RF_BLOCKi_13_Q_reg_23_inst : DFF_X1 port map( D => n3541, CK => CLK
                           , Q => n_3313, QN => 
                           DataPath_RF_bus_reg_dataout_183_port);
   DataPath_RF_BLOCKi_14_Q_reg_23_inst : DFF_X1 port map( D => n3579, CK => CLK
                           , Q => n_3314, QN => 
                           DataPath_RF_bus_reg_dataout_215_port);
   DataPath_RF_BLOCKi_15_Q_reg_23_inst : DFF_X1 port map( D => n3617, CK => CLK
                           , Q => n_3315, QN => 
                           DataPath_RF_bus_reg_dataout_247_port);
   DataPath_RF_BLOCKi_16_Q_reg_23_inst : DFF_X1 port map( D => n3655, CK => CLK
                           , Q => n_3316, QN => 
                           DataPath_RF_bus_reg_dataout_279_port);
   DataPath_RF_BLOCKi_17_Q_reg_23_inst : DFF_X1 port map( D => n3692, CK => CLK
                           , Q => n_3317, QN => 
                           DataPath_RF_bus_reg_dataout_311_port);
   DataPath_RF_BLOCKi_18_Q_reg_23_inst : DFF_X1 port map( D => n3729, CK => CLK
                           , Q => n_3318, QN => 
                           DataPath_RF_bus_reg_dataout_343_port);
   DataPath_RF_BLOCKi_19_Q_reg_23_inst : DFF_X1 port map( D => n3766, CK => CLK
                           , Q => n_3319, QN => 
                           DataPath_RF_bus_reg_dataout_375_port);
   DataPath_RF_BLOCKi_20_Q_reg_23_inst : DFF_X1 port map( D => n3801, CK => CLK
                           , Q => n_3320, QN => 
                           DataPath_RF_bus_reg_dataout_407_port);
   DataPath_RF_BLOCKi_21_Q_reg_23_inst : DFF_X1 port map( D => n3836, CK => CLK
                           , Q => n_3321, QN => 
                           DataPath_RF_bus_reg_dataout_439_port);
   DataPath_RF_BLOCKi_22_Q_reg_23_inst : DFF_X1 port map( D => n3871, CK => CLK
                           , Q => n_3322, QN => 
                           DataPath_RF_bus_reg_dataout_471_port);
   DataPath_RF_BLOCKi_23_Q_reg_23_inst : DFF_X1 port map( D => n3914, CK => CLK
                           , Q => n_3323, QN => 
                           DataPath_RF_bus_reg_dataout_503_port);
   DataPath_RF_BLOCKi_24_Q_reg_23_inst : DFF_X1 port map( D => n3982, CK => CLK
                           , Q => n_3324, QN => 
                           DataPath_RF_bus_reg_dataout_535_port);
   DataPath_RF_BLOCKi_25_Q_reg_23_inst : DFF_X1 port map( D => n4042, CK => CLK
                           , Q => n_3325, QN => 
                           DataPath_RF_bus_reg_dataout_567_port);
   DataPath_RF_BLOCKi_26_Q_reg_23_inst : DFF_X1 port map( D => n4077, CK => CLK
                           , Q => n_3326, QN => 
                           DataPath_RF_bus_reg_dataout_599_port);
   DataPath_RF_BLOCKi_27_Q_reg_23_inst : DFF_X1 port map( D => n4112, CK => CLK
                           , Q => n_3327, QN => 
                           DataPath_RF_bus_reg_dataout_631_port);
   DataPath_RF_BLOCKi_28_Q_reg_23_inst : DFF_X1 port map( D => n4147, CK => CLK
                           , Q => n_3328, QN => 
                           DataPath_RF_bus_reg_dataout_663_port);
   DataPath_RF_BLOCKi_29_Q_reg_23_inst : DFF_X1 port map( D => n4182, CK => CLK
                           , Q => n_3329, QN => 
                           DataPath_RF_bus_reg_dataout_695_port);
   DataPath_RF_BLOCKi_30_Q_reg_23_inst : DFF_X1 port map( D => n4217, CK => CLK
                           , Q => n_3330, QN => 
                           DataPath_RF_bus_reg_dataout_727_port);
   DataPath_RF_BLOCKi_31_Q_reg_23_inst : DFF_X1 port map( D => n4252, CK => CLK
                           , Q => n_3331, QN => 
                           DataPath_RF_bus_reg_dataout_759_port);
   DataPath_RF_BLOCKi_32_Q_reg_23_inst : DFF_X1 port map( D => n4287, CK => CLK
                           , Q => n_3332, QN => 
                           DataPath_RF_bus_reg_dataout_791_port);
   DataPath_RF_BLOCKi_33_Q_reg_23_inst : DFF_X1 port map( D => n4322, CK => CLK
                           , Q => n_3333, QN => 
                           DataPath_RF_bus_reg_dataout_823_port);
   DataPath_RF_BLOCKi_34_Q_reg_23_inst : DFF_X1 port map( D => n4357, CK => CLK
                           , Q => n_3334, QN => 
                           DataPath_RF_bus_reg_dataout_855_port);
   DataPath_RF_BLOCKi_35_Q_reg_23_inst : DFF_X1 port map( D => n4392, CK => CLK
                           , Q => n_3335, QN => 
                           DataPath_RF_bus_reg_dataout_887_port);
   DataPath_RF_BLOCKi_36_Q_reg_23_inst : DFF_X1 port map( D => n4427, CK => CLK
                           , Q => n_3336, QN => 
                           DataPath_RF_bus_reg_dataout_919_port);
   DataPath_RF_BLOCKi_37_Q_reg_23_inst : DFF_X1 port map( D => n4462, CK => CLK
                           , Q => n_3337, QN => 
                           DataPath_RF_bus_reg_dataout_951_port);
   DataPath_RF_BLOCKi_38_Q_reg_23_inst : DFF_X1 port map( D => n4497, CK => CLK
                           , Q => n_3338, QN => 
                           DataPath_RF_bus_reg_dataout_983_port);
   DataPath_RF_BLOCKi_39_Q_reg_23_inst : DFF_X1 port map( D => n4532, CK => CLK
                           , Q => n_3339, QN => 
                           DataPath_RF_bus_reg_dataout_1015_port);
   DataPath_RF_BLOCKi_40_Q_reg_23_inst : DFF_X1 port map( D => n4575, CK => CLK
                           , Q => n_3340, QN => 
                           DataPath_RF_bus_reg_dataout_1047_port);
   DataPath_RF_BLOCKi_41_Q_reg_23_inst : DFF_X1 port map( D => n4635, CK => CLK
                           , Q => n_3341, QN => 
                           DataPath_RF_bus_reg_dataout_1079_port);
   DataPath_RF_BLOCKi_42_Q_reg_23_inst : DFF_X1 port map( D => n4670, CK => CLK
                           , Q => n_3342, QN => 
                           DataPath_RF_bus_reg_dataout_1111_port);
   DataPath_RF_BLOCKi_43_Q_reg_23_inst : DFF_X1 port map( D => n4705, CK => CLK
                           , Q => n_3343, QN => 
                           DataPath_RF_bus_reg_dataout_1143_port);
   DataPath_RF_BLOCKi_44_Q_reg_23_inst : DFF_X1 port map( D => n4740, CK => CLK
                           , Q => n_3344, QN => 
                           DataPath_RF_bus_reg_dataout_1175_port);
   DataPath_RF_BLOCKi_45_Q_reg_23_inst : DFF_X1 port map( D => n4775, CK => CLK
                           , Q => n_3345, QN => 
                           DataPath_RF_bus_reg_dataout_1207_port);
   DataPath_RF_BLOCKi_46_Q_reg_23_inst : DFF_X1 port map( D => n4810, CK => CLK
                           , Q => n_3346, QN => 
                           DataPath_RF_bus_reg_dataout_1239_port);
   DataPath_RF_BLOCKi_47_Q_reg_23_inst : DFF_X1 port map( D => n4845, CK => CLK
                           , Q => n_3347, QN => 
                           DataPath_RF_bus_reg_dataout_1271_port);
   DataPath_RF_BLOCKi_48_Q_reg_23_inst : DFF_X1 port map( D => n4880, CK => CLK
                           , Q => n_3348, QN => 
                           DataPath_RF_bus_reg_dataout_1303_port);
   DataPath_RF_BLOCKi_49_Q_reg_23_inst : DFF_X1 port map( D => n4915, CK => CLK
                           , Q => n_3349, QN => 
                           DataPath_RF_bus_reg_dataout_1335_port);
   DataPath_RF_BLOCKi_50_Q_reg_23_inst : DFF_X1 port map( D => n4950, CK => CLK
                           , Q => n_3350, QN => 
                           DataPath_RF_bus_reg_dataout_1367_port);
   DataPath_RF_BLOCKi_51_Q_reg_23_inst : DFF_X1 port map( D => n4985, CK => CLK
                           , Q => n_3351, QN => 
                           DataPath_RF_bus_reg_dataout_1399_port);
   DataPath_RF_BLOCKi_52_Q_reg_23_inst : DFF_X1 port map( D => n5020, CK => CLK
                           , Q => n_3352, QN => 
                           DataPath_RF_bus_reg_dataout_1431_port);
   DataPath_RF_BLOCKi_53_Q_reg_23_inst : DFF_X1 port map( D => n5055, CK => CLK
                           , Q => n_3353, QN => 
                           DataPath_RF_bus_reg_dataout_1463_port);
   DataPath_RF_BLOCKi_54_Q_reg_23_inst : DFF_X1 port map( D => n5090, CK => CLK
                           , Q => n_3354, QN => 
                           DataPath_RF_bus_reg_dataout_1495_port);
   DataPath_RF_BLOCKi_55_Q_reg_23_inst : DFF_X1 port map( D => n5125, CK => CLK
                           , Q => n_3355, QN => 
                           DataPath_RF_bus_reg_dataout_1527_port);
   DataPath_RF_BLOCKi_56_Q_reg_23_inst : DFF_X1 port map( D => n5168, CK => CLK
                           , Q => n_3356, QN => 
                           DataPath_RF_bus_reg_dataout_1559_port);
   DataPath_RF_BLOCKi_57_Q_reg_23_inst : DFF_X1 port map( D => n5227, CK => CLK
                           , Q => n_3357, QN => 
                           DataPath_RF_bus_reg_dataout_1591_port);
   DataPath_RF_BLOCKi_58_Q_reg_23_inst : DFF_X1 port map( D => n5263, CK => CLK
                           , Q => n_3358, QN => 
                           DataPath_RF_bus_reg_dataout_1623_port);
   DataPath_RF_BLOCKi_59_Q_reg_23_inst : DFF_X1 port map( D => n5298, CK => CLK
                           , Q => n_3359, QN => 
                           DataPath_RF_bus_reg_dataout_1655_port);
   DataPath_RF_BLOCKi_60_Q_reg_23_inst : DFF_X1 port map( D => n5333, CK => CLK
                           , Q => n_3360, QN => 
                           DataPath_RF_bus_reg_dataout_1687_port);
   DataPath_RF_BLOCKi_61_Q_reg_23_inst : DFF_X1 port map( D => n5368, CK => CLK
                           , Q => n_3361, QN => 
                           DataPath_RF_bus_reg_dataout_1719_port);
   DataPath_RF_BLOCKi_62_Q_reg_23_inst : DFF_X1 port map( D => n5403, CK => CLK
                           , Q => n_3362, QN => 
                           DataPath_RF_bus_reg_dataout_1751_port);
   DataPath_RF_BLOCKi_63_Q_reg_23_inst : DFF_X1 port map( D => n5438, CK => CLK
                           , Q => n_3363, QN => 
                           DataPath_RF_bus_reg_dataout_1783_port);
   DataPath_RF_BLOCKi_64_Q_reg_23_inst : DFF_X1 port map( D => n5473, CK => CLK
                           , Q => n_3364, QN => 
                           DataPath_RF_bus_reg_dataout_1815_port);
   DataPath_RF_BLOCKi_65_Q_reg_23_inst : DFF_X1 port map( D => n5508, CK => CLK
                           , Q => n_3365, QN => 
                           DataPath_RF_bus_reg_dataout_1847_port);
   DataPath_RF_BLOCKi_66_Q_reg_23_inst : DFF_X1 port map( D => n5543, CK => CLK
                           , Q => n_3366, QN => 
                           DataPath_RF_bus_reg_dataout_1879_port);
   DataPath_RF_BLOCKi_67_Q_reg_23_inst : DFF_X1 port map( D => n5578, CK => CLK
                           , Q => n_3367, QN => 
                           DataPath_RF_bus_reg_dataout_1911_port);
   DataPath_RF_BLOCKi_68_Q_reg_23_inst : DFF_X1 port map( D => n5617, CK => CLK
                           , Q => n_3368, QN => 
                           DataPath_RF_bus_reg_dataout_1943_port);
   DataPath_RF_BLOCKi_69_Q_reg_23_inst : DFF_X1 port map( D => n5654, CK => CLK
                           , Q => n_3369, QN => 
                           DataPath_RF_bus_reg_dataout_1975_port);
   DataPath_RF_BLOCKi_70_Q_reg_23_inst : DFF_X1 port map( D => n5691, CK => CLK
                           , Q => n_3370, QN => 
                           DataPath_RF_bus_reg_dataout_2007_port);
   DataPath_RF_BLOCKi_71_Q_reg_23_inst : DFF_X1 port map( D => n5728, CK => CLK
                           , Q => n_3371, QN => 
                           DataPath_RF_bus_reg_dataout_2039_port);
   DataPath_RF_BLOCKi_83_Q_reg_23_inst : DFF_X1 port map( D => n932, CK => CLK,
                           Q => n_3372, QN => 
                           DataPath_RF_bus_reg_dataout_2423_port);
   DataPath_RF_BLOCKi_84_Q_reg_23_inst : DFF_X1 port map( D => n978, CK => CLK,
                           Q => n_3373, QN => 
                           DataPath_RF_bus_reg_dataout_2455_port);
   DataPath_RF_BLOCKi_85_Q_reg_23_inst : DFF_X1 port map( D => n1015, CK => CLK
                           , Q => n_3374, QN => 
                           DataPath_RF_bus_reg_dataout_2487_port);
   DataPath_RF_BLOCKi_86_Q_reg_23_inst : DFF_X1 port map( D => n1052, CK => CLK
                           , Q => n_3375, QN => 
                           DataPath_RF_bus_reg_dataout_2519_port);
   DataPath_RF_BLOCKi_87_Q_reg_23_inst : DFF_X1 port map( D => n1089, CK => CLK
                           , Q => n_3376, QN => 
                           DataPath_RF_bus_reg_dataout_2551_port);
   DataPath_RF_BLOCKi_72_Q_reg_23_inst : DFF_X1 port map( D => n5765, CK => CLK
                           , Q => n_3377, QN => 
                           DataPath_RF_bus_reg_dataout_2071_port);
   DataPath_RF_BLOCKi_73_Q_reg_23_inst : DFF_X1 port map( D => n5804, CK => CLK
                           , Q => n_3378, QN => 
                           DataPath_RF_bus_reg_dataout_2103_port);
   DataPath_RF_BLOCKi_74_Q_reg_23_inst : DFF_X1 port map( D => n5840, CK => CLK
                           , Q => n_3379, QN => 
                           DataPath_RF_bus_reg_dataout_2135_port);
   DataPath_RF_BLOCKi_75_Q_reg_23_inst : DFF_X1 port map( D => n5876, CK => CLK
                           , Q => n_3380, QN => 
                           DataPath_RF_bus_reg_dataout_2167_port);
   DataPath_RF_BLOCKi_76_Q_reg_23_inst : DFF_X1 port map( D => n5912, CK => CLK
                           , Q => n_3381, QN => 
                           DataPath_RF_bus_reg_dataout_2199_port);
   DataPath_RF_BLOCKi_77_Q_reg_23_inst : DFF_X1 port map( D => n5948, CK => CLK
                           , Q => n_3382, QN => 
                           DataPath_RF_bus_reg_dataout_2231_port);
   DataPath_RF_BLOCKi_78_Q_reg_23_inst : DFF_X1 port map( D => n5984, CK => CLK
                           , Q => n_3383, QN => 
                           DataPath_RF_bus_reg_dataout_2263_port);
   DataPath_RF_BLOCKi_79_Q_reg_23_inst : DFF_X1 port map( D => n6020, CK => CLK
                           , Q => n_3384, QN => 
                           DataPath_RF_bus_reg_dataout_2295_port);
   DataPath_RF_BLOCKi_80_Q_reg_23_inst : DFF_X1 port map( D => n6057, CK => CLK
                           , Q => n_3385, QN => 
                           DataPath_RF_bus_reg_dataout_2327_port);
   DataPath_RF_BLOCKi_81_Q_reg_23_inst : DFF_X1 port map( D => n6093, CK => CLK
                           , Q => n_3386, QN => 
                           DataPath_RF_bus_reg_dataout_2359_port);
   DataPath_RF_BLOCKi_82_Q_reg_23_inst : DFF_X1 port map( D => n6127, CK => CLK
                           , Q => n_3387, QN => 
                           DataPath_RF_bus_reg_dataout_2391_port);
   DataPath_REG_ALU_OUT_Q_reg_24_inst : DFF_X1 port map( D => n6999, CK => CLK,
                           Q => DRAM_ADDRESS_24_port, QN => n510);
   DataPath_REG_MEM_ALUOUT_Q_reg_24_inst : DFF_X1 port map( D => n1125, CK => 
                           CLK, Q => n_3388, QN => 
                           DataPath_i_REG_MEM_ALUOUT_24_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_24_inst : DFF_X1 port map( D => n6775, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_56_port,
                           QN => n623);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_24_inst : DFF_X1 port map( D => n6807, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_88_port,
                           QN => n655);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_24_inst : DFF_X1 port map( D => n6839, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_120_port
                           , QN => n687);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_24_inst : DFF_X1 port map( D => n6871, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_152_port
                           , QN => n719);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_24_inst : DFF_X1 port map( D => n6903, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_184_port
                           , QN => n751);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_24_inst : DFF_X1 port map( D => n6935, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_216_port
                           , QN => n783);
   DataPath_RF_BLOCKi_8_Q_reg_24_inst : DFF_X1 port map( D => n3324, CK => CLK,
                           Q => n_3389, QN => 
                           DataPath_RF_bus_reg_dataout_24_port);
   DataPath_RF_BLOCKi_9_Q_reg_24_inst : DFF_X1 port map( D => n3388, CK => CLK,
                           Q => n_3390, QN => 
                           DataPath_RF_bus_reg_dataout_56_port);
   DataPath_RF_BLOCKi_10_Q_reg_24_inst : DFF_X1 port map( D => n3426, CK => CLK
                           , Q => n_3391, QN => 
                           DataPath_RF_bus_reg_dataout_88_port);
   DataPath_RF_BLOCKi_11_Q_reg_24_inst : DFF_X1 port map( D => n3464, CK => CLK
                           , Q => n_3392, QN => 
                           DataPath_RF_bus_reg_dataout_120_port);
   DataPath_RF_BLOCKi_12_Q_reg_24_inst : DFF_X1 port map( D => n3502, CK => CLK
                           , Q => n_3393, QN => 
                           DataPath_RF_bus_reg_dataout_152_port);
   DataPath_RF_BLOCKi_13_Q_reg_24_inst : DFF_X1 port map( D => n3540, CK => CLK
                           , Q => n_3394, QN => 
                           DataPath_RF_bus_reg_dataout_184_port);
   DataPath_RF_BLOCKi_14_Q_reg_24_inst : DFF_X1 port map( D => n3578, CK => CLK
                           , Q => n_3395, QN => 
                           DataPath_RF_bus_reg_dataout_216_port);
   DataPath_RF_BLOCKi_15_Q_reg_24_inst : DFF_X1 port map( D => n3616, CK => CLK
                           , Q => n_3396, QN => 
                           DataPath_RF_bus_reg_dataout_248_port);
   DataPath_RF_BLOCKi_16_Q_reg_24_inst : DFF_X1 port map( D => n3654, CK => CLK
                           , Q => n_3397, QN => 
                           DataPath_RF_bus_reg_dataout_280_port);
   DataPath_RF_BLOCKi_17_Q_reg_24_inst : DFF_X1 port map( D => n3691, CK => CLK
                           , Q => n_3398, QN => 
                           DataPath_RF_bus_reg_dataout_312_port);
   DataPath_RF_BLOCKi_18_Q_reg_24_inst : DFF_X1 port map( D => n3728, CK => CLK
                           , Q => n_3399, QN => 
                           DataPath_RF_bus_reg_dataout_344_port);
   DataPath_RF_BLOCKi_19_Q_reg_24_inst : DFF_X1 port map( D => n3765, CK => CLK
                           , Q => n_3400, QN => 
                           DataPath_RF_bus_reg_dataout_376_port);
   DataPath_RF_BLOCKi_20_Q_reg_24_inst : DFF_X1 port map( D => n3800, CK => CLK
                           , Q => n_3401, QN => 
                           DataPath_RF_bus_reg_dataout_408_port);
   DataPath_RF_BLOCKi_21_Q_reg_24_inst : DFF_X1 port map( D => n3835, CK => CLK
                           , Q => n_3402, QN => 
                           DataPath_RF_bus_reg_dataout_440_port);
   DataPath_RF_BLOCKi_22_Q_reg_24_inst : DFF_X1 port map( D => n3870, CK => CLK
                           , Q => n_3403, QN => 
                           DataPath_RF_bus_reg_dataout_472_port);
   DataPath_RF_BLOCKi_23_Q_reg_24_inst : DFF_X1 port map( D => n3912, CK => CLK
                           , Q => n_3404, QN => 
                           DataPath_RF_bus_reg_dataout_504_port);
   DataPath_RF_BLOCKi_24_Q_reg_24_inst : DFF_X1 port map( D => n3980, CK => CLK
                           , Q => n_3405, QN => 
                           DataPath_RF_bus_reg_dataout_536_port);
   DataPath_RF_BLOCKi_25_Q_reg_24_inst : DFF_X1 port map( D => n4041, CK => CLK
                           , Q => n_3406, QN => 
                           DataPath_RF_bus_reg_dataout_568_port);
   DataPath_RF_BLOCKi_26_Q_reg_24_inst : DFF_X1 port map( D => n4076, CK => CLK
                           , Q => n_3407, QN => 
                           DataPath_RF_bus_reg_dataout_600_port);
   DataPath_RF_BLOCKi_27_Q_reg_24_inst : DFF_X1 port map( D => n4111, CK => CLK
                           , Q => n_3408, QN => 
                           DataPath_RF_bus_reg_dataout_632_port);
   DataPath_RF_BLOCKi_28_Q_reg_24_inst : DFF_X1 port map( D => n4146, CK => CLK
                           , Q => n_3409, QN => 
                           DataPath_RF_bus_reg_dataout_664_port);
   DataPath_RF_BLOCKi_29_Q_reg_24_inst : DFF_X1 port map( D => n4181, CK => CLK
                           , Q => n_3410, QN => 
                           DataPath_RF_bus_reg_dataout_696_port);
   DataPath_RF_BLOCKi_30_Q_reg_24_inst : DFF_X1 port map( D => n4216, CK => CLK
                           , Q => n_3411, QN => 
                           DataPath_RF_bus_reg_dataout_728_port);
   DataPath_RF_BLOCKi_31_Q_reg_24_inst : DFF_X1 port map( D => n4251, CK => CLK
                           , Q => n_3412, QN => 
                           DataPath_RF_bus_reg_dataout_760_port);
   DataPath_RF_BLOCKi_32_Q_reg_24_inst : DFF_X1 port map( D => n4286, CK => CLK
                           , Q => n_3413, QN => 
                           DataPath_RF_bus_reg_dataout_792_port);
   DataPath_RF_BLOCKi_33_Q_reg_24_inst : DFF_X1 port map( D => n4321, CK => CLK
                           , Q => n_3414, QN => 
                           DataPath_RF_bus_reg_dataout_824_port);
   DataPath_RF_BLOCKi_34_Q_reg_24_inst : DFF_X1 port map( D => n4356, CK => CLK
                           , Q => n_3415, QN => 
                           DataPath_RF_bus_reg_dataout_856_port);
   DataPath_RF_BLOCKi_35_Q_reg_24_inst : DFF_X1 port map( D => n4391, CK => CLK
                           , Q => n_3416, QN => 
                           DataPath_RF_bus_reg_dataout_888_port);
   DataPath_RF_BLOCKi_36_Q_reg_24_inst : DFF_X1 port map( D => n4426, CK => CLK
                           , Q => n_3417, QN => 
                           DataPath_RF_bus_reg_dataout_920_port);
   DataPath_RF_BLOCKi_37_Q_reg_24_inst : DFF_X1 port map( D => n4461, CK => CLK
                           , Q => n_3418, QN => 
                           DataPath_RF_bus_reg_dataout_952_port);
   DataPath_RF_BLOCKi_38_Q_reg_24_inst : DFF_X1 port map( D => n4496, CK => CLK
                           , Q => n_3419, QN => 
                           DataPath_RF_bus_reg_dataout_984_port);
   DataPath_RF_BLOCKi_39_Q_reg_24_inst : DFF_X1 port map( D => n4531, CK => CLK
                           , Q => n_3420, QN => 
                           DataPath_RF_bus_reg_dataout_1016_port);
   DataPath_RF_BLOCKi_40_Q_reg_24_inst : DFF_X1 port map( D => n4573, CK => CLK
                           , Q => n_3421, QN => 
                           DataPath_RF_bus_reg_dataout_1048_port);
   DataPath_RF_BLOCKi_41_Q_reg_24_inst : DFF_X1 port map( D => n4634, CK => CLK
                           , Q => n_3422, QN => 
                           DataPath_RF_bus_reg_dataout_1080_port);
   DataPath_RF_BLOCKi_42_Q_reg_24_inst : DFF_X1 port map( D => n4669, CK => CLK
                           , Q => n_3423, QN => 
                           DataPath_RF_bus_reg_dataout_1112_port);
   DataPath_RF_BLOCKi_43_Q_reg_24_inst : DFF_X1 port map( D => n4704, CK => CLK
                           , Q => n_3424, QN => 
                           DataPath_RF_bus_reg_dataout_1144_port);
   DataPath_RF_BLOCKi_44_Q_reg_24_inst : DFF_X1 port map( D => n4739, CK => CLK
                           , Q => n_3425, QN => 
                           DataPath_RF_bus_reg_dataout_1176_port);
   DataPath_RF_BLOCKi_45_Q_reg_24_inst : DFF_X1 port map( D => n4774, CK => CLK
                           , Q => n_3426, QN => 
                           DataPath_RF_bus_reg_dataout_1208_port);
   DataPath_RF_BLOCKi_46_Q_reg_24_inst : DFF_X1 port map( D => n4809, CK => CLK
                           , Q => n_3427, QN => 
                           DataPath_RF_bus_reg_dataout_1240_port);
   DataPath_RF_BLOCKi_47_Q_reg_24_inst : DFF_X1 port map( D => n4844, CK => CLK
                           , Q => n_3428, QN => 
                           DataPath_RF_bus_reg_dataout_1272_port);
   DataPath_RF_BLOCKi_48_Q_reg_24_inst : DFF_X1 port map( D => n4879, CK => CLK
                           , Q => n_3429, QN => 
                           DataPath_RF_bus_reg_dataout_1304_port);
   DataPath_RF_BLOCKi_49_Q_reg_24_inst : DFF_X1 port map( D => n4914, CK => CLK
                           , Q => n_3430, QN => 
                           DataPath_RF_bus_reg_dataout_1336_port);
   DataPath_RF_BLOCKi_50_Q_reg_24_inst : DFF_X1 port map( D => n4949, CK => CLK
                           , Q => n_3431, QN => 
                           DataPath_RF_bus_reg_dataout_1368_port);
   DataPath_RF_BLOCKi_51_Q_reg_24_inst : DFF_X1 port map( D => n4984, CK => CLK
                           , Q => n_3432, QN => 
                           DataPath_RF_bus_reg_dataout_1400_port);
   DataPath_RF_BLOCKi_52_Q_reg_24_inst : DFF_X1 port map( D => n5019, CK => CLK
                           , Q => n_3433, QN => 
                           DataPath_RF_bus_reg_dataout_1432_port);
   DataPath_RF_BLOCKi_53_Q_reg_24_inst : DFF_X1 port map( D => n5054, CK => CLK
                           , Q => n_3434, QN => 
                           DataPath_RF_bus_reg_dataout_1464_port);
   DataPath_RF_BLOCKi_54_Q_reg_24_inst : DFF_X1 port map( D => n5089, CK => CLK
                           , Q => n_3435, QN => 
                           DataPath_RF_bus_reg_dataout_1496_port);
   DataPath_RF_BLOCKi_55_Q_reg_24_inst : DFF_X1 port map( D => n5124, CK => CLK
                           , Q => n_3436, QN => 
                           DataPath_RF_bus_reg_dataout_1528_port);
   DataPath_RF_BLOCKi_56_Q_reg_24_inst : DFF_X1 port map( D => n5166, CK => CLK
                           , Q => n_3437, QN => 
                           DataPath_RF_bus_reg_dataout_1560_port);
   DataPath_RF_BLOCKi_57_Q_reg_24_inst : DFF_X1 port map( D => n5226, CK => CLK
                           , Q => n_3438, QN => 
                           DataPath_RF_bus_reg_dataout_1592_port);
   DataPath_RF_BLOCKi_58_Q_reg_24_inst : DFF_X1 port map( D => n5262, CK => CLK
                           , Q => n_3439, QN => 
                           DataPath_RF_bus_reg_dataout_1624_port);
   DataPath_RF_BLOCKi_59_Q_reg_24_inst : DFF_X1 port map( D => n5297, CK => CLK
                           , Q => n_3440, QN => 
                           DataPath_RF_bus_reg_dataout_1656_port);
   DataPath_RF_BLOCKi_60_Q_reg_24_inst : DFF_X1 port map( D => n5332, CK => CLK
                           , Q => n_3441, QN => 
                           DataPath_RF_bus_reg_dataout_1688_port);
   DataPath_RF_BLOCKi_61_Q_reg_24_inst : DFF_X1 port map( D => n5367, CK => CLK
                           , Q => n_3442, QN => 
                           DataPath_RF_bus_reg_dataout_1720_port);
   DataPath_RF_BLOCKi_62_Q_reg_24_inst : DFF_X1 port map( D => n5402, CK => CLK
                           , Q => n_3443, QN => 
                           DataPath_RF_bus_reg_dataout_1752_port);
   DataPath_RF_BLOCKi_63_Q_reg_24_inst : DFF_X1 port map( D => n5437, CK => CLK
                           , Q => n_3444, QN => 
                           DataPath_RF_bus_reg_dataout_1784_port);
   DataPath_RF_BLOCKi_64_Q_reg_24_inst : DFF_X1 port map( D => n5472, CK => CLK
                           , Q => n_3445, QN => 
                           DataPath_RF_bus_reg_dataout_1816_port);
   DataPath_RF_BLOCKi_65_Q_reg_24_inst : DFF_X1 port map( D => n5507, CK => CLK
                           , Q => n_3446, QN => 
                           DataPath_RF_bus_reg_dataout_1848_port);
   DataPath_RF_BLOCKi_66_Q_reg_24_inst : DFF_X1 port map( D => n5542, CK => CLK
                           , Q => n_3447, QN => 
                           DataPath_RF_bus_reg_dataout_1880_port);
   DataPath_RF_BLOCKi_67_Q_reg_24_inst : DFF_X1 port map( D => n5577, CK => CLK
                           , Q => n_3448, QN => 
                           DataPath_RF_bus_reg_dataout_1912_port);
   DataPath_RF_BLOCKi_68_Q_reg_24_inst : DFF_X1 port map( D => n5616, CK => CLK
                           , Q => n_3449, QN => 
                           DataPath_RF_bus_reg_dataout_1944_port);
   DataPath_RF_BLOCKi_69_Q_reg_24_inst : DFF_X1 port map( D => n5653, CK => CLK
                           , Q => n_3450, QN => 
                           DataPath_RF_bus_reg_dataout_1976_port);
   DataPath_RF_BLOCKi_70_Q_reg_24_inst : DFF_X1 port map( D => n5690, CK => CLK
                           , Q => n_3451, QN => 
                           DataPath_RF_bus_reg_dataout_2008_port);
   DataPath_RF_BLOCKi_71_Q_reg_24_inst : DFF_X1 port map( D => n5727, CK => CLK
                           , Q => n_3452, QN => 
                           DataPath_RF_bus_reg_dataout_2040_port);
   DataPath_RF_BLOCKi_83_Q_reg_24_inst : DFF_X1 port map( D => n930, CK => CLK,
                           Q => n_3453, QN => 
                           DataPath_RF_bus_reg_dataout_2424_port);
   DataPath_RF_BLOCKi_84_Q_reg_24_inst : DFF_X1 port map( D => n977, CK => CLK,
                           Q => n_3454, QN => 
                           DataPath_RF_bus_reg_dataout_2456_port);
   DataPath_RF_BLOCKi_85_Q_reg_24_inst : DFF_X1 port map( D => n1014, CK => CLK
                           , Q => n_3455, QN => 
                           DataPath_RF_bus_reg_dataout_2488_port);
   DataPath_RF_BLOCKi_86_Q_reg_24_inst : DFF_X1 port map( D => n1051, CK => CLK
                           , Q => n_3456, QN => 
                           DataPath_RF_bus_reg_dataout_2520_port);
   DataPath_RF_BLOCKi_87_Q_reg_24_inst : DFF_X1 port map( D => n1088, CK => CLK
                           , Q => n_3457, QN => 
                           DataPath_RF_bus_reg_dataout_2552_port);
   DataPath_RF_BLOCKi_72_Q_reg_24_inst : DFF_X1 port map( D => n5764, CK => CLK
                           , Q => n_3458, QN => 
                           DataPath_RF_bus_reg_dataout_2072_port);
   DataPath_RF_BLOCKi_73_Q_reg_24_inst : DFF_X1 port map( D => n5803, CK => CLK
                           , Q => n_3459, QN => 
                           DataPath_RF_bus_reg_dataout_2104_port);
   DataPath_RF_BLOCKi_74_Q_reg_24_inst : DFF_X1 port map( D => n5839, CK => CLK
                           , Q => n_3460, QN => 
                           DataPath_RF_bus_reg_dataout_2136_port);
   DataPath_RF_BLOCKi_75_Q_reg_24_inst : DFF_X1 port map( D => n5875, CK => CLK
                           , Q => n_3461, QN => 
                           DataPath_RF_bus_reg_dataout_2168_port);
   DataPath_RF_BLOCKi_76_Q_reg_24_inst : DFF_X1 port map( D => n5911, CK => CLK
                           , Q => n_3462, QN => 
                           DataPath_RF_bus_reg_dataout_2200_port);
   DataPath_RF_BLOCKi_77_Q_reg_24_inst : DFF_X1 port map( D => n5947, CK => CLK
                           , Q => n_3463, QN => 
                           DataPath_RF_bus_reg_dataout_2232_port);
   DataPath_RF_BLOCKi_78_Q_reg_24_inst : DFF_X1 port map( D => n5983, CK => CLK
                           , Q => n_3464, QN => 
                           DataPath_RF_bus_reg_dataout_2264_port);
   DataPath_RF_BLOCKi_79_Q_reg_24_inst : DFF_X1 port map( D => n6019, CK => CLK
                           , Q => n_3465, QN => 
                           DataPath_RF_bus_reg_dataout_2296_port);
   DataPath_RF_BLOCKi_80_Q_reg_24_inst : DFF_X1 port map( D => n6056, CK => CLK
                           , Q => n_3466, QN => 
                           DataPath_RF_bus_reg_dataout_2328_port);
   DataPath_RF_BLOCKi_81_Q_reg_24_inst : DFF_X1 port map( D => n6092, CK => CLK
                           , Q => n_3467, QN => 
                           DataPath_RF_bus_reg_dataout_2360_port);
   DataPath_RF_BLOCKi_82_Q_reg_24_inst : DFF_X1 port map( D => n6126, CK => CLK
                           , Q => n_3468, QN => 
                           DataPath_RF_bus_reg_dataout_2392_port);
   DataPath_REG_ALU_OUT_Q_reg_26_inst : DFF_X1 port map( D => n6997, CK => CLK,
                           Q => DRAM_ADDRESS_26_port, QN => n511);
   DataPath_REG_MEM_ALUOUT_Q_reg_26_inst : DFF_X1 port map( D => n1123, CK => 
                           CLK, Q => n_3469, QN => 
                           DataPath_i_REG_MEM_ALUOUT_26_port);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_26_inst : DFF_X1 port map( D => n6837, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_122_port
                           , QN => n689);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_26_inst : DFF_X1 port map( D => n6869, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_154_port
                           , QN => n721);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_26_inst : DFF_X1 port map( D => n6933, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_218_port
                           , QN => n785);
   DataPath_RF_BLOCKi_8_Q_reg_26_inst : DFF_X1 port map( D => n3320, CK => CLK,
                           Q => n_3470, QN => 
                           DataPath_RF_bus_reg_dataout_26_port);
   DataPath_RF_BLOCKi_9_Q_reg_26_inst : DFF_X1 port map( D => n3386, CK => CLK,
                           Q => n_3471, QN => 
                           DataPath_RF_bus_reg_dataout_58_port);
   DataPath_RF_BLOCKi_10_Q_reg_26_inst : DFF_X1 port map( D => n3424, CK => CLK
                           , Q => n_3472, QN => 
                           DataPath_RF_bus_reg_dataout_90_port);
   DataPath_RF_BLOCKi_11_Q_reg_26_inst : DFF_X1 port map( D => n3462, CK => CLK
                           , Q => n_3473, QN => 
                           DataPath_RF_bus_reg_dataout_122_port);
   DataPath_RF_BLOCKi_12_Q_reg_26_inst : DFF_X1 port map( D => n3500, CK => CLK
                           , Q => n_3474, QN => 
                           DataPath_RF_bus_reg_dataout_154_port);
   DataPath_RF_BLOCKi_13_Q_reg_26_inst : DFF_X1 port map( D => n3538, CK => CLK
                           , Q => n_3475, QN => 
                           DataPath_RF_bus_reg_dataout_186_port);
   DataPath_RF_BLOCKi_14_Q_reg_26_inst : DFF_X1 port map( D => n3576, CK => CLK
                           , Q => n_3476, QN => 
                           DataPath_RF_bus_reg_dataout_218_port);
   DataPath_RF_BLOCKi_15_Q_reg_26_inst : DFF_X1 port map( D => n3614, CK => CLK
                           , Q => n_3477, QN => 
                           DataPath_RF_bus_reg_dataout_250_port);
   DataPath_RF_BLOCKi_16_Q_reg_26_inst : DFF_X1 port map( D => n3652, CK => CLK
                           , Q => n_3478, QN => 
                           DataPath_RF_bus_reg_dataout_282_port);
   DataPath_RF_BLOCKi_17_Q_reg_26_inst : DFF_X1 port map( D => n3689, CK => CLK
                           , Q => n_3479, QN => 
                           DataPath_RF_bus_reg_dataout_314_port);
   DataPath_RF_BLOCKi_18_Q_reg_26_inst : DFF_X1 port map( D => n3726, CK => CLK
                           , Q => n_3480, QN => 
                           DataPath_RF_bus_reg_dataout_346_port);
   DataPath_RF_BLOCKi_19_Q_reg_26_inst : DFF_X1 port map( D => n3763, CK => CLK
                           , Q => n_3481, QN => 
                           DataPath_RF_bus_reg_dataout_378_port);
   DataPath_RF_BLOCKi_20_Q_reg_26_inst : DFF_X1 port map( D => n3798, CK => CLK
                           , Q => n_3482, QN => 
                           DataPath_RF_bus_reg_dataout_410_port);
   DataPath_RF_BLOCKi_21_Q_reg_26_inst : DFF_X1 port map( D => n3833, CK => CLK
                           , Q => n_3483, QN => 
                           DataPath_RF_bus_reg_dataout_442_port);
   DataPath_RF_BLOCKi_22_Q_reg_26_inst : DFF_X1 port map( D => n3868, CK => CLK
                           , Q => n_3484, QN => 
                           DataPath_RF_bus_reg_dataout_474_port);
   DataPath_RF_BLOCKi_23_Q_reg_26_inst : DFF_X1 port map( D => n3908, CK => CLK
                           , Q => n_3485, QN => 
                           DataPath_RF_bus_reg_dataout_506_port);
   DataPath_RF_BLOCKi_24_Q_reg_26_inst : DFF_X1 port map( D => n3976, CK => CLK
                           , Q => n_3486, QN => 
                           DataPath_RF_bus_reg_dataout_538_port);
   DataPath_RF_BLOCKi_25_Q_reg_26_inst : DFF_X1 port map( D => n4039, CK => CLK
                           , Q => n_3487, QN => 
                           DataPath_RF_bus_reg_dataout_570_port);
   DataPath_RF_BLOCKi_26_Q_reg_26_inst : DFF_X1 port map( D => n4074, CK => CLK
                           , Q => n_3488, QN => 
                           DataPath_RF_bus_reg_dataout_602_port);
   DataPath_RF_BLOCKi_27_Q_reg_26_inst : DFF_X1 port map( D => n4109, CK => CLK
                           , Q => n_3489, QN => 
                           DataPath_RF_bus_reg_dataout_634_port);
   DataPath_RF_BLOCKi_28_Q_reg_26_inst : DFF_X1 port map( D => n4144, CK => CLK
                           , Q => n_3490, QN => 
                           DataPath_RF_bus_reg_dataout_666_port);
   DataPath_RF_BLOCKi_29_Q_reg_26_inst : DFF_X1 port map( D => n4179, CK => CLK
                           , Q => n_3491, QN => 
                           DataPath_RF_bus_reg_dataout_698_port);
   DataPath_RF_BLOCKi_30_Q_reg_26_inst : DFF_X1 port map( D => n4214, CK => CLK
                           , Q => n_3492, QN => 
                           DataPath_RF_bus_reg_dataout_730_port);
   DataPath_RF_BLOCKi_31_Q_reg_26_inst : DFF_X1 port map( D => n4249, CK => CLK
                           , Q => n_3493, QN => 
                           DataPath_RF_bus_reg_dataout_762_port);
   DataPath_RF_BLOCKi_32_Q_reg_26_inst : DFF_X1 port map( D => n4284, CK => CLK
                           , Q => n_3494, QN => 
                           DataPath_RF_bus_reg_dataout_794_port);
   DataPath_RF_BLOCKi_33_Q_reg_26_inst : DFF_X1 port map( D => n4319, CK => CLK
                           , Q => n_3495, QN => 
                           DataPath_RF_bus_reg_dataout_826_port);
   DataPath_RF_BLOCKi_34_Q_reg_26_inst : DFF_X1 port map( D => n4354, CK => CLK
                           , Q => n_3496, QN => 
                           DataPath_RF_bus_reg_dataout_858_port);
   DataPath_RF_BLOCKi_35_Q_reg_26_inst : DFF_X1 port map( D => n4389, CK => CLK
                           , Q => n_3497, QN => 
                           DataPath_RF_bus_reg_dataout_890_port);
   DataPath_RF_BLOCKi_36_Q_reg_26_inst : DFF_X1 port map( D => n4424, CK => CLK
                           , Q => n_3498, QN => 
                           DataPath_RF_bus_reg_dataout_922_port);
   DataPath_RF_BLOCKi_37_Q_reg_26_inst : DFF_X1 port map( D => n4459, CK => CLK
                           , Q => n_3499, QN => 
                           DataPath_RF_bus_reg_dataout_954_port);
   DataPath_RF_BLOCKi_38_Q_reg_26_inst : DFF_X1 port map( D => n4494, CK => CLK
                           , Q => n_3500, QN => 
                           DataPath_RF_bus_reg_dataout_986_port);
   DataPath_RF_BLOCKi_39_Q_reg_26_inst : DFF_X1 port map( D => n4529, CK => CLK
                           , Q => n_3501, QN => 
                           DataPath_RF_bus_reg_dataout_1018_port);
   DataPath_RF_BLOCKi_40_Q_reg_26_inst : DFF_X1 port map( D => n4569, CK => CLK
                           , Q => n_3502, QN => 
                           DataPath_RF_bus_reg_dataout_1050_port);
   DataPath_RF_BLOCKi_41_Q_reg_26_inst : DFF_X1 port map( D => n4632, CK => CLK
                           , Q => n_3503, QN => 
                           DataPath_RF_bus_reg_dataout_1082_port);
   DataPath_RF_BLOCKi_42_Q_reg_26_inst : DFF_X1 port map( D => n4667, CK => CLK
                           , Q => n_3504, QN => 
                           DataPath_RF_bus_reg_dataout_1114_port);
   DataPath_RF_BLOCKi_43_Q_reg_26_inst : DFF_X1 port map( D => n4702, CK => CLK
                           , Q => n_3505, QN => 
                           DataPath_RF_bus_reg_dataout_1146_port);
   DataPath_RF_BLOCKi_44_Q_reg_26_inst : DFF_X1 port map( D => n4737, CK => CLK
                           , Q => n_3506, QN => 
                           DataPath_RF_bus_reg_dataout_1178_port);
   DataPath_RF_BLOCKi_45_Q_reg_26_inst : DFF_X1 port map( D => n4772, CK => CLK
                           , Q => n_3507, QN => 
                           DataPath_RF_bus_reg_dataout_1210_port);
   DataPath_RF_BLOCKi_46_Q_reg_26_inst : DFF_X1 port map( D => n4807, CK => CLK
                           , Q => n_3508, QN => 
                           DataPath_RF_bus_reg_dataout_1242_port);
   DataPath_RF_BLOCKi_47_Q_reg_26_inst : DFF_X1 port map( D => n4842, CK => CLK
                           , Q => n_3509, QN => 
                           DataPath_RF_bus_reg_dataout_1274_port);
   DataPath_RF_BLOCKi_48_Q_reg_26_inst : DFF_X1 port map( D => n4877, CK => CLK
                           , Q => n_3510, QN => 
                           DataPath_RF_bus_reg_dataout_1306_port);
   DataPath_RF_BLOCKi_49_Q_reg_26_inst : DFF_X1 port map( D => n4912, CK => CLK
                           , Q => n_3511, QN => 
                           DataPath_RF_bus_reg_dataout_1338_port);
   DataPath_RF_BLOCKi_50_Q_reg_26_inst : DFF_X1 port map( D => n4947, CK => CLK
                           , Q => n_3512, QN => 
                           DataPath_RF_bus_reg_dataout_1370_port);
   DataPath_RF_BLOCKi_51_Q_reg_26_inst : DFF_X1 port map( D => n4982, CK => CLK
                           , Q => n_3513, QN => 
                           DataPath_RF_bus_reg_dataout_1402_port);
   DataPath_RF_BLOCKi_52_Q_reg_26_inst : DFF_X1 port map( D => n5017, CK => CLK
                           , Q => n_3514, QN => 
                           DataPath_RF_bus_reg_dataout_1434_port);
   DataPath_RF_BLOCKi_53_Q_reg_26_inst : DFF_X1 port map( D => n5052, CK => CLK
                           , Q => n_3515, QN => 
                           DataPath_RF_bus_reg_dataout_1466_port);
   DataPath_RF_BLOCKi_54_Q_reg_26_inst : DFF_X1 port map( D => n5087, CK => CLK
                           , Q => n_3516, QN => 
                           DataPath_RF_bus_reg_dataout_1498_port);
   DataPath_RF_BLOCKi_55_Q_reg_26_inst : DFF_X1 port map( D => n5122, CK => CLK
                           , Q => n_3517, QN => 
                           DataPath_RF_bus_reg_dataout_1530_port);
   DataPath_RF_BLOCKi_56_Q_reg_26_inst : DFF_X1 port map( D => n5162, CK => CLK
                           , Q => n_3518, QN => 
                           DataPath_RF_bus_reg_dataout_1562_port);
   DataPath_RF_BLOCKi_57_Q_reg_26_inst : DFF_X1 port map( D => n5224, CK => CLK
                           , Q => n_3519, QN => 
                           DataPath_RF_bus_reg_dataout_1594_port);
   DataPath_RF_BLOCKi_58_Q_reg_26_inst : DFF_X1 port map( D => n5260, CK => CLK
                           , Q => n_3520, QN => 
                           DataPath_RF_bus_reg_dataout_1626_port);
   DataPath_RF_BLOCKi_59_Q_reg_26_inst : DFF_X1 port map( D => n5295, CK => CLK
                           , Q => n_3521, QN => 
                           DataPath_RF_bus_reg_dataout_1658_port);
   DataPath_RF_BLOCKi_60_Q_reg_26_inst : DFF_X1 port map( D => n5330, CK => CLK
                           , Q => n_3522, QN => 
                           DataPath_RF_bus_reg_dataout_1690_port);
   DataPath_RF_BLOCKi_61_Q_reg_26_inst : DFF_X1 port map( D => n5365, CK => CLK
                           , Q => n_3523, QN => 
                           DataPath_RF_bus_reg_dataout_1722_port);
   DataPath_RF_BLOCKi_62_Q_reg_26_inst : DFF_X1 port map( D => n5400, CK => CLK
                           , Q => n_3524, QN => 
                           DataPath_RF_bus_reg_dataout_1754_port);
   DataPath_RF_BLOCKi_63_Q_reg_26_inst : DFF_X1 port map( D => n5435, CK => CLK
                           , Q => n_3525, QN => 
                           DataPath_RF_bus_reg_dataout_1786_port);
   DataPath_RF_BLOCKi_64_Q_reg_26_inst : DFF_X1 port map( D => n5470, CK => CLK
                           , Q => n_3526, QN => 
                           DataPath_RF_bus_reg_dataout_1818_port);
   DataPath_RF_BLOCKi_65_Q_reg_26_inst : DFF_X1 port map( D => n5505, CK => CLK
                           , Q => n_3527, QN => 
                           DataPath_RF_bus_reg_dataout_1850_port);
   DataPath_RF_BLOCKi_66_Q_reg_26_inst : DFF_X1 port map( D => n5540, CK => CLK
                           , Q => n_3528, QN => 
                           DataPath_RF_bus_reg_dataout_1882_port);
   DataPath_RF_BLOCKi_67_Q_reg_26_inst : DFF_X1 port map( D => n5575, CK => CLK
                           , Q => n_3529, QN => 
                           DataPath_RF_bus_reg_dataout_1914_port);
   DataPath_RF_BLOCKi_68_Q_reg_26_inst : DFF_X1 port map( D => n5614, CK => CLK
                           , Q => n_3530, QN => 
                           DataPath_RF_bus_reg_dataout_1946_port);
   DataPath_RF_BLOCKi_69_Q_reg_26_inst : DFF_X1 port map( D => n5651, CK => CLK
                           , Q => n_3531, QN => 
                           DataPath_RF_bus_reg_dataout_1978_port);
   DataPath_RF_BLOCKi_70_Q_reg_26_inst : DFF_X1 port map( D => n5688, CK => CLK
                           , Q => n_3532, QN => 
                           DataPath_RF_bus_reg_dataout_2010_port);
   DataPath_RF_BLOCKi_71_Q_reg_26_inst : DFF_X1 port map( D => n5725, CK => CLK
                           , Q => n_3533, QN => 
                           DataPath_RF_bus_reg_dataout_2042_port);
   DataPath_RF_BLOCKi_83_Q_reg_26_inst : DFF_X1 port map( D => n926, CK => CLK,
                           Q => n_3534, QN => 
                           DataPath_RF_bus_reg_dataout_2426_port);
   DataPath_RF_BLOCKi_84_Q_reg_26_inst : DFF_X1 port map( D => n975, CK => CLK,
                           Q => n_3535, QN => 
                           DataPath_RF_bus_reg_dataout_2458_port);
   DataPath_RF_BLOCKi_85_Q_reg_26_inst : DFF_X1 port map( D => n1012, CK => CLK
                           , Q => n_3536, QN => 
                           DataPath_RF_bus_reg_dataout_2490_port);
   DataPath_RF_BLOCKi_86_Q_reg_26_inst : DFF_X1 port map( D => n1049, CK => CLK
                           , Q => n_3537, QN => 
                           DataPath_RF_bus_reg_dataout_2522_port);
   DataPath_RF_BLOCKi_87_Q_reg_26_inst : DFF_X1 port map( D => n1086, CK => CLK
                           , Q => n_3538, QN => 
                           DataPath_RF_bus_reg_dataout_2554_port);
   DataPath_RF_BLOCKi_72_Q_reg_26_inst : DFF_X1 port map( D => n5762, CK => CLK
                           , Q => n_3539, QN => 
                           DataPath_RF_bus_reg_dataout_2074_port);
   DataPath_RF_BLOCKi_73_Q_reg_26_inst : DFF_X1 port map( D => n5801, CK => CLK
                           , Q => n_3540, QN => 
                           DataPath_RF_bus_reg_dataout_2106_port);
   DataPath_RF_BLOCKi_74_Q_reg_26_inst : DFF_X1 port map( D => n5837, CK => CLK
                           , Q => n_3541, QN => 
                           DataPath_RF_bus_reg_dataout_2138_port);
   DataPath_RF_BLOCKi_75_Q_reg_26_inst : DFF_X1 port map( D => n5873, CK => CLK
                           , Q => n_3542, QN => 
                           DataPath_RF_bus_reg_dataout_2170_port);
   DataPath_RF_BLOCKi_76_Q_reg_26_inst : DFF_X1 port map( D => n5909, CK => CLK
                           , Q => n_3543, QN => 
                           DataPath_RF_bus_reg_dataout_2202_port);
   DataPath_RF_BLOCKi_77_Q_reg_26_inst : DFF_X1 port map( D => n5945, CK => CLK
                           , Q => n_3544, QN => 
                           DataPath_RF_bus_reg_dataout_2234_port);
   DataPath_RF_BLOCKi_78_Q_reg_26_inst : DFF_X1 port map( D => n5981, CK => CLK
                           , Q => n_3545, QN => 
                           DataPath_RF_bus_reg_dataout_2266_port);
   DataPath_RF_BLOCKi_79_Q_reg_26_inst : DFF_X1 port map( D => n6017, CK => CLK
                           , Q => n_3546, QN => 
                           DataPath_RF_bus_reg_dataout_2298_port);
   DataPath_RF_BLOCKi_80_Q_reg_26_inst : DFF_X1 port map( D => n6054, CK => CLK
                           , Q => n_3547, QN => 
                           DataPath_RF_bus_reg_dataout_2330_port);
   DataPath_RF_BLOCKi_81_Q_reg_26_inst : DFF_X1 port map( D => n6090, CK => CLK
                           , Q => n_3548, QN => 
                           DataPath_RF_bus_reg_dataout_2362_port);
   DataPath_RF_BLOCKi_82_Q_reg_26_inst : DFF_X1 port map( D => n6124, CK => CLK
                           , Q => n_3549, QN => 
                           DataPath_RF_bus_reg_dataout_2394_port);
   DataPath_REG_ALU_OUT_Q_reg_27_inst : DFF_X1 port map( D => n6996, CK => CLK,
                           Q => DRAM_ADDRESS_27_port, QN => n512);
   DataPath_REG_MEM_ALUOUT_Q_reg_27_inst : DFF_X1 port map( D => n1122, CK => 
                           CLK, Q => n_3550, QN => 
                           DataPath_i_REG_MEM_ALUOUT_27_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_27_inst : DFF_X1 port map( D => n6772, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_59_port,
                           QN => n626);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_27_inst : DFF_X1 port map( D => n6804, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_91_port,
                           QN => n658);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_27_inst : DFF_X1 port map( D => n6836, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_123_port
                           , QN => n690);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_27_inst : DFF_X1 port map( D => n6868, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_155_port
                           , QN => n722);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_27_inst : DFF_X1 port map( D => n6900, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_187_port
                           , QN => n754);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_27_inst : DFF_X1 port map( D => n6932, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_219_port
                           , QN => n786);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_27_inst : DFF_X1 port map( D => n6964, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_251_port
                           , QN => n818);
   DataPath_RF_BLOCKi_8_Q_reg_27_inst : DFF_X1 port map( D => n3318, CK => CLK,
                           Q => n_3551, QN => 
                           DataPath_RF_bus_reg_dataout_27_port);
   DataPath_RF_BLOCKi_9_Q_reg_27_inst : DFF_X1 port map( D => n3385, CK => CLK,
                           Q => n_3552, QN => 
                           DataPath_RF_bus_reg_dataout_59_port);
   DataPath_RF_BLOCKi_10_Q_reg_27_inst : DFF_X1 port map( D => n3423, CK => CLK
                           , Q => n_3553, QN => 
                           DataPath_RF_bus_reg_dataout_91_port);
   DataPath_RF_BLOCKi_11_Q_reg_27_inst : DFF_X1 port map( D => n3461, CK => CLK
                           , Q => n_3554, QN => 
                           DataPath_RF_bus_reg_dataout_123_port);
   DataPath_RF_BLOCKi_12_Q_reg_27_inst : DFF_X1 port map( D => n3499, CK => CLK
                           , Q => n_3555, QN => 
                           DataPath_RF_bus_reg_dataout_155_port);
   DataPath_RF_BLOCKi_13_Q_reg_27_inst : DFF_X1 port map( D => n3537, CK => CLK
                           , Q => n_3556, QN => 
                           DataPath_RF_bus_reg_dataout_187_port);
   DataPath_RF_BLOCKi_14_Q_reg_27_inst : DFF_X1 port map( D => n3575, CK => CLK
                           , Q => n_3557, QN => 
                           DataPath_RF_bus_reg_dataout_219_port);
   DataPath_RF_BLOCKi_15_Q_reg_27_inst : DFF_X1 port map( D => n3613, CK => CLK
                           , Q => n_3558, QN => 
                           DataPath_RF_bus_reg_dataout_251_port);
   DataPath_RF_BLOCKi_16_Q_reg_27_inst : DFF_X1 port map( D => n3651, CK => CLK
                           , Q => n_3559, QN => 
                           DataPath_RF_bus_reg_dataout_283_port);
   DataPath_RF_BLOCKi_17_Q_reg_27_inst : DFF_X1 port map( D => n3688, CK => CLK
                           , Q => n_3560, QN => 
                           DataPath_RF_bus_reg_dataout_315_port);
   DataPath_RF_BLOCKi_18_Q_reg_27_inst : DFF_X1 port map( D => n3725, CK => CLK
                           , Q => n_3561, QN => 
                           DataPath_RF_bus_reg_dataout_347_port);
   DataPath_RF_BLOCKi_19_Q_reg_27_inst : DFF_X1 port map( D => n3762, CK => CLK
                           , Q => n_3562, QN => 
                           DataPath_RF_bus_reg_dataout_379_port);
   DataPath_RF_BLOCKi_20_Q_reg_27_inst : DFF_X1 port map( D => n3797, CK => CLK
                           , Q => n_3563, QN => 
                           DataPath_RF_bus_reg_dataout_411_port);
   DataPath_RF_BLOCKi_21_Q_reg_27_inst : DFF_X1 port map( D => n3832, CK => CLK
                           , Q => n_3564, QN => 
                           DataPath_RF_bus_reg_dataout_443_port);
   DataPath_RF_BLOCKi_22_Q_reg_27_inst : DFF_X1 port map( D => n3867, CK => CLK
                           , Q => n_3565, QN => 
                           DataPath_RF_bus_reg_dataout_475_port);
   DataPath_RF_BLOCKi_23_Q_reg_27_inst : DFF_X1 port map( D => n3906, CK => CLK
                           , Q => n_3566, QN => 
                           DataPath_RF_bus_reg_dataout_507_port);
   DataPath_RF_BLOCKi_24_Q_reg_27_inst : DFF_X1 port map( D => n3974, CK => CLK
                           , Q => n_3567, QN => 
                           DataPath_RF_bus_reg_dataout_539_port);
   DataPath_RF_BLOCKi_25_Q_reg_27_inst : DFF_X1 port map( D => n4038, CK => CLK
                           , Q => n_3568, QN => 
                           DataPath_RF_bus_reg_dataout_571_port);
   DataPath_RF_BLOCKi_26_Q_reg_27_inst : DFF_X1 port map( D => n4073, CK => CLK
                           , Q => n_3569, QN => 
                           DataPath_RF_bus_reg_dataout_603_port);
   DataPath_RF_BLOCKi_27_Q_reg_27_inst : DFF_X1 port map( D => n4108, CK => CLK
                           , Q => n_3570, QN => 
                           DataPath_RF_bus_reg_dataout_635_port);
   DataPath_RF_BLOCKi_28_Q_reg_27_inst : DFF_X1 port map( D => n4143, CK => CLK
                           , Q => n_3571, QN => 
                           DataPath_RF_bus_reg_dataout_667_port);
   DataPath_RF_BLOCKi_29_Q_reg_27_inst : DFF_X1 port map( D => n4178, CK => CLK
                           , Q => n_3572, QN => 
                           DataPath_RF_bus_reg_dataout_699_port);
   DataPath_RF_BLOCKi_30_Q_reg_27_inst : DFF_X1 port map( D => n4213, CK => CLK
                           , Q => n_3573, QN => 
                           DataPath_RF_bus_reg_dataout_731_port);
   DataPath_RF_BLOCKi_31_Q_reg_27_inst : DFF_X1 port map( D => n4248, CK => CLK
                           , Q => n_3574, QN => 
                           DataPath_RF_bus_reg_dataout_763_port);
   DataPath_RF_BLOCKi_32_Q_reg_27_inst : DFF_X1 port map( D => n4283, CK => CLK
                           , Q => n_3575, QN => 
                           DataPath_RF_bus_reg_dataout_795_port);
   DataPath_RF_BLOCKi_33_Q_reg_27_inst : DFF_X1 port map( D => n4318, CK => CLK
                           , Q => n_3576, QN => 
                           DataPath_RF_bus_reg_dataout_827_port);
   DataPath_RF_BLOCKi_34_Q_reg_27_inst : DFF_X1 port map( D => n4353, CK => CLK
                           , Q => n_3577, QN => 
                           DataPath_RF_bus_reg_dataout_859_port);
   DataPath_RF_BLOCKi_35_Q_reg_27_inst : DFF_X1 port map( D => n4388, CK => CLK
                           , Q => n_3578, QN => 
                           DataPath_RF_bus_reg_dataout_891_port);
   DataPath_RF_BLOCKi_36_Q_reg_27_inst : DFF_X1 port map( D => n4423, CK => CLK
                           , Q => n_3579, QN => 
                           DataPath_RF_bus_reg_dataout_923_port);
   DataPath_RF_BLOCKi_37_Q_reg_27_inst : DFF_X1 port map( D => n4458, CK => CLK
                           , Q => n_3580, QN => 
                           DataPath_RF_bus_reg_dataout_955_port);
   DataPath_RF_BLOCKi_38_Q_reg_27_inst : DFF_X1 port map( D => n4493, CK => CLK
                           , Q => n_3581, QN => 
                           DataPath_RF_bus_reg_dataout_987_port);
   DataPath_RF_BLOCKi_39_Q_reg_27_inst : DFF_X1 port map( D => n4528, CK => CLK
                           , Q => n_3582, QN => 
                           DataPath_RF_bus_reg_dataout_1019_port);
   DataPath_RF_BLOCKi_40_Q_reg_27_inst : DFF_X1 port map( D => n4567, CK => CLK
                           , Q => n_3583, QN => 
                           DataPath_RF_bus_reg_dataout_1051_port);
   DataPath_RF_BLOCKi_41_Q_reg_27_inst : DFF_X1 port map( D => n4631, CK => CLK
                           , Q => n_3584, QN => 
                           DataPath_RF_bus_reg_dataout_1083_port);
   DataPath_RF_BLOCKi_42_Q_reg_27_inst : DFF_X1 port map( D => n4666, CK => CLK
                           , Q => n_3585, QN => 
                           DataPath_RF_bus_reg_dataout_1115_port);
   DataPath_RF_BLOCKi_43_Q_reg_27_inst : DFF_X1 port map( D => n4701, CK => CLK
                           , Q => n_3586, QN => 
                           DataPath_RF_bus_reg_dataout_1147_port);
   DataPath_RF_BLOCKi_44_Q_reg_27_inst : DFF_X1 port map( D => n4736, CK => CLK
                           , Q => n_3587, QN => 
                           DataPath_RF_bus_reg_dataout_1179_port);
   DataPath_RF_BLOCKi_45_Q_reg_27_inst : DFF_X1 port map( D => n4771, CK => CLK
                           , Q => n_3588, QN => 
                           DataPath_RF_bus_reg_dataout_1211_port);
   DataPath_RF_BLOCKi_46_Q_reg_27_inst : DFF_X1 port map( D => n4806, CK => CLK
                           , Q => n_3589, QN => 
                           DataPath_RF_bus_reg_dataout_1243_port);
   DataPath_RF_BLOCKi_47_Q_reg_27_inst : DFF_X1 port map( D => n4841, CK => CLK
                           , Q => n_3590, QN => 
                           DataPath_RF_bus_reg_dataout_1275_port);
   DataPath_RF_BLOCKi_48_Q_reg_27_inst : DFF_X1 port map( D => n4876, CK => CLK
                           , Q => n_3591, QN => 
                           DataPath_RF_bus_reg_dataout_1307_port);
   DataPath_RF_BLOCKi_49_Q_reg_27_inst : DFF_X1 port map( D => n4911, CK => CLK
                           , Q => n_3592, QN => 
                           DataPath_RF_bus_reg_dataout_1339_port);
   DataPath_RF_BLOCKi_50_Q_reg_27_inst : DFF_X1 port map( D => n4946, CK => CLK
                           , Q => n_3593, QN => 
                           DataPath_RF_bus_reg_dataout_1371_port);
   DataPath_RF_BLOCKi_51_Q_reg_27_inst : DFF_X1 port map( D => n4981, CK => CLK
                           , Q => n_3594, QN => 
                           DataPath_RF_bus_reg_dataout_1403_port);
   DataPath_RF_BLOCKi_52_Q_reg_27_inst : DFF_X1 port map( D => n5016, CK => CLK
                           , Q => n_3595, QN => 
                           DataPath_RF_bus_reg_dataout_1435_port);
   DataPath_RF_BLOCKi_53_Q_reg_27_inst : DFF_X1 port map( D => n5051, CK => CLK
                           , Q => n_3596, QN => 
                           DataPath_RF_bus_reg_dataout_1467_port);
   DataPath_RF_BLOCKi_54_Q_reg_27_inst : DFF_X1 port map( D => n5086, CK => CLK
                           , Q => n_3597, QN => 
                           DataPath_RF_bus_reg_dataout_1499_port);
   DataPath_RF_BLOCKi_55_Q_reg_27_inst : DFF_X1 port map( D => n5121, CK => CLK
                           , Q => n_3598, QN => 
                           DataPath_RF_bus_reg_dataout_1531_port);
   DataPath_RF_BLOCKi_56_Q_reg_27_inst : DFF_X1 port map( D => n5160, CK => CLK
                           , Q => n_3599, QN => 
                           DataPath_RF_bus_reg_dataout_1563_port);
   DataPath_RF_BLOCKi_57_Q_reg_27_inst : DFF_X1 port map( D => n5223, CK => CLK
                           , Q => n_3600, QN => 
                           DataPath_RF_bus_reg_dataout_1595_port);
   DataPath_RF_BLOCKi_58_Q_reg_27_inst : DFF_X1 port map( D => n5259, CK => CLK
                           , Q => n_3601, QN => 
                           DataPath_RF_bus_reg_dataout_1627_port);
   DataPath_RF_BLOCKi_59_Q_reg_27_inst : DFF_X1 port map( D => n5294, CK => CLK
                           , Q => n_3602, QN => 
                           DataPath_RF_bus_reg_dataout_1659_port);
   DataPath_RF_BLOCKi_60_Q_reg_27_inst : DFF_X1 port map( D => n5329, CK => CLK
                           , Q => n_3603, QN => 
                           DataPath_RF_bus_reg_dataout_1691_port);
   DataPath_RF_BLOCKi_61_Q_reg_27_inst : DFF_X1 port map( D => n5364, CK => CLK
                           , Q => n_3604, QN => 
                           DataPath_RF_bus_reg_dataout_1723_port);
   DataPath_RF_BLOCKi_62_Q_reg_27_inst : DFF_X1 port map( D => n5399, CK => CLK
                           , Q => n_3605, QN => 
                           DataPath_RF_bus_reg_dataout_1755_port);
   DataPath_RF_BLOCKi_63_Q_reg_27_inst : DFF_X1 port map( D => n5434, CK => CLK
                           , Q => n_3606, QN => 
                           DataPath_RF_bus_reg_dataout_1787_port);
   DataPath_RF_BLOCKi_64_Q_reg_27_inst : DFF_X1 port map( D => n5469, CK => CLK
                           , Q => n_3607, QN => 
                           DataPath_RF_bus_reg_dataout_1819_port);
   DataPath_RF_BLOCKi_65_Q_reg_27_inst : DFF_X1 port map( D => n5504, CK => CLK
                           , Q => n_3608, QN => 
                           DataPath_RF_bus_reg_dataout_1851_port);
   DataPath_RF_BLOCKi_66_Q_reg_27_inst : DFF_X1 port map( D => n5539, CK => CLK
                           , Q => n_3609, QN => 
                           DataPath_RF_bus_reg_dataout_1883_port);
   DataPath_RF_BLOCKi_67_Q_reg_27_inst : DFF_X1 port map( D => n5574, CK => CLK
                           , Q => n_3610, QN => 
                           DataPath_RF_bus_reg_dataout_1915_port);
   DataPath_RF_BLOCKi_68_Q_reg_27_inst : DFF_X1 port map( D => n5613, CK => CLK
                           , Q => n_3611, QN => 
                           DataPath_RF_bus_reg_dataout_1947_port);
   DataPath_RF_BLOCKi_69_Q_reg_27_inst : DFF_X1 port map( D => n5650, CK => CLK
                           , Q => n_3612, QN => 
                           DataPath_RF_bus_reg_dataout_1979_port);
   DataPath_RF_BLOCKi_70_Q_reg_27_inst : DFF_X1 port map( D => n5687, CK => CLK
                           , Q => n_3613, QN => 
                           DataPath_RF_bus_reg_dataout_2011_port);
   DataPath_RF_BLOCKi_71_Q_reg_27_inst : DFF_X1 port map( D => n5724, CK => CLK
                           , Q => n_3614, QN => 
                           DataPath_RF_bus_reg_dataout_2043_port);
   DataPath_RF_BLOCKi_83_Q_reg_27_inst : DFF_X1 port map( D => n924, CK => CLK,
                           Q => n_3615, QN => 
                           DataPath_RF_bus_reg_dataout_2427_port);
   DataPath_RF_BLOCKi_84_Q_reg_27_inst : DFF_X1 port map( D => n974, CK => CLK,
                           Q => n_3616, QN => 
                           DataPath_RF_bus_reg_dataout_2459_port);
   DataPath_RF_BLOCKi_85_Q_reg_27_inst : DFF_X1 port map( D => n1011, CK => CLK
                           , Q => n_3617, QN => 
                           DataPath_RF_bus_reg_dataout_2491_port);
   DataPath_RF_BLOCKi_86_Q_reg_27_inst : DFF_X1 port map( D => n1048, CK => CLK
                           , Q => n_3618, QN => 
                           DataPath_RF_bus_reg_dataout_2523_port);
   DataPath_RF_BLOCKi_87_Q_reg_27_inst : DFF_X1 port map( D => n1085, CK => CLK
                           , Q => n_3619, QN => 
                           DataPath_RF_bus_reg_dataout_2555_port);
   DataPath_RF_BLOCKi_72_Q_reg_27_inst : DFF_X1 port map( D => n5761, CK => CLK
                           , Q => n_3620, QN => 
                           DataPath_RF_bus_reg_dataout_2075_port);
   DataPath_RF_BLOCKi_73_Q_reg_27_inst : DFF_X1 port map( D => n5800, CK => CLK
                           , Q => n_3621, QN => 
                           DataPath_RF_bus_reg_dataout_2107_port);
   DataPath_RF_BLOCKi_74_Q_reg_27_inst : DFF_X1 port map( D => n5836, CK => CLK
                           , Q => n_3622, QN => 
                           DataPath_RF_bus_reg_dataout_2139_port);
   DataPath_RF_BLOCKi_75_Q_reg_27_inst : DFF_X1 port map( D => n5872, CK => CLK
                           , Q => n_3623, QN => 
                           DataPath_RF_bus_reg_dataout_2171_port);
   DataPath_RF_BLOCKi_76_Q_reg_27_inst : DFF_X1 port map( D => n5908, CK => CLK
                           , Q => n_3624, QN => 
                           DataPath_RF_bus_reg_dataout_2203_port);
   DataPath_RF_BLOCKi_77_Q_reg_27_inst : DFF_X1 port map( D => n5944, CK => CLK
                           , Q => n_3625, QN => 
                           DataPath_RF_bus_reg_dataout_2235_port);
   DataPath_RF_BLOCKi_78_Q_reg_27_inst : DFF_X1 port map( D => n5980, CK => CLK
                           , Q => n_3626, QN => 
                           DataPath_RF_bus_reg_dataout_2267_port);
   DataPath_RF_BLOCKi_79_Q_reg_27_inst : DFF_X1 port map( D => n6016, CK => CLK
                           , Q => n_3627, QN => 
                           DataPath_RF_bus_reg_dataout_2299_port);
   DataPath_RF_BLOCKi_80_Q_reg_27_inst : DFF_X1 port map( D => n6053, CK => CLK
                           , Q => n_3628, QN => 
                           DataPath_RF_bus_reg_dataout_2331_port);
   DataPath_RF_BLOCKi_81_Q_reg_27_inst : DFF_X1 port map( D => n6089, CK => CLK
                           , Q => n_3629, QN => 
                           DataPath_RF_bus_reg_dataout_2363_port);
   DataPath_RF_BLOCKi_82_Q_reg_27_inst : DFF_X1 port map( D => n6123, CK => CLK
                           , Q => n_3630, QN => 
                           DataPath_RF_bus_reg_dataout_2395_port);
   DataPath_REG_ALU_OUT_Q_reg_28_inst : DFF_X1 port map( D => n6995, CK => CLK,
                           Q => DRAM_ADDRESS_28_port, QN => n513);
   DataPath_REG_MEM_ALUOUT_Q_reg_28_inst : DFF_X1 port map( D => n1121, CK => 
                           CLK, Q => n_3631, QN => 
                           DataPath_i_REG_MEM_ALUOUT_28_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_28_inst : DFF_X1 port map( D => n6771, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_60_port,
                           QN => n627);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_28_inst : DFF_X1 port map( D => n6803, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_92_port,
                           QN => n659);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_28_inst : DFF_X1 port map( D => n6835, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_124_port
                           , QN => n691);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_28_inst : DFF_X1 port map( D => n6867, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_156_port
                           , QN => n723);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_28_inst : DFF_X1 port map( D => n6899, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_188_port
                           , QN => n755);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_28_inst : DFF_X1 port map( D => n6931, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_220_port
                           , QN => n787);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_28_inst : DFF_X1 port map( D => n6963, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_252_port
                           , QN => n819);
   DataPath_RF_BLOCKi_8_Q_reg_28_inst : DFF_X1 port map( D => n3316, CK => CLK,
                           Q => n_3632, QN => 
                           DataPath_RF_bus_reg_dataout_28_port);
   DataPath_RF_BLOCKi_9_Q_reg_28_inst : DFF_X1 port map( D => n3384, CK => CLK,
                           Q => n_3633, QN => 
                           DataPath_RF_bus_reg_dataout_60_port);
   DataPath_RF_BLOCKi_10_Q_reg_28_inst : DFF_X1 port map( D => n3422, CK => CLK
                           , Q => n_3634, QN => 
                           DataPath_RF_bus_reg_dataout_92_port);
   DataPath_RF_BLOCKi_11_Q_reg_28_inst : DFF_X1 port map( D => n3460, CK => CLK
                           , Q => n_3635, QN => 
                           DataPath_RF_bus_reg_dataout_124_port);
   DataPath_RF_BLOCKi_12_Q_reg_28_inst : DFF_X1 port map( D => n3498, CK => CLK
                           , Q => n_3636, QN => 
                           DataPath_RF_bus_reg_dataout_156_port);
   DataPath_RF_BLOCKi_13_Q_reg_28_inst : DFF_X1 port map( D => n3536, CK => CLK
                           , Q => n_3637, QN => 
                           DataPath_RF_bus_reg_dataout_188_port);
   DataPath_RF_BLOCKi_14_Q_reg_28_inst : DFF_X1 port map( D => n3574, CK => CLK
                           , Q => n_3638, QN => 
                           DataPath_RF_bus_reg_dataout_220_port);
   DataPath_RF_BLOCKi_15_Q_reg_28_inst : DFF_X1 port map( D => n3612, CK => CLK
                           , Q => n_3639, QN => 
                           DataPath_RF_bus_reg_dataout_252_port);
   DataPath_RF_BLOCKi_16_Q_reg_28_inst : DFF_X1 port map( D => n3650, CK => CLK
                           , Q => n_3640, QN => 
                           DataPath_RF_bus_reg_dataout_284_port);
   DataPath_RF_BLOCKi_17_Q_reg_28_inst : DFF_X1 port map( D => n3687, CK => CLK
                           , Q => n_3641, QN => 
                           DataPath_RF_bus_reg_dataout_316_port);
   DataPath_RF_BLOCKi_18_Q_reg_28_inst : DFF_X1 port map( D => n3724, CK => CLK
                           , Q => n_3642, QN => 
                           DataPath_RF_bus_reg_dataout_348_port);
   DataPath_RF_BLOCKi_19_Q_reg_28_inst : DFF_X1 port map( D => n3761, CK => CLK
                           , Q => n_3643, QN => 
                           DataPath_RF_bus_reg_dataout_380_port);
   DataPath_RF_BLOCKi_20_Q_reg_28_inst : DFF_X1 port map( D => n3796, CK => CLK
                           , Q => n_3644, QN => 
                           DataPath_RF_bus_reg_dataout_412_port);
   DataPath_RF_BLOCKi_21_Q_reg_28_inst : DFF_X1 port map( D => n3831, CK => CLK
                           , Q => n_3645, QN => 
                           DataPath_RF_bus_reg_dataout_444_port);
   DataPath_RF_BLOCKi_22_Q_reg_28_inst : DFF_X1 port map( D => n3866, CK => CLK
                           , Q => n_3646, QN => 
                           DataPath_RF_bus_reg_dataout_476_port);
   DataPath_RF_BLOCKi_23_Q_reg_28_inst : DFF_X1 port map( D => n3904, CK => CLK
                           , Q => n_3647, QN => 
                           DataPath_RF_bus_reg_dataout_508_port);
   DataPath_RF_BLOCKi_24_Q_reg_28_inst : DFF_X1 port map( D => n3972, CK => CLK
                           , Q => n_3648, QN => 
                           DataPath_RF_bus_reg_dataout_540_port);
   DataPath_RF_BLOCKi_25_Q_reg_28_inst : DFF_X1 port map( D => n4037, CK => CLK
                           , Q => n_3649, QN => 
                           DataPath_RF_bus_reg_dataout_572_port);
   DataPath_RF_BLOCKi_26_Q_reg_28_inst : DFF_X1 port map( D => n4072, CK => CLK
                           , Q => n_3650, QN => 
                           DataPath_RF_bus_reg_dataout_604_port);
   DataPath_RF_BLOCKi_27_Q_reg_28_inst : DFF_X1 port map( D => n4107, CK => CLK
                           , Q => n_3651, QN => 
                           DataPath_RF_bus_reg_dataout_636_port);
   DataPath_RF_BLOCKi_28_Q_reg_28_inst : DFF_X1 port map( D => n4142, CK => CLK
                           , Q => n_3652, QN => 
                           DataPath_RF_bus_reg_dataout_668_port);
   DataPath_RF_BLOCKi_29_Q_reg_28_inst : DFF_X1 port map( D => n4177, CK => CLK
                           , Q => n_3653, QN => 
                           DataPath_RF_bus_reg_dataout_700_port);
   DataPath_RF_BLOCKi_30_Q_reg_28_inst : DFF_X1 port map( D => n4212, CK => CLK
                           , Q => n_3654, QN => 
                           DataPath_RF_bus_reg_dataout_732_port);
   DataPath_RF_BLOCKi_31_Q_reg_28_inst : DFF_X1 port map( D => n4247, CK => CLK
                           , Q => n_3655, QN => 
                           DataPath_RF_bus_reg_dataout_764_port);
   DataPath_RF_BLOCKi_32_Q_reg_28_inst : DFF_X1 port map( D => n4282, CK => CLK
                           , Q => n_3656, QN => 
                           DataPath_RF_bus_reg_dataout_796_port);
   DataPath_RF_BLOCKi_33_Q_reg_28_inst : DFF_X1 port map( D => n4317, CK => CLK
                           , Q => n_3657, QN => 
                           DataPath_RF_bus_reg_dataout_828_port);
   DataPath_RF_BLOCKi_34_Q_reg_28_inst : DFF_X1 port map( D => n4352, CK => CLK
                           , Q => n_3658, QN => 
                           DataPath_RF_bus_reg_dataout_860_port);
   DataPath_RF_BLOCKi_35_Q_reg_28_inst : DFF_X1 port map( D => n4387, CK => CLK
                           , Q => n_3659, QN => 
                           DataPath_RF_bus_reg_dataout_892_port);
   DataPath_RF_BLOCKi_36_Q_reg_28_inst : DFF_X1 port map( D => n4422, CK => CLK
                           , Q => n_3660, QN => 
                           DataPath_RF_bus_reg_dataout_924_port);
   DataPath_RF_BLOCKi_37_Q_reg_28_inst : DFF_X1 port map( D => n4457, CK => CLK
                           , Q => n_3661, QN => 
                           DataPath_RF_bus_reg_dataout_956_port);
   DataPath_RF_BLOCKi_38_Q_reg_28_inst : DFF_X1 port map( D => n4492, CK => CLK
                           , Q => n_3662, QN => 
                           DataPath_RF_bus_reg_dataout_988_port);
   DataPath_RF_BLOCKi_39_Q_reg_28_inst : DFF_X1 port map( D => n4527, CK => CLK
                           , Q => n_3663, QN => 
                           DataPath_RF_bus_reg_dataout_1020_port);
   DataPath_RF_BLOCKi_40_Q_reg_28_inst : DFF_X1 port map( D => n4565, CK => CLK
                           , Q => n_3664, QN => 
                           DataPath_RF_bus_reg_dataout_1052_port);
   DataPath_RF_BLOCKi_41_Q_reg_28_inst : DFF_X1 port map( D => n4630, CK => CLK
                           , Q => n_3665, QN => 
                           DataPath_RF_bus_reg_dataout_1084_port);
   DataPath_RF_BLOCKi_42_Q_reg_28_inst : DFF_X1 port map( D => n4665, CK => CLK
                           , Q => n_3666, QN => 
                           DataPath_RF_bus_reg_dataout_1116_port);
   DataPath_RF_BLOCKi_43_Q_reg_28_inst : DFF_X1 port map( D => n4700, CK => CLK
                           , Q => n_3667, QN => 
                           DataPath_RF_bus_reg_dataout_1148_port);
   DataPath_RF_BLOCKi_44_Q_reg_28_inst : DFF_X1 port map( D => n4735, CK => CLK
                           , Q => n_3668, QN => 
                           DataPath_RF_bus_reg_dataout_1180_port);
   DataPath_RF_BLOCKi_45_Q_reg_28_inst : DFF_X1 port map( D => n4770, CK => CLK
                           , Q => n_3669, QN => 
                           DataPath_RF_bus_reg_dataout_1212_port);
   DataPath_RF_BLOCKi_46_Q_reg_28_inst : DFF_X1 port map( D => n4805, CK => CLK
                           , Q => n_3670, QN => 
                           DataPath_RF_bus_reg_dataout_1244_port);
   DataPath_RF_BLOCKi_47_Q_reg_28_inst : DFF_X1 port map( D => n4840, CK => CLK
                           , Q => n_3671, QN => 
                           DataPath_RF_bus_reg_dataout_1276_port);
   DataPath_RF_BLOCKi_48_Q_reg_28_inst : DFF_X1 port map( D => n4875, CK => CLK
                           , Q => n_3672, QN => 
                           DataPath_RF_bus_reg_dataout_1308_port);
   DataPath_RF_BLOCKi_49_Q_reg_28_inst : DFF_X1 port map( D => n4910, CK => CLK
                           , Q => n_3673, QN => 
                           DataPath_RF_bus_reg_dataout_1340_port);
   DataPath_RF_BLOCKi_50_Q_reg_28_inst : DFF_X1 port map( D => n4945, CK => CLK
                           , Q => n_3674, QN => 
                           DataPath_RF_bus_reg_dataout_1372_port);
   DataPath_RF_BLOCKi_51_Q_reg_28_inst : DFF_X1 port map( D => n4980, CK => CLK
                           , Q => n_3675, QN => 
                           DataPath_RF_bus_reg_dataout_1404_port);
   DataPath_RF_BLOCKi_52_Q_reg_28_inst : DFF_X1 port map( D => n5015, CK => CLK
                           , Q => n_3676, QN => 
                           DataPath_RF_bus_reg_dataout_1436_port);
   DataPath_RF_BLOCKi_53_Q_reg_28_inst : DFF_X1 port map( D => n5050, CK => CLK
                           , Q => n_3677, QN => 
                           DataPath_RF_bus_reg_dataout_1468_port);
   DataPath_RF_BLOCKi_54_Q_reg_28_inst : DFF_X1 port map( D => n5085, CK => CLK
                           , Q => n_3678, QN => 
                           DataPath_RF_bus_reg_dataout_1500_port);
   DataPath_RF_BLOCKi_55_Q_reg_28_inst : DFF_X1 port map( D => n5120, CK => CLK
                           , Q => n_3679, QN => 
                           DataPath_RF_bus_reg_dataout_1532_port);
   DataPath_RF_BLOCKi_56_Q_reg_28_inst : DFF_X1 port map( D => n5158, CK => CLK
                           , Q => n_3680, QN => 
                           DataPath_RF_bus_reg_dataout_1564_port);
   DataPath_RF_BLOCKi_57_Q_reg_28_inst : DFF_X1 port map( D => n5222, CK => CLK
                           , Q => n_3681, QN => 
                           DataPath_RF_bus_reg_dataout_1596_port);
   DataPath_RF_BLOCKi_58_Q_reg_28_inst : DFF_X1 port map( D => n5258, CK => CLK
                           , Q => n_3682, QN => 
                           DataPath_RF_bus_reg_dataout_1628_port);
   DataPath_RF_BLOCKi_59_Q_reg_28_inst : DFF_X1 port map( D => n5293, CK => CLK
                           , Q => n_3683, QN => 
                           DataPath_RF_bus_reg_dataout_1660_port);
   DataPath_RF_BLOCKi_60_Q_reg_28_inst : DFF_X1 port map( D => n5328, CK => CLK
                           , Q => n_3684, QN => 
                           DataPath_RF_bus_reg_dataout_1692_port);
   DataPath_RF_BLOCKi_61_Q_reg_28_inst : DFF_X1 port map( D => n5363, CK => CLK
                           , Q => n_3685, QN => 
                           DataPath_RF_bus_reg_dataout_1724_port);
   DataPath_RF_BLOCKi_62_Q_reg_28_inst : DFF_X1 port map( D => n5398, CK => CLK
                           , Q => n_3686, QN => 
                           DataPath_RF_bus_reg_dataout_1756_port);
   DataPath_RF_BLOCKi_63_Q_reg_28_inst : DFF_X1 port map( D => n5433, CK => CLK
                           , Q => n_3687, QN => 
                           DataPath_RF_bus_reg_dataout_1788_port);
   DataPath_RF_BLOCKi_64_Q_reg_28_inst : DFF_X1 port map( D => n5468, CK => CLK
                           , Q => n_3688, QN => 
                           DataPath_RF_bus_reg_dataout_1820_port);
   DataPath_RF_BLOCKi_65_Q_reg_28_inst : DFF_X1 port map( D => n5503, CK => CLK
                           , Q => n_3689, QN => 
                           DataPath_RF_bus_reg_dataout_1852_port);
   DataPath_RF_BLOCKi_66_Q_reg_28_inst : DFF_X1 port map( D => n5538, CK => CLK
                           , Q => n_3690, QN => 
                           DataPath_RF_bus_reg_dataout_1884_port);
   DataPath_RF_BLOCKi_67_Q_reg_28_inst : DFF_X1 port map( D => n5573, CK => CLK
                           , Q => n_3691, QN => 
                           DataPath_RF_bus_reg_dataout_1916_port);
   DataPath_RF_BLOCKi_68_Q_reg_28_inst : DFF_X1 port map( D => n5612, CK => CLK
                           , Q => n_3692, QN => 
                           DataPath_RF_bus_reg_dataout_1948_port);
   DataPath_RF_BLOCKi_69_Q_reg_28_inst : DFF_X1 port map( D => n5649, CK => CLK
                           , Q => n_3693, QN => 
                           DataPath_RF_bus_reg_dataout_1980_port);
   DataPath_RF_BLOCKi_70_Q_reg_28_inst : DFF_X1 port map( D => n5686, CK => CLK
                           , Q => n_3694, QN => 
                           DataPath_RF_bus_reg_dataout_2012_port);
   DataPath_RF_BLOCKi_71_Q_reg_28_inst : DFF_X1 port map( D => n5723, CK => CLK
                           , Q => n_3695, QN => 
                           DataPath_RF_bus_reg_dataout_2044_port);
   DataPath_RF_BLOCKi_83_Q_reg_28_inst : DFF_X1 port map( D => n922, CK => CLK,
                           Q => n_3696, QN => 
                           DataPath_RF_bus_reg_dataout_2428_port);
   DataPath_RF_BLOCKi_84_Q_reg_28_inst : DFF_X1 port map( D => n973, CK => CLK,
                           Q => n_3697, QN => 
                           DataPath_RF_bus_reg_dataout_2460_port);
   DataPath_RF_BLOCKi_85_Q_reg_28_inst : DFF_X1 port map( D => n1010, CK => CLK
                           , Q => n_3698, QN => 
                           DataPath_RF_bus_reg_dataout_2492_port);
   DataPath_RF_BLOCKi_86_Q_reg_28_inst : DFF_X1 port map( D => n1047, CK => CLK
                           , Q => n_3699, QN => 
                           DataPath_RF_bus_reg_dataout_2524_port);
   DataPath_RF_BLOCKi_87_Q_reg_28_inst : DFF_X1 port map( D => n1084, CK => CLK
                           , Q => n_3700, QN => 
                           DataPath_RF_bus_reg_dataout_2556_port);
   DataPath_RF_BLOCKi_72_Q_reg_28_inst : DFF_X1 port map( D => n5760, CK => CLK
                           , Q => n_3701, QN => 
                           DataPath_RF_bus_reg_dataout_2076_port);
   DataPath_RF_BLOCKi_73_Q_reg_28_inst : DFF_X1 port map( D => n5799, CK => CLK
                           , Q => n_3702, QN => 
                           DataPath_RF_bus_reg_dataout_2108_port);
   DataPath_RF_BLOCKi_74_Q_reg_28_inst : DFF_X1 port map( D => n5835, CK => CLK
                           , Q => n_3703, QN => 
                           DataPath_RF_bus_reg_dataout_2140_port);
   DataPath_RF_BLOCKi_75_Q_reg_28_inst : DFF_X1 port map( D => n5871, CK => CLK
                           , Q => n_3704, QN => 
                           DataPath_RF_bus_reg_dataout_2172_port);
   DataPath_RF_BLOCKi_76_Q_reg_28_inst : DFF_X1 port map( D => n5907, CK => CLK
                           , Q => n_3705, QN => 
                           DataPath_RF_bus_reg_dataout_2204_port);
   DataPath_RF_BLOCKi_77_Q_reg_28_inst : DFF_X1 port map( D => n5943, CK => CLK
                           , Q => n_3706, QN => 
                           DataPath_RF_bus_reg_dataout_2236_port);
   DataPath_RF_BLOCKi_78_Q_reg_28_inst : DFF_X1 port map( D => n5979, CK => CLK
                           , Q => n_3707, QN => 
                           DataPath_RF_bus_reg_dataout_2268_port);
   DataPath_RF_BLOCKi_79_Q_reg_28_inst : DFF_X1 port map( D => n6015, CK => CLK
                           , Q => n_3708, QN => 
                           DataPath_RF_bus_reg_dataout_2300_port);
   DataPath_RF_BLOCKi_80_Q_reg_28_inst : DFF_X1 port map( D => n6052, CK => CLK
                           , Q => n_3709, QN => 
                           DataPath_RF_bus_reg_dataout_2332_port);
   DataPath_RF_BLOCKi_81_Q_reg_28_inst : DFF_X1 port map( D => n6088, CK => CLK
                           , Q => n_3710, QN => 
                           DataPath_RF_bus_reg_dataout_2364_port);
   DataPath_RF_BLOCKi_82_Q_reg_28_inst : DFF_X1 port map( D => n6122, CK => CLK
                           , Q => n_3711, QN => 
                           DataPath_RF_bus_reg_dataout_2396_port);
   DataPath_REG_ALU_OUT_Q_reg_30_inst : DFF_X1 port map( D => n6993, CK => CLK,
                           Q => DRAM_ADDRESS_30_port, QN => n514);
   DataPath_REG_MEM_ALUOUT_Q_reg_30_inst : DFF_X1 port map( D => n1119, CK => 
                           CLK, Q => n_3712, QN => 
                           DataPath_i_REG_MEM_ALUOUT_30_port);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_30_inst : DFF_X1 port map( D => n6769, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_62_port,
                           QN => n629);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_30_inst : DFF_X1 port map( D => n6801, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_94_port,
                           QN => n661);
   DataPath_RF_BLOCK_GLOB_3_Q_reg_30_inst : DFF_X1 port map( D => n6833, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_126_port
                           , QN => n693);
   DataPath_RF_BLOCK_GLOB_4_Q_reg_30_inst : DFF_X1 port map( D => n6865, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_158_port
                           , QN => n725);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_30_inst : DFF_X1 port map( D => n6897, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_190_port
                           , QN => n757);
   DataPath_RF_BLOCK_GLOB_6_Q_reg_30_inst : DFF_X1 port map( D => n6929, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_222_port
                           , QN => n789);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_30_inst : DFF_X1 port map( D => n6961, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_254_port
                           , QN => n821);
   DataPath_RF_BLOCKi_8_Q_reg_30_inst : DFF_X1 port map( D => n3312, CK => CLK,
                           Q => n_3713, QN => 
                           DataPath_RF_bus_reg_dataout_30_port);
   DataPath_RF_BLOCKi_9_Q_reg_30_inst : DFF_X1 port map( D => n3382, CK => CLK,
                           Q => n_3714, QN => 
                           DataPath_RF_bus_reg_dataout_62_port);
   DataPath_RF_BLOCKi_10_Q_reg_30_inst : DFF_X1 port map( D => n3420, CK => CLK
                           , Q => n_3715, QN => 
                           DataPath_RF_bus_reg_dataout_94_port);
   DataPath_RF_BLOCKi_11_Q_reg_30_inst : DFF_X1 port map( D => n3458, CK => CLK
                           , Q => n_3716, QN => 
                           DataPath_RF_bus_reg_dataout_126_port);
   DataPath_RF_BLOCKi_12_Q_reg_30_inst : DFF_X1 port map( D => n3496, CK => CLK
                           , Q => n_3717, QN => 
                           DataPath_RF_bus_reg_dataout_158_port);
   DataPath_RF_BLOCKi_13_Q_reg_30_inst : DFF_X1 port map( D => n3534, CK => CLK
                           , Q => n_3718, QN => 
                           DataPath_RF_bus_reg_dataout_190_port);
   DataPath_RF_BLOCKi_14_Q_reg_30_inst : DFF_X1 port map( D => n3572, CK => CLK
                           , Q => n_3719, QN => 
                           DataPath_RF_bus_reg_dataout_222_port);
   DataPath_RF_BLOCKi_15_Q_reg_30_inst : DFF_X1 port map( D => n3610, CK => CLK
                           , Q => n_3720, QN => 
                           DataPath_RF_bus_reg_dataout_254_port);
   DataPath_RF_BLOCKi_16_Q_reg_30_inst : DFF_X1 port map( D => n3648, CK => CLK
                           , Q => n_3721, QN => 
                           DataPath_RF_bus_reg_dataout_286_port);
   DataPath_RF_BLOCKi_17_Q_reg_30_inst : DFF_X1 port map( D => n3685, CK => CLK
                           , Q => n_3722, QN => 
                           DataPath_RF_bus_reg_dataout_318_port);
   DataPath_RF_BLOCKi_18_Q_reg_30_inst : DFF_X1 port map( D => n3722, CK => CLK
                           , Q => n_3723, QN => 
                           DataPath_RF_bus_reg_dataout_350_port);
   DataPath_RF_BLOCKi_19_Q_reg_30_inst : DFF_X1 port map( D => n3759, CK => CLK
                           , Q => n_3724, QN => 
                           DataPath_RF_bus_reg_dataout_382_port);
   DataPath_RF_BLOCKi_20_Q_reg_30_inst : DFF_X1 port map( D => n3794, CK => CLK
                           , Q => n_3725, QN => 
                           DataPath_RF_bus_reg_dataout_414_port);
   DataPath_RF_BLOCKi_21_Q_reg_30_inst : DFF_X1 port map( D => n3829, CK => CLK
                           , Q => n_3726, QN => 
                           DataPath_RF_bus_reg_dataout_446_port);
   DataPath_RF_BLOCKi_22_Q_reg_30_inst : DFF_X1 port map( D => n3864, CK => CLK
                           , Q => n_3727, QN => 
                           DataPath_RF_bus_reg_dataout_478_port);
   DataPath_RF_BLOCKi_23_Q_reg_30_inst : DFF_X1 port map( D => n3900, CK => CLK
                           , Q => n_3728, QN => 
                           DataPath_RF_bus_reg_dataout_510_port);
   DataPath_RF_BLOCKi_24_Q_reg_30_inst : DFF_X1 port map( D => n3968, CK => CLK
                           , Q => n_3729, QN => 
                           DataPath_RF_bus_reg_dataout_542_port);
   DataPath_RF_BLOCKi_25_Q_reg_30_inst : DFF_X1 port map( D => n4035, CK => CLK
                           , Q => n_3730, QN => 
                           DataPath_RF_bus_reg_dataout_574_port);
   DataPath_RF_BLOCKi_26_Q_reg_30_inst : DFF_X1 port map( D => n4070, CK => CLK
                           , Q => n_3731, QN => 
                           DataPath_RF_bus_reg_dataout_606_port);
   DataPath_RF_BLOCKi_27_Q_reg_30_inst : DFF_X1 port map( D => n4105, CK => CLK
                           , Q => n_3732, QN => 
                           DataPath_RF_bus_reg_dataout_638_port);
   DataPath_RF_BLOCKi_28_Q_reg_30_inst : DFF_X1 port map( D => n4140, CK => CLK
                           , Q => n_3733, QN => 
                           DataPath_RF_bus_reg_dataout_670_port);
   DataPath_RF_BLOCKi_29_Q_reg_30_inst : DFF_X1 port map( D => n4175, CK => CLK
                           , Q => n_3734, QN => 
                           DataPath_RF_bus_reg_dataout_702_port);
   DataPath_RF_BLOCKi_30_Q_reg_30_inst : DFF_X1 port map( D => n4210, CK => CLK
                           , Q => n_3735, QN => 
                           DataPath_RF_bus_reg_dataout_734_port);
   DataPath_RF_BLOCKi_31_Q_reg_30_inst : DFF_X1 port map( D => n4245, CK => CLK
                           , Q => n_3736, QN => 
                           DataPath_RF_bus_reg_dataout_766_port);
   DataPath_RF_BLOCKi_32_Q_reg_30_inst : DFF_X1 port map( D => n4280, CK => CLK
                           , Q => n_3737, QN => 
                           DataPath_RF_bus_reg_dataout_798_port);
   DataPath_RF_BLOCKi_33_Q_reg_30_inst : DFF_X1 port map( D => n4315, CK => CLK
                           , Q => n_3738, QN => 
                           DataPath_RF_bus_reg_dataout_830_port);
   DataPath_RF_BLOCKi_34_Q_reg_30_inst : DFF_X1 port map( D => n4350, CK => CLK
                           , Q => n_3739, QN => 
                           DataPath_RF_bus_reg_dataout_862_port);
   DataPath_RF_BLOCKi_35_Q_reg_30_inst : DFF_X1 port map( D => n4385, CK => CLK
                           , Q => n_3740, QN => 
                           DataPath_RF_bus_reg_dataout_894_port);
   DataPath_RF_BLOCKi_36_Q_reg_30_inst : DFF_X1 port map( D => n4420, CK => CLK
                           , Q => n_3741, QN => 
                           DataPath_RF_bus_reg_dataout_926_port);
   DataPath_RF_BLOCKi_37_Q_reg_30_inst : DFF_X1 port map( D => n4455, CK => CLK
                           , Q => n_3742, QN => 
                           DataPath_RF_bus_reg_dataout_958_port);
   DataPath_RF_BLOCKi_38_Q_reg_30_inst : DFF_X1 port map( D => n4490, CK => CLK
                           , Q => n_3743, QN => 
                           DataPath_RF_bus_reg_dataout_990_port);
   DataPath_RF_BLOCKi_39_Q_reg_30_inst : DFF_X1 port map( D => n4525, CK => CLK
                           , Q => n_3744, QN => 
                           DataPath_RF_bus_reg_dataout_1022_port);
   DataPath_RF_BLOCKi_40_Q_reg_30_inst : DFF_X1 port map( D => n4561, CK => CLK
                           , Q => n_3745, QN => 
                           DataPath_RF_bus_reg_dataout_1054_port);
   DataPath_RF_BLOCKi_41_Q_reg_30_inst : DFF_X1 port map( D => n4628, CK => CLK
                           , Q => n_3746, QN => 
                           DataPath_RF_bus_reg_dataout_1086_port);
   DataPath_RF_BLOCKi_42_Q_reg_30_inst : DFF_X1 port map( D => n4663, CK => CLK
                           , Q => n_3747, QN => 
                           DataPath_RF_bus_reg_dataout_1118_port);
   DataPath_RF_BLOCKi_43_Q_reg_30_inst : DFF_X1 port map( D => n4698, CK => CLK
                           , Q => n_3748, QN => 
                           DataPath_RF_bus_reg_dataout_1150_port);
   DataPath_RF_BLOCKi_44_Q_reg_30_inst : DFF_X1 port map( D => n4733, CK => CLK
                           , Q => n_3749, QN => 
                           DataPath_RF_bus_reg_dataout_1182_port);
   DataPath_RF_BLOCKi_45_Q_reg_30_inst : DFF_X1 port map( D => n4768, CK => CLK
                           , Q => n_3750, QN => 
                           DataPath_RF_bus_reg_dataout_1214_port);
   DataPath_RF_BLOCKi_46_Q_reg_30_inst : DFF_X1 port map( D => n4803, CK => CLK
                           , Q => n_3751, QN => 
                           DataPath_RF_bus_reg_dataout_1246_port);
   DataPath_RF_BLOCKi_47_Q_reg_30_inst : DFF_X1 port map( D => n4838, CK => CLK
                           , Q => n_3752, QN => 
                           DataPath_RF_bus_reg_dataout_1278_port);
   DataPath_RF_BLOCKi_48_Q_reg_30_inst : DFF_X1 port map( D => n4873, CK => CLK
                           , Q => n_3753, QN => 
                           DataPath_RF_bus_reg_dataout_1310_port);
   DataPath_RF_BLOCKi_49_Q_reg_30_inst : DFF_X1 port map( D => n4908, CK => CLK
                           , Q => n_3754, QN => 
                           DataPath_RF_bus_reg_dataout_1342_port);
   DataPath_RF_BLOCKi_50_Q_reg_30_inst : DFF_X1 port map( D => n4943, CK => CLK
                           , Q => n_3755, QN => 
                           DataPath_RF_bus_reg_dataout_1374_port);
   DataPath_RF_BLOCKi_51_Q_reg_30_inst : DFF_X1 port map( D => n4978, CK => CLK
                           , Q => n_3756, QN => 
                           DataPath_RF_bus_reg_dataout_1406_port);
   DataPath_RF_BLOCKi_52_Q_reg_30_inst : DFF_X1 port map( D => n5013, CK => CLK
                           , Q => n_3757, QN => 
                           DataPath_RF_bus_reg_dataout_1438_port);
   DataPath_RF_BLOCKi_53_Q_reg_30_inst : DFF_X1 port map( D => n5048, CK => CLK
                           , Q => n_3758, QN => 
                           DataPath_RF_bus_reg_dataout_1470_port);
   DataPath_RF_BLOCKi_54_Q_reg_30_inst : DFF_X1 port map( D => n5083, CK => CLK
                           , Q => n_3759, QN => 
                           DataPath_RF_bus_reg_dataout_1502_port);
   DataPath_RF_BLOCKi_55_Q_reg_30_inst : DFF_X1 port map( D => n5118, CK => CLK
                           , Q => n_3760, QN => 
                           DataPath_RF_bus_reg_dataout_1534_port);
   DataPath_RF_BLOCKi_56_Q_reg_30_inst : DFF_X1 port map( D => n5154, CK => CLK
                           , Q => n_3761, QN => 
                           DataPath_RF_bus_reg_dataout_1566_port);
   DataPath_RF_BLOCKi_57_Q_reg_30_inst : DFF_X1 port map( D => n5220, CK => CLK
                           , Q => n_3762, QN => 
                           DataPath_RF_bus_reg_dataout_1598_port);
   DataPath_RF_BLOCKi_58_Q_reg_30_inst : DFF_X1 port map( D => n5256, CK => CLK
                           , Q => n_3763, QN => 
                           DataPath_RF_bus_reg_dataout_1630_port);
   DataPath_RF_BLOCKi_59_Q_reg_30_inst : DFF_X1 port map( D => n5291, CK => CLK
                           , Q => n_3764, QN => 
                           DataPath_RF_bus_reg_dataout_1662_port);
   DataPath_RF_BLOCKi_60_Q_reg_30_inst : DFF_X1 port map( D => n5326, CK => CLK
                           , Q => n_3765, QN => 
                           DataPath_RF_bus_reg_dataout_1694_port);
   DataPath_RF_BLOCKi_61_Q_reg_30_inst : DFF_X1 port map( D => n5361, CK => CLK
                           , Q => n_3766, QN => 
                           DataPath_RF_bus_reg_dataout_1726_port);
   DataPath_RF_BLOCKi_62_Q_reg_30_inst : DFF_X1 port map( D => n5396, CK => CLK
                           , Q => n_3767, QN => 
                           DataPath_RF_bus_reg_dataout_1758_port);
   DataPath_RF_BLOCKi_63_Q_reg_30_inst : DFF_X1 port map( D => n5431, CK => CLK
                           , Q => n_3768, QN => 
                           DataPath_RF_bus_reg_dataout_1790_port);
   DataPath_RF_BLOCKi_64_Q_reg_30_inst : DFF_X1 port map( D => n5466, CK => CLK
                           , Q => n_3769, QN => 
                           DataPath_RF_bus_reg_dataout_1822_port);
   DataPath_RF_BLOCKi_65_Q_reg_30_inst : DFF_X1 port map( D => n5501, CK => CLK
                           , Q => n_3770, QN => 
                           DataPath_RF_bus_reg_dataout_1854_port);
   DataPath_RF_BLOCKi_66_Q_reg_30_inst : DFF_X1 port map( D => n5536, CK => CLK
                           , Q => n_3771, QN => 
                           DataPath_RF_bus_reg_dataout_1886_port);
   DataPath_RF_BLOCKi_67_Q_reg_30_inst : DFF_X1 port map( D => n5571, CK => CLK
                           , Q => n_3772, QN => 
                           DataPath_RF_bus_reg_dataout_1918_port);
   DataPath_RF_BLOCKi_68_Q_reg_30_inst : DFF_X1 port map( D => n5610, CK => CLK
                           , Q => n_3773, QN => 
                           DataPath_RF_bus_reg_dataout_1950_port);
   DataPath_RF_BLOCKi_69_Q_reg_30_inst : DFF_X1 port map( D => n5647, CK => CLK
                           , Q => n_3774, QN => 
                           DataPath_RF_bus_reg_dataout_1982_port);
   DataPath_RF_BLOCKi_70_Q_reg_30_inst : DFF_X1 port map( D => n5684, CK => CLK
                           , Q => n_3775, QN => 
                           DataPath_RF_bus_reg_dataout_2014_port);
   DataPath_RF_BLOCKi_71_Q_reg_30_inst : DFF_X1 port map( D => n5721, CK => CLK
                           , Q => n_3776, QN => 
                           DataPath_RF_bus_reg_dataout_2046_port);
   DataPath_RF_BLOCKi_83_Q_reg_30_inst : DFF_X1 port map( D => n918, CK => CLK,
                           Q => n_3777, QN => 
                           DataPath_RF_bus_reg_dataout_2430_port);
   DataPath_RF_BLOCKi_84_Q_reg_30_inst : DFF_X1 port map( D => n971, CK => CLK,
                           Q => n_3778, QN => 
                           DataPath_RF_bus_reg_dataout_2462_port);
   DataPath_RF_BLOCKi_85_Q_reg_30_inst : DFF_X1 port map( D => n1008, CK => CLK
                           , Q => n_3779, QN => 
                           DataPath_RF_bus_reg_dataout_2494_port);
   DataPath_RF_BLOCKi_86_Q_reg_30_inst : DFF_X1 port map( D => n1045, CK => CLK
                           , Q => n_3780, QN => 
                           DataPath_RF_bus_reg_dataout_2526_port);
   DataPath_RF_BLOCKi_87_Q_reg_30_inst : DFF_X1 port map( D => n1082, CK => CLK
                           , Q => n_3781, QN => 
                           DataPath_RF_bus_reg_dataout_2558_port);
   DataPath_RF_BLOCKi_72_Q_reg_30_inst : DFF_X1 port map( D => n5758, CK => CLK
                           , Q => n_3782, QN => 
                           DataPath_RF_bus_reg_dataout_2078_port);
   DataPath_RF_BLOCKi_73_Q_reg_30_inst : DFF_X1 port map( D => n5797, CK => CLK
                           , Q => n_3783, QN => 
                           DataPath_RF_bus_reg_dataout_2110_port);
   DataPath_RF_BLOCKi_74_Q_reg_30_inst : DFF_X1 port map( D => n5833, CK => CLK
                           , Q => n_3784, QN => 
                           DataPath_RF_bus_reg_dataout_2142_port);
   DataPath_RF_BLOCKi_75_Q_reg_30_inst : DFF_X1 port map( D => n5869, CK => CLK
                           , Q => n_3785, QN => 
                           DataPath_RF_bus_reg_dataout_2174_port);
   DataPath_RF_BLOCKi_76_Q_reg_30_inst : DFF_X1 port map( D => n5905, CK => CLK
                           , Q => n_3786, QN => 
                           DataPath_RF_bus_reg_dataout_2206_port);
   DataPath_RF_BLOCKi_77_Q_reg_30_inst : DFF_X1 port map( D => n5941, CK => CLK
                           , Q => n_3787, QN => 
                           DataPath_RF_bus_reg_dataout_2238_port);
   DataPath_RF_BLOCKi_78_Q_reg_30_inst : DFF_X1 port map( D => n5977, CK => CLK
                           , Q => n_3788, QN => 
                           DataPath_RF_bus_reg_dataout_2270_port);
   DataPath_RF_BLOCKi_79_Q_reg_30_inst : DFF_X1 port map( D => n6013, CK => CLK
                           , Q => n_3789, QN => 
                           DataPath_RF_bus_reg_dataout_2302_port);
   DataPath_RF_BLOCKi_80_Q_reg_30_inst : DFF_X1 port map( D => n6050, CK => CLK
                           , Q => n_3790, QN => 
                           DataPath_RF_bus_reg_dataout_2334_port);
   DataPath_RF_BLOCKi_81_Q_reg_30_inst : DFF_X1 port map( D => n6086, CK => CLK
                           , Q => n_3791, QN => 
                           DataPath_RF_bus_reg_dataout_2366_port);
   DataPath_RF_BLOCKi_82_Q_reg_30_inst : DFF_X1 port map( D => n6120, CK => CLK
                           , Q => n_3792, QN => 
                           DataPath_RF_bus_reg_dataout_2398_port);
   DataPath_RF_BLOCKi_8_Q_reg_7_inst : DFF_X1 port map( D => n3358, CK => CLK, 
                           Q => n_3793, QN => 
                           DataPath_RF_bus_reg_dataout_7_port);
   DataPath_RF_BLOCKi_9_Q_reg_7_inst : DFF_X1 port map( D => n3405, CK => CLK, 
                           Q => n_3794, QN => 
                           DataPath_RF_bus_reg_dataout_39_port);
   DataPath_RF_BLOCKi_10_Q_reg_7_inst : DFF_X1 port map( D => n3443, CK => CLK,
                           Q => n_3795, QN => 
                           DataPath_RF_bus_reg_dataout_71_port);
   DataPath_RF_BLOCKi_11_Q_reg_7_inst : DFF_X1 port map( D => n3481, CK => CLK,
                           Q => n_3796, QN => 
                           DataPath_RF_bus_reg_dataout_103_port);
   DataPath_RF_BLOCKi_12_Q_reg_7_inst : DFF_X1 port map( D => n3519, CK => CLK,
                           Q => n_3797, QN => 
                           DataPath_RF_bus_reg_dataout_135_port);
   DataPath_RF_BLOCKi_13_Q_reg_7_inst : DFF_X1 port map( D => n3557, CK => CLK,
                           Q => n_3798, QN => 
                           DataPath_RF_bus_reg_dataout_167_port);
   DataPath_RF_BLOCKi_14_Q_reg_7_inst : DFF_X1 port map( D => n3595, CK => CLK,
                           Q => n_3799, QN => 
                           DataPath_RF_bus_reg_dataout_199_port);
   DataPath_RF_BLOCKi_15_Q_reg_7_inst : DFF_X1 port map( D => n3633, CK => CLK,
                           Q => n_3800, QN => 
                           DataPath_RF_bus_reg_dataout_231_port);
   DataPath_RF_BLOCKi_16_Q_reg_7_inst : DFF_X1 port map( D => n3671, CK => CLK,
                           Q => n_3801, QN => 
                           DataPath_RF_bus_reg_dataout_263_port);
   DataPath_RF_BLOCKi_17_Q_reg_7_inst : DFF_X1 port map( D => n3708, CK => CLK,
                           Q => n_3802, QN => 
                           DataPath_RF_bus_reg_dataout_295_port);
   DataPath_RF_BLOCKi_18_Q_reg_7_inst : DFF_X1 port map( D => n3745, CK => CLK,
                           Q => n_3803, QN => 
                           DataPath_RF_bus_reg_dataout_327_port);
   DataPath_RF_BLOCKi_19_Q_reg_7_inst : DFF_X1 port map( D => n3782, CK => CLK,
                           Q => n_3804, QN => 
                           DataPath_RF_bus_reg_dataout_359_port);
   DataPath_RF_BLOCKi_20_Q_reg_7_inst : DFF_X1 port map( D => n3817, CK => CLK,
                           Q => n_3805, QN => 
                           DataPath_RF_bus_reg_dataout_391_port);
   DataPath_RF_BLOCKi_21_Q_reg_7_inst : DFF_X1 port map( D => n3852, CK => CLK,
                           Q => n_3806, QN => 
                           DataPath_RF_bus_reg_dataout_423_port);
   DataPath_RF_BLOCKi_22_Q_reg_7_inst : DFF_X1 port map( D => n3887, CK => CLK,
                           Q => n_3807, QN => 
                           DataPath_RF_bus_reg_dataout_455_port);
   DataPath_RF_BLOCKi_23_Q_reg_7_inst : DFF_X1 port map( D => n3946, CK => CLK,
                           Q => n_3808, QN => 
                           DataPath_RF_bus_reg_dataout_487_port);
   DataPath_RF_BLOCKi_24_Q_reg_7_inst : DFF_X1 port map( D => n4014, CK => CLK,
                           Q => n_3809, QN => 
                           DataPath_RF_bus_reg_dataout_519_port);
   DataPath_RF_BLOCKi_25_Q_reg_7_inst : DFF_X1 port map( D => n4058, CK => CLK,
                           Q => n_3810, QN => 
                           DataPath_RF_bus_reg_dataout_551_port);
   DataPath_RF_BLOCKi_26_Q_reg_7_inst : DFF_X1 port map( D => n4093, CK => CLK,
                           Q => n_3811, QN => 
                           DataPath_RF_bus_reg_dataout_583_port);
   DataPath_RF_BLOCKi_27_Q_reg_7_inst : DFF_X1 port map( D => n4128, CK => CLK,
                           Q => n_3812, QN => 
                           DataPath_RF_bus_reg_dataout_615_port);
   DataPath_RF_BLOCKi_28_Q_reg_7_inst : DFF_X1 port map( D => n4163, CK => CLK,
                           Q => n_3813, QN => 
                           DataPath_RF_bus_reg_dataout_647_port);
   DataPath_RF_BLOCKi_29_Q_reg_7_inst : DFF_X1 port map( D => n4198, CK => CLK,
                           Q => n_3814, QN => 
                           DataPath_RF_bus_reg_dataout_679_port);
   DataPath_RF_BLOCKi_30_Q_reg_7_inst : DFF_X1 port map( D => n4233, CK => CLK,
                           Q => n_3815, QN => 
                           DataPath_RF_bus_reg_dataout_711_port);
   DataPath_RF_BLOCKi_31_Q_reg_7_inst : DFF_X1 port map( D => n4268, CK => CLK,
                           Q => n_3816, QN => 
                           DataPath_RF_bus_reg_dataout_743_port);
   DataPath_RF_BLOCKi_32_Q_reg_7_inst : DFF_X1 port map( D => n4303, CK => CLK,
                           Q => n_3817, QN => 
                           DataPath_RF_bus_reg_dataout_775_port);
   DataPath_RF_BLOCKi_33_Q_reg_7_inst : DFF_X1 port map( D => n4338, CK => CLK,
                           Q => n_3818, QN => 
                           DataPath_RF_bus_reg_dataout_807_port);
   DataPath_RF_BLOCKi_34_Q_reg_7_inst : DFF_X1 port map( D => n4373, CK => CLK,
                           Q => n_3819, QN => 
                           DataPath_RF_bus_reg_dataout_839_port);
   DataPath_RF_BLOCKi_35_Q_reg_7_inst : DFF_X1 port map( D => n4408, CK => CLK,
                           Q => n_3820, QN => 
                           DataPath_RF_bus_reg_dataout_871_port);
   DataPath_RF_BLOCKi_36_Q_reg_7_inst : DFF_X1 port map( D => n4443, CK => CLK,
                           Q => n_3821, QN => 
                           DataPath_RF_bus_reg_dataout_903_port);
   DataPath_RF_BLOCKi_37_Q_reg_7_inst : DFF_X1 port map( D => n4478, CK => CLK,
                           Q => n_3822, QN => 
                           DataPath_RF_bus_reg_dataout_935_port);
   DataPath_RF_BLOCKi_38_Q_reg_7_inst : DFF_X1 port map( D => n4513, CK => CLK,
                           Q => n_3823, QN => 
                           DataPath_RF_bus_reg_dataout_967_port);
   DataPath_RF_BLOCKi_39_Q_reg_7_inst : DFF_X1 port map( D => n4548, CK => CLK,
                           Q => n_3824, QN => 
                           DataPath_RF_bus_reg_dataout_999_port);
   DataPath_RF_BLOCKi_40_Q_reg_7_inst : DFF_X1 port map( D => n4607, CK => CLK,
                           Q => n_3825, QN => 
                           DataPath_RF_bus_reg_dataout_1031_port);
   DataPath_RF_BLOCKi_41_Q_reg_7_inst : DFF_X1 port map( D => n4651, CK => CLK,
                           Q => n_3826, QN => 
                           DataPath_RF_bus_reg_dataout_1063_port);
   DataPath_RF_BLOCKi_42_Q_reg_7_inst : DFF_X1 port map( D => n4686, CK => CLK,
                           Q => n_3827, QN => 
                           DataPath_RF_bus_reg_dataout_1095_port);
   DataPath_RF_BLOCKi_43_Q_reg_7_inst : DFF_X1 port map( D => n4721, CK => CLK,
                           Q => n_3828, QN => 
                           DataPath_RF_bus_reg_dataout_1127_port);
   DataPath_RF_BLOCKi_44_Q_reg_7_inst : DFF_X1 port map( D => n4756, CK => CLK,
                           Q => n_3829, QN => 
                           DataPath_RF_bus_reg_dataout_1159_port);
   DataPath_RF_BLOCKi_45_Q_reg_7_inst : DFF_X1 port map( D => n4791, CK => CLK,
                           Q => n_3830, QN => 
                           DataPath_RF_bus_reg_dataout_1191_port);
   DataPath_RF_BLOCKi_46_Q_reg_7_inst : DFF_X1 port map( D => n4826, CK => CLK,
                           Q => n_3831, QN => 
                           DataPath_RF_bus_reg_dataout_1223_port);
   DataPath_RF_BLOCKi_47_Q_reg_7_inst : DFF_X1 port map( D => n4861, CK => CLK,
                           Q => n_3832, QN => 
                           DataPath_RF_bus_reg_dataout_1255_port);
   DataPath_RF_BLOCKi_48_Q_reg_7_inst : DFF_X1 port map( D => n4896, CK => CLK,
                           Q => n_3833, QN => 
                           DataPath_RF_bus_reg_dataout_1287_port);
   DataPath_RF_BLOCKi_49_Q_reg_7_inst : DFF_X1 port map( D => n4931, CK => CLK,
                           Q => n_3834, QN => 
                           DataPath_RF_bus_reg_dataout_1319_port);
   DataPath_RF_BLOCKi_50_Q_reg_7_inst : DFF_X1 port map( D => n4966, CK => CLK,
                           Q => n_3835, QN => 
                           DataPath_RF_bus_reg_dataout_1351_port);
   DataPath_RF_BLOCKi_51_Q_reg_7_inst : DFF_X1 port map( D => n5001, CK => CLK,
                           Q => n_3836, QN => 
                           DataPath_RF_bus_reg_dataout_1383_port);
   DataPath_RF_BLOCKi_52_Q_reg_7_inst : DFF_X1 port map( D => n5036, CK => CLK,
                           Q => n_3837, QN => 
                           DataPath_RF_bus_reg_dataout_1415_port);
   DataPath_RF_BLOCKi_53_Q_reg_7_inst : DFF_X1 port map( D => n5071, CK => CLK,
                           Q => n_3838, QN => 
                           DataPath_RF_bus_reg_dataout_1447_port);
   DataPath_RF_BLOCKi_54_Q_reg_7_inst : DFF_X1 port map( D => n5106, CK => CLK,
                           Q => n_3839, QN => 
                           DataPath_RF_bus_reg_dataout_1479_port);
   DataPath_RF_BLOCKi_55_Q_reg_7_inst : DFF_X1 port map( D => n5141, CK => CLK,
                           Q => n_3840, QN => 
                           DataPath_RF_bus_reg_dataout_1511_port);
   DataPath_RF_BLOCKi_56_Q_reg_7_inst : DFF_X1 port map( D => n5200, CK => CLK,
                           Q => n_3841, QN => 
                           DataPath_RF_bus_reg_dataout_1543_port);
   DataPath_RF_BLOCKi_57_Q_reg_7_inst : DFF_X1 port map( D => n5243, CK => CLK,
                           Q => n_3842, QN => 
                           DataPath_RF_bus_reg_dataout_1575_port);
   DataPath_RF_BLOCKi_58_Q_reg_7_inst : DFF_X1 port map( D => n5279, CK => CLK,
                           Q => n_3843, QN => 
                           DataPath_RF_bus_reg_dataout_1607_port);
   DataPath_RF_BLOCKi_59_Q_reg_7_inst : DFF_X1 port map( D => n5314, CK => CLK,
                           Q => n_3844, QN => 
                           DataPath_RF_bus_reg_dataout_1639_port);
   DataPath_RF_BLOCKi_60_Q_reg_7_inst : DFF_X1 port map( D => n5349, CK => CLK,
                           Q => n_3845, QN => 
                           DataPath_RF_bus_reg_dataout_1671_port);
   DataPath_RF_BLOCKi_61_Q_reg_7_inst : DFF_X1 port map( D => n5384, CK => CLK,
                           Q => n_3846, QN => 
                           DataPath_RF_bus_reg_dataout_1703_port);
   DataPath_RF_BLOCKi_62_Q_reg_7_inst : DFF_X1 port map( D => n5419, CK => CLK,
                           Q => n_3847, QN => 
                           DataPath_RF_bus_reg_dataout_1735_port);
   DataPath_RF_BLOCKi_63_Q_reg_7_inst : DFF_X1 port map( D => n5454, CK => CLK,
                           Q => n_3848, QN => 
                           DataPath_RF_bus_reg_dataout_1767_port);
   DataPath_RF_BLOCKi_64_Q_reg_7_inst : DFF_X1 port map( D => n5489, CK => CLK,
                           Q => n_3849, QN => 
                           DataPath_RF_bus_reg_dataout_1799_port);
   DataPath_RF_BLOCKi_65_Q_reg_7_inst : DFF_X1 port map( D => n5524, CK => CLK,
                           Q => n_3850, QN => 
                           DataPath_RF_bus_reg_dataout_1831_port);
   DataPath_RF_BLOCKi_66_Q_reg_7_inst : DFF_X1 port map( D => n5559, CK => CLK,
                           Q => n_3851, QN => 
                           DataPath_RF_bus_reg_dataout_1863_port);
   DataPath_RF_BLOCKi_67_Q_reg_7_inst : DFF_X1 port map( D => n5594, CK => CLK,
                           Q => n_3852, QN => 
                           DataPath_RF_bus_reg_dataout_1895_port);
   DataPath_RF_BLOCKi_68_Q_reg_7_inst : DFF_X1 port map( D => n5633, CK => CLK,
                           Q => n_3853, QN => 
                           DataPath_RF_bus_reg_dataout_1927_port);
   DataPath_RF_BLOCKi_69_Q_reg_7_inst : DFF_X1 port map( D => n5670, CK => CLK,
                           Q => n_3854, QN => 
                           DataPath_RF_bus_reg_dataout_1959_port);
   DataPath_RF_BLOCKi_70_Q_reg_7_inst : DFF_X1 port map( D => n5707, CK => CLK,
                           Q => n_3855, QN => 
                           DataPath_RF_bus_reg_dataout_1991_port);
   DataPath_RF_BLOCKi_71_Q_reg_7_inst : DFF_X1 port map( D => n5744, CK => CLK,
                           Q => n_3856, QN => 
                           DataPath_RF_bus_reg_dataout_2023_port);
   DataPath_RF_BLOCKi_82_Q_reg_7_inst : DFF_X1 port map( D => n898, CK => CLK, 
                           Q => n_3857, QN => 
                           DataPath_RF_bus_reg_dataout_2375_port);
   DataPath_RF_BLOCKi_83_Q_reg_7_inst : DFF_X1 port map( D => n956, CK => CLK, 
                           Q => n_3858, QN => 
                           DataPath_RF_bus_reg_dataout_2407_port);
   DataPath_RF_BLOCKi_84_Q_reg_7_inst : DFF_X1 port map( D => n994, CK => CLK, 
                           Q => n_3859, QN => 
                           DataPath_RF_bus_reg_dataout_2439_port);
   DataPath_RF_BLOCKi_85_Q_reg_7_inst : DFF_X1 port map( D => n1031, CK => CLK,
                           Q => n_3860, QN => 
                           DataPath_RF_bus_reg_dataout_2471_port);
   DataPath_RF_BLOCKi_86_Q_reg_7_inst : DFF_X1 port map( D => n1068, CK => CLK,
                           Q => n_3861, QN => 
                           DataPath_RF_bus_reg_dataout_2503_port);
   DataPath_RF_BLOCKi_87_Q_reg_7_inst : DFF_X1 port map( D => n1105, CK => CLK,
                           Q => n_3862, QN => 
                           DataPath_RF_bus_reg_dataout_2535_port);
   DataPath_RF_BLOCKi_72_Q_reg_7_inst : DFF_X1 port map( D => n5781, CK => CLK,
                           Q => n_3863, QN => 
                           DataPath_RF_bus_reg_dataout_2055_port);
   DataPath_RF_BLOCKi_73_Q_reg_7_inst : DFF_X1 port map( D => n5820, CK => CLK,
                           Q => n_3864, QN => 
                           DataPath_RF_bus_reg_dataout_2087_port);
   DataPath_RF_BLOCKi_74_Q_reg_7_inst : DFF_X1 port map( D => n5856, CK => CLK,
                           Q => n_3865, QN => 
                           DataPath_RF_bus_reg_dataout_2119_port);
   DataPath_RF_BLOCKi_75_Q_reg_7_inst : DFF_X1 port map( D => n5892, CK => CLK,
                           Q => n_3866, QN => 
                           DataPath_RF_bus_reg_dataout_2151_port);
   DataPath_RF_BLOCKi_76_Q_reg_7_inst : DFF_X1 port map( D => n5928, CK => CLK,
                           Q => n_3867, QN => 
                           DataPath_RF_bus_reg_dataout_2183_port);
   DataPath_RF_BLOCKi_77_Q_reg_7_inst : DFF_X1 port map( D => n5964, CK => CLK,
                           Q => n_3868, QN => 
                           DataPath_RF_bus_reg_dataout_2215_port);
   DataPath_RF_BLOCKi_78_Q_reg_7_inst : DFF_X1 port map( D => n6000, CK => CLK,
                           Q => n_3869, QN => 
                           DataPath_RF_bus_reg_dataout_2247_port);
   DataPath_RF_BLOCKi_79_Q_reg_7_inst : DFF_X1 port map( D => n6036, CK => CLK,
                           Q => n_3870, QN => 
                           DataPath_RF_bus_reg_dataout_2279_port);
   DataPath_RF_BLOCKi_80_Q_reg_7_inst : DFF_X1 port map( D => n6073, CK => CLK,
                           Q => n_3871, QN => 
                           DataPath_RF_bus_reg_dataout_2311_port);
   DataPath_RF_BLOCKi_81_Q_reg_7_inst : DFF_X1 port map( D => n6109, CK => CLK,
                           Q => n_3872, QN => 
                           DataPath_RF_bus_reg_dataout_2343_port);
   DataPath_RF_CWP_Q_reg_0_inst : DFF_X2 port map( D => n7074, CK => CLK, Q => 
                           DataPath_RF_c_win_0_port, QN => n8191);
   DataPath_RF_CWP_Q_reg_1_inst : DFF_X2 port map( D => n7073, CK => CLK, Q => 
                           DataPath_RF_c_win_1_port, QN => n8333);
   CU_I_CW_MEM_reg_DRAM_RE_inst : DFF_X2 port map( D => n7096, CK => CLK, Q => 
                           i_DATAMEM_RM, QN => n8293);
   IR_reg_30_inst : DFFS_X1 port map( D => n7119, CK => CLK, SN => n8574, Q => 
                           n8237, QN => n161);
   IR_reg_31_inst : DFFS_X1 port map( D => n8391, CK => CLK, SN => n8575, Q => 
                           n159, QN => n8586);
   DataPath_WRF_CUhw_curr_state_reg_1_inst : DFF_X1 port map( D => 
                           DataPath_WRF_CUhw_N145, CK => CLK, Q => n8230, QN =>
                           n466);
   CU_I_aluOpcode1_reg_2_inst : DFF_X2 port map( D => n7093, CK => CLK, Q => 
                           i_ALU_OP_2_port, QN => n8188);
   DataPath_WRF_CUhw_curr_addr_reg_29_inst : DFF_X1 port map( D => n8395, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_29_port, QN =>
                           n_3873);
   DataPath_WRF_CUhw_curr_addr_reg_30_inst : DFF_X1 port map( D => n8394, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_30_port, QN =>
                           n_3874);
   PC_reg_28_inst : DFFS_X1 port map( D => n8392, CK => CLK, SN => n8581, Q => 
                           n10281, QN => IRAM_ADDRESS_28_port);
   PC_reg_29_inst : DFFS_X1 port map( D => n7190, CK => CLK, SN => n8575, Q => 
                           n10275, QN => IRAM_ADDRESS_29_port);
   IR_reg_22_inst : DFFR_X1 port map( D => n7126, CK => CLK, RN => n8581, Q => 
                           n8302, QN => n171);
   PC_reg_10_inst : DFFR_X1 port map( D => n7051, CK => CLK, RN => n8577, Q => 
                           IRAM_ADDRESS_10_port, QN => n8314);
   PC_reg_23_inst : DFFR_X1 port map( D => n7038, CK => CLK, RN => n8572, Q => 
                           IRAM_ADDRESS_23_port, QN => n8289);
   PC_reg_4_inst : DFFR_X1 port map( D => n7057, CK => CLK, RN => n8579, Q => 
                           IRAM_ADDRESS_4_port, QN => n8313);
   PC_reg_11_inst : DFFR_X1 port map( D => n7050, CK => CLK, RN => n8571, Q => 
                           IRAM_ADDRESS_11_port, QN => n8312);
   intadd_0_U6 : NOR2_X1 port map( A1 => intadd_0_B_3_port, A2 => 
                           IRAM_ADDRESS_4_port, ZN => intadd_0_n6);
   intadd_0_U7 : NAND2_X1 port map( A1 => intadd_0_B_3_port, A2 => 
                           IRAM_ADDRESS_4_port, ZN => intadd_0_n7);
   intadd_1_U28 : NOR2_X1 port map( A1 => intadd_1_B_0_port, A2 => 
                           IRAM_ADDRESS_10_port, ZN => intadd_1_n21);
   intadd_1_U20 : NOR2_X1 port map( A1 => intadd_1_B_1_port, A2 => 
                           IRAM_ADDRESS_11_port, ZN => intadd_1_n16);
   intadd_1_U16 : NOR2_X1 port map( A1 => intadd_1_n21, A2 => intadd_1_n16, ZN 
                           => intadd_1_n14);
   intadd_1_U29 : NAND2_X1 port map( A1 => intadd_1_B_0_port, A2 => 
                           IRAM_ADDRESS_10_port, ZN => intadd_1_n22);
   intadd_1_U21 : NAND2_X1 port map( A1 => intadd_1_B_1_port, A2 => 
                           IRAM_ADDRESS_11_port, ZN => intadd_1_n17);
   intadd_1_U17 : OAI21_X1 port map( B1 => intadd_1_n16, B2 => intadd_1_n22, A 
                           => intadd_1_n17, ZN => intadd_1_n15);
   intadd_1_U13 : NAND2_X1 port map( A1 => intadd_1_B_2_port, A2 => 
                           IRAM_ADDRESS_12_port, ZN => intadd_1_n12);
   intadd_1_U10 : NAND2_X1 port map( A1 => n8222, A2 => intadd_1_n12, ZN => 
                           intadd_1_n1);
   intadd_1_U18 : NAND2_X1 port map( A1 => intadd_1_n26, A2 => intadd_1_n17, ZN
                           => intadd_1_n2);
   intadd_1_U26 : NAND2_X1 port map( A1 => intadd_1_n27, A2 => intadd_1_n22, ZN
                           => intadd_1_n3);
   intadd_0_U18 : NAND2_X1 port map( A1 => intadd_0_n23, A2 => intadd_0_n15, ZN
                           => intadd_0_n3);
   intadd_0_U16 : XOR2_X1 port map( A => intadd_0_n16, B => intadd_0_n3, Z => 
                           intadd_0_SUM_1_port);
   intadd_0_U12 : NAND2_X1 port map( A1 => intadd_0_n22, A2 => intadd_0_n12, ZN
                           => intadd_0_n2);
   intadd_0_U4 : NAND2_X1 port map( A1 => intadd_0_n21, A2 => intadd_0_n7, ZN 
                           => intadd_0_n1);
   DP_OP_1091J1_126_6973_U29 : FA_X1 port map( A => DP_OP_1091J1_126_6973_n31, 
                           B => DataPath_WRF_CUhw_curr_addr_4_port, CI => 
                           DP_OP_1091J1_126_6973_n29, CO => 
                           DP_OP_1091J1_126_6973_n28, S => C620_DATA2_4);
   DP_OP_1091J1_126_6973_U28 : FA_X1 port map( A => DP_OP_1091J1_126_6973_n31, 
                           B => DataPath_WRF_CUhw_curr_addr_5_port, CI => 
                           DP_OP_1091J1_126_6973_n28, CO => 
                           DP_OP_1091J1_126_6973_n27, S => C620_DATA2_5);
   DP_OP_1091J1_126_6973_U27 : FA_X1 port map( A => DP_OP_1091J1_126_6973_n31, 
                           B => DataPath_WRF_CUhw_curr_addr_6_port, CI => 
                           DP_OP_1091J1_126_6973_n27, CO => 
                           DP_OP_1091J1_126_6973_n26, S => C620_DATA2_6);
   DP_OP_1091J1_126_6973_U26 : FA_X1 port map( A => DP_OP_1091J1_126_6973_n31, 
                           B => DataPath_WRF_CUhw_curr_addr_7_port, CI => 
                           DP_OP_1091J1_126_6973_n26, CO => 
                           DP_OP_1091J1_126_6973_n25, S => C620_DATA2_7);
   DP_OP_1091J1_126_6973_U21 : FA_X1 port map( A => DP_OP_1091J1_126_6973_n31, 
                           B => DataPath_WRF_CUhw_curr_addr_12_port, CI => 
                           DP_OP_1091J1_126_6973_n21, CO => 
                           DP_OP_1091J1_126_6973_n20, S => C620_DATA2_12);
   DP_OP_1091J1_126_6973_U16 : FA_X1 port map( A => DP_OP_1091J1_126_6973_n31, 
                           B => DataPath_WRF_CUhw_curr_addr_17_port, CI => 
                           DP_OP_1091J1_126_6973_n16, CO => 
                           DP_OP_1091J1_126_6973_n15, S => C620_DATA2_17);
   DP_OP_1091J1_126_6973_U15 : FA_X1 port map( A => DP_OP_1091J1_126_6973_n31, 
                           B => DataPath_WRF_CUhw_curr_addr_18_port, CI => 
                           DP_OP_1091J1_126_6973_n15, CO => 
                           DP_OP_1091J1_126_6973_n14, S => C620_DATA2_18);
   DP_OP_751_130_6421_U208 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n26, B 
                           => n8167, ZN => DataPath_ALUhw_i_Q_EXTENDED_34_port)
                           ;
   DP_OP_751_130_6421_U212 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n166, 
                           A2 => DP_OP_751_130_6421_n167, ZN => 
                           DP_OP_751_130_6421_n26);
   DP_OP_751_130_6421_U185 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n23, B 
                           => DP_OP_751_130_6421_n154, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_37_port);
   DP_OP_751_130_6421_U156 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n19, B 
                           => DP_OP_751_130_6421_n138, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_41_port);
   DP_OP_751_130_6421_U161 : NAND2_X1 port map( A1 => n8160, A2 => 
                           DP_OP_751_130_6421_n137, ZN => 
                           DP_OP_751_130_6421_n19);
   DP_OP_751_130_6421_U148 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n18, B 
                           => DP_OP_751_130_6421_n132, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_42_port);
   DP_OP_751_130_6421_U152 : NAND2_X1 port map( A1 => n8166, A2 => 
                           DP_OP_751_130_6421_n131, ZN => 
                           DP_OP_751_130_6421_n18);
   DP_OP_751_130_6421_U142 : XOR2_X1 port map( A => DP_OP_751_130_6421_n17, B 
                           => DP_OP_751_130_6421_n127, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_43_port);
   DP_OP_751_130_6421_U144 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n190, 
                           A2 => DP_OP_751_130_6421_n126, ZN => 
                           DP_OP_751_130_6421_n17);
   DP_OP_751_130_6421_U193 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n24, B 
                           => DP_OP_751_130_6421_n160, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_36_port);
   DP_OP_751_130_6421_U198 : NAND2_X1 port map( A1 => n8162, A2 => 
                           DP_OP_751_130_6421_n159, ZN => 
                           DP_OP_751_130_6421_n24);
   DP_OP_751_130_6421_U134 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n16, B 
                           => DP_OP_751_130_6421_n124, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_44_port);
   DP_OP_751_130_6421_U138 : NAND2_X1 port map( A1 => n8163, A2 => 
                           DP_OP_751_130_6421_n123, ZN => 
                           DP_OP_751_130_6421_n16);
   DP_OP_751_130_6421_U167 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n193, 
                           A2 => DP_OP_751_130_6421_n140, ZN => 
                           DP_OP_751_130_6421_n20);
   DP_OP_751_130_6421_U120 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n14, B 
                           => n7699, ZN => DataPath_ALUhw_i_Q_EXTENDED_46_port)
                           ;
   DP_OP_751_130_6421_U124 : NAND2_X1 port map( A1 => n8168, A2 => 
                           DP_OP_751_130_6421_n115, ZN => 
                           DP_OP_751_130_6421_n14);
   DP_OP_751_130_6421_U113 : XOR2_X1 port map( A => DP_OP_751_130_6421_n13, B 
                           => DP_OP_751_130_6421_n111, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_47_port);
   DP_OP_751_130_6421_U116 : NAND2_X1 port map( A1 => n8150, A2 => 
                           DP_OP_751_130_6421_n110, ZN => 
                           DP_OP_751_130_6421_n13);
   DP_OP_751_130_6421_U89 : NAND2_X1 port map( A1 => n8165, A2 => 
                           DP_OP_751_130_6421_n95, ZN => DP_OP_751_130_6421_n9)
                           ;
   DP_OP_751_130_6421_U93 : XOR2_X1 port map( A => DP_OP_751_130_6421_n10, B =>
                           DP_OP_751_130_6421_n99, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_50_port);
   DP_OP_751_130_6421_U95 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n183, 
                           A2 => DP_OP_751_130_6421_n98, ZN => 
                           DP_OP_751_130_6421_n10);
   DP_OP_751_130_6421_U81 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n181, 
                           A2 => DP_OP_751_130_6421_n90, ZN => 
                           DP_OP_751_130_6421_n8);
   DP_OP_751_130_6421_U56 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n5, B =>
                           n7950, ZN => DataPath_ALUhw_i_Q_EXTENDED_55_port);
   DP_OP_751_130_6421_U61 : NAND2_X1 port map( A1 => n8159, A2 => 
                           DP_OP_751_130_6421_n79, ZN => DP_OP_751_130_6421_n5)
                           ;
   DP_OP_751_130_6421_U65 : XOR2_X1 port map( A => DP_OP_751_130_6421_n6, B => 
                           n7922, Z => DataPath_ALUhw_i_Q_EXTENDED_54_port);
   DP_OP_751_130_6421_U67 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n179, 
                           A2 => DP_OP_751_130_6421_n82, ZN => 
                           DP_OP_751_130_6421_n6);
   DP_OP_751_130_6421_U48 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n4, B =>
                           n7925, ZN => DataPath_ALUhw_i_Q_EXTENDED_56_port);
   DP_OP_751_130_6421_U52 : NAND2_X1 port map( A1 => n8158, A2 => 
                           DP_OP_751_130_6421_n73, ZN => DP_OP_751_130_6421_n4)
                           ;
   DP_OP_751_130_6421_U41 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n268, 
                           A2 => DP_OP_751_130_6421_n366, ZN => 
                           DP_OP_751_130_6421_n63);
   DP_OP_751_130_6421_U55 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n574, 
                           A2 => DP_OP_751_130_6421_n672, ZN => 
                           DP_OP_751_130_6421_n73);
   DP_OP_751_130_6421_U64 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n674, 
                           A2 => DP_OP_751_130_6421_n675, ZN => 
                           DP_OP_751_130_6421_n79);
   DP_OP_751_130_6421_U70 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n676, 
                           A2 => DP_OP_751_130_6421_n774, ZN => 
                           DP_OP_751_130_6421_n82);
   DP_OP_751_130_6421_U69 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n676, A2
                           => DP_OP_751_130_6421_n774, ZN => 
                           DP_OP_751_130_6421_n81);
   DP_OP_751_130_6421_U84 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n778, 
                           A2 => DP_OP_751_130_6421_n876, ZN => 
                           DP_OP_751_130_6421_n90);
   DP_OP_751_130_6421_U83 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n778, A2
                           => DP_OP_751_130_6421_n876, ZN => 
                           DP_OP_751_130_6421_n89);
   DP_OP_751_130_6421_U647 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_20_port, B => 
                           DP_OP_751_130_6421_n813, Z => 
                           DP_OP_751_130_6421_n812);
   DP_OP_751_130_6421_U716 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_19_port, B => n8149, Z
                           => DP_OP_751_130_6421_n913);
   DP_OP_751_130_6421_U98 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n880, 
                           A2 => DP_OP_751_130_6421_n978, ZN => 
                           DP_OP_751_130_6421_n98);
   DP_OP_751_130_6421_U112 : NAND2_X1 port map( A1 => n7187, A2 => 
                           DP_OP_751_130_6421_n1080, ZN => 
                           DP_OP_751_130_6421_n106);
   DP_OP_751_130_6421_U119 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1082,
                           A2 => DP_OP_751_130_6421_n1083, ZN => 
                           DP_OP_751_130_6421_n110);
   DP_OP_751_130_6421_U856 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_15_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1117);
   DP_OP_751_130_6421_U787 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_16_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1016);
   DP_OP_751_130_6421_U121 : AOI21_X1 port map( B1 => n8168, B2 => 
                           DP_OP_751_130_6421_n116, A => 
                           DP_OP_751_130_6421_n113, ZN => 
                           DP_OP_751_130_6421_n111);
   DP_OP_751_130_6421_U127 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1084,
                           A2 => DP_OP_751_130_6421_n1182, ZN => 
                           DP_OP_751_130_6421_n115);
   DP_OP_751_130_6421_U133 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1184,
                           A2 => DP_OP_751_130_6421_n1185, ZN => 
                           DP_OP_751_130_6421_n118);
   DP_OP_751_130_6421_U132 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n1184, 
                           A2 => DP_OP_751_130_6421_n1185, ZN => 
                           DP_OP_751_130_6421_n117);
   DP_OP_751_130_6421_U147 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1286,
                           A2 => DP_OP_751_130_6421_n1287, ZN => 
                           DP_OP_751_130_6421_n126);
   DP_OP_751_130_6421_U146 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n1286, 
                           A2 => DP_OP_751_130_6421_n1287, ZN => 
                           DP_OP_751_130_6421_n125);
   DP_OP_751_130_6421_U155 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1288,
                           A2 => DP_OP_751_130_6421_n1386, ZN => 
                           DP_OP_751_130_6421_n131);
   DP_OP_751_130_6421_U164 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1388,
                           A2 => DP_OP_751_130_6421_n1389, ZN => 
                           DP_OP_751_130_6421_n137);
   DP_OP_751_130_6421_U170 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1390,
                           A2 => DP_OP_751_130_6421_n1488, ZN => 
                           DP_OP_751_130_6421_n140);
   DP_OP_751_130_6421_U178 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1490,
                           A2 => DP_OP_751_130_6421_n1491, ZN => 
                           DP_OP_751_130_6421_n145);
   DP_OP_751_130_6421_U184 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1492,
                           A2 => DP_OP_751_130_6421_n1590, ZN => 
                           DP_OP_751_130_6421_n148);
   DP_OP_751_130_6421_U192 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1592,
                           A2 => DP_OP_751_130_6421_n1593, ZN => 
                           DP_OP_751_130_6421_n153);
   DP_OP_751_130_6421_U201 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1594,
                           A2 => DP_OP_751_130_6421_n1692, ZN => 
                           DP_OP_751_130_6421_n159);
   DP_OP_751_130_6421_U203 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n161, 
                           B2 => DP_OP_751_130_6421_n163, A => 
                           DP_OP_751_130_6421_n162, ZN => 
                           DP_OP_751_130_6421_n160);
   DP_OP_751_130_6421_U207 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1694,
                           A2 => DP_OP_751_130_6421_n1695, ZN => 
                           DP_OP_751_130_6421_n162);
   DP_OP_751_130_6421_U209 : AOI21_X1 port map( B1 => DP_OP_751_130_6421_n166, 
                           B2 => n8167, A => DP_OP_751_130_6421_n165, ZN => 
                           DP_OP_751_130_6421_n163);
   DP_OP_751_130_6421_U215 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1696,
                           A2 => DP_OP_751_130_6421_n1762, ZN => 
                           DP_OP_751_130_6421_n167);
   DP_OP_751_130_6421_U228 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1765,
                           A2 => n7998, ZN => DP_OP_751_130_6421_n174);
   DP_OP_751_130_6421_U206 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n1694, 
                           A2 => DP_OP_751_130_6421_n1695, ZN => 
                           DP_OP_751_130_6421_n161);
   DP_OP_751_130_6421_U1278 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_1_3_port, B => n8146, Z 
                           => DP_OP_751_130_6421_n1695);
   DP_OP_751_130_6421_U183 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n1492, 
                           A2 => DP_OP_751_130_6421_n1590, ZN => 
                           DP_OP_751_130_6421_n147);
   DP_OP_751_130_6421_U1206 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_5_port, B => n7775, Z 
                           => DP_OP_751_130_6421_n1627);
   DP_OP_751_130_6421_U1309 : MUX2_X1 port map( A => DP_OP_751_130_6421_n1795, 
                           B => DataPath_ALUhw_MULT_mux_out_0_4_port, S => 
                           n8148, Z => DP_OP_751_130_6421_n1760);
   DP_OP_751_130_6421_U1137 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_6_port, B => n7797, Z 
                           => DP_OP_751_130_6421_n1526);
   DP_OP_751_130_6421_U169 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n1390, 
                           A2 => DP_OP_751_130_6421_n1488, ZN => 
                           DP_OP_751_130_6421_n139);
   DP_OP_751_130_6421_U1136 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_7_port, B => n7797, Z 
                           => DP_OP_751_130_6421_n1525);
   DP_OP_751_130_6421_U1205 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_6_port, B => n7775, Z 
                           => DP_OP_751_130_6421_n1626);
   DP_OP_751_130_6421_U1308 : MUX2_X1 port map( A => DP_OP_751_130_6421_n1794, 
                           B => DataPath_ALUhw_MULT_mux_out_0_5_port, S => 
                           n8147, Z => DP_OP_751_130_6421_n1759);
   DP_OP_751_130_6421_U1276 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_1_5_port, B => n8146, Z 
                           => DP_OP_751_130_6421_n1729);
   DP_OP_751_130_6421_U1066 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_9_port, B => n7792, Z 
                           => DP_OP_751_130_6421_n1423);
   DP_OP_751_130_6421_U1135 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_8_port, B => n7797, Z 
                           => DP_OP_751_130_6421_n1524);
   DP_OP_751_130_6421_U1204 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_7_port, B => n7775, Z 
                           => DP_OP_751_130_6421_n1625);
   DP_OP_751_130_6421_U996 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_11_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1321);
   DP_OP_751_130_6421_U1065 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_10_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1422);
   DP_OP_751_130_6421_U1134 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_9_port, B => n7797, Z 
                           => DP_OP_751_130_6421_n1523);
   DP_OP_751_130_6421_U1203 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_8_port, B => n7775, Z 
                           => DP_OP_751_130_6421_n1624);
   DP_OP_751_130_6421_U927 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_12_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1220);
   DP_OP_751_130_6421_U925 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_14_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1218);
   DP_OP_751_130_6421_U994 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_13_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1319);
   DP_OP_751_130_6421_U926 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_13_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1219);
   DP_OP_751_130_6421_U1063 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_12_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1420);
   DP_OP_751_130_6421_U995 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_12_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1320);
   DP_OP_751_130_6421_U1132 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_11_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1521);
   DP_OP_751_130_6421_U1064 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_11_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1421);
   DP_OP_751_130_6421_U1201 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_10_port, B => n7775, Z
                           => DP_OP_751_130_6421_n1622);
   DP_OP_751_130_6421_U1133 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_10_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1522);
   DP_OP_751_130_6421_U1202 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_9_port, B => n7775, Z 
                           => DP_OP_751_130_6421_n1623);
   DP_OP_751_130_6421_U1305 : MUX2_X1 port map( A => DP_OP_751_130_6421_n1791, 
                           B => DataPath_ALUhw_MULT_mux_out_0_8_port, S => 
                           n8147, Z => DP_OP_751_130_6421_n1756);
   DP_OP_751_130_6421_U1273 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_1_8_port, B => n8146, Z 
                           => DP_OP_751_130_6421_n1726);
   DP_OP_751_130_6421_U857 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_14_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1118);
   DP_OP_751_130_6421_U97 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n880, A2
                           => DP_OP_751_130_6421_n978, ZN => 
                           DP_OP_751_130_6421_n97);
   DP_OP_751_130_6421_U785 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_18_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1014);
   DP_OP_751_130_6421_U854 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_17_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1115);
   DP_OP_751_130_6421_U786 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_17_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1015);
   DP_OP_751_130_6421_U923 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_16_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1216);
   DP_OP_751_130_6421_U855 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_16_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1116);
   DP_OP_751_130_6421_U992 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_15_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1317);
   DP_OP_751_130_6421_U924 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_15_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1217);
   DP_OP_751_130_6421_U1061 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_14_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1418);
   DP_OP_751_130_6421_U993 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_14_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1318);
   DP_OP_751_130_6421_U1130 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_13_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1519);
   DP_OP_751_130_6421_U1062 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_13_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1419);
   DP_OP_751_130_6421_U1199 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_12_port, B => n7775, Z
                           => DP_OP_751_130_6421_n1620);
   DP_OP_751_130_6421_U1131 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_12_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1520);
   DP_OP_751_130_6421_U1200 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_11_port, B => n7775, Z
                           => DP_OP_751_130_6421_n1621);
   DP_OP_751_130_6421_U1271 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_1_10_port, B => n8146, Z
                           => DP_OP_751_130_6421_n1724);
   DP_OP_751_130_6421_U646 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_21_port, B => 
                           DP_OP_751_130_6421_n813, Z => 
                           DP_OP_751_130_6421_n811);
   DP_OP_751_130_6421_U715 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_20_port, B => n8149, Z
                           => DP_OP_751_130_6421_n912);
   DP_OP_751_130_6421_U784 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_19_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1013);
   DP_OP_751_130_6421_U853 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_18_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1114);
   DP_OP_751_130_6421_U922 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_17_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1215);
   DP_OP_751_130_6421_U991 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_16_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1316);
   DP_OP_751_130_6421_U1060 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_15_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1417);
   DP_OP_751_130_6421_U1129 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_14_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1518);
   DP_OP_751_130_6421_U1198 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_13_port, B => n7775, Z
                           => DP_OP_751_130_6421_n1619);
   DP_OP_751_130_6421_U577 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_22_port, B => 
                           DP_OP_751_130_6421_n711, Z => 
                           DP_OP_751_130_6421_n710);
   DP_OP_751_130_6421_U576 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_23_port, B => 
                           DP_OP_751_130_6421_n711, Z => 
                           DP_OP_751_130_6421_n709);
   DP_OP_751_130_6421_U645 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_22_port, B => 
                           DP_OP_751_130_6421_n813, Z => 
                           DP_OP_751_130_6421_n810);
   DP_OP_751_130_6421_U714 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_21_port, B => n8149, Z
                           => DP_OP_751_130_6421_n911);
   DP_OP_751_130_6421_U783 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_20_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1012);
   DP_OP_751_130_6421_U852 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_19_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1113);
   DP_OP_751_130_6421_U921 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_18_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1214);
   DP_OP_751_130_6421_U990 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_17_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1315);
   DP_OP_751_130_6421_U1059 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_16_port, B => n8144, Z
                           => DP_OP_751_130_6421_n1416);
   DP_OP_751_130_6421_U1128 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_15_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1517);
   DP_OP_751_130_6421_U1197 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_14_port, B => n7775, Z
                           => DP_OP_751_130_6421_n1618);
   DP_OP_751_130_6421_U507 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_24_port, B => n7817, 
                           Z => DP_OP_751_130_6421_n608);
   DP_OP_751_130_6421_U506 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_25_port, B => n7817, 
                           Z => DP_OP_751_130_6421_n607);
   DP_OP_751_130_6421_U575 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_24_port, B => 
                           DP_OP_751_130_6421_n711, Z => 
                           DP_OP_751_130_6421_n708);
   DP_OP_751_130_6421_U644 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_23_port, B => 
                           DP_OP_751_130_6421_n813, Z => 
                           DP_OP_751_130_6421_n809);
   DP_OP_751_130_6421_U713 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_22_port, B => n8149, Z
                           => DP_OP_751_130_6421_n910);
   DP_OP_751_130_6421_U782 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_21_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1011);
   DP_OP_751_130_6421_U851 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_20_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1112);
   DP_OP_751_130_6421_U920 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_19_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1213);
   DP_OP_751_130_6421_U989 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_18_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1314);
   DP_OP_751_130_6421_U1058 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_17_port, B => n8144, Z
                           => DP_OP_751_130_6421_n1415);
   DP_OP_751_130_6421_U1127 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_16_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1516);
   DP_OP_751_130_6421_U1196 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_15_port, B => n7775, Z
                           => DP_OP_751_130_6421_n1617);
   DP_OP_751_130_6421_U1299 : MUX2_X1 port map( A => DP_OP_751_130_6421_n1785, 
                           B => DataPath_ALUhw_MULT_mux_out_0_14_port, S => 
                           n8147, Z => DP_OP_751_130_6421_n1750);
   DP_OP_751_130_6421_U437 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_13_26_port, B => 
                           DP_OP_751_130_6421_n507, Z => 
                           DP_OP_751_130_6421_n506);
   DP_OP_751_130_6421_U436 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_13_27_port, B => 
                           DP_OP_751_130_6421_n507, Z => 
                           DP_OP_751_130_6421_n505);
   DP_OP_751_130_6421_U505 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_26_port, B => n7817, 
                           Z => DP_OP_751_130_6421_n606);
   DP_OP_751_130_6421_U643 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_24_port, B => 
                           DP_OP_751_130_6421_n813, Z => 
                           DP_OP_751_130_6421_n808);
   DP_OP_751_130_6421_U712 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_23_port, B => n8149, Z
                           => DP_OP_751_130_6421_n909);
   DP_OP_751_130_6421_U781 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_22_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1010);
   DP_OP_751_130_6421_U850 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_21_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1111);
   DP_OP_751_130_6421_U919 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_20_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1212);
   DP_OP_751_130_6421_U988 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_19_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1313);
   DP_OP_751_130_6421_U1057 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_18_port, B => n8144, Z
                           => DP_OP_751_130_6421_n1414);
   DP_OP_751_130_6421_U1126 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_17_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1515);
   DP_OP_751_130_6421_U367 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_14_28_port, B => 
                           DP_OP_751_130_6421_n405, Z => 
                           DP_OP_751_130_6421_n404);
   DP_OP_751_130_6421_U366 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_14_29_port, B => 
                           DP_OP_751_130_6421_n405, Z => 
                           DP_OP_751_130_6421_n403);
   DP_OP_751_130_6421_U435 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_13_28_port, B => 
                           DP_OP_751_130_6421_n507, Z => 
                           DP_OP_751_130_6421_n504);
   DP_OP_751_130_6421_U504 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_27_port, B => n7817, 
                           Z => DP_OP_751_130_6421_n605);
   DP_OP_751_130_6421_U573 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_26_port, B => 
                           DP_OP_751_130_6421_n711, Z => 
                           DP_OP_751_130_6421_n706);
   DP_OP_751_130_6421_U642 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_25_port, B => 
                           DP_OP_751_130_6421_n813, Z => 
                           DP_OP_751_130_6421_n807);
   DP_OP_751_130_6421_U711 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_24_port, B => n8149, Z
                           => DP_OP_751_130_6421_n908);
   DP_OP_751_130_6421_U780 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_23_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1009);
   DP_OP_751_130_6421_U849 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_22_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1110);
   DP_OP_751_130_6421_U918 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_21_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1211);
   DP_OP_751_130_6421_U987 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_20_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1312);
   DP_OP_751_130_6421_U1056 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_19_port, B => n8144, Z
                           => DP_OP_751_130_6421_n1413);
   DP_OP_751_130_6421_U1125 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_18_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1514);
   DP_OP_751_130_6421_U1297 : MUX2_X1 port map( A => DP_OP_751_130_6421_n1783, 
                           B => DataPath_ALUhw_MULT_mux_out_0_16_port, S => 
                           n8147, Z => DP_OP_751_130_6421_n1748);
   DP_OP_751_130_6421_U297 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_15_30_port, B => n7816, 
                           Z => DP_OP_751_130_6421_n302);
   DP_OP_751_130_6421_U1282 : MUX2_X1 port map( A => DP_OP_751_130_6421_n1768, 
                           B => DataPath_ALUhw_MULT_mux_out_0_31_port, S => 
                           n8147, Z => DP_OP_751_130_6421_n1733);
   DP_OP_751_130_6421_U1250 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_1_31_port, B => n8146, Z
                           => DP_OP_751_130_6421_n1703);
   DP_OP_751_130_6421_U1180 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_31_port, B => n8145, Z
                           => DP_OP_751_130_6421_n1601);
   DP_OP_751_130_6421_U1112 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_31_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1501);
   DP_OP_751_130_6421_U1044 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_31_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1401);
   DP_OP_751_130_6421_U976 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_31_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1301);
   DP_OP_751_130_6421_U908 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_31_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1201);
   DP_OP_751_130_6421_U840 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_31_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1101);
   DP_OP_751_130_6421_U772 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_31_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1001);
   DP_OP_751_130_6421_U704 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_31_port, B => n8149, Z
                           => DP_OP_751_130_6421_n901);
   DP_OP_751_130_6421_U636 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_31_port, B => 
                           DP_OP_751_130_6421_n813, Z => 
                           DP_OP_751_130_6421_n801);
   DP_OP_751_130_6421_U568 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_31_port, B => 
                           DP_OP_751_130_6421_n711, Z => 
                           DP_OP_751_130_6421_n701);
   DP_OP_751_130_6421_U500 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_31_port, B => n7817, 
                           Z => DP_OP_751_130_6421_n601);
   DP_OP_751_130_6421_U432 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_13_31_port, B => 
                           DP_OP_751_130_6421_n507, Z => 
                           DP_OP_751_130_6421_n501);
   DP_OP_751_130_6421_U364 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_14_31_port, B => 
                           DP_OP_751_130_6421_n405, Z => 
                           DP_OP_751_130_6421_n401);
   DP_OP_751_130_6421_U296 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_15_31_port, B => n7816, 
                           Z => DP_OP_751_130_6421_n301);
   DP_OP_751_130_6421_U1181 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_30_port, B => n8145, Z
                           => DP_OP_751_130_6421_n1602);
   DP_OP_751_130_6421_U1113 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_30_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1502);
   DP_OP_751_130_6421_U1045 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_30_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1402);
   DP_OP_751_130_6421_U977 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_30_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1302);
   DP_OP_751_130_6421_U909 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_30_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1202);
   DP_OP_751_130_6421_U841 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_30_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1102);
   DP_OP_751_130_6421_U773 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_30_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1002);
   DP_OP_751_130_6421_U705 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_30_port, B => n8149, Z
                           => DP_OP_751_130_6421_n902);
   DP_OP_751_130_6421_U637 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_30_port, B => 
                           DP_OP_751_130_6421_n813, Z => 
                           DP_OP_751_130_6421_n802);
   DP_OP_751_130_6421_U569 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_30_port, B => 
                           DP_OP_751_130_6421_n711, Z => 
                           DP_OP_751_130_6421_n702);
   DP_OP_751_130_6421_U501 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_30_port, B => n7817, 
                           Z => DP_OP_751_130_6421_n602);
   DP_OP_751_130_6421_U433 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_13_30_port, B => 
                           DP_OP_751_130_6421_n507, Z => 
                           DP_OP_751_130_6421_n502);
   DP_OP_751_130_6421_U365 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_14_30_port, B => n7821, 
                           Z => DP_OP_751_130_6421_n402);
   DP_OP_751_130_6421_U1284 : MUX2_X1 port map( A => DP_OP_751_130_6421_n1770, 
                           B => DataPath_ALUhw_MULT_mux_out_0_29_port, S => 
                           n8148, Z => DP_OP_751_130_6421_n1735);
   DP_OP_751_130_6421_U1182 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_29_port, B => n8145, Z
                           => DP_OP_751_130_6421_n1603);
   DP_OP_751_130_6421_U1114 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_29_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1503);
   DP_OP_751_130_6421_U1046 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_29_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1403);
   DP_OP_751_130_6421_U978 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_29_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1303);
   DP_OP_751_130_6421_U910 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_29_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1203);
   DP_OP_751_130_6421_U842 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_29_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1103);
   DP_OP_751_130_6421_U774 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_29_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1003);
   DP_OP_751_130_6421_U706 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_29_port, B => n8149, Z
                           => DP_OP_751_130_6421_n903);
   DP_OP_751_130_6421_U638 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_29_port, B => 
                           DP_OP_751_130_6421_n813, Z => 
                           DP_OP_751_130_6421_n803);
   DP_OP_751_130_6421_U570 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_29_port, B => 
                           DP_OP_751_130_6421_n711, Z => 
                           DP_OP_751_130_6421_n703);
   DP_OP_751_130_6421_U502 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_29_port, B => n7817, 
                           Z => DP_OP_751_130_6421_n603);
   DP_OP_751_130_6421_U434 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_13_29_port, B => 
                           DP_OP_751_130_6421_n507, Z => 
                           DP_OP_751_130_6421_n503);
   DP_OP_751_130_6421_U1183 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_28_port, B => n8145, Z
                           => DP_OP_751_130_6421_n1604);
   DP_OP_751_130_6421_U1115 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_28_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1504);
   DP_OP_751_130_6421_U1047 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_28_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1404);
   DP_OP_751_130_6421_U979 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_28_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1304);
   DP_OP_751_130_6421_U911 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_28_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1204);
   DP_OP_751_130_6421_U843 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_28_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1104);
   DP_OP_751_130_6421_U775 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_28_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1004);
   DP_OP_751_130_6421_U707 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_28_port, B => n8149, Z
                           => DP_OP_751_130_6421_n904);
   DP_OP_751_130_6421_U639 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_28_port, B => 
                           DP_OP_751_130_6421_n813, Z => 
                           DP_OP_751_130_6421_n804);
   DP_OP_751_130_6421_U571 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_28_port, B => 
                           DP_OP_751_130_6421_n711, Z => 
                           DP_OP_751_130_6421_n704);
   DP_OP_751_130_6421_U503 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_12_28_port, B => n7817, 
                           Z => DP_OP_751_130_6421_n604);
   DP_OP_751_130_6421_U1286 : MUX2_X1 port map( A => DP_OP_751_130_6421_n1772, 
                           B => DataPath_ALUhw_MULT_mux_out_0_27_port, S => 
                           n8147, Z => DP_OP_751_130_6421_n1737);
   DP_OP_751_130_6421_U1116 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_27_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1505);
   DP_OP_751_130_6421_U1048 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_27_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1405);
   DP_OP_751_130_6421_U980 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_27_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1305);
   DP_OP_751_130_6421_U912 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_27_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1205);
   DP_OP_751_130_6421_U844 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_27_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1105);
   DP_OP_751_130_6421_U776 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_27_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1005);
   DP_OP_751_130_6421_U708 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_27_port, B => n8149, Z
                           => DP_OP_751_130_6421_n905);
   DP_OP_751_130_6421_U640 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_27_port, B => 
                           DP_OP_751_130_6421_n813, Z => 
                           DP_OP_751_130_6421_n805);
   DP_OP_751_130_6421_U572 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_11_27_port, B => 
                           DP_OP_751_130_6421_n711, Z => 
                           DP_OP_751_130_6421_n705);
   DP_OP_751_130_6421_U1117 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_26_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1506);
   DP_OP_751_130_6421_U1049 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_26_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1406);
   DP_OP_751_130_6421_U981 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_26_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1306);
   DP_OP_751_130_6421_U913 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_26_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1206);
   DP_OP_751_130_6421_U845 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_26_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1106);
   DP_OP_751_130_6421_U777 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_26_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1006);
   DP_OP_751_130_6421_U709 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_26_port, B => n8149, Z
                           => DP_OP_751_130_6421_n906);
   DP_OP_751_130_6421_U641 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_10_26_port, B => 
                           DP_OP_751_130_6421_n813, Z => 
                           DP_OP_751_130_6421_n806);
   DP_OP_751_130_6421_U1288 : MUX2_X1 port map( A => DP_OP_751_130_6421_n1774, 
                           B => DataPath_ALUhw_MULT_mux_out_0_25_port, S => 
                           n8147, Z => DP_OP_751_130_6421_n1739);
   DP_OP_751_130_6421_U1050 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_25_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1407);
   DP_OP_751_130_6421_U982 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_25_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1307);
   DP_OP_751_130_6421_U914 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_25_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1207);
   DP_OP_751_130_6421_U846 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_25_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1107);
   DP_OP_751_130_6421_U778 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_25_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1007);
   DP_OP_751_130_6421_U710 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_9_25_port, B => n8149, Z
                           => DP_OP_751_130_6421_n907);
   DP_OP_751_130_6421_U1187 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_24_port, B => n8145, Z
                           => DP_OP_751_130_6421_n1608);
   DP_OP_751_130_6421_U1119 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_24_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1508);
   DP_OP_751_130_6421_U1051 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_24_port, B => n7792, Z
                           => DP_OP_751_130_6421_n1408);
   DP_OP_751_130_6421_U983 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_24_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1308);
   DP_OP_751_130_6421_U847 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_24_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1108);
   DP_OP_751_130_6421_U779 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_8_24_port, B => 
                           DP_OP_751_130_6421_n1017, Z => 
                           DP_OP_751_130_6421_n1008);
   DP_OP_751_130_6421_U1188 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_23_port, B => n8145, Z
                           => DP_OP_751_130_6421_n1609);
   DP_OP_751_130_6421_U1120 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_23_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1509);
   DP_OP_751_130_6421_U1052 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_23_port, B => n8144, Z
                           => DP_OP_751_130_6421_n1409);
   DP_OP_751_130_6421_U984 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_23_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1309);
   DP_OP_751_130_6421_U916 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_23_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1209);
   DP_OP_751_130_6421_U848 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_7_23_port, B => n7793, Z
                           => DP_OP_751_130_6421_n1109);
   DP_OP_751_130_6421_U1291 : MUX2_X1 port map( A => DP_OP_751_130_6421_n1777, 
                           B => DataPath_ALUhw_MULT_mux_out_0_22_port, S => 
                           n8147, Z => DP_OP_751_130_6421_n1742);
   DP_OP_751_130_6421_U1121 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_22_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1510);
   DP_OP_751_130_6421_U985 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_22_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1310);
   DP_OP_751_130_6421_U917 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_6_22_port, B => 
                           DP_OP_751_130_6421_n1221, Z => 
                           DP_OP_751_130_6421_n1210);
   DP_OP_751_130_6421_U1122 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_21_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1511);
   DP_OP_751_130_6421_U1054 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_21_port, B => n8144, Z
                           => DP_OP_751_130_6421_n1411);
   DP_OP_751_130_6421_U986 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_5_21_port, B => 
                           DP_OP_751_130_6421_n1323, Z => 
                           DP_OP_751_130_6421_n1311);
   DP_OP_751_130_6421_U1191 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_20_port, B => n8145, Z
                           => DP_OP_751_130_6421_n1612);
   DP_OP_751_130_6421_U1123 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_20_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1512);
   DP_OP_751_130_6421_U1055 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_4_20_port, B => n8144, Z
                           => DP_OP_751_130_6421_n1412);
   DP_OP_751_130_6421_U1192 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_19_port, B => n7775, Z
                           => DP_OP_751_130_6421_n1613);
   DP_OP_751_130_6421_U1124 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_3_19_port, B => n7797, Z
                           => DP_OP_751_130_6421_n1513);
   DP_OP_751_130_6421_U1193 : XOR2_X1 port map( A => 
                           DataPath_ALUhw_MULT_mux_out_2_18_port, B => n7775, Z
                           => DP_OP_751_130_6421_n1614);
   DP_OP_751_130_6421_U1242 : HA_X1 port map( A => DP_OP_751_130_6421_n1729, B 
                           => DP_OP_751_130_6421_n1759, CO => 
                           DP_OP_751_130_6421_n1689, S => 
                           DP_OP_751_130_6421_n1690);
   DP_OP_751_130_6421_U1239 : HA_X1 port map( A => DP_OP_751_130_6421_n1726, B 
                           => DP_OP_751_130_6421_n1756, CO => 
                           DP_OP_751_130_6421_n1683, S => 
                           DP_OP_751_130_6421_n1684);
   DP_OP_751_130_6421_U1233 : HA_X1 port map( A => DP_OP_751_130_6421_n1720, B 
                           => DP_OP_751_130_6421_n1750, CO => 
                           DP_OP_751_130_6421_n1671, S => 
                           DP_OP_751_130_6421_n1672);
   DP_OP_751_130_6421_U1228 : HA_X1 port map( A => DP_OP_751_130_6421_n1715, B 
                           => DP_OP_751_130_6421_n1745, CO => 
                           DP_OP_751_130_6421_n1661, S => 
                           DP_OP_751_130_6421_n1662);
   DP_OP_751_130_6421_U1218 : HA_X1 port map( A => DP_OP_751_130_6421_n1705, B 
                           => DP_OP_751_130_6421_n1735, CO => 
                           DP_OP_751_130_6421_n1641, S => 
                           DP_OP_751_130_6421_n1642);
   DP_OP_751_130_6421_U1172 : FA_X1 port map( A => DP_OP_751_130_6421_n1691, B 
                           => DP_OP_751_130_6421_n1627, CI => 
                           DP_OP_751_130_6421_n1690, CO => 
                           DP_OP_751_130_6421_n1591, S => 
                           DP_OP_751_130_6421_n1592);
   DP_OP_751_130_6421_U1171 : FA_X1 port map( A => DP_OP_751_130_6421_n1689, B 
                           => DP_OP_751_130_6421_n1626, CI => 
                           DP_OP_751_130_6421_n1688, CO => 
                           DP_OP_751_130_6421_n1589, S => 
                           DP_OP_751_130_6421_n1590);
   DP_OP_751_130_6421_U1170 : FA_X1 port map( A => DP_OP_751_130_6421_n1687, B 
                           => DP_OP_751_130_6421_n1625, CI => 
                           DP_OP_751_130_6421_n1686, CO => 
                           DP_OP_751_130_6421_n1587, S => 
                           DP_OP_751_130_6421_n1588);
   DP_OP_751_130_6421_U1169 : FA_X1 port map( A => DP_OP_751_130_6421_n1685, B 
                           => DP_OP_751_130_6421_n1624, CI => 
                           DP_OP_751_130_6421_n1684, CO => 
                           DP_OP_751_130_6421_n1585, S => 
                           DP_OP_751_130_6421_n1586);
   DP_OP_751_130_6421_U1168 : FA_X1 port map( A => DP_OP_751_130_6421_n1683, B 
                           => DP_OP_751_130_6421_n1623, CI => 
                           DP_OP_751_130_6421_n1682, CO => 
                           DP_OP_751_130_6421_n1583, S => 
                           DP_OP_751_130_6421_n1584);
   DP_OP_751_130_6421_U1167 : FA_X1 port map( A => DP_OP_751_130_6421_n1681, B 
                           => DP_OP_751_130_6421_n1622, CI => 
                           DP_OP_751_130_6421_n1680, CO => 
                           DP_OP_751_130_6421_n1581, S => 
                           DP_OP_751_130_6421_n1582);
   DP_OP_751_130_6421_U1166 : FA_X1 port map( A => n7189, B => 
                           DP_OP_751_130_6421_n1621, CI => 
                           DP_OP_751_130_6421_n1678, CO => 
                           DP_OP_751_130_6421_n1579, S => 
                           DP_OP_751_130_6421_n1580);
   DP_OP_751_130_6421_U1165 : FA_X1 port map( A => DP_OP_751_130_6421_n1677, B 
                           => DP_OP_751_130_6421_n1620, CI => 
                           DP_OP_751_130_6421_n1676, CO => 
                           DP_OP_751_130_6421_n1577, S => 
                           DP_OP_751_130_6421_n1578);
   DP_OP_751_130_6421_U1164 : FA_X1 port map( A => DP_OP_751_130_6421_n1675, B 
                           => DP_OP_751_130_6421_n1619, CI => 
                           DP_OP_751_130_6421_n1674, CO => 
                           DP_OP_751_130_6421_n1575, S => 
                           DP_OP_751_130_6421_n1576);
   DP_OP_751_130_6421_U1163 : FA_X1 port map( A => DP_OP_751_130_6421_n1673, B 
                           => DP_OP_751_130_6421_n1618, CI => 
                           DP_OP_751_130_6421_n1672, CO => 
                           DP_OP_751_130_6421_n1573, S => 
                           DP_OP_751_130_6421_n1574);
   DP_OP_751_130_6421_U1162 : FA_X1 port map( A => DP_OP_751_130_6421_n1671, B 
                           => DP_OP_751_130_6421_n1617, CI => 
                           DP_OP_751_130_6421_n1670, CO => 
                           DP_OP_751_130_6421_n1571, S => 
                           DP_OP_751_130_6421_n1572);
   DP_OP_751_130_6421_U1161 : FA_X1 port map( A => DP_OP_751_130_6421_n1669, B 
                           => DP_OP_751_130_6421_n1616, CI => 
                           DP_OP_751_130_6421_n1668, CO => 
                           DP_OP_751_130_6421_n1569, S => 
                           DP_OP_751_130_6421_n1570);
   DP_OP_751_130_6421_U1159 : FA_X1 port map( A => DP_OP_751_130_6421_n1665, B 
                           => DP_OP_751_130_6421_n1614, CI => 
                           DP_OP_751_130_6421_n1664, CO => 
                           DP_OP_751_130_6421_n1565, S => 
                           DP_OP_751_130_6421_n1566);
   DP_OP_751_130_6421_U1158 : FA_X1 port map( A => DP_OP_751_130_6421_n1663, B 
                           => DP_OP_751_130_6421_n1613, CI => 
                           DP_OP_751_130_6421_n1662, CO => 
                           DP_OP_751_130_6421_n1563, S => 
                           DP_OP_751_130_6421_n1564);
   DP_OP_751_130_6421_U1157 : FA_X1 port map( A => DP_OP_751_130_6421_n1661, B 
                           => DP_OP_751_130_6421_n1612, CI => 
                           DP_OP_751_130_6421_n1660, CO => 
                           DP_OP_751_130_6421_n1561, S => 
                           DP_OP_751_130_6421_n1562);
   DP_OP_751_130_6421_U1154 : FA_X1 port map( A => DP_OP_751_130_6421_n1609, B 
                           => DP_OP_751_130_6421_n1655, CI => 
                           DP_OP_751_130_6421_n1654, CO => 
                           DP_OP_751_130_6421_n1555, S => 
                           DP_OP_751_130_6421_n1556);
   DP_OP_751_130_6421_U1153 : FA_X1 port map( A => DP_OP_751_130_6421_n1608, B 
                           => DP_OP_751_130_6421_n1653, CI => 
                           DP_OP_751_130_6421_n1652, CO => 
                           DP_OP_751_130_6421_n1553, S => 
                           DP_OP_751_130_6421_n1554);
   DP_OP_751_130_6421_U1150 : FA_X1 port map( A => DP_OP_751_130_6421_n1647, B 
                           => DP_OP_751_130_6421_n1605, CI => 
                           DP_OP_751_130_6421_n1646, CO => 
                           DP_OP_751_130_6421_n1547, S => 
                           DP_OP_751_130_6421_n1548);
   DP_OP_751_130_6421_U1149 : FA_X1 port map( A => DP_OP_751_130_6421_n1645, B 
                           => DP_OP_751_130_6421_n1604, CI => 
                           DP_OP_751_130_6421_n1644, CO => 
                           DP_OP_751_130_6421_n1545, S => 
                           DP_OP_751_130_6421_n1546);
   DP_OP_751_130_6421_U1147 : FA_X1 port map( A => DP_OP_751_130_6421_n1641, B 
                           => DP_OP_751_130_6421_n1602, CI => 
                           DP_OP_751_130_6421_n1640, CO => 
                           DP_OP_751_130_6421_n1541, S => 
                           DP_OP_751_130_6421_n1542);
   DP_OP_751_130_6421_U1146 : FA_X1 port map( A => DP_OP_751_130_6421_n1639, B 
                           => DP_OP_751_130_6421_n1601, CI => 
                           DP_OP_751_130_6421_n1638, CO => n_3875, S => 
                           DP_OP_751_130_6421_n1540);
   DP_OP_751_130_6421_U1103 : FA_X1 port map( A => DP_OP_751_130_6421_n1526, B 
                           => n7797, CI => DP_OP_751_130_6421_n1591, CO => 
                           DP_OP_751_130_6421_n1491, S => 
                           DP_OP_751_130_6421_n1492);
   DP_OP_751_130_6421_U1102 : FA_X1 port map( A => DP_OP_751_130_6421_n1589, B 
                           => DP_OP_751_130_6421_n1525, CI => 
                           DP_OP_751_130_6421_n1588, CO => 
                           DP_OP_751_130_6421_n1489, S => 
                           DP_OP_751_130_6421_n1490);
   DP_OP_751_130_6421_U1101 : FA_X1 port map( A => DP_OP_751_130_6421_n1587, B 
                           => DP_OP_751_130_6421_n1524, CI => 
                           DP_OP_751_130_6421_n1586, CO => 
                           DP_OP_751_130_6421_n1487, S => 
                           DP_OP_751_130_6421_n1488);
   DP_OP_751_130_6421_U1100 : FA_X1 port map( A => DP_OP_751_130_6421_n1585, B 
                           => DP_OP_751_130_6421_n1523, CI => 
                           DP_OP_751_130_6421_n1584, CO => 
                           DP_OP_751_130_6421_n1485, S => 
                           DP_OP_751_130_6421_n1486);
   DP_OP_751_130_6421_U1099 : FA_X1 port map( A => DP_OP_751_130_6421_n1583, B 
                           => DP_OP_751_130_6421_n1522, CI => 
                           DP_OP_751_130_6421_n1582, CO => 
                           DP_OP_751_130_6421_n1483, S => 
                           DP_OP_751_130_6421_n1484);
   DP_OP_751_130_6421_U1098 : FA_X1 port map( A => DP_OP_751_130_6421_n1581, B 
                           => DP_OP_751_130_6421_n1521, CI => 
                           DP_OP_751_130_6421_n1580, CO => 
                           DP_OP_751_130_6421_n1481, S => 
                           DP_OP_751_130_6421_n1482);
   DP_OP_751_130_6421_U1097 : FA_X1 port map( A => DP_OP_751_130_6421_n1579, B 
                           => DP_OP_751_130_6421_n1520, CI => 
                           DP_OP_751_130_6421_n1578, CO => 
                           DP_OP_751_130_6421_n1479, S => 
                           DP_OP_751_130_6421_n1480);
   DP_OP_751_130_6421_U1096 : FA_X1 port map( A => DP_OP_751_130_6421_n1577, B 
                           => DP_OP_751_130_6421_n1519, CI => 
                           DP_OP_751_130_6421_n1576, CO => 
                           DP_OP_751_130_6421_n1477, S => 
                           DP_OP_751_130_6421_n1478);
   DP_OP_751_130_6421_U1095 : FA_X1 port map( A => DP_OP_751_130_6421_n1575, B 
                           => DP_OP_751_130_6421_n1518, CI => 
                           DP_OP_751_130_6421_n1574, CO => 
                           DP_OP_751_130_6421_n1475, S => 
                           DP_OP_751_130_6421_n1476);
   DP_OP_751_130_6421_U1094 : FA_X1 port map( A => DP_OP_751_130_6421_n1573, B 
                           => DP_OP_751_130_6421_n1517, CI => 
                           DP_OP_751_130_6421_n1572, CO => 
                           DP_OP_751_130_6421_n1473, S => 
                           DP_OP_751_130_6421_n1474);
   DP_OP_751_130_6421_U1093 : FA_X1 port map( A => DP_OP_751_130_6421_n1571, B 
                           => DP_OP_751_130_6421_n1516, CI => 
                           DP_OP_751_130_6421_n1570, CO => 
                           DP_OP_751_130_6421_n1471, S => 
                           DP_OP_751_130_6421_n1472);
   DP_OP_751_130_6421_U1091 : FA_X1 port map( A => DP_OP_751_130_6421_n1567, B 
                           => DP_OP_751_130_6421_n1514, CI => 
                           DP_OP_751_130_6421_n1566, CO => 
                           DP_OP_751_130_6421_n1467, S => 
                           DP_OP_751_130_6421_n1468);
   DP_OP_751_130_6421_U1090 : FA_X1 port map( A => DP_OP_751_130_6421_n1565, B 
                           => DP_OP_751_130_6421_n1513, CI => 
                           DP_OP_751_130_6421_n1564, CO => 
                           DP_OP_751_130_6421_n1465, S => 
                           DP_OP_751_130_6421_n1466);
   DP_OP_751_130_6421_U1089 : FA_X1 port map( A => DP_OP_751_130_6421_n1563, B 
                           => DP_OP_751_130_6421_n1512, CI => 
                           DP_OP_751_130_6421_n1562, CO => 
                           DP_OP_751_130_6421_n1463, S => 
                           DP_OP_751_130_6421_n1464);
   DP_OP_751_130_6421_U1087 : FA_X1 port map( A => DP_OP_751_130_6421_n1559, B 
                           => DP_OP_751_130_6421_n1510, CI => 
                           DP_OP_751_130_6421_n1558, CO => 
                           DP_OP_751_130_6421_n1459, S => 
                           DP_OP_751_130_6421_n1460);
   DP_OP_751_130_6421_U1086 : FA_X1 port map( A => DP_OP_751_130_6421_n1557, B 
                           => DP_OP_751_130_6421_n1509, CI => 
                           DP_OP_751_130_6421_n1556, CO => 
                           DP_OP_751_130_6421_n1457, S => 
                           DP_OP_751_130_6421_n1458);
   DP_OP_751_130_6421_U1085 : FA_X1 port map( A => DP_OP_751_130_6421_n1555, B 
                           => DP_OP_751_130_6421_n1508, CI => 
                           DP_OP_751_130_6421_n1554, CO => 
                           DP_OP_751_130_6421_n1455, S => 
                           DP_OP_751_130_6421_n1456);
   DP_OP_751_130_6421_U1083 : FA_X1 port map( A => DP_OP_751_130_6421_n1551, B 
                           => DP_OP_751_130_6421_n1506, CI => 
                           DP_OP_751_130_6421_n1550, CO => 
                           DP_OP_751_130_6421_n1451, S => 
                           DP_OP_751_130_6421_n1452);
   DP_OP_751_130_6421_U1081 : FA_X1 port map( A => DP_OP_751_130_6421_n1547, B 
                           => DP_OP_751_130_6421_n1504, CI => 
                           DP_OP_751_130_6421_n1546, CO => 
                           DP_OP_751_130_6421_n1447, S => 
                           DP_OP_751_130_6421_n1448);
   DP_OP_751_130_6421_U1079 : FA_X1 port map( A => DP_OP_751_130_6421_n1543, B 
                           => DP_OP_751_130_6421_n1502, CI => 
                           DP_OP_751_130_6421_n1542, CO => 
                           DP_OP_751_130_6421_n1443, S => 
                           DP_OP_751_130_6421_n1444);
   DP_OP_751_130_6421_U1078 : FA_X1 port map( A => DP_OP_751_130_6421_n1541, B 
                           => DP_OP_751_130_6421_n1501, CI => 
                           DP_OP_751_130_6421_n1540, CO => n_3876, S => 
                           DP_OP_751_130_6421_n1442);
   DP_OP_751_130_6421_U1032 : FA_X1 port map( A => DP_OP_751_130_6421_n1487, B 
                           => DP_OP_751_130_6421_n1423, CI => 
                           DP_OP_751_130_6421_n1486, CO => 
                           DP_OP_751_130_6421_n1387, S => 
                           DP_OP_751_130_6421_n1388);
   DP_OP_751_130_6421_U1031 : FA_X1 port map( A => DP_OP_751_130_6421_n1485, B 
                           => DP_OP_751_130_6421_n1422, CI => 
                           DP_OP_751_130_6421_n1484, CO => 
                           DP_OP_751_130_6421_n1385, S => 
                           DP_OP_751_130_6421_n1386);
   DP_OP_751_130_6421_U1030 : FA_X1 port map( A => DP_OP_751_130_6421_n1483, B 
                           => DP_OP_751_130_6421_n1421, CI => 
                           DP_OP_751_130_6421_n1482, CO => 
                           DP_OP_751_130_6421_n1383, S => 
                           DP_OP_751_130_6421_n1384);
   DP_OP_751_130_6421_U1029 : FA_X1 port map( A => DP_OP_751_130_6421_n1481, B 
                           => DP_OP_751_130_6421_n1420, CI => 
                           DP_OP_751_130_6421_n1480, CO => 
                           DP_OP_751_130_6421_n1381, S => 
                           DP_OP_751_130_6421_n1382);
   DP_OP_751_130_6421_U1028 : FA_X1 port map( A => DP_OP_751_130_6421_n1479, B 
                           => DP_OP_751_130_6421_n1419, CI => 
                           DP_OP_751_130_6421_n1478, CO => 
                           DP_OP_751_130_6421_n1379, S => 
                           DP_OP_751_130_6421_n1380);
   DP_OP_751_130_6421_U1027 : FA_X1 port map( A => DP_OP_751_130_6421_n1477, B 
                           => DP_OP_751_130_6421_n1418, CI => 
                           DP_OP_751_130_6421_n1476, CO => 
                           DP_OP_751_130_6421_n1377, S => 
                           DP_OP_751_130_6421_n1378);
   DP_OP_751_130_6421_U1026 : FA_X1 port map( A => DP_OP_751_130_6421_n1475, B 
                           => DP_OP_751_130_6421_n1417, CI => 
                           DP_OP_751_130_6421_n1474, CO => 
                           DP_OP_751_130_6421_n1375, S => 
                           DP_OP_751_130_6421_n1376);
   DP_OP_751_130_6421_U1025 : FA_X1 port map( A => DP_OP_751_130_6421_n1473, B 
                           => DP_OP_751_130_6421_n1416, CI => 
                           DP_OP_751_130_6421_n1472, CO => 
                           DP_OP_751_130_6421_n1373, S => 
                           DP_OP_751_130_6421_n1374);
   DP_OP_751_130_6421_U1024 : FA_X1 port map( A => DP_OP_751_130_6421_n1471, B 
                           => DP_OP_751_130_6421_n1415, CI => 
                           DP_OP_751_130_6421_n1470, CO => 
                           DP_OP_751_130_6421_n1371, S => 
                           DP_OP_751_130_6421_n1372);
   DP_OP_751_130_6421_U1023 : FA_X1 port map( A => DP_OP_751_130_6421_n1469, B 
                           => DP_OP_751_130_6421_n1414, CI => 
                           DP_OP_751_130_6421_n1468, CO => 
                           DP_OP_751_130_6421_n1369, S => 
                           DP_OP_751_130_6421_n1370);
   DP_OP_751_130_6421_U1022 : FA_X1 port map( A => DP_OP_751_130_6421_n1467, B 
                           => DP_OP_751_130_6421_n1413, CI => 
                           DP_OP_751_130_6421_n1466, CO => 
                           DP_OP_751_130_6421_n1367, S => 
                           DP_OP_751_130_6421_n1368);
   DP_OP_751_130_6421_U1021 : FA_X1 port map( A => DP_OP_751_130_6421_n1465, B 
                           => DP_OP_751_130_6421_n1412, CI => 
                           DP_OP_751_130_6421_n1464, CO => 
                           DP_OP_751_130_6421_n1365, S => 
                           DP_OP_751_130_6421_n1366);
   DP_OP_751_130_6421_U1020 : FA_X1 port map( A => DP_OP_751_130_6421_n1463, B 
                           => DP_OP_751_130_6421_n1411, CI => 
                           DP_OP_751_130_6421_n1462, CO => 
                           DP_OP_751_130_6421_n1363, S => 
                           DP_OP_751_130_6421_n1364);
   DP_OP_751_130_6421_U1016 : FA_X1 port map( A => DP_OP_751_130_6421_n1455, B 
                           => DP_OP_751_130_6421_n1407, CI => 
                           DP_OP_751_130_6421_n1454, CO => 
                           DP_OP_751_130_6421_n1355, S => 
                           DP_OP_751_130_6421_n1356);
   DP_OP_751_130_6421_U1013 : FA_X1 port map( A => DP_OP_751_130_6421_n1449, B 
                           => DP_OP_751_130_6421_n1404, CI => 
                           DP_OP_751_130_6421_n1448, CO => 
                           DP_OP_751_130_6421_n1349, S => 
                           DP_OP_751_130_6421_n1350);
   DP_OP_751_130_6421_U1011 : FA_X1 port map( A => DP_OP_751_130_6421_n1445, B 
                           => DP_OP_751_130_6421_n1402, CI => 
                           DP_OP_751_130_6421_n1444, CO => 
                           DP_OP_751_130_6421_n1345, S => 
                           DP_OP_751_130_6421_n1346);
   DP_OP_751_130_6421_U1010 : FA_X1 port map( A => DP_OP_751_130_6421_n1443, B 
                           => DP_OP_751_130_6421_n1401, CI => 
                           DP_OP_751_130_6421_n1442, CO => n_3877, S => 
                           DP_OP_751_130_6421_n1344);
   DP_OP_751_130_6421_U962 : FA_X1 port map( A => DP_OP_751_130_6421_n1385, B 
                           => DP_OP_751_130_6421_n1321, CI => 
                           DP_OP_751_130_6421_n1384, CO => 
                           DP_OP_751_130_6421_n1285, S => 
                           DP_OP_751_130_6421_n1286);
   DP_OP_751_130_6421_U961 : FA_X1 port map( A => DP_OP_751_130_6421_n1383, B 
                           => DP_OP_751_130_6421_n1320, CI => 
                           DP_OP_751_130_6421_n1382, CO => 
                           DP_OP_751_130_6421_n1283, S => 
                           DP_OP_751_130_6421_n1284);
   DP_OP_751_130_6421_U960 : FA_X1 port map( A => DP_OP_751_130_6421_n1381, B 
                           => DP_OP_751_130_6421_n1319, CI => 
                           DP_OP_751_130_6421_n1380, CO => 
                           DP_OP_751_130_6421_n1281, S => 
                           DP_OP_751_130_6421_n1282);
   DP_OP_751_130_6421_U959 : FA_X1 port map( A => DP_OP_751_130_6421_n1379, B 
                           => DP_OP_751_130_6421_n1318, CI => 
                           DP_OP_751_130_6421_n1378, CO => 
                           DP_OP_751_130_6421_n1279, S => 
                           DP_OP_751_130_6421_n1280);
   DP_OP_751_130_6421_U958 : FA_X1 port map( A => DP_OP_751_130_6421_n1377, B 
                           => DP_OP_751_130_6421_n1317, CI => 
                           DP_OP_751_130_6421_n1376, CO => 
                           DP_OP_751_130_6421_n1277, S => 
                           DP_OP_751_130_6421_n1278);
   DP_OP_751_130_6421_U957 : FA_X1 port map( A => DP_OP_751_130_6421_n1375, B 
                           => DP_OP_751_130_6421_n1316, CI => 
                           DP_OP_751_130_6421_n1374, CO => 
                           DP_OP_751_130_6421_n1275, S => 
                           DP_OP_751_130_6421_n1276);
   DP_OP_751_130_6421_U956 : FA_X1 port map( A => DP_OP_751_130_6421_n1373, B 
                           => DP_OP_751_130_6421_n1315, CI => 
                           DP_OP_751_130_6421_n1372, CO => 
                           DP_OP_751_130_6421_n1273, S => 
                           DP_OP_751_130_6421_n1274);
   DP_OP_751_130_6421_U955 : FA_X1 port map( A => DP_OP_751_130_6421_n1371, B 
                           => DP_OP_751_130_6421_n1314, CI => 
                           DP_OP_751_130_6421_n1370, CO => 
                           DP_OP_751_130_6421_n1271, S => 
                           DP_OP_751_130_6421_n1272);
   DP_OP_751_130_6421_U954 : FA_X1 port map( A => DP_OP_751_130_6421_n1369, B 
                           => DP_OP_751_130_6421_n1313, CI => 
                           DP_OP_751_130_6421_n1368, CO => 
                           DP_OP_751_130_6421_n1269, S => 
                           DP_OP_751_130_6421_n1270);
   DP_OP_751_130_6421_U953 : FA_X1 port map( A => DP_OP_751_130_6421_n1367, B 
                           => DP_OP_751_130_6421_n1312, CI => 
                           DP_OP_751_130_6421_n1366, CO => 
                           DP_OP_751_130_6421_n1267, S => 
                           DP_OP_751_130_6421_n1268);
   DP_OP_751_130_6421_U952 : FA_X1 port map( A => DP_OP_751_130_6421_n1365, B 
                           => DP_OP_751_130_6421_n1311, CI => 
                           DP_OP_751_130_6421_n1364, CO => 
                           DP_OP_751_130_6421_n1265, S => 
                           DP_OP_751_130_6421_n1266);
   DP_OP_751_130_6421_U951 : FA_X1 port map( A => DP_OP_751_130_6421_n1363, B 
                           => DP_OP_751_130_6421_n1310, CI => 
                           DP_OP_751_130_6421_n1362, CO => 
                           DP_OP_751_130_6421_n1263, S => 
                           DP_OP_751_130_6421_n1264);
   DP_OP_751_130_6421_U950 : FA_X1 port map( A => DP_OP_751_130_6421_n1361, B 
                           => DP_OP_751_130_6421_n1309, CI => 
                           DP_OP_751_130_6421_n1360, CO => 
                           DP_OP_751_130_6421_n1261, S => 
                           DP_OP_751_130_6421_n1262);
   DP_OP_751_130_6421_U948 : FA_X1 port map( A => DP_OP_751_130_6421_n1357, B 
                           => DP_OP_751_130_6421_n1307, CI => 
                           DP_OP_751_130_6421_n1356, CO => 
                           DP_OP_751_130_6421_n1257, S => 
                           DP_OP_751_130_6421_n1258);
   DP_OP_751_130_6421_U947 : FA_X1 port map( A => DP_OP_751_130_6421_n1355, B 
                           => DP_OP_751_130_6421_n1306, CI => 
                           DP_OP_751_130_6421_n1354, CO => 
                           DP_OP_751_130_6421_n1255, S => 
                           DP_OP_751_130_6421_n1256);
   DP_OP_751_130_6421_U944 : FA_X1 port map( A => DP_OP_751_130_6421_n1349, B 
                           => DP_OP_751_130_6421_n1303, CI => 
                           DP_OP_751_130_6421_n1348, CO => 
                           DP_OP_751_130_6421_n1249, S => 
                           DP_OP_751_130_6421_n1250);
   DP_OP_751_130_6421_U942 : FA_X1 port map( A => DP_OP_751_130_6421_n1345, B 
                           => DP_OP_751_130_6421_n1301, CI => 
                           DP_OP_751_130_6421_n1344, CO => n_3878, S => 
                           DP_OP_751_130_6421_n1246);
   DP_OP_751_130_6421_U893 : FA_X1 port map( A => DP_OP_751_130_6421_n1220, B 
                           => DP_OP_751_130_6421_n1221, CI => 
                           DP_OP_751_130_6421_n1285, CO => 
                           DP_OP_751_130_6421_n1185, S => 
                           DP_OP_751_130_6421_n1186);
   DP_OP_751_130_6421_U892 : FA_X1 port map( A => DP_OP_751_130_6421_n1283, B 
                           => DP_OP_751_130_6421_n1219, CI => 
                           DP_OP_751_130_6421_n1282, CO => 
                           DP_OP_751_130_6421_n1183, S => 
                           DP_OP_751_130_6421_n1184);
   DP_OP_751_130_6421_U890 : FA_X1 port map( A => DP_OP_751_130_6421_n1279, B 
                           => DP_OP_751_130_6421_n1217, CI => 
                           DP_OP_751_130_6421_n1278, CO => 
                           DP_OP_751_130_6421_n1179, S => 
                           DP_OP_751_130_6421_n1180);
   DP_OP_751_130_6421_U889 : FA_X1 port map( A => DP_OP_751_130_6421_n1277, B 
                           => DP_OP_751_130_6421_n1216, CI => 
                           DP_OP_751_130_6421_n1276, CO => 
                           DP_OP_751_130_6421_n1177, S => 
                           DP_OP_751_130_6421_n1178);
   DP_OP_751_130_6421_U888 : FA_X1 port map( A => DP_OP_751_130_6421_n1275, B 
                           => DP_OP_751_130_6421_n1215, CI => 
                           DP_OP_751_130_6421_n1274, CO => 
                           DP_OP_751_130_6421_n1175, S => 
                           DP_OP_751_130_6421_n1176);
   DP_OP_751_130_6421_U887 : FA_X1 port map( A => DP_OP_751_130_6421_n1273, B 
                           => DP_OP_751_130_6421_n1214, CI => 
                           DP_OP_751_130_6421_n1272, CO => 
                           DP_OP_751_130_6421_n1173, S => 
                           DP_OP_751_130_6421_n1174);
   DP_OP_751_130_6421_U886 : FA_X1 port map( A => DP_OP_751_130_6421_n1271, B 
                           => DP_OP_751_130_6421_n1213, CI => 
                           DP_OP_751_130_6421_n1270, CO => 
                           DP_OP_751_130_6421_n1171, S => 
                           DP_OP_751_130_6421_n1172);
   DP_OP_751_130_6421_U885 : FA_X1 port map( A => DP_OP_751_130_6421_n1269, B 
                           => DP_OP_751_130_6421_n1212, CI => 
                           DP_OP_751_130_6421_n1268, CO => 
                           DP_OP_751_130_6421_n1169, S => 
                           DP_OP_751_130_6421_n1170);
   DP_OP_751_130_6421_U884 : FA_X1 port map( A => DP_OP_751_130_6421_n1267, B 
                           => DP_OP_751_130_6421_n1211, CI => 
                           DP_OP_751_130_6421_n1266, CO => 
                           DP_OP_751_130_6421_n1167, S => 
                           DP_OP_751_130_6421_n1168);
   DP_OP_751_130_6421_U882 : FA_X1 port map( A => DP_OP_751_130_6421_n1263, B 
                           => DP_OP_751_130_6421_n1209, CI => 
                           DP_OP_751_130_6421_n1262, CO => 
                           DP_OP_751_130_6421_n1163, S => 
                           DP_OP_751_130_6421_n1164);
   DP_OP_751_130_6421_U880 : FA_X1 port map( A => DP_OP_751_130_6421_n1259, B 
                           => DP_OP_751_130_6421_n1207, CI => 
                           DP_OP_751_130_6421_n1258, CO => 
                           DP_OP_751_130_6421_n1159, S => 
                           DP_OP_751_130_6421_n1160);
   DP_OP_751_130_6421_U879 : FA_X1 port map( A => DP_OP_751_130_6421_n1257, B 
                           => DP_OP_751_130_6421_n1206, CI => 
                           DP_OP_751_130_6421_n1256, CO => 
                           DP_OP_751_130_6421_n1157, S => 
                           DP_OP_751_130_6421_n1158);
   DP_OP_751_130_6421_U877 : FA_X1 port map( A => DP_OP_751_130_6421_n1253, B 
                           => DP_OP_751_130_6421_n1204, CI => 
                           DP_OP_751_130_6421_n1252, CO => 
                           DP_OP_751_130_6421_n1153, S => 
                           DP_OP_751_130_6421_n1154);
   DP_OP_751_130_6421_U876 : FA_X1 port map( A => DP_OP_751_130_6421_n1251, B 
                           => DP_OP_751_130_6421_n1203, CI => 
                           DP_OP_751_130_6421_n1250, CO => 
                           DP_OP_751_130_6421_n1151, S => 
                           DP_OP_751_130_6421_n1152);
   DP_OP_751_130_6421_U875 : FA_X1 port map( A => DP_OP_751_130_6421_n1249, B 
                           => DP_OP_751_130_6421_n1202, CI => 
                           DP_OP_751_130_6421_n1248, CO => 
                           DP_OP_751_130_6421_n1149, S => 
                           DP_OP_751_130_6421_n1150);
   DP_OP_751_130_6421_U874 : FA_X1 port map( A => DP_OP_751_130_6421_n1247, B 
                           => DP_OP_751_130_6421_n1201, CI => 
                           DP_OP_751_130_6421_n1246, CO => n_3879, S => 
                           DP_OP_751_130_6421_n1148);
   DP_OP_751_130_6421_U823 : FA_X1 port map( A => DP_OP_751_130_6421_n1118, B 
                           => n7793, CI => DP_OP_751_130_6421_n1183, CO => 
                           DP_OP_751_130_6421_n1083, S => 
                           DP_OP_751_130_6421_n1084);
   DP_OP_751_130_6421_U822 : FA_X1 port map( A => DP_OP_751_130_6421_n1181, B 
                           => DP_OP_751_130_6421_n1117, CI => 
                           DP_OP_751_130_6421_n1180, CO => 
                           DP_OP_751_130_6421_n1081, S => 
                           DP_OP_751_130_6421_n1082);
   DP_OP_751_130_6421_U821 : FA_X1 port map( A => DP_OP_751_130_6421_n1179, B 
                           => DP_OP_751_130_6421_n1116, CI => 
                           DP_OP_751_130_6421_n1178, CO => 
                           DP_OP_751_130_6421_n1079, S => 
                           DP_OP_751_130_6421_n1080);
   DP_OP_751_130_6421_U820 : FA_X1 port map( A => DP_OP_751_130_6421_n1177, B 
                           => DP_OP_751_130_6421_n1115, CI => 
                           DP_OP_751_130_6421_n1176, CO => 
                           DP_OP_751_130_6421_n1077, S => 
                           DP_OP_751_130_6421_n1078);
   DP_OP_751_130_6421_U819 : FA_X1 port map( A => DP_OP_751_130_6421_n1175, B 
                           => DP_OP_751_130_6421_n1114, CI => 
                           DP_OP_751_130_6421_n1174, CO => 
                           DP_OP_751_130_6421_n1075, S => 
                           DP_OP_751_130_6421_n1076);
   DP_OP_751_130_6421_U818 : FA_X1 port map( A => DP_OP_751_130_6421_n1173, B 
                           => DP_OP_751_130_6421_n1113, CI => 
                           DP_OP_751_130_6421_n1172, CO => 
                           DP_OP_751_130_6421_n1073, S => 
                           DP_OP_751_130_6421_n1074);
   DP_OP_751_130_6421_U817 : FA_X1 port map( A => DP_OP_751_130_6421_n1171, B 
                           => DP_OP_751_130_6421_n1112, CI => 
                           DP_OP_751_130_6421_n1170, CO => 
                           DP_OP_751_130_6421_n1071, S => 
                           DP_OP_751_130_6421_n1072);
   DP_OP_751_130_6421_U816 : FA_X1 port map( A => DP_OP_751_130_6421_n1169, B 
                           => DP_OP_751_130_6421_n1111, CI => 
                           DP_OP_751_130_6421_n1168, CO => 
                           DP_OP_751_130_6421_n1069, S => 
                           DP_OP_751_130_6421_n1070);
   DP_OP_751_130_6421_U814 : FA_X1 port map( A => DP_OP_751_130_6421_n1165, B 
                           => DP_OP_751_130_6421_n1109, CI => 
                           DP_OP_751_130_6421_n1164, CO => 
                           DP_OP_751_130_6421_n1065, S => 
                           DP_OP_751_130_6421_n1066);
   DP_OP_751_130_6421_U812 : FA_X1 port map( A => DP_OP_751_130_6421_n1161, B 
                           => DP_OP_751_130_6421_n1107, CI => 
                           DP_OP_751_130_6421_n1160, CO => 
                           DP_OP_751_130_6421_n1061, S => 
                           DP_OP_751_130_6421_n1062);
   DP_OP_751_130_6421_U811 : FA_X1 port map( A => DP_OP_751_130_6421_n1159, B 
                           => DP_OP_751_130_6421_n1106, CI => 
                           DP_OP_751_130_6421_n1158, CO => 
                           DP_OP_751_130_6421_n1059, S => 
                           DP_OP_751_130_6421_n1060);
   DP_OP_751_130_6421_U810 : FA_X1 port map( A => DP_OP_751_130_6421_n1157, B 
                           => DP_OP_751_130_6421_n1105, CI => 
                           DP_OP_751_130_6421_n1156, CO => 
                           DP_OP_751_130_6421_n1057, S => 
                           DP_OP_751_130_6421_n1058);
   DP_OP_751_130_6421_U808 : FA_X1 port map( A => DP_OP_751_130_6421_n1153, B 
                           => DP_OP_751_130_6421_n1103, CI => 
                           DP_OP_751_130_6421_n1152, CO => 
                           DP_OP_751_130_6421_n1053, S => 
                           DP_OP_751_130_6421_n1054);
   DP_OP_751_130_6421_U807 : FA_X1 port map( A => DP_OP_751_130_6421_n1151, B 
                           => DP_OP_751_130_6421_n1102, CI => 
                           DP_OP_751_130_6421_n1150, CO => 
                           DP_OP_751_130_6421_n1051, S => 
                           DP_OP_751_130_6421_n1052);
   DP_OP_751_130_6421_U806 : FA_X1 port map( A => DP_OP_751_130_6421_n1149, B 
                           => DP_OP_751_130_6421_n1101, CI => 
                           DP_OP_751_130_6421_n1148, CO => n_3880, S => 
                           DP_OP_751_130_6421_n1050);
   DP_OP_751_130_6421_U752 : FA_X1 port map( A => DP_OP_751_130_6421_n1079, B 
                           => DP_OP_751_130_6421_n1015, CI => 
                           DP_OP_751_130_6421_n1078, CO => 
                           DP_OP_751_130_6421_n979, S => 
                           DP_OP_751_130_6421_n980);
   DP_OP_751_130_6421_U751 : FA_X1 port map( A => DP_OP_751_130_6421_n1077, B 
                           => DP_OP_751_130_6421_n1014, CI => 
                           DP_OP_751_130_6421_n1076, CO => 
                           DP_OP_751_130_6421_n977, S => 
                           DP_OP_751_130_6421_n978);
   DP_OP_751_130_6421_U750 : FA_X1 port map( A => DP_OP_751_130_6421_n1075, B 
                           => DP_OP_751_130_6421_n1013, CI => 
                           DP_OP_751_130_6421_n1074, CO => 
                           DP_OP_751_130_6421_n975, S => 
                           DP_OP_751_130_6421_n976);
   DP_OP_751_130_6421_U749 : FA_X1 port map( A => DP_OP_751_130_6421_n1073, B 
                           => DP_OP_751_130_6421_n1012, CI => 
                           DP_OP_751_130_6421_n1072, CO => 
                           DP_OP_751_130_6421_n973, S => 
                           DP_OP_751_130_6421_n974);
   DP_OP_751_130_6421_U748 : FA_X1 port map( A => DP_OP_751_130_6421_n1071, B 
                           => DP_OP_751_130_6421_n1011, CI => 
                           DP_OP_751_130_6421_n1070, CO => 
                           DP_OP_751_130_6421_n971, S => 
                           DP_OP_751_130_6421_n972);
   DP_OP_751_130_6421_U747 : FA_X1 port map( A => DP_OP_751_130_6421_n1069, B 
                           => DP_OP_751_130_6421_n1010, CI => 
                           DP_OP_751_130_6421_n1068, CO => 
                           DP_OP_751_130_6421_n969, S => 
                           DP_OP_751_130_6421_n970);
   DP_OP_751_130_6421_U746 : FA_X1 port map( A => DP_OP_751_130_6421_n1067, B 
                           => DP_OP_751_130_6421_n1009, CI => 
                           DP_OP_751_130_6421_n1066, CO => 
                           DP_OP_751_130_6421_n967, S => 
                           DP_OP_751_130_6421_n968);
   DP_OP_751_130_6421_U744 : FA_X1 port map( A => DP_OP_751_130_6421_n1063, B 
                           => DP_OP_751_130_6421_n1007, CI => 
                           DP_OP_751_130_6421_n1062, CO => 
                           DP_OP_751_130_6421_n963, S => 
                           DP_OP_751_130_6421_n964);
   DP_OP_751_130_6421_U743 : FA_X1 port map( A => DP_OP_751_130_6421_n1061, B 
                           => DP_OP_751_130_6421_n1006, CI => 
                           DP_OP_751_130_6421_n1060, CO => 
                           DP_OP_751_130_6421_n961, S => 
                           DP_OP_751_130_6421_n962);
   DP_OP_751_130_6421_U742 : FA_X1 port map( A => DP_OP_751_130_6421_n1059, B 
                           => DP_OP_751_130_6421_n1005, CI => 
                           DP_OP_751_130_6421_n1058, CO => 
                           DP_OP_751_130_6421_n959, S => 
                           DP_OP_751_130_6421_n960);
   DP_OP_751_130_6421_U741 : FA_X1 port map( A => DP_OP_751_130_6421_n1057, B 
                           => DP_OP_751_130_6421_n1004, CI => 
                           DP_OP_751_130_6421_n1056, CO => 
                           DP_OP_751_130_6421_n957, S => 
                           DP_OP_751_130_6421_n958);
   DP_OP_751_130_6421_U738 : FA_X1 port map( A => DP_OP_751_130_6421_n1051, B 
                           => DP_OP_751_130_6421_n1001, CI => 
                           DP_OP_751_130_6421_n1050, CO => n_3881, S => 
                           DP_OP_751_130_6421_n952);
   DP_OP_751_130_6421_U682 : FA_X1 port map( A => DP_OP_751_130_6421_n977, B =>
                           DP_OP_751_130_6421_n913, CI => 
                           DP_OP_751_130_6421_n976, CO => 
                           DP_OP_751_130_6421_n877, S => 
                           DP_OP_751_130_6421_n878);
   DP_OP_751_130_6421_U681 : FA_X1 port map( A => DP_OP_751_130_6421_n975, B =>
                           DP_OP_751_130_6421_n912, CI => 
                           DP_OP_751_130_6421_n974, CO => 
                           DP_OP_751_130_6421_n875, S => 
                           DP_OP_751_130_6421_n876);
   DP_OP_751_130_6421_U680 : FA_X1 port map( A => DP_OP_751_130_6421_n973, B =>
                           DP_OP_751_130_6421_n911, CI => 
                           DP_OP_751_130_6421_n972, CO => 
                           DP_OP_751_130_6421_n873, S => 
                           DP_OP_751_130_6421_n874);
   DP_OP_751_130_6421_U679 : FA_X1 port map( A => DP_OP_751_130_6421_n971, B =>
                           DP_OP_751_130_6421_n910, CI => 
                           DP_OP_751_130_6421_n970, CO => 
                           DP_OP_751_130_6421_n871, S => 
                           DP_OP_751_130_6421_n872);
   DP_OP_751_130_6421_U677 : FA_X1 port map( A => DP_OP_751_130_6421_n967, B =>
                           DP_OP_751_130_6421_n908, CI => 
                           DP_OP_751_130_6421_n966, CO => 
                           DP_OP_751_130_6421_n867, S => 
                           DP_OP_751_130_6421_n868);
   DP_OP_751_130_6421_U676 : FA_X1 port map( A => DP_OP_751_130_6421_n965, B =>
                           DP_OP_751_130_6421_n907, CI => 
                           DP_OP_751_130_6421_n964, CO => 
                           DP_OP_751_130_6421_n865, S => 
                           DP_OP_751_130_6421_n866);
   DP_OP_751_130_6421_U675 : FA_X1 port map( A => DP_OP_751_130_6421_n963, B =>
                           DP_OP_751_130_6421_n906, CI => 
                           DP_OP_751_130_6421_n962, CO => 
                           DP_OP_751_130_6421_n863, S => 
                           DP_OP_751_130_6421_n864);
   DP_OP_751_130_6421_U674 : FA_X1 port map( A => DP_OP_751_130_6421_n961, B =>
                           DP_OP_751_130_6421_n905, CI => 
                           DP_OP_751_130_6421_n960, CO => 
                           DP_OP_751_130_6421_n861, S => 
                           DP_OP_751_130_6421_n862);
   DP_OP_751_130_6421_U673 : FA_X1 port map( A => DP_OP_751_130_6421_n959, B =>
                           DP_OP_751_130_6421_n904, CI => 
                           DP_OP_751_130_6421_n958, CO => 
                           DP_OP_751_130_6421_n859, S => 
                           DP_OP_751_130_6421_n860);
   DP_OP_751_130_6421_U672 : FA_X1 port map( A => DP_OP_751_130_6421_n957, B =>
                           DP_OP_751_130_6421_n903, CI => 
                           DP_OP_751_130_6421_n956, CO => 
                           DP_OP_751_130_6421_n857, S => 
                           DP_OP_751_130_6421_n858);
   DP_OP_751_130_6421_U670 : FA_X1 port map( A => DP_OP_751_130_6421_n953, B =>
                           DP_OP_751_130_6421_n901, CI => 
                           DP_OP_751_130_6421_n952, CO => n_3882, S => 
                           DP_OP_751_130_6421_n854);
   DP_OP_751_130_6421_U612 : FA_X1 port map( A => DP_OP_751_130_6421_n875, B =>
                           DP_OP_751_130_6421_n811, CI => 
                           DP_OP_751_130_6421_n874, CO => 
                           DP_OP_751_130_6421_n775, S => 
                           DP_OP_751_130_6421_n776);
   DP_OP_751_130_6421_U611 : FA_X1 port map( A => DP_OP_751_130_6421_n873, B =>
                           DP_OP_751_130_6421_n810, CI => 
                           DP_OP_751_130_6421_n872, CO => 
                           DP_OP_751_130_6421_n773, S => 
                           DP_OP_751_130_6421_n774);
   DP_OP_751_130_6421_U609 : FA_X1 port map( A => DP_OP_751_130_6421_n869, B =>
                           DP_OP_751_130_6421_n808, CI => 
                           DP_OP_751_130_6421_n868, CO => 
                           DP_OP_751_130_6421_n769, S => 
                           DP_OP_751_130_6421_n770);
   DP_OP_751_130_6421_U608 : FA_X1 port map( A => DP_OP_751_130_6421_n867, B =>
                           DP_OP_751_130_6421_n807, CI => 
                           DP_OP_751_130_6421_n866, CO => 
                           DP_OP_751_130_6421_n767, S => 
                           DP_OP_751_130_6421_n768);
   DP_OP_751_130_6421_U607 : FA_X1 port map( A => DP_OP_751_130_6421_n865, B =>
                           DP_OP_751_130_6421_n806, CI => 
                           DP_OP_751_130_6421_n864, CO => 
                           DP_OP_751_130_6421_n765, S => 
                           DP_OP_751_130_6421_n766);
   DP_OP_751_130_6421_U606 : FA_X1 port map( A => DP_OP_751_130_6421_n863, B =>
                           DP_OP_751_130_6421_n805, CI => 
                           DP_OP_751_130_6421_n862, CO => 
                           DP_OP_751_130_6421_n763, S => 
                           DP_OP_751_130_6421_n764);
   DP_OP_751_130_6421_U605 : FA_X1 port map( A => DP_OP_751_130_6421_n861, B =>
                           DP_OP_751_130_6421_n804, CI => 
                           DP_OP_751_130_6421_n860, CO => 
                           DP_OP_751_130_6421_n761, S => 
                           DP_OP_751_130_6421_n762);
   DP_OP_751_130_6421_U604 : FA_X1 port map( A => DP_OP_751_130_6421_n859, B =>
                           DP_OP_751_130_6421_n803, CI => 
                           DP_OP_751_130_6421_n858, CO => 
                           DP_OP_751_130_6421_n759, S => 
                           DP_OP_751_130_6421_n760);
   DP_OP_751_130_6421_U602 : FA_X1 port map( A => DP_OP_751_130_6421_n855, B =>
                           DP_OP_751_130_6421_n801, CI => 
                           DP_OP_751_130_6421_n854, CO => n_3883, S => 
                           DP_OP_751_130_6421_n756);
   DP_OP_751_130_6421_U542 : FA_X1 port map( A => DP_OP_751_130_6421_n773, B =>
                           DP_OP_751_130_6421_n709, CI => 
                           DP_OP_751_130_6421_n772, CO => 
                           DP_OP_751_130_6421_n673, S => 
                           DP_OP_751_130_6421_n674);
   DP_OP_751_130_6421_U541 : FA_X1 port map( A => DP_OP_751_130_6421_n771, B =>
                           DP_OP_751_130_6421_n708, CI => 
                           DP_OP_751_130_6421_n770, CO => 
                           DP_OP_751_130_6421_n671, S => 
                           DP_OP_751_130_6421_n672);
   DP_OP_751_130_6421_U539 : FA_X1 port map( A => DP_OP_751_130_6421_n767, B =>
                           DP_OP_751_130_6421_n706, CI => 
                           DP_OP_751_130_6421_n766, CO => 
                           DP_OP_751_130_6421_n667, S => 
                           DP_OP_751_130_6421_n668);
   DP_OP_751_130_6421_U538 : FA_X1 port map( A => DP_OP_751_130_6421_n765, B =>
                           DP_OP_751_130_6421_n705, CI => 
                           DP_OP_751_130_6421_n764, CO => 
                           DP_OP_751_130_6421_n665, S => 
                           DP_OP_751_130_6421_n666);
   DP_OP_751_130_6421_U537 : FA_X1 port map( A => DP_OP_751_130_6421_n763, B =>
                           DP_OP_751_130_6421_n704, CI => 
                           DP_OP_751_130_6421_n762, CO => 
                           DP_OP_751_130_6421_n663, S => 
                           DP_OP_751_130_6421_n664);
   DP_OP_751_130_6421_U536 : FA_X1 port map( A => DP_OP_751_130_6421_n761, B =>
                           DP_OP_751_130_6421_n703, CI => 
                           DP_OP_751_130_6421_n760, CO => 
                           DP_OP_751_130_6421_n661, S => 
                           DP_OP_751_130_6421_n662);
   DP_OP_751_130_6421_U535 : FA_X1 port map( A => DP_OP_751_130_6421_n759, B =>
                           DP_OP_751_130_6421_n702, CI => 
                           DP_OP_751_130_6421_n758, CO => 
                           DP_OP_751_130_6421_n659, S => 
                           DP_OP_751_130_6421_n660);
   DP_OP_751_130_6421_U534 : FA_X1 port map( A => DP_OP_751_130_6421_n757, B =>
                           DP_OP_751_130_6421_n701, CI => 
                           DP_OP_751_130_6421_n756, CO => n_3884, S => 
                           DP_OP_751_130_6421_n658);
   DP_OP_751_130_6421_U472 : FA_X1 port map( A => DP_OP_751_130_6421_n671, B =>
                           DP_OP_751_130_6421_n607, CI => 
                           DP_OP_751_130_6421_n670, CO => 
                           DP_OP_751_130_6421_n571, S => 
                           DP_OP_751_130_6421_n572);
   DP_OP_751_130_6421_U471 : FA_X1 port map( A => DP_OP_751_130_6421_n669, B =>
                           DP_OP_751_130_6421_n606, CI => 
                           DP_OP_751_130_6421_n668, CO => 
                           DP_OP_751_130_6421_n569, S => 
                           DP_OP_751_130_6421_n570);
   DP_OP_751_130_6421_U470 : FA_X1 port map( A => DP_OP_751_130_6421_n667, B =>
                           DP_OP_751_130_6421_n605, CI => 
                           DP_OP_751_130_6421_n666, CO => 
                           DP_OP_751_130_6421_n567, S => 
                           DP_OP_751_130_6421_n568);
   DP_OP_751_130_6421_U469 : FA_X1 port map( A => DP_OP_751_130_6421_n665, B =>
                           DP_OP_751_130_6421_n604, CI => 
                           DP_OP_751_130_6421_n664, CO => 
                           DP_OP_751_130_6421_n565, S => 
                           DP_OP_751_130_6421_n566);
   DP_OP_751_130_6421_U468 : FA_X1 port map( A => DP_OP_751_130_6421_n663, B =>
                           DP_OP_751_130_6421_n603, CI => 
                           DP_OP_751_130_6421_n662, CO => 
                           DP_OP_751_130_6421_n563, S => 
                           DP_OP_751_130_6421_n564);
   DP_OP_751_130_6421_U467 : FA_X1 port map( A => DP_OP_751_130_6421_n661, B =>
                           DP_OP_751_130_6421_n602, CI => 
                           DP_OP_751_130_6421_n660, CO => 
                           DP_OP_751_130_6421_n561, S => 
                           DP_OP_751_130_6421_n562);
   DP_OP_751_130_6421_U466 : FA_X1 port map( A => DP_OP_751_130_6421_n659, B =>
                           DP_OP_751_130_6421_n601, CI => 
                           DP_OP_751_130_6421_n658, CO => n_3885, S => 
                           DP_OP_751_130_6421_n560);
   DP_OP_751_130_6421_U402 : FA_X1 port map( A => DP_OP_751_130_6421_n505, B =>
                           DP_OP_751_130_6421_n569, CI => 
                           DP_OP_751_130_6421_n568, CO => 
                           DP_OP_751_130_6421_n469, S => 
                           DP_OP_751_130_6421_n470);
   DP_OP_751_130_6421_U401 : FA_X1 port map( A => DP_OP_751_130_6421_n567, B =>
                           DP_OP_751_130_6421_n504, CI => 
                           DP_OP_751_130_6421_n566, CO => 
                           DP_OP_751_130_6421_n467, S => 
                           DP_OP_751_130_6421_n468);
   DP_OP_751_130_6421_U399 : FA_X1 port map( A => DP_OP_751_130_6421_n563, B =>
                           DP_OP_751_130_6421_n502, CI => 
                           DP_OP_751_130_6421_n562, CO => 
                           DP_OP_751_130_6421_n463, S => 
                           DP_OP_751_130_6421_n464);
   DP_OP_751_130_6421_U398 : FA_X1 port map( A => DP_OP_751_130_6421_n561, B =>
                           DP_OP_751_130_6421_n501, CI => 
                           DP_OP_751_130_6421_n560, CO => n_3886, S => 
                           DP_OP_751_130_6421_n462);
   DP_OP_751_130_6421_U331 : FA_X1 port map( A => DP_OP_751_130_6421_n465, B =>
                           DP_OP_751_130_6421_n402, CI => 
                           DP_OP_751_130_6421_n464, CO => 
                           DP_OP_751_130_6421_n365, S => 
                           DP_OP_751_130_6421_n366);
   IR_reg_26_inst : DFFS_X1 port map( D => n7123, CK => CLK, SN => n8579, Q => 
                           IR_26_port, QN => n8223);
   DataPath_REG_ALU_OUT_Q_reg_31_inst : DFF_X1 port map( D => n6992, CK => CLK,
                           Q => DRAM_ADDRESS_31_port, QN => n515);
   intadd_0_U21 : NAND2_X1 port map( A1 => intadd_0_B_1_port, A2 => 
                           IRAM_ADDRESS_2_port, ZN => intadd_0_n15);
   intadd_0_U20 : NOR2_X1 port map( A1 => intadd_0_B_1_port, A2 => 
                           IRAM_ADDRESS_2_port, ZN => intadd_0_n14);
   CU_I_CW_EX_reg_MUXB_SEL_inst : DFF_X1 port map( D => n7086, CK => CLK, Q => 
                           n8193, QN => n8221);
   DataPath_WRF_CUhw_curr_addr_reg_2_inst : DFF_X1 port map( D => n7649, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_2_port, QN => 
                           n_3887);
   DataPath_WRF_CUhw_curr_addr_reg_3_inst : DFF_X1 port map( D => n7648, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_3_port, QN => 
                           n8129);
   DataPath_WRF_CUhw_curr_addr_reg_4_inst : DFF_X1 port map( D => n7647, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_4_port, QN => 
                           n_3888);
   DataPath_WRF_CUhw_curr_addr_reg_5_inst : DFF_X1 port map( D => n7646, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_5_port, QN => 
                           n_3889);
   DataPath_WRF_CUhw_curr_addr_reg_6_inst : DFF_X1 port map( D => n7645, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_6_port, QN => 
                           n_3890);
   DataPath_WRF_CUhw_curr_addr_reg_7_inst : DFF_X1 port map( D => n7644, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_7_port, QN => 
                           n_3891);
   DataPath_WRF_CUhw_curr_addr_reg_8_inst : DFF_X1 port map( D => n7643, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_8_port, QN => 
                           n_3892);
   DataPath_WRF_CUhw_curr_addr_reg_10_inst : DFF_X1 port map( D => n7642, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_10_port, QN =>
                           n_3893);
   DataPath_WRF_CUhw_curr_addr_reg_9_inst : DFF_X1 port map( D => n7641, CK => 
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_9_port, QN => 
                           n_3894);
   DataPath_WRF_CUhw_curr_addr_reg_11_inst : DFF_X1 port map( D => n7640, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_11_port, QN =>
                           n_3895);
   DataPath_WRF_CUhw_curr_addr_reg_12_inst : DFF_X1 port map( D => n7639, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_12_port, QN =>
                           n_3896);
   DataPath_WRF_CUhw_curr_addr_reg_13_inst : DFF_X1 port map( D => n7638, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_13_port, QN =>
                           n_3897);
   DataPath_WRF_CUhw_curr_addr_reg_14_inst : DFF_X1 port map( D => n7637, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_14_port, QN =>
                           n_3898);
   DataPath_WRF_CUhw_curr_addr_reg_15_inst : DFF_X1 port map( D => n7636, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_15_port, QN =>
                           n_3899);
   DataPath_WRF_CUhw_curr_addr_reg_16_inst : DFF_X1 port map( D => n7635, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_16_port, QN =>
                           n_3900);
   DataPath_WRF_CUhw_curr_addr_reg_17_inst : DFF_X1 port map( D => n7634, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_17_port, QN =>
                           n_3901);
   DataPath_WRF_CUhw_curr_addr_reg_18_inst : DFF_X1 port map( D => n7633, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_18_port, QN =>
                           n_3902);
   DataPath_WRF_CUhw_curr_addr_reg_19_inst : DFF_X1 port map( D => n7632, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_19_port, QN =>
                           n_3903);
   DataPath_WRF_CUhw_curr_addr_reg_20_inst : DFF_X1 port map( D => n7631, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_20_port, QN =>
                           n_3904);
   DataPath_WRF_CUhw_curr_addr_reg_21_inst : DFF_X1 port map( D => n7630, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_21_port, QN =>
                           n_3905);
   DataPath_WRF_CUhw_curr_addr_reg_22_inst : DFF_X1 port map( D => n7629, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_22_port, QN =>
                           n_3906);
   DataPath_WRF_CUhw_curr_addr_reg_23_inst : DFF_X1 port map( D => n7628, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_23_port, QN =>
                           n_3907);
   DataPath_WRF_CUhw_curr_addr_reg_24_inst : DFF_X1 port map( D => n7627, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_24_port, QN =>
                           n_3908);
   DataPath_WRF_CUhw_curr_addr_reg_28_inst : DFF_X1 port map( D => n7626, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_28_port, QN =>
                           n8110);
   DataPath_WRF_CUhw_curr_addr_reg_25_inst : DFF_X1 port map( D => n7625, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_25_port, QN =>
                           n_3909);
   DataPath_WRF_CUhw_curr_addr_reg_27_inst : DFF_X1 port map( D => n7624, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_27_port, QN =>
                           n_3910);
   DataPath_WRF_CUhw_curr_addr_reg_26_inst : DFF_X1 port map( D => n7623, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_26_port, QN =>
                           n_3911);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_0_inst : DFF_X1 port map( D => 
                           n7165, CK => CLK, Q => n_3912, QN => n541);
   DataPath_WRF_CUhw_curr_data_reg_22_inst : DFF_X1 port map( D => n3215, CK =>
                           CLK, Q => n_3913, QN => 
                           DataPath_WRF_CUhw_curr_data_22_port);
   DataPath_WRF_CUhw_curr_data_reg_21_inst : DFF_X1 port map( D => n3216, CK =>
                           CLK, Q => n_3914, QN => 
                           DataPath_WRF_CUhw_curr_data_21_port);
   DataPath_WRF_CUhw_curr_data_reg_18_inst : DFF_X1 port map( D => n3219, CK =>
                           CLK, Q => n_3915, QN => 
                           DataPath_WRF_CUhw_curr_data_18_port);
   DataPath_WRF_CUhw_curr_data_reg_14_inst : DFF_X1 port map( D => n3223, CK =>
                           CLK, Q => n_3916, QN => 
                           DataPath_WRF_CUhw_curr_data_14_port);
   DataPath_WRF_CUhw_curr_data_reg_13_inst : DFF_X1 port map( D => n3224, CK =>
                           CLK, Q => n_3917, QN => 
                           DataPath_WRF_CUhw_curr_data_13_port);
   DataPath_WRF_CUhw_curr_data_reg_12_inst : DFF_X1 port map( D => n3225, CK =>
                           CLK, Q => n_3918, QN => 
                           DataPath_WRF_CUhw_curr_data_12_port);
   DataPath_WRF_CUhw_curr_data_reg_11_inst : DFF_X1 port map( D => n3226, CK =>
                           CLK, Q => n_3919, QN => 
                           DataPath_WRF_CUhw_curr_data_11_port);
   DataPath_WRF_CUhw_curr_data_reg_10_inst : DFF_X1 port map( D => n3227, CK =>
                           CLK, Q => n_3920, QN => 
                           DataPath_WRF_CUhw_curr_data_10_port);
   DataPath_WRF_CUhw_curr_data_reg_8_inst : DFF_X1 port map( D => n3229, CK => 
                           CLK, Q => n_3921, QN => 
                           DataPath_WRF_CUhw_curr_data_8_port);
   DataPath_WRF_CUhw_curr_data_reg_6_inst : DFF_X1 port map( D => n3231, CK => 
                           CLK, Q => n_3922, QN => 
                           DataPath_WRF_CUhw_curr_data_6_port);
   DataPath_WRF_CUhw_curr_data_reg_1_inst : DFF_X1 port map( D => n3236, CK => 
                           CLK, Q => n_3923, QN => 
                           DataPath_WRF_CUhw_curr_data_1_port);
   DataPath_WRF_CUhw_curr_data_reg_26_inst : DFF_X1 port map( D => n3211, CK =>
                           CLK, Q => n_3924, QN => 
                           DataPath_WRF_CUhw_curr_data_26_port);
   DataPath_WRF_CUhw_curr_data_reg_7_inst : DFF_X1 port map( D => n3230, CK => 
                           CLK, Q => n_3925, QN => 
                           DataPath_WRF_CUhw_curr_data_7_port);
   DataPath_WRF_CUhw_curr_data_reg_4_inst : DFF_X1 port map( D => n3233, CK => 
                           CLK, Q => n_3926, QN => 
                           DataPath_WRF_CUhw_curr_data_4_port);
   DataPath_WRF_CUhw_curr_data_reg_3_inst : DFF_X1 port map( D => n3234, CK => 
                           CLK, Q => n_3927, QN => 
                           DataPath_WRF_CUhw_curr_data_3_port);
   DataPath_WRF_CUhw_curr_data_reg_2_inst : DFF_X1 port map( D => n3235, CK => 
                           CLK, Q => n_3928, QN => 
                           DataPath_WRF_CUhw_curr_data_2_port);
   DataPath_WRF_CUhw_curr_data_reg_0_inst : DFF_X1 port map( D => n3237, CK => 
                           CLK, Q => n_3929, QN => 
                           DataPath_WRF_CUhw_curr_data_0_port);
   DataPath_WRF_CUhw_curr_data_reg_20_inst : DFF_X1 port map( D => n3217, CK =>
                           CLK, Q => n_3930, QN => 
                           DataPath_WRF_CUhw_curr_data_20_port);
   DataPath_WRF_CUhw_curr_data_reg_29_inst : DFF_X1 port map( D => n3208, CK =>
                           CLK, Q => n_3931, QN => 
                           DataPath_WRF_CUhw_curr_data_29_port);
   DataPath_WRF_CUhw_curr_data_reg_31_inst : DFF_X1 port map( D => n3204, CK =>
                           CLK, Q => n_3932, QN => 
                           DataPath_WRF_CUhw_curr_data_31_port);
   DataPath_WRF_CUhw_curr_data_reg_30_inst : DFF_X1 port map( D => n3207, CK =>
                           CLK, Q => n_3933, QN => 
                           DataPath_WRF_CUhw_curr_data_30_port);
   DataPath_WRF_CUhw_curr_data_reg_28_inst : DFF_X1 port map( D => n3209, CK =>
                           CLK, Q => n_3934, QN => 
                           DataPath_WRF_CUhw_curr_data_28_port);
   DataPath_WRF_CUhw_curr_data_reg_19_inst : DFF_X1 port map( D => n3218, CK =>
                           CLK, Q => n_3935, QN => 
                           DataPath_WRF_CUhw_curr_data_19_port);
   DataPath_WRF_CUhw_curr_data_reg_17_inst : DFF_X1 port map( D => n3220, CK =>
                           CLK, Q => n_3936, QN => 
                           DataPath_WRF_CUhw_curr_data_17_port);
   DataPath_WRF_CUhw_curr_data_reg_16_inst : DFF_X1 port map( D => n3221, CK =>
                           CLK, Q => n_3937, QN => 
                           DataPath_WRF_CUhw_curr_data_16_port);
   DataPath_WRF_CUhw_curr_data_reg_27_inst : DFF_X1 port map( D => n3210, CK =>
                           CLK, Q => n_3938, QN => 
                           DataPath_WRF_CUhw_curr_data_27_port);
   DataPath_WRF_CUhw_curr_data_reg_15_inst : DFF_X1 port map( D => n3222, CK =>
                           CLK, Q => n_3939, QN => 
                           DataPath_WRF_CUhw_curr_data_15_port);
   DataPath_WRF_CUhw_curr_data_reg_9_inst : DFF_X1 port map( D => n3228, CK => 
                           CLK, Q => n_3940, QN => 
                           DataPath_WRF_CUhw_curr_data_9_port);
   DataPath_WRF_CUhw_curr_data_reg_5_inst : DFF_X1 port map( D => n3232, CK => 
                           CLK, Q => n_3941, QN => 
                           DataPath_WRF_CUhw_curr_data_5_port);
   DataPath_WRF_CUhw_curr_data_reg_25_inst : DFF_X1 port map( D => n3212, CK =>
                           CLK, Q => n_3942, QN => 
                           DataPath_WRF_CUhw_curr_data_25_port);
   DataPath_WRF_CUhw_curr_data_reg_24_inst : DFF_X1 port map( D => n3213, CK =>
                           CLK, Q => n_3943, QN => 
                           DataPath_WRF_CUhw_curr_data_24_port);
   DataPath_WRF_CUhw_curr_data_reg_23_inst : DFF_X1 port map( D => n3214, CK =>
                           CLK, Q => n_3944, QN => 
                           DataPath_WRF_CUhw_curr_data_23_port);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_1_inst : DFF_X1 port map( D => 
                           n7164, CK => CLK, Q => n_3945, QN => n542);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_3_inst : DFF_X1 port map( D => 
                           n7162, CK => CLK, Q => n_3946, QN => n544);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_5_inst : DFF_X1 port map( D => 
                           n7160, CK => CLK, Q => n_3947, QN => n546);
   DataPath_RF_PUSH_ADDRGEN_curr_state_reg_1_inst : DFF_X1 port map( D => n90, 
                           CK => CLK, Q => n_3948, QN => n838);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_7_inst : DFF_X1 port map( D => 
                           n7158, CK => CLK, Q => n_3949, QN => n548);
   CU_I_unsigned_2_reg : DFF_X1 port map( D => n7083, CK => CLK, Q => n_3950, 
                           QN => n212);
   CU_I_unsigned_1_reg : DFF_X1 port map( D => n7084, CK => CLK, Q => n_3951, 
                           QN => n213);
   CU_I_i_SPILL_delay_reg : DFF_X1 port map( D => CU_I_N318, CK => CLK, Q => 
                           n_3952, QN => n8272);
   DataPath_REG_IN2_Q_reg_6_inst : DFF_X1 port map( D => n7026, CK => CLK, Q =>
                           n_3953, QN => n486);
   DataPath_RF_POP_ADDRGEN_curr_state_reg_0_inst : DFF_X1 port map( D => n7063,
                           CK => CLK, Q => n_3954, QN => n866);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_9_inst : DFF_X1 port map( D => 
                           n7156, CK => CLK, Q => n_3955, QN => n550);
   CU_I_sel_alu_setcmp_1_reg : DFF_X1 port map( D => n7087, CK => CLK, Q => 
                           n_3956, QN => n217);
   CU_I_setcmp_1_reg_2_inst : DFF_X1 port map( D => n7088, CK => CLK, Q => 
                           n_3957, QN => n219);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_14_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N60, CK => CLK, Q => n_3958
                           , QN => n8310);
   DataPath_WRF_CUhw_curr_state_reg_0_inst : DFF_X1 port map( D => n99, CK => 
                           CLK, Q => n_3959, QN => n465);
   CU_I_CW_MEM_reg_WB_MUX_SEL_inst : DFF_X1 port map( D => n2832, CK => CLK, Q 
                           => n_3960, QN => CU_I_CW_MEM_WB_MUX_SEL_port);
   CU_I_CW_MEM_reg_WB_EN_inst : DFF_X1 port map( D => n2833, CK => CLK, Q => 
                           n_3961, QN => CU_I_CW_MEM_WB_EN_port);
   CU_I_CW_EX_reg_WB_MUX_SEL_inst : DFF_X1 port map( D => n2838, CK => CLK, Q 
                           => n_3962, QN => CU_I_CW_EX_WB_MUX_SEL_port);
   CU_I_CW_EX_reg_WB_EN_inst : DFF_X1 port map( D => n2839, CK => CLK, Q => 
                           n_3963, QN => CU_I_CW_EX_WB_EN_port);
   DataPath_REG_IN2_Q_reg_5_inst : DFF_X1 port map( D => n2380, CK => CLK, Q =>
                           n_3964, QN => DataPath_i_PIPLIN_IN2_5_port);
   DataPath_REG_IN1_Q_reg_14_inst : DFF_X1 port map( D => n2842, CK => CLK, Q 
                           => n_3965, QN => DataPath_i_PIPLIN_IN1_14_port);
   DataPath_REG_IN1_Q_reg_13_inst : DFF_X1 port map( D => n2843, CK => CLK, Q 
                           => n_3966, QN => DataPath_i_PIPLIN_IN1_13_port);
   DataPath_REG_IN1_Q_reg_12_inst : DFF_X1 port map( D => n2844, CK => CLK, Q 
                           => n_3967, QN => DataPath_i_PIPLIN_IN1_12_port);
   DataPath_REG_IN1_Q_reg_10_inst : DFF_X1 port map( D => n2846, CK => CLK, Q 
                           => n_3968, QN => DataPath_i_PIPLIN_IN1_10_port);
   DataPath_REG_IN1_Q_reg_8_inst : DFF_X1 port map( D => n2848, CK => CLK, Q =>
                           n_3969, QN => DataPath_i_PIPLIN_IN1_8_port);
   DataPath_REG_IN1_Q_reg_3_inst : DFF_X1 port map( D => n2853, CK => CLK, Q =>
                           n_3970, QN => DataPath_i_PIPLIN_IN1_3_port);
   DataPath_REG_IN1_Q_reg_1_inst : DFF_X1 port map( D => n2858, CK => CLK, Q =>
                           n_3971, QN => DataPath_i_PIPLIN_IN1_1_port);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_11_inst : DFF_X1 port map( D => 
                           n7154, CK => CLK, Q => n_3972, QN => n552);
   DataPath_REG_B_Q_reg_23_inst : DFF_X1 port map( D => n2740, CK => CLK, Q => 
                           n9102, QN => DataPath_i_PIPLIN_B_23_port);
   DataPath_REG_B_Q_reg_21_inst : DFF_X1 port map( D => n2742, CK => CLK, Q => 
                           n9097, QN => DataPath_i_PIPLIN_B_21_port);
   DataPath_REG_A_Q_reg_30_inst : DFF_X1 port map( D => n3239, CK => CLK, Q => 
                           n_3973, QN => DataPath_i_PIPLIN_A_30_port);
   IR_reg_1_inst : DFFS_X1 port map( D => n10411, CK => CLK, SN => n8573, Q => 
                           n10160, QN => IR_1_port);
   IR_reg_29_inst : DFFS_X1 port map( D => n10414, CK => CLK, SN => n8572, Q =>
                           n8281, QN => IR_29_port);
   IR_reg_27_inst : DFFR_X1 port map( D => n7122, CK => CLK, RN => n8570, Q => 
                           n10149, QN => n167);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_15_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N61, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_15_port, QN => 
                           n8203);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_4_inst : DFF_X1 port map( D => 
                           n11710, CK => CLK, Q => n8266, QN => 
                           DECODEhw_i_tickcounter_4_port);
   DataPath_RF_PUSH_ADDRGEN_curr_addr_reg_0_inst : DFF_X1 port map( D => 
                           DataPath_RF_PUSH_ADDRGEN_N46, CK => CLK, Q => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, QN => 
                           n8325);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_0_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N46, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_0_port, QN => 
                           n8327);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_15_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N61, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_15_port, QN => 
                           n8291);
   DataPath_RF_SWP_Q_reg_0_inst : DFF_X1 port map( D => n7068, CK => CLK, Q => 
                           DataPath_RF_c_swin_0_port, QN => n8242);
   DataPath_REG_B_Q_reg_6_inst : DFF_X1 port map( D => n7080, CK => CLK, Q => 
                           n8320, QN => n477);
   DataPath_RF_SWP_Q_reg_4_inst : DFF_X1 port map( D => n7064, CK => CLK, Q => 
                           DataPath_RF_c_swin_4_port, QN => n8334);
   DataPath_RF_SWP_Q_reg_2_inst : DFF_X1 port map( D => n7066, CK => CLK, Q => 
                           DataPath_RF_c_swin_2_port, QN => n825);
   DataPath_RF_SWP_Q_reg_1_inst : DFF_X1 port map( D => n7067, CK => CLK, Q => 
                           DataPath_RF_c_swin_1_port, QN => n824);
   DataPath_RF_SWP_Q_reg_3_inst : DFF_X1 port map( D => n7065, CK => CLK, Q => 
                           DataPath_RF_c_swin_3_port, QN => n826);
   DataPath_REG_B_Q_reg_13_inst : DFF_X1 port map( D => n7077, CK => CLK, Q => 
                           DataPath_i_PIPLIN_B_13_port, QN => n8324);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_8_inst : DFF_X1 port map( D => n6823, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_72_port,
                           QN => n639);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_7_inst : DFF_X1 port map( D => n6824, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_71_port,
                           QN => n638);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_6_inst : DFF_X1 port map( D => n6825, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_70_port,
                           QN => n637);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_5_inst : DFF_X1 port map( D => n6826, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_69_port,
                           QN => n636);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_4_inst : DFF_X1 port map( D => n6827, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_68_port,
                           QN => n635);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_3_inst : DFF_X1 port map( D => n6828, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_67_port,
                           QN => n634);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_2_inst : DFF_X1 port map( D => n6829, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_66_port,
                           QN => n633);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_1_inst : DFF_X1 port map( D => n6830, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_65_port,
                           QN => n632);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_0_inst : DFF_X1 port map( D => n6831, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_64_port,
                           QN => n631);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_8_inst : DFF_X1 port map( D => n6983, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_232_port
                           , QN => n799);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_7_inst : DFF_X1 port map( D => n6984, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_231_port
                           , QN => n798);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_6_inst : DFF_X1 port map( D => n6985, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_230_port
                           , QN => n797);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_5_inst : DFF_X1 port map( D => n6986, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_229_port
                           , QN => n796);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_4_inst : DFF_X1 port map( D => n6987, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_228_port
                           , QN => n795);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_3_inst : DFF_X1 port map( D => n6988, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_227_port
                           , QN => n794);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_2_inst : DFF_X1 port map( D => n6989, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_226_port
                           , QN => n793);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_1_inst : DFF_X1 port map( D => n6990, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_225_port
                           , QN => n792);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_0_inst : DFF_X1 port map( D => n6991, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_224_port
                           , QN => n791);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_14_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N60, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_14_port, QN => 
                           n8211);
   DataPath_RF_POP_ADDRGEN_curr_addr_reg_8_inst : DFF_X1 port map( D => 
                           DataPath_RF_POP_ADDRGEN_N54, CK => CLK, Q => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_8_port, QN => 
                           n8308);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_22_inst : DFF_X1 port map( D => n6969, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_246_port
                           , QN => n813);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_22_inst : DFF_X1 port map( D => n6809, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_86_port,
                           QN => n653);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_26_inst : DFF_X1 port map( D => n6965, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_250_port
                           , QN => n817);
   DataPath_RF_BLOCK_GLOB_2_Q_reg_26_inst : DFF_X1 port map( D => n6805, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_90_port,
                           QN => n657);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_26_inst : DFF_X1 port map( D => n6901, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_186_port
                           , QN => n753);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_22_inst : DFF_X1 port map( D => n6905, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_182_port
                           , QN => n749);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_10_inst : DFF_X1 port map( D => n6917, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_170_port
                           , QN => n737);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_8_inst : DFF_X1 port map( D => n6919, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_168_port
                           , QN => n735);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_7_inst : DFF_X1 port map( D => n6920, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_167_port
                           , QN => n734);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_6_inst : DFF_X1 port map( D => n6921, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_166_port
                           , QN => n733);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_5_inst : DFF_X1 port map( D => n6922, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_165_port
                           , QN => n732);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_4_inst : DFF_X1 port map( D => n6923, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_164_port
                           , QN => n731);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_3_inst : DFF_X1 port map( D => n6924, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_163_port
                           , QN => n730);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_2_inst : DFF_X1 port map( D => n6925, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_162_port
                           , QN => n729);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_1_inst : DFF_X1 port map( D => n6926, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_161_port
                           , QN => n728);
   DataPath_RF_BLOCK_GLOB_5_Q_reg_0_inst : DFF_X1 port map( D => n6927, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_160_port
                           , QN => n727);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_26_inst : DFF_X1 port map( D => n6773, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_58_port,
                           QN => n625);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_22_inst : DFF_X1 port map( D => n6777, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_54_port,
                           QN => n621);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_10_inst : DFF_X1 port map( D => n6789, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_42_port,
                           QN => n609);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_8_inst : DFF_X1 port map( D => n6791, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_40_port,
                           QN => n607);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_7_inst : DFF_X1 port map( D => n6792, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_39_port,
                           QN => n606);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_6_inst : DFF_X1 port map( D => n6793, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_38_port,
                           QN => n605);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_5_inst : DFF_X1 port map( D => n6794, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_37_port,
                           QN => n604);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_4_inst : DFF_X1 port map( D => n6795, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_36_port,
                           QN => n603);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_3_inst : DFF_X1 port map( D => n6796, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_35_port,
                           QN => n602);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_2_inst : DFF_X1 port map( D => n6797, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_34_port,
                           QN => n601);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_1_inst : DFF_X1 port map( D => n6798, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_33_port,
                           QN => n600);
   DataPath_RF_BLOCK_GLOB_1_Q_reg_0_inst : DFF_X1 port map( D => n6799, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_32_port,
                           QN => n599);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_25_inst : DFF_X1 port map( D => n6966, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_249_port
                           , QN => n816);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_24_inst : DFF_X1 port map( D => n6967, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_248_port
                           , QN => n815);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_23_inst : DFF_X1 port map( D => n6968, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_247_port
                           , QN => n814);
   DataPath_RF_BLOCK_GLOB_7_Q_reg_9_inst : DFF_X1 port map( D => n6982, CK => 
                           CLK, Q => DataPath_RF_bus_complete_win_data_233_port
                           , QN => n800);
   DECODEhw_HALF_ADDER_COUNTER_REG_TICK_Q_reg_2_inst : DFF_X1 port map( D => 
                           n11707, CK => CLK, Q => n_3974, QN => 
                           DECODEhw_i_tickcounter_2_port);
   PC_reg_30_inst : DFFR_X1 port map( D => n7031, CK => CLK, RN => n8570, Q => 
                           IRAM_ADDRESS_30_port, QN => n8003);
   PC_reg_31_inst : DFFR_X1 port map( D => n7030, CK => CLK, RN => n8570, Q => 
                           IRAM_ADDRESS_31_port, QN => n8048);
   DataPath_RF_CWP_Q_reg_2_inst : DFF_X2 port map( D => n7072, CK => CLK, Q => 
                           DataPath_RF_c_win_2_port, QN => n575);
   DataPath_RF_CWP_Q_reg_4_inst : DFF_X2 port map( D => n7070, CK => CLK, Q => 
                           DataPath_RF_c_win_4_port, QN => n8219);
   DataPath_RF_CWP_Q_reg_3_inst : DFF_X1 port map( D => n7071, CK => CLK, Q => 
                           DataPath_RF_c_win_3_port, QN => n576);
   IR_reg_6_inst : DFFR_X1 port map( D => n40, CK => CLK, RN => n8571, Q => 
                           IR_6_port, QN => n8228);
   DataPath_WRF_CUhw_curr_addr_reg_31_inst : DFF_X1 port map( D => n8393, CK =>
                           CLK, Q => DataPath_WRF_CUhw_curr_addr_31_port, QN =>
                           n_3975);
   U7551 : OAI33_X1 port map( A1 => n7425, A2 => n7423, A3 => n7424, B1 => 
                           n10317, B2 => n8386, B3 => n10315, ZN => n7426);
   U7552 : CLKBUF_X3 port map( A => n9061, Z => n8441);
   U7553 : CLKBUF_X3 port map( A => n9061, Z => n8440);
   U7554 : CLKBUF_X3 port map( A => n9061, Z => n8442);
   U7555 : BUF_X1 port map( A => DP_OP_751_130_6421_n982, Z => n7187);
   U7556 : XOR2_X1 port map( A => n7912, B => n7837, Z => n7188);
   U7557 : CLKBUF_X3 port map( A => n9062, Z => n8432);
   U7558 : CLKBUF_X1 port map( A => n7309, Z => n7981);
   U7559 : BUF_X2 port map( A => n9059, Z => n7750);
   U7560 : CLKBUF_X3 port map( A => n9062, Z => n8429);
   U7561 : NAND2_X2 port map( A1 => DataPath_i_PIPLIN_A_18_port, A2 => n8555, 
                           ZN => n9495);
   U7562 : AND2_X1 port map( A1 => DP_OP_751_130_6421_n1724, A2 => 
                           DP_OP_751_130_6421_n1754, ZN => n7189);
   U7563 : AND2_X1 port map( A1 => n7597, A2 => n10277, ZN => n7190);
   U7564 : BUF_X2 port map( A => n9239, Z => n7795);
   U7565 : BUF_X2 port map( A => n8193, Z => n7929);
   U7566 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1651, A2 => 
                           DP_OP_751_130_6421_n1607, ZN => n7956);
   U7567 : BUF_X2 port map( A => n7795, Z => n7823);
   U7568 : BUF_X2 port map( A => n10032, Z => n8427);
   U7569 : BUF_X2 port map( A => n9069, Z => n7616);
   U7570 : NAND2_X1 port map( A1 => n8599, A2 => n8600, ZN => n10238);
   U7571 : BUF_X2 port map( A => n8556, Z => n7617);
   U7572 : BUF_X1 port map( A => n10261, Z => n7604);
   U7573 : AND2_X1 port map( A1 => n10242, A2 => IRAM_ADDRESS_16_port, ZN => 
                           n7728);
   U7574 : BUF_X2 port map( A => n7749, Z => n7880);
   U7575 : OR2_X1 port map( A1 => n7779, A2 => 
                           DataPath_WRF_CUhw_curr_addr_2_port, ZN => n8131);
   U7576 : INV_X1 port map( A => n8069, ZN => n8136);
   U7577 : BUF_X1 port map( A => n9806, Z => n7893);
   U7578 : BUF_X1 port map( A => n9197, Z => n7897);
   U7579 : BUF_X1 port map( A => n8004, Z => n7974);
   U7580 : INV_X1 port map( A => n7728, ZN => n10334);
   U7581 : BUF_X1 port map( A => n167, Z => n7752);
   U7582 : INV_X1 port map( A => n7691, ZN => DP_OP_751_130_6421_n95);
   U7583 : AOI22_X1 port map( A1 => n8136, A2 => DataPath_i_PIPLIN_B_14_port, 
                           B1 => DataPath_i_PIPLIN_IN2_14_port, B2 => n8137, ZN
                           => n7191);
   U7584 : INV_X1 port map( A => n7191, ZN => n9807);
   U7585 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n106, A2 => n8151, ZN =>
                           n7192);
   U7586 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n111, B2 => 
                           DP_OP_751_130_6421_n109, A => 
                           DP_OP_751_130_6421_n110, ZN => n7193);
   U7587 : XNOR2_X1 port map( A => n7193, B => n7192, ZN => n7194);
   U7588 : OR2_X1 port map( A1 => n10051, A2 => n10048, ZN => n7195);
   U7589 : AOI22_X1 port map( A1 => n8438, A2 => n10088, B1 => n10033, B2 => 
                           n8439, ZN => n7196);
   U7590 : OAI221_X1 port map( B1 => n8439, B2 => n10035, C1 => n8438, C2 => 
                           n10088, A => n9754, ZN => n7197);
   U7591 : OAI21_X1 port map( B1 => n7196, B2 => n9754, A => n7197, ZN => n7198
                           );
   U7592 : AOI21_X1 port map( B1 => n10052, B2 => n7195, A => n7198, ZN => 
                           n7199);
   U7593 : OAI21_X1 port map( B1 => n10055, B2 => n7195, A => n7199, ZN => 
                           n7200);
   U7594 : AOI21_X1 port map( B1 => n10094, B2 => n7194, A => n7200, ZN => 
                           n7201);
   U7595 : AOI22_X1 port map( A1 => n10062, A2 => n10117, B1 => n10120, B2 => 
                           n10063, ZN => n7202);
   U7596 : AOI22_X1 port map( A1 => n10064, A2 => n10112, B1 => n10110, B2 => 
                           n10065, ZN => n7203);
   U7597 : OAI211_X1 port map( C1 => n10067, C2 => n10002, A => n7202, B => 
                           n7203, ZN => n7204);
   U7598 : OAI22_X1 port map( A1 => n10057, A2 => n10106, B1 => n10058, B2 => 
                           n10066, ZN => n7205);
   U7599 : OAI22_X1 port map( A1 => n10060, A2 => n10046, B1 => n10039, B2 => 
                           n10104, ZN => n7206);
   U7600 : NOR3_X1 port map( A1 => n7204, A2 => n7205, A3 => n7206, ZN => n7207
                           );
   U7601 : OAI222_X1 port map( A1 => n11885, A2 => n7201, B1 => n11884, B2 => 
                           n504, C1 => n7207, C2 => n11881, ZN => n7007);
   U7602 : OAI22_X1 port map( A1 => n7726, A2 => n8405, B1 => n9753, B2 => 
                           n8134, ZN => DataPath_ALUhw_MULT_mux_out_0_17_port);
   U7603 : AOI22_X1 port map( A1 => n8148, A2 => 
                           DataPath_ALUhw_MULT_mux_out_0_9_port, B1 => 
                           DP_OP_751_130_6421_n1790, B2 => n7998, ZN => n7208);
   U7604 : OAI22_X1 port map( A1 => n8430, A2 => n9248, B1 => n9239, B2 => 
                           n8442, ZN => n7209);
   U7605 : XNOR2_X1 port map( A => n8146, B => n7209, ZN => n7210);
   U7606 : NOR2_X1 port map( A1 => n7208, A2 => n7210, ZN => 
                           DP_OP_751_130_6421_n1681);
   U7607 : XOR2_X1 port map( A => n7208, B => n7210, Z => 
                           DP_OP_751_130_6421_n1682);
   U7608 : AOI22_X1 port map( A1 => n8562, A2 => n9754, B1 => 
                           DP_OP_751_130_6421_n1017, B2 => 
                           DP_OP_751_130_6421_n1119, ZN => n7211);
   U7609 : OAI21_X1 port map( B1 => n9754, B2 => DP_OP_751_130_6421_n1017, A =>
                           n7211, ZN => n9088);
   U7610 : NAND2_X1 port map( A1 => n9727, A2 => n10103, ZN => n7212);
   U7611 : AOI21_X1 port map( B1 => n7212, B2 => n9728, A => n9732, ZN => n7213
                           );
   U7612 : AOI21_X1 port map( B1 => n9731, B2 => n7788, A => n7213, ZN => n7214
                           );
   U7613 : NAND2_X1 port map( A1 => n9725, A2 => n9724, ZN => n7215);
   U7614 : OAI21_X1 port map( B1 => n7215, B2 => n9726, A => n7214, ZN => n7216
                           );
   U7615 : AOI21_X1 port map( B1 => n9730, B2 => n9729, A => n7216, ZN => 
                           n10067);
   U7616 : NAND2_X1 port map( A1 => n7897, A2 => n8146, ZN => n7217);
   U7617 : NAND2_X1 port map( A1 => n10036, A2 => n7217, ZN => n7218);
   U7618 : OAI221_X1 port map( B1 => n7217, B2 => n10035, C1 => n7897, C2 => 
                           n8146, A => n7218, ZN => n7219);
   U7619 : INV_X1 port map( A => DP_OP_751_130_6421_n162, ZN => n7220);
   U7620 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n161, A2 => n7220, ZN => 
                           n7221);
   U7621 : XNOR2_X1 port map( A => n8398, B => n9201, ZN => n7222);
   U7622 : INV_X1 port map( A => n10427, ZN => n7223);
   U7623 : OAI21_X1 port map( B1 => n7223, B2 => n11856, A => n9198, ZN => 
                           n7224);
   U7624 : XNOR2_X1 port map( A => n7224, B => n7222, ZN => n7225);
   U7625 : NAND2_X1 port map( A1 => n10427, A2 => n11857, ZN => n7226);
   U7626 : OAI21_X1 port map( B1 => n7222, B2 => n7226, A => n11858, ZN => 
                           n7227);
   U7627 : AOI222_X1 port map( A1 => n7225, A2 => n7227, B1 => n7225, B2 => 
                           n7226, C1 => n7227, C2 => n11859, ZN => n7228);
   U7628 : XNOR2_X1 port map( A => n7221, B => DP_OP_751_130_6421_n163, ZN => 
                           n7229);
   U7629 : AOI21_X1 port map( B1 => n7229, B2 => n10094, A => n7228, ZN => 
                           n7230);
   U7630 : NAND3_X1 port map( A1 => n10033, A2 => n8398, A3 => n7774, ZN => 
                           n7231);
   U7631 : NAND3_X1 port map( A1 => n7219, A2 => n7230, A3 => n7231, ZN => 
                           n7232);
   U7632 : OAI22_X1 port map( A1 => n10001, A2 => n9977, B1 => n9185, B2 => 
                           n10104, ZN => n7233);
   U7633 : OAI22_X1 port map( A1 => n9885, A2 => n10038, B1 => n9975, B2 => 
                           n10002, ZN => n7234);
   U7634 : AOI211_X1 port map( C1 => n10430, C2 => n11866, A => n7233, B => 
                           n7234, ZN => n7235);
   U7635 : AOI22_X1 port map( A1 => n9247, A2 => n10120, B1 => n10113, B2 => 
                           n9888, ZN => n7236);
   U7636 : AOI22_X1 port map( A1 => n9972, A2 => n10116, B1 => n10117, B2 => 
                           n9890, ZN => n7237);
   U7637 : NAND3_X1 port map( A1 => n7235, A2 => n7236, A3 => n7237, ZN => 
                           n7238);
   U7638 : AOI222_X1 port map( A1 => n7232, A2 => n10429, B1 => 
                           DRAM_ADDRESS_3_port, B2 => n7791, C1 => n7238, C2 =>
                           n10428, ZN => n2119);
   U7639 : AND2_X1 port map( A1 => n8572, A2 => 
                           DataPath_RF_internal_out2_19_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N23);
   U7640 : AND2_X1 port map( A1 => n8572, A2 => 
                           DataPath_RF_internal_out1_29_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N33);
   U7641 : OAI22_X1 port map( A1 => n8134, A2 => n9122, B1 => n7726, B2 => 
                           n9844, ZN => n7239);
   U7642 : XOR2_X1 port map( A => n8148, B => n7239, Z => n7240);
   U7643 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_11_port, B => 
                           n8146, ZN => n7241);
   U7644 : NOR2_X1 port map( A1 => n7240, A2 => n7241, ZN => 
                           DP_OP_751_130_6421_n1677);
   U7645 : XOR2_X1 port map( A => n7240, B => n7241, Z => 
                           DP_OP_751_130_6421_n1678);
   U7646 : INV_X1 port map( A => n7693, ZN => n7242);
   U7647 : NAND2_X1 port map( A1 => n8164, A2 => n7242, ZN => n7243);
   U7648 : XNOR2_X1 port map( A => n7918, B => n7243, ZN => n7244);
   U7649 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n813, A2 => n9962, ZN =>
                           n7245);
   U7650 : OAI22_X1 port map( A1 => DP_OP_751_130_6421_n813, A2 => n9962, B1 =>
                           n10035, B2 => n7245, ZN => n7246);
   U7651 : NAND3_X1 port map( A1 => n9961, A2 => n10033, A3 => n7794, ZN => 
                           n7247);
   U7652 : OAI221_X1 port map( B1 => n7246, B2 => n10036, C1 => n7246, C2 => 
                           n7245, A => n7247, ZN => n7248);
   U7653 : INV_X1 port map( A => n9957, ZN => n7249);
   U7654 : OAI22_X1 port map( A1 => n9959, A2 => n9958, B1 => n9960, B2 => 
                           n7249, ZN => n7250);
   U7655 : AOI22_X1 port map( A1 => n9965, A2 => n7250, B1 => n9964, B2 => 
                           n9963, ZN => n7251);
   U7656 : OAI21_X1 port map( B1 => n9965, B2 => n9966, A => n7251, ZN => n7252
                           );
   U7657 : AOI211_X1 port map( C1 => n10094, C2 => n7244, A => n7248, B => 
                           n7252, ZN => n7253);
   U7658 : AOI22_X1 port map( A1 => n9967, A2 => n10430, B1 => n10121, B2 => 
                           n10062, ZN => n7254);
   U7659 : AOI22_X1 port map( A1 => n10042, A2 => n10045, B1 => n10113, B2 => 
                           n10065, ZN => n7255);
   U7660 : OAI211_X1 port map( C1 => n9968, C2 => n10046, A => n7254, B => 
                           n7255, ZN => n7256);
   U7661 : OAI22_X1 port map( A1 => n10061, A2 => n10059, B1 => n10057, B2 => 
                           n10038, ZN => n7257);
   U7662 : OAI22_X1 port map( A1 => n7810, A2 => n9977, B1 => n9969, B2 => 
                           n10056, ZN => n7258);
   U7663 : NOR3_X1 port map( A1 => n7256, A2 => n7257, A3 => n7258, ZN => n7259
                           );
   U7664 : OAI222_X1 port map( A1 => n8329, A2 => n11884, B1 => n11880, B2 => 
                           n7253, C1 => n7259, C2 => n11881, ZN => n7002);
   U7665 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_29_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N33);
   U7666 : AND2_X1 port map( A1 => n8580, A2 => 
                           DataPath_RF_internal_out1_19_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N23);
   U7667 : NAND2_X1 port map( A1 => n9056, A2 => n9011, ZN => n7260);
   U7668 : AOI21_X1 port map( B1 => n11868, B2 => n9137, A => n7260, ZN => 
                           n9347);
   U7669 : OAI22_X1 port map( A1 => n8134, A2 => n9168, B1 => n7726, B2 => 
                           n8399, ZN => n7261);
   U7670 : XNOR2_X1 port map( A => n8148, B => n7261, ZN => n7262);
   U7671 : AND2_X1 port map( A1 => n7262, A2 => DP_OP_751_130_6421_n1698, ZN =>
                           DP_OP_751_130_6421_n1697);
   U7672 : XOR2_X1 port map( A => n7262, B => DP_OP_751_130_6421_n1698, Z => 
                           DP_OP_751_130_6421_n1694);
   U7673 : AOI22_X1 port map( A1 => n8136, A2 => DataPath_i_PIPLIN_B_12_port, 
                           B1 => DataPath_i_PIPLIN_IN2_12_port, B2 => n8069, ZN
                           => n7263);
   U7674 : INV_X1 port map( A => n7263, ZN => n9823);
   U7675 : NAND3_X1 port map( A1 => n7788, A2 => n7806, A3 => n7805, ZN => 
                           n7264);
   U7676 : NAND2_X1 port map( A1 => n9548, A2 => n10103, ZN => n7265);
   U7677 : OAI211_X1 port map( C1 => n9544, C2 => n7982, A => n7264, B => n7265
                           , ZN => n7266);
   U7678 : AOI21_X1 port map( B1 => n8438, B2 => n9657, A => n7266, ZN => n7267
                           );
   U7679 : OAI21_X1 port map( B1 => n8189, B2 => n9379, A => n9531, ZN => n7268
                           );
   U7680 : NAND3_X1 port map( A1 => n9549, A2 => n9724, A3 => n7268, ZN => 
                           n7269);
   U7681 : OAI211_X1 port map( C1 => n9264, C2 => n9246, A => n7267, B => n7269
                           , ZN => n9972);
   U7682 : AND2_X1 port map( A1 => n8576, A2 => 
                           DataPath_RF_internal_out2_17_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N21);
   U7683 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out1_18_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N22);
   U7684 : OAI22_X1 port map( A1 => n8431, A2 => n9986, B1 => n8441, B2 => 
                           n9188, ZN => n7270);
   U7685 : XNOR2_X1 port map( A => n8146, B => n7270, ZN => n7271);
   U7686 : OAI22_X1 port map( A1 => n7756, A2 => n9239, B1 => n7726, B2 => 
                           n9248, ZN => n7272);
   U7687 : XOR2_X1 port map( A => n8148, B => n7272, Z => n7273);
   U7688 : XOR2_X1 port map( A => n7271, B => n7273, Z => 
                           DP_OP_751_130_6421_n1686);
   U7689 : NOR2_X1 port map( A1 => n7271, A2 => n7273, ZN => 
                           DP_OP_751_130_6421_n1685);
   U7690 : NAND2_X1 port map( A1 => n7794, A2 => n9637, ZN => n7274);
   U7691 : OAI221_X1 port map( B1 => n9601, B2 => n7794, C1 => n9637, C2 => 
                           DP_OP_751_130_6421_n711, A => n7274, ZN => n9104);
   U7692 : INV_X1 port map( A => n9179, ZN => n7275);
   U7693 : AOI21_X1 port map( B1 => n8398, B2 => i_ALU_OP_2_port, A => n7275, 
                           ZN => n9702);
   U7694 : NAND2_X1 port map( A1 => n7851, A2 => n7849, ZN => n7276);
   U7695 : NAND2_X1 port map( A1 => intadd_1_n6, A2 => n10345, ZN => n7277);
   U7696 : NAND3_X1 port map( A1 => n7277, A2 => n10344, A3 => n7276, ZN => 
                           n7610);
   U7697 : AOI22_X1 port map( A1 => n8136, A2 => DataPath_i_PIPLIN_B_20_port, 
                           B1 => DataPath_i_PIPLIN_IN2_20_port, B2 => n8137, ZN
                           => n7278);
   U7698 : INV_X1 port map( A => n7278, ZN => n9651);
   U7699 : INV_X1 port map( A => n10097, ZN => n7279);
   U7700 : AOI222_X1 port map( A1 => n9730, A2 => n7279, B1 => n10103, B2 => 
                           n9244, C1 => n7788, C2 => n9243, ZN => n7280);
   U7701 : OR2_X1 port map( A1 => n9583, A2 => n9585, ZN => n7281);
   U7702 : AOI22_X1 port map( A1 => n9245, A2 => n9582, B1 => n7789, B2 => 
                           n7281, ZN => n7282);
   U7703 : OAI211_X1 port map( C1 => n7353, C2 => n9246, A => n7280, B => n7282
                           , ZN => n10043);
   U7704 : NAND3_X1 port map( A1 => n163, A2 => n8601, A3 => n7752, ZN => n7283
                           );
   U7705 : NAND3_X1 port map( A1 => n8602, A2 => n10392, A3 => n7283, ZN => 
                           n7284);
   U7706 : AOI211_X1 port map( C1 => n159, C2 => n7962, A => n10222, B => n7284
                           , ZN => n7285);
   U7707 : NOR2_X1 port map( A1 => n11753, A2 => n7285, ZN => n10434);
   U7708 : XNOR2_X1 port map( A => n9148, B => n9147, ZN => n7286);
   U7709 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n170, B2 => 
                           DP_OP_751_130_6421_n172, A => n10094, ZN => n7287);
   U7710 : AOI21_X1 port map( B1 => DP_OP_751_130_6421_n170, B2 => 
                           DP_OP_751_130_6421_n172, A => n7287, ZN => n7288);
   U7711 : NAND3_X1 port map( A1 => n9137, A2 => n10035, A3 => n7998, ZN => 
                           n7289);
   U7712 : NAND3_X1 port map( A1 => n10033, A2 => n8148, A3 => n9133, ZN => 
                           n7290);
   U7713 : AOI21_X1 port map( B1 => n7998, B2 => n9137, A => n10036, ZN => 
                           n7291);
   U7714 : OAI21_X1 port map( B1 => n7998, B2 => n9137, A => n7291, ZN => n7292
                           );
   U7715 : AOI21_X1 port map( B1 => n9149, B2 => n9132, A => n11859, ZN => 
                           n7293);
   U7716 : OAI21_X1 port map( B1 => n9149, B2 => n9132, A => n7293, ZN => n7294
                           );
   U7717 : NAND4_X1 port map( A1 => n7289, A2 => n7290, A3 => n7292, A4 => 
                           n7294, ZN => n7295);
   U7718 : AOI211_X1 port map( C1 => n11858, C2 => n7286, A => n7288, B => 
                           n7295, ZN => n7296);
   U7719 : OAI22_X1 port map( A1 => n9976, A2 => n9977, B1 => n9134, B2 => 
                           n10104, ZN => n7297);
   U7720 : OAI22_X1 port map( A1 => n9135, A2 => n10038, B1 => n9185, B2 => 
                           n10002, ZN => n7298);
   U7721 : OAI22_X1 port map( A1 => n9884, A2 => n10056, B1 => n9885, B2 => 
                           n10046, ZN => n7299);
   U7722 : OAI22_X1 port map( A1 => n10106, A2 => n10001, B1 => n10066, B2 => 
                           n9153, ZN => n7300);
   U7723 : NOR2_X1 port map( A1 => n7299, A2 => n7300, ZN => n7301);
   U7724 : OAI21_X1 port map( B1 => n9975, B2 => n10059, A => n7301, ZN => 
                           n7302);
   U7725 : NOR3_X1 port map( A1 => n7297, A2 => n7298, A3 => n7302, ZN => n7303
                           );
   U7726 : OAI222_X1 port map( A1 => n11880, A2 => n7296, B1 => n11884, B2 => 
                           n495, C1 => n7303, C2 => n11881, ZN => n7019);
   U7727 : AND2_X1 port map( A1 => n8578, A2 => 
                           DataPath_RF_internal_out2_18_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N22);
   U7728 : AND2_X1 port map( A1 => n8576, A2 => 
                           DataPath_RF_internal_out1_17_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N21);
   U7729 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1709, B => 
                           DP_OP_751_130_6421_n1739, Z => n7958);
   U7730 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1351, B2 => 
                           DP_OP_751_130_6421_n1304, A => 
                           DP_OP_751_130_6421_n1350, ZN => n7831);
   U7731 : OAI22_X1 port map( A1 => n8440, A2 => n8398, B1 => n8432, B2 => 
                           n9188, ZN => n7304);
   U7732 : XNOR2_X1 port map( A => n8146, B => n7304, ZN => n7305);
   U7733 : OAI22_X1 port map( A1 => n7750, A2 => n9986, B1 => n7726, B2 => 
                           n9239, ZN => n7306);
   U7734 : XOR2_X1 port map( A => n8148, B => n7306, Z => n7307);
   U7735 : NOR2_X1 port map( A1 => n7305, A2 => n7307, ZN => 
                           DP_OP_751_130_6421_n1687);
   U7736 : XOR2_X1 port map( A => n7305, B => n7307, Z => 
                           DP_OP_751_130_6421_n1688);
   U7737 : NAND4_X1 port map( A1 => n10128, A2 => IR_26_port, A3 => n8354, A4 
                           => n10440, ZN => n8240);
   U7738 : AOI22_X1 port map( A1 => n9935, A2 => n9518, B1 => 
                           DP_OP_751_130_6421_n507, B2 => n7817, ZN => n7308);
   U7739 : OAI21_X1 port map( B1 => n9518, B2 => DP_OP_751_130_6421_n507, A => 
                           n7308, ZN => n9113);
   U7740 : AOI22_X1 port map( A1 => n8225, A2 => DataPath_i_PIPLIN_IN1_14_port,
                           B1 => n8555, B2 => DataPath_i_PIPLIN_A_14_port, ZN 
                           => n7309);
   U7741 : INV_X1 port map( A => n7309, ZN => n9806);
   U7742 : OAI221_X1 port map( B1 => n9243, B2 => n9283, C1 => n9243, C2 => 
                           n11853, A => n7789, ZN => n7310);
   U7743 : OAI211_X1 port map( C1 => n10081, C2 => n8566, A => n9242, B => 
                           n9708, ZN => n7311);
   U7744 : AOI22_X1 port map( A1 => n7898, A2 => n9547, B1 => n9283, B2 => 
                           n9047, ZN => n7312);
   U7745 : NAND2_X1 port map( A1 => n9586, A2 => n9244, ZN => n7313);
   U7746 : NAND3_X1 port map( A1 => n7313, A2 => n7312, A3 => n7311, ZN => 
                           n7314);
   U7747 : AOI21_X1 port map( B1 => n9582, B2 => n9045, A => n7314, ZN => n7315
                           );
   U7748 : NAND2_X1 port map( A1 => n9585, A2 => n9542, ZN => n7316);
   U7749 : NAND3_X1 port map( A1 => n7316, A2 => n7315, A3 => n7310, ZN => 
                           n9247);
   U7750 : INV_X1 port map( A => n10271, ZN => n7317);
   U7751 : NAND2_X1 port map( A1 => n10279, A2 => n7317, ZN => n7318);
   U7752 : XNOR2_X1 port map( A => n10280, B => n7318, ZN => n7319);
   U7753 : OAI22_X1 port map( A1 => n10281, A2 => n10367, B1 => n7757, B2 => 
                           n7319, ZN => n7320);
   U7754 : AOI21_X1 port map( B1 => i_RD1_28_port, B2 => n10418, A => n7320, ZN
                           => n8392);
   U7755 : AOI22_X1 port map( A1 => n10064, A2 => n10110, B1 => n10430, B2 => 
                           n10042, ZN => n7321);
   U7756 : AOI22_X1 port map( A1 => n10121, A2 => n10043, B1 => n10044, B2 => 
                           n10045, ZN => n7322);
   U7757 : OAI211_X1 port map( C1 => n10067, C2 => n10046, A => n7321, B => 
                           n7322, ZN => n7323);
   U7758 : OAI22_X1 port map( A1 => n10039, A2 => n10038, B1 => n10058, B2 => 
                           n10059, ZN => n7324);
   U7759 : OAI22_X1 port map( A1 => n10040, A2 => n10066, B1 => n10041, B2 => 
                           n10056, ZN => n7325);
   U7760 : NOR3_X1 port map( A1 => n7323, A2 => n7324, A3 => n7325, ZN => n7326
                           );
   U7761 : INV_X1 port map( A => DP_OP_751_130_6421_n118, ZN => n7327);
   U7762 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n117, A2 => n7327, ZN => 
                           n7328);
   U7763 : XNOR2_X1 port map( A => n7328, B => DP_OP_751_130_6421_n119, ZN => 
                           n7329);
   U7764 : NAND2_X1 port map( A1 => n10031, A2 => n10030, ZN => n7330);
   U7765 : AOI21_X1 port map( B1 => n10029, B2 => n10028, A => n7330, ZN => 
                           n7331);
   U7766 : INV_X1 port map( A => n10026, ZN => n7332);
   U7767 : AOI21_X1 port map( B1 => n10028, B2 => n10027, A => n7332, ZN => 
                           n7333);
   U7768 : NAND2_X1 port map( A1 => n10034, A2 => DP_OP_751_130_6421_n1221, ZN 
                           => n7334);
   U7769 : NAND2_X1 port map( A1 => n10036, A2 => n7334, ZN => n7335);
   U7770 : OAI221_X1 port map( B1 => n7334, B2 => n10035, C1 => n10034, C2 => 
                           DP_OP_751_130_6421_n1221, A => n7335, ZN => n7336);
   U7771 : NAND3_X1 port map( A1 => n8227, A2 => n10033, A3 => n8428, ZN => 
                           n7337);
   U7772 : OAI211_X1 port map( C1 => n10037, C2 => n7333, A => n7336, B => 
                           n7337, ZN => n7338);
   U7773 : AOI211_X1 port map( C1 => n10094, C2 => n7329, A => n7331, B => 
                           n7338, ZN => n7339);
   U7774 : OAI222_X1 port map( A1 => n8330, A2 => n11884, B1 => n7326, B2 => 
                           n11881, C1 => n11880, C2 => n7339, ZN => n7010);
   U7775 : AND2_X1 port map( A1 => n8570, A2 => 
                           DataPath_RF_internal_out2_15_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N19);
   U7776 : AND2_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_internal_out1_16_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N20);
   U7777 : OAI22_X1 port map( A1 => n7751, A2 => n9913, B1 => n7726, B2 => 
                           n9619, ZN => n7340);
   U7778 : XNOR2_X1 port map( A => n8147, B => n7340, ZN => 
                           DP_OP_751_130_6421_n1734);
   U7779 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1713, B => 
                           DP_OP_751_130_6421_n1743, Z => 
                           DP_OP_751_130_6421_n1658);
   U7780 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1155, B2 => 
                           DP_OP_751_130_6421_n1104, A => 
                           DP_OP_751_130_6421_n1154, ZN => n7341);
   U7781 : OAI21_X1 port map( B1 => n7342, B2 => n7343, A => n7341, ZN => 
                           DP_OP_751_130_6421_n1055);
   U7782 : INV_X1 port map( A => DP_OP_751_130_6421_n1104, ZN => n7342);
   U7783 : INV_X1 port map( A => DP_OP_751_130_6421_n1155, ZN => n7343);
   U7784 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1456, B => 
                           DP_OP_751_130_6421_n1408, ZN => n7344);
   U7785 : XNOR2_X1 port map( A => n7344, B => DP_OP_751_130_6421_n1457, ZN => 
                           DP_OP_751_130_6421_n1358);
   U7786 : NAND3_X1 port map( A1 => n8354, A2 => n8272, A3 => n8587, ZN => 
                           n7345);
   U7787 : NOR2_X1 port map( A1 => i_BUSY_WINDOW, A2 => n7345, ZN => n8358);
   U7788 : OAI22_X1 port map( A1 => n8431, A2 => n9168, B1 => n7620, B2 => 
                           n9133, ZN => n7346);
   U7789 : XNOR2_X1 port map( A => n8146, B => n7346, ZN => n7347);
   U7790 : NOR2_X1 port map( A1 => n8446, A2 => n9130, ZN => n7348);
   U7791 : XNOR2_X1 port map( A => n7347, B => n7348, ZN => 
                           DP_OP_751_130_6421_n1594);
   U7792 : INV_X1 port map( A => n7348, ZN => n7349);
   U7793 : AOI22_X1 port map( A1 => n7348, A2 => n7347, B1 => n7772, B2 => 
                           n7349, ZN => DP_OP_751_130_6421_n1593);
   U7794 : NAND2_X1 port map( A1 => n7617, A2 => DataPath_i_PIPLIN_A_0_port, ZN
                           => n7350);
   U7795 : OAI21_X1 port map( B1 => n8557, B2 => n8262, A => n7350, ZN => n9060
                           );
   U7796 : INV_X1 port map( A => n9332, ZN => n7351);
   U7797 : OAI21_X1 port map( B1 => n7714, B2 => n9531, A => n7351, ZN => n9221
                           );
   U7798 : INV_X1 port map( A => n9761, ZN => n7352);
   U7799 : NAND2_X1 port map( A1 => n9758, A2 => n7352, ZN => n9140);
   U7800 : AOI22_X1 port map( A1 => n7983, A2 => n7809, B1 => i_ALU_OP_2_port, 
                           B2 => n9602, ZN => n7353);
   U7801 : INV_X1 port map( A => n7353, ZN => n9283);
   U7802 : OAI21_X1 port map( B1 => n8188, B2 => n7913, A => n9157, ZN => n7354
                           );
   U7803 : INV_X1 port map( A => n7354, ZN => n9507);
   U7804 : NOR2_X1 port map( A1 => n7929, A2 => n8248, ZN => n7355);
   U7805 : AOI21_X1 port map( B1 => n7929, B2 => DataPath_i_PIPLIN_IN2_11_port,
                           A => n7355, ZN => n7803);
   U7806 : NAND2_X1 port map( A1 => n8197, A2 => n9126, ZN => n7356);
   U7807 : NAND2_X1 port map( A1 => n11870, A2 => i_ALU_OP_3_port, ZN => n7357)
                           ;
   U7808 : NAND4_X1 port map( A1 => i_ALU_OP_1_port, A2 => n8292, A3 => n7356, 
                           A4 => n7357, ZN => n10036);
   U7809 : AOI22_X1 port map( A1 => n10062, A2 => n10110, B1 => n10112, B2 => 
                           n10063, ZN => n7358);
   U7810 : AOI22_X1 port map( A1 => n10064, A2 => n10121, B1 => n10116, B2 => 
                           n10065, ZN => n7359);
   U7811 : OAI211_X1 port map( C1 => n10067, C2 => n10066, A => n7358, B => 
                           n7359, ZN => n7360);
   U7812 : OAI22_X1 port map( A1 => n10057, A2 => n10056, B1 => n10058, B2 => 
                           n10104, ZN => n7361);
   U7813 : OAI22_X1 port map( A1 => n10060, A2 => n10059, B1 => n10061, B2 => 
                           n10106, ZN => n7362);
   U7814 : NOR3_X1 port map( A1 => n7360, A2 => n7361, A3 => n7362, ZN => n7363
                           );
   U7815 : OAI21_X1 port map( B1 => n10050, B2 => n10051, A => n10049, ZN => 
                           n7364);
   U7816 : INV_X1 port map( A => DP_OP_751_130_6421_n103, ZN => n7365);
   U7817 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n111, B2 => n8152, A => 
                           n8154, ZN => n7366);
   U7818 : NOR2_X1 port map( A1 => n7365, A2 => n8155, ZN => n7367);
   U7819 : OAI21_X1 port map( B1 => n7366, B2 => n7367, A => n10094, ZN => 
                           n7368);
   U7820 : AOI21_X1 port map( B1 => n7366, B2 => n7367, A => n7368, ZN => n7369
                           );
   U7821 : OAI21_X1 port map( B1 => n10050, B2 => n10048, A => n10047, ZN => 
                           n7370);
   U7822 : XNOR2_X1 port map( A => n8405, B => DP_OP_751_130_6421_n1017, ZN => 
                           n7371);
   U7823 : NOR3_X1 port map( A1 => n8563, A2 => n8405, A3 => n10084, ZN => 
                           n7372);
   U7824 : NOR3_X1 port map( A1 => n7924, A2 => DP_OP_751_130_6421_n1017, A3 =>
                           n10082, ZN => n7373);
   U7825 : AOI211_X1 port map( C1 => n10088, C2 => n7371, A => n7372, B => 
                           n7373, ZN => n7374);
   U7826 : OAI21_X1 port map( B1 => n10055, B2 => n7370, A => n7374, ZN => 
                           n7375);
   U7827 : AOI211_X1 port map( C1 => n10052, C2 => n7364, A => n7369, B => 
                           n7375, ZN => n7376);
   U7828 : OAI222_X1 port map( A1 => n8331, A2 => n11884, B1 => n7363, B2 => 
                           n11881, C1 => n11880, C2 => n7376, ZN => n7006);
   U7829 : INV_X1 port map( A => i_RD1_22_port, ZN => n7377);
   U7830 : XOR2_X1 port map( A => n10310, B => n8274, Z => n7378);
   U7831 : NAND2_X1 port map( A1 => n10313, A2 => n10311, ZN => n7379);
   U7832 : OAI22_X1 port map( A1 => n7379, A2 => n10312, B1 => n10313, B2 => 
                           n7378, ZN => n7380);
   U7833 : OAI222_X1 port map( A1 => n7377, A2 => n11845, B1 => n7380, B2 => 
                           n7757, C1 => n10367, C2 => n8274, ZN => n7039);
   U7834 : AND2_X1 port map( A1 => n8578, A2 => 
                           DataPath_RF_internal_out2_16_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N20);
   U7835 : AND2_X1 port map( A1 => n8573, A2 => 
                           DataPath_RF_internal_out1_15_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N19);
   U7836 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1708, B => 
                           DP_OP_751_130_6421_n1738, Z => n7934);
   U7837 : XOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_17_port, B => 
                           n7774, Z => n7381);
   U7838 : AOI22_X1 port map( A1 => n8148, A2 => 
                           DataPath_ALUhw_MULT_mux_out_0_17_port, B1 => 
                           DP_OP_751_130_6421_n1782, B2 => n7837, ZN => n7382);
   U7839 : NOR2_X1 port map( A1 => n7381, A2 => n7382, ZN => 
                           DP_OP_751_130_6421_n1665);
   U7840 : XOR2_X1 port map( A => n7381, B => n7382, Z => 
                           DP_OP_751_130_6421_n1666);
   U7841 : OAI22_X1 port map( A1 => n9822, A2 => n7750, B1 => n7726, B2 => 
                           n10032, ZN => n7383);
   U7842 : XOR2_X1 port map( A => n8147, B => n7383, Z => n7384);
   U7843 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_13_port, B => 
                           n8146, ZN => n7385);
   U7844 : NOR2_X1 port map( A1 => n7384, A2 => n7385, ZN => 
                           DP_OP_751_130_6421_n1673);
   U7845 : XOR2_X1 port map( A => n7384, B => n7385, Z => 
                           DP_OP_751_130_6421_n1674);
   U7846 : OAI22_X1 port map( A1 => n7756, A2 => n8404, B1 => n7726, B2 => 
                           n7800, ZN => n7386);
   U7847 : XNOR2_X1 port map( A => n8148, B => n7386, ZN => 
                           DP_OP_751_130_6421_n1754);
   U7848 : OAI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n31, B2 => 
                           DataPath_WRF_CUhw_curr_addr_26_port, A => n7868, ZN 
                           => n7387);
   U7849 : AOI21_X1 port map( B1 => n8033, B2 => n7869, A => n7387, ZN => n7867
                           );
   U7850 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n507, B2 => 
                           DP_OP_751_130_6421_n506, A => 
                           DP_OP_751_130_6421_n571, ZN => n7388);
   U7851 : OAI21_X1 port map( B1 => n7389, B2 => n9461, A => n7388, ZN => 
                           DP_OP_751_130_6421_n471);
   U7852 : INV_X1 port map( A => DP_OP_751_130_6421_n506, ZN => n7389);
   U7853 : NOR2_X1 port map( A1 => n8454, A2 => n9130, ZN => n7390);
   U7854 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1387, B => n7390, Z => 
                           DP_OP_751_130_6421_n1288);
   U7855 : NOR2_X1 port map( A1 => n8454, A2 => n9130, ZN => n7391);
   U7856 : MUX2_X1 port map( A => DP_OP_751_130_6421_n1323, B => 
                           DP_OP_751_130_6421_n1387, S => n7391, Z => 
                           DP_OP_751_130_6421_n1287);
   U7857 : NOR2_X1 port map( A1 => n9130, A2 => n7771, ZN => n7392);
   U7858 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1489, B => n7392, Z => 
                           DP_OP_751_130_6421_n1390);
   U7859 : NOR2_X1 port map( A1 => n9130, A2 => n7771, ZN => n7393);
   U7860 : MUX2_X1 port map( A => n7792, B => DP_OP_751_130_6421_n1489, S => 
                           n7393, Z => DP_OP_751_130_6421_n1389);
   U7861 : OAI21_X1 port map( B1 => n9240, B2 => n8188, A => n9220, ZN => n9362
                           );
   U7862 : OAI22_X1 port map( A1 => n8566, A2 => n7824, B1 => n9137, B2 => 
                           n7809, ZN => n9764);
   U7863 : OAI21_X1 port map( B1 => n7983, B2 => i_ALU_OP_2_port, A => n9242, 
                           ZN => n10097);
   U7864 : OAI21_X1 port map( B1 => n7827, B2 => n8188, A => n9229, ZN => n9670
                           );
   U7865 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n160, A2 => n8162, ZN =>
                           n7394);
   U7866 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n159, A2 => n7394, ZN =>
                           DP_OP_751_130_6421_n154);
   U7867 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_IN2_13_port, A2 => n8069,
                           B1 => DataPath_i_PIPLIN_B_13_port, B2 => n8136, ZN 
                           => n8227);
   U7868 : INV_X1 port map( A => n10441, ZN => n7395);
   U7869 : NAND2_X1 port map( A1 => IR_26_port, A2 => n8051, ZN => n7396);
   U7870 : OAI222_X1 port map( A1 => n10441, A2 => n10392, B1 => n10441, B2 => 
                           n10377, C1 => n7395, C2 => n7396, ZN => n8592);
   U7871 : AOI22_X1 port map( A1 => n8283, A2 => i_SEL_LGET_0_port, B1 => 
                           i_SEL_LGET_1_port, B2 => n493, ZN => n7397);
   U7872 : AOI22_X1 port map( A1 => i_SEL_LGET_0_port, A2 => n492, B1 => n7397,
                           B2 => n8319, ZN => n7398);
   U7873 : NOR2_X1 port map( A1 => n493, A2 => n219, ZN => n7399);
   U7874 : OAI221_X1 port map( B1 => n492, B2 => n7399, C1 => n8319, C2 => 
                           n8332, A => n8283, ZN => n7400);
   U7875 : NAND2_X1 port map( A1 => n219, A2 => n7398, ZN => n7401);
   U7876 : AOI21_X1 port map( B1 => n7401, B2 => n7400, A => n217, ZN => n7402)
                           ;
   U7877 : AOI211_X1 port map( C1 => n11878, C2 => n10036, A => n9130, B => 
                           n8020, ZN => n7403);
   U7878 : OAI21_X1 port map( B1 => n11858, B2 => n10088, A => n7596, ZN => 
                           n7404);
   U7879 : AOI221_X1 port map( B1 => n8020, B2 => n7404, C1 => n10082, C2 => 
                           n7404, A => n9060, ZN => n7405);
   U7880 : AOI211_X1 port map( C1 => n10035, C2 => 
                           DataPath_ALUhw_MULT_mux_out_0_0_port, A => n7403, B 
                           => n7405, ZN => n7406);
   U7881 : OAI211_X1 port map( C1 => n7998, C2 => DP_OP_751_130_6421_n1765, A 
                           => n10094, B => DP_OP_751_130_6421_n174, ZN => n7407
                           );
   U7882 : OAI211_X1 port map( C1 => n11859, C2 => n9149, A => n7406, B => 
                           n7407, ZN => n7408);
   U7883 : AOI22_X1 port map( A1 => n7796, A2 => n7402, B1 => n10429, B2 => 
                           n7408, ZN => n7409);
   U7884 : OAI22_X1 port map( A1 => n9135, A2 => n10059, B1 => n9975, B2 => 
                           n10046, ZN => n7410);
   U7885 : NOR2_X1 port map( A1 => n9885, A2 => n9977, ZN => n7411);
   U7886 : OAI21_X1 port map( B1 => n8438, B2 => n9548, A => n9586, ZN => n7412
                           );
   U7887 : OAI21_X1 port map( B1 => n9130, B2 => n9505, A => n7412, ZN => n7413
                           );
   U7888 : AOI21_X1 port map( B1 => n7806, B2 => n7789, A => n9708, ZN => n7414
                           );
   U7889 : AOI21_X1 port map( B1 => n11853, B2 => n7789, A => n9047, ZN => 
                           n7415);
   U7890 : OAI22_X1 port map( A1 => n9528, A2 => n7414, B1 => n9264, B2 => 
                           n7415, ZN => n7416);
   U7891 : AOI211_X1 port map( C1 => n9550, C2 => n9045, A => n7413, B => n7416
                           , ZN => n7417);
   U7892 : OAI22_X1 port map( A1 => n10104, A2 => n7417, B1 => n9134, B2 => 
                           n10066, ZN => n7418);
   U7893 : AOI211_X1 port map( C1 => n9150, C2 => n10112, A => n7411, B => 
                           n7418, ZN => n7419);
   U7894 : AOI22_X1 port map( A1 => n9972, A2 => n10430, B1 => n10117, B2 => 
                           n9247, ZN => n7420);
   U7895 : OAI211_X1 port map( C1 => n9153, C2 => n10002, A => n7419, B => 
                           n7420, ZN => n7421);
   U7896 : OAI21_X1 port map( B1 => n7410, B2 => n7421, A => n10428, ZN => 
                           n7422);
   U7897 : OAI211_X1 port map( C1 => n494, C2 => n11884, A => n7409, B => n7422
                           , ZN => n7020);
   U7898 : XOR2_X1 port map( A => n8275, B => n10316, Z => n7423);
   U7899 : INV_X1 port map( A => n10317, ZN => n7424);
   n7425 <= '0';
   U7901 : OAI222_X1 port map( A1 => n7426, A2 => n7757, B1 => n8275, B2 => 
                           n10367, C1 => n10318, C2 => n11845, ZN => n7040);
   U7902 : AND2_X1 port map( A1 => n8570, A2 => 
                           DataPath_RF_internal_out2_13_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N17);
   U7903 : AND2_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_internal_out1_14_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N18);
   U7904 : XOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_15_port, B => 
                           n7774, Z => n7427);
   U7905 : OAI22_X1 port map( A1 => n7751, A2 => n7309, B1 => n7726, B2 => 
                           n9784, ZN => n7428);
   U7906 : XOR2_X1 port map( A => n8148, B => n7428, Z => n7429);
   U7907 : XOR2_X1 port map( A => n7427, B => n7429, Z => 
                           DP_OP_751_130_6421_n1670);
   U7908 : NOR2_X1 port map( A1 => n7427, A2 => n7429, ZN => 
                           DP_OP_751_130_6421_n1669);
   U7909 : INV_X1 port map( A => DP_OP_751_130_6421_n1459, ZN => n7430);
   U7910 : INV_X1 port map( A => DP_OP_751_130_6421_n1409, ZN => n7431);
   U7911 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1409, B2 => 
                           DP_OP_751_130_6421_n1459, A => 
                           DP_OP_751_130_6421_n1458, ZN => n7432);
   U7912 : OAI21_X1 port map( B1 => n7430, B2 => n7431, A => n7432, ZN => 
                           DP_OP_751_130_6421_n1359);
   U7913 : INV_X1 port map( A => DP_OP_751_130_6421_n1055, ZN => n7433);
   U7914 : INV_X1 port map( A => DP_OP_751_130_6421_n1003, ZN => n7434);
   U7915 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1003, B2 => 
                           DP_OP_751_130_6421_n1055, A => 
                           DP_OP_751_130_6421_n1054, ZN => n7435);
   U7916 : OAI21_X1 port map( B1 => n7433, B2 => n7434, A => n7435, ZN => 
                           DP_OP_751_130_6421_n955);
   U7917 : OAI22_X1 port map( A1 => n9822, A2 => n9081, B1 => n7770, B2 => 
                           n8401, ZN => n7436);
   U7918 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1221, B => n7436, Z => 
                           DP_OP_751_130_6421_n1208);
   U7919 : NAND2_X1 port map( A1 => n9461, A2 => n9441, ZN => n7437);
   U7920 : OAI221_X1 port map( B1 => n9914, B2 => n9461, C1 => n9441, C2 => 
                           DP_OP_751_130_6421_n405, A => n7437, ZN => n9117);
   U7921 : INV_X1 port map( A => n10436, ZN => n7438);
   U7922 : NOR4_X1 port map( A1 => n11996, A2 => n8593, A3 => n11993, A4 => 
                           n7438, ZN => n8378);
   U7923 : INV_X1 port map( A => n8996, ZN => n7439);
   U7924 : AOI21_X1 port map( B1 => n7897, B2 => n11861, A => n7439, ZN => 
                           n9477);
   U7925 : OAI211_X1 port map( C1 => n7809, C2 => n7875, A => n11879, B => 
                           n9369, ZN => n7440);
   U7926 : INV_X1 port map( A => n7440, ZN => n9428);
   U7927 : AOI22_X2 port map( A1 => n7618, A2 => DataPath_i_PIPLIN_A_8_port, B1
                           => DataPath_i_PIPLIN_IN1_8_port, B2 => n8225, ZN => 
                           n8435);
   U7928 : OAI22_X1 port map( A1 => n8134, A2 => n9133, B1 => n7726, B2 => 
                           n9168, ZN => n7441);
   U7929 : XNOR2_X1 port map( A => n8148, B => n7441, ZN => 
                           DP_OP_751_130_6421_n1762);
   U7930 : INV_X1 port map( A => DP_OP_751_130_6421_n877, ZN => n7442);
   U7931 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n877, B2 => 
                           DP_OP_751_130_6421_n813, A => 
                           DP_OP_751_130_6421_n812, ZN => n7443);
   U7932 : OAI21_X1 port map( B1 => n7794, B2 => n7442, A => n7443, ZN => 
                           DP_OP_751_130_6421_n777);
   U7933 : INV_X1 port map( A => DP_OP_751_130_6421_n1016, ZN => n7444);
   U7934 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1017, B2 => 
                           DP_OP_751_130_6421_n1016, A => 
                           DP_OP_751_130_6421_n1081, ZN => n7445);
   U7935 : OAI21_X1 port map( B1 => n7444, B2 => n8563, A => n7445, ZN => 
                           DP_OP_751_130_6421_n981);
   U7936 : OR3_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_25_port, A3 => n7871, ZN
                           => n7868);
   U7937 : OAI21_X1 port map( B1 => n8107, B2 => n8109, A => 
                           DP_OP_1091J1_126_6973_n6, ZN => n7446);
   U7938 : NAND3_X1 port map( A1 => n8104, A2 => n8105, A3 => n7446, ZN => 
                           n7447);
   U7939 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_29_port, ZN => n7448);
   U7940 : XNOR2_X1 port map( A => n7448, B => n7447, ZN => C620_DATA2_29);
   U7941 : INV_X1 port map( A => DP_OP_751_130_6421_n123, ZN => n7449);
   U7942 : AOI21_X1 port map( B1 => DP_OP_751_130_6421_n124, B2 => n8163, A => 
                           n7449, ZN => DP_OP_751_130_6421_n119);
   U7943 : NOR2_X1 port map( A1 => n9249, A2 => n9248, ZN => n9259);
   U7944 : NAND2_X1 port map( A1 => n8222, A2 => intadd_1_n15, ZN => n7450);
   U7945 : NAND2_X1 port map( A1 => intadd_1_n12, A2 => n7450, ZN => 
                           intadd_1_n6);
   U7946 : NOR2_X1 port map( A1 => n9250, A2 => n9252, ZN => n7451);
   U7947 : XOR2_X1 port map( A => n7451, B => n11862, Z => n7452);
   U7948 : NOR2_X1 port map( A1 => n9251, A2 => n7451, ZN => n7453);
   U7949 : AOI211_X1 port map( C1 => n9251, C2 => n7451, A => n9993, B => n7453
                           , ZN => n7454);
   U7950 : AOI22_X1 port map( A1 => n7795, A2 => n10088, B1 => n10035, B2 => 
                           n9240, ZN => n7455);
   U7951 : INV_X1 port map( A => DP_OP_751_130_6421_n148, ZN => n7456);
   U7952 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n147, A2 => n7456, ZN => 
                           n7457);
   U7953 : XNOR2_X1 port map( A => n7457, B => DP_OP_751_130_6421_n149, ZN => 
                           n7458);
   U7954 : AOI22_X1 port map( A1 => n9889, A2 => n10112, B1 => n10113, B2 => 
                           n9247, ZN => n7459);
   U7955 : OAI22_X1 port map( A1 => n10040, A2 => n10106, B1 => n9868, B2 => 
                           n9977, ZN => n7460);
   U7956 : OAI22_X1 port map( A1 => n9884, A2 => n10002, B1 => n9267, B2 => 
                           n10056, ZN => n7461);
   U7957 : AOI211_X1 port map( C1 => n10045, C2 => n9971, A => n7460, B => 
                           n7461, ZN => n7462);
   U7958 : AOI22_X1 port map( A1 => n11866, A2 => n10116, B1 => n10120, B2 => 
                           n9890, ZN => n7463);
   U7959 : NAND3_X1 port map( A1 => n7459, A2 => n7462, A3 => n7463, ZN => 
                           n7464);
   U7960 : AOI22_X1 port map( A1 => n10094, A2 => n7458, B1 => n9897, B2 => 
                           n7464, ZN => n7465);
   U7961 : OAI221_X1 port map( B1 => n9240, B2 => n10033, C1 => n7795, C2 => 
                           n10088, A => n9241, ZN => n7466);
   U7962 : OAI211_X1 port map( C1 => n7455, C2 => n9241, A => n7465, B => n7466
                           , ZN => n7467);
   U7963 : AOI211_X1 port map( C1 => n10426, C2 => n7452, A => n7454, B => 
                           n7467, ZN => n7468);
   U7964 : OAI22_X1 port map( A1 => n11885, A2 => n7468, B1 => n497, B2 => 
                           n11884, ZN => n7016);
   U7965 : INV_X1 port map( A => n10230, ZN => n7469);
   U7966 : NOR3_X1 port map( A1 => n10229, A2 => n8281, A3 => n7469, ZN => n143
                           );
   U7967 : INV_X1 port map( A => n10324, ZN => n7470);
   U7968 : OAI21_X1 port map( B1 => n10339, B2 => n8236, A => n7470, ZN => 
                           n7471);
   U7969 : XOR2_X1 port map( A => n10325, B => n7471, Z => n7472);
   U7970 : AOI22_X1 port map( A1 => n10417, A2 => IRAM_ADDRESS_19_port, B1 => 
                           i_RD1_19_port, B2 => n10418, ZN => n7473);
   U7971 : OAI21_X1 port map( B1 => n7757, B2 => n7472, A => n7473, ZN => n7042
                           );
   U7972 : AND2_X1 port map( A1 => n8574, A2 => 
                           DataPath_RF_internal_out2_14_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N18);
   U7973 : AND2_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_internal_out1_13_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N17);
   U7974 : INV_X1 port map( A => DP_OP_751_130_6421_n1714, ZN => n7474);
   U7975 : NOR2_X1 port map( A1 => n7908, A2 => n7474, ZN => 
                           DP_OP_751_130_6421_n1659);
   U7976 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1703, B => 
                           DP_OP_751_130_6421_n1733, Z => 
                           DP_OP_751_130_6421_n1638);
   U7977 : OAI22_X1 port map( A1 => n7771, A2 => n7981, B1 => n8452, B2 => 
                           n8428, ZN => n7475);
   U7978 : XOR2_X1 port map( A => n8144, B => n7475, Z => 
                           DP_OP_751_130_6421_n1410);
   U7979 : AOI22_X1 port map( A1 => n8148, A2 => 
                           DataPath_ALUhw_MULT_mux_out_0_12_port, B1 => 
                           DP_OP_751_130_6421_n1787, B2 => n7837, ZN => n7476);
   U7980 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_12_port, B => 
                           n8146, ZN => n7477);
   U7981 : NOR2_X1 port map( A1 => n7476, A2 => n7477, ZN => 
                           DP_OP_751_130_6421_n1675);
   U7982 : XOR2_X1 port map( A => n7476, B => n7477, Z => 
                           DP_OP_751_130_6421_n1676);
   U7983 : NAND2_X1 port map( A1 => n10475, A2 => n10482, ZN => n7478);
   U7984 : OAI21_X1 port map( B1 => n7478, B2 => n10478, A => n10479, ZN => 
                           n10480);
   U7985 : AOI22_X1 port map( A1 => n825, A2 => DataPath_RF_c_win_0_port, B1 =>
                           n824, B2 => DataPath_RF_c_win_4_port, ZN => n8220);
   U7986 : INV_X1 port map( A => DP_OP_751_130_6421_n467, ZN => n7479);
   U7987 : INV_X1 port map( A => DP_OP_751_130_6421_n403, ZN => n7480);
   U7988 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n467, B2 => 
                           DP_OP_751_130_6421_n403, A => 
                           DP_OP_751_130_6421_n466, ZN => n7481);
   U7989 : OAI21_X1 port map( B1 => n7479, B2 => n7480, A => n7481, ZN => 
                           DP_OP_751_130_6421_n367);
   U7990 : OAI22_X1 port map( A1 => n9105, A2 => n8399, B1 => n9104, B2 => 
                           n9168, ZN => n7482);
   U7991 : XOR2_X1 port map( A => DP_OP_751_130_6421_n711, B => n7482, Z => 
                           DP_OP_751_130_6421_n707);
   U7992 : AOI22_X1 port map( A1 => n7803, A2 => n9823, B1 => 
                           DP_OP_751_130_6421_n1221, B2 => 
                           DP_OP_751_130_6421_n1323, ZN => n7483);
   U7993 : OAI21_X1 port map( B1 => n9823, B2 => DP_OP_751_130_6421_n1221, A =>
                           n7483, ZN => n9080);
   U7994 : AOI21_X1 port map( B1 => IRAM_ADDRESS_20_port, B2 => n10319, A => 
                           n7936, ZN => n7859);
   U7995 : INV_X1 port map( A => n8175, ZN => n7484);
   U7996 : AOI221_X1 port map( B1 => DataPath_WRF_CUhw_curr_addr_29_port, B2 =>
                           DataPath_WRF_CUhw_curr_addr_30_port, C1 => n7484, C2
                           => DataPath_WRF_CUhw_curr_addr_30_port, A => 
                           DP_OP_1091J1_126_6973_n31, ZN => n7485);
   U7997 : INV_X1 port map( A => n8170, ZN => n7486);
   U7998 : NAND2_X1 port map( A1 => n7485, A2 => n7486, ZN => n8132);
   U7999 : OAI21_X1 port map( B1 => n9656, B2 => n11869, A => n9373, ZN => 
                           n9426);
   U8000 : INV_X1 port map( A => n8431, ZN => n7487);
   U8001 : AOI21_X1 port map( B1 => n9060, B2 => n7487, A => n7774, ZN => 
                           DP_OP_751_130_6421_n1698);
   U8002 : AND2_X1 port map( A1 => n9060, A2 => n7487, ZN => 
                           DP_OP_751_130_6421_n1696);
   U8003 : INV_X1 port map( A => n8982, ZN => n7488);
   U8004 : AOI21_X1 port map( B1 => n7913, B2 => n11861, A => n7488, ZN => 
                           n9494);
   U8005 : AOI21_X1 port map( B1 => n7824, B2 => n7809, A => n9351, ZN => n7489
                           );
   U8006 : INV_X1 port map( A => n7489, ZN => n9348);
   U8007 : INV_X1 port map( A => n7869, ZN => n7490);
   U8008 : AOI22_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_26_port, B1 => n7867, B2
                           => n7490, ZN => n7865);
   U8009 : NAND2_X1 port map( A1 => n9531, A2 => n9544, ZN => n7491);
   U8010 : OAI211_X1 port map( C1 => n11879, C2 => n7805, A => n10103, B => 
                           n7491, ZN => n7492);
   U8011 : NOR2_X1 port map( A1 => n9264, A2 => n9658, ZN => n7493);
   U8012 : OAI22_X1 port map( A1 => n9531, A2 => n9546, B1 => n9704, B2 => 
                           n7493, ZN => n7494);
   U8013 : OAI221_X1 port map( B1 => n9586, B2 => n9548, C1 => n9586, C2 => 
                           n7788, A => n9549, ZN => n7495);
   U8014 : NAND3_X1 port map( A1 => n7492, A2 => n7494, A3 => n7495, ZN => 
                           n7496);
   U8015 : AOI21_X1 port map( B1 => n9550, B2 => n9730, A => n7496, ZN => 
                           n10039);
   U8016 : NOR2_X1 port map( A1 => n8250, A2 => n7929, ZN => n7497);
   U8017 : AOI21_X1 port map( B1 => DataPath_i_PIPLIN_IN2_17_port, B2 => n8137,
                           A => n7497, ZN => n8563);
   U8018 : AOI22_X1 port map( A1 => n7853, A2 => n8921, B1 => n7852, B2 => 
                           n8920, ZN => n7498);
   U8019 : INV_X1 port map( A => n7849, ZN => n7499);
   U8020 : NAND2_X1 port map( A1 => n7498, A2 => n7499, ZN => intadd_1_n23);
   U8021 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_2_port, Z => n7500);
   U8022 : OAI21_X1 port map( B1 => n7601, B2 => n7500, A => n10443, ZN => 
                           n7501);
   U8023 : AOI21_X1 port map( B1 => n7601, B2 => n7500, A => n7501, ZN => 
                           DRAMRF_ADDRESS_2_port);
   U8024 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_25_port, Z => n7502);
   U8025 : NAND2_X1 port map( A1 => n8032, A2 => n7872, ZN => n7503);
   U8026 : OAI21_X1 port map( B1 => n7502, B2 => n7503, A => n10443, ZN => 
                           n7504);
   U8027 : AOI21_X1 port map( B1 => n7502, B2 => n7503, A => n7504, ZN => 
                           DRAMRF_ADDRESS_25_port);
   U8028 : AOI22_X1 port map( A1 => n8136, A2 => DataPath_i_PIPLIN_B_10_port, 
                           B1 => DataPath_i_PIPLIN_IN2_10_port, B2 => n8069, ZN
                           => n7505);
   U8029 : INV_X1 port map( A => n7505, ZN => n9872);
   U8030 : NOR2_X1 port map( A1 => n7898, A2 => DP_OP_751_130_6421_n1527, ZN =>
                           n7506);
   U8031 : AOI21_X1 port map( B1 => DP_OP_751_130_6421_n1527, B2 => n7898, A =>
                           n7506, ZN => n7507);
   U8032 : AOI22_X1 port map( A1 => n9247, A2 => n10045, B1 => n10121, B2 => 
                           n9889, ZN => n7508);
   U8033 : NAND2_X1 port map( A1 => n10120, A2 => n11866, ZN => n7509);
   U8034 : OAI21_X1 port map( B1 => n9868, B2 => n10046, A => n7509, ZN => 
                           n7510);
   U8035 : AOI21_X1 port map( B1 => n9865, B2 => n10117, A => n7510, ZN => 
                           n7511);
   U8036 : AOI22_X1 port map( A1 => n10430, A2 => n10043, B1 => n10110, B2 => 
                           n10044, ZN => n7512);
   U8037 : AOI22_X1 port map( A1 => n10112, A2 => n9890, B1 => n10113, B2 => 
                           n9972, ZN => n7513);
   U8038 : NAND4_X1 port map( A1 => n7508, A2 => n7511, A3 => n7512, A4 => 
                           n7513, ZN => n7514);
   U8039 : AOI222_X1 port map( A1 => n10088, A2 => n7507, B1 => n7506, B2 => 
                           n10033, C1 => n7514, C2 => n9897, ZN => n7515);
   U8040 : NAND2_X1 port map( A1 => n8161, A2 => DP_OP_751_130_6421_n145, ZN =>
                           n7516);
   U8041 : XNOR2_X1 port map( A => n7516, B => DP_OP_751_130_6421_n146, ZN => 
                           n7517);
   U8042 : INV_X1 port map( A => n9258, ZN => n7518);
   U8043 : NOR2_X1 port map( A1 => n9259, A2 => n7518, ZN => n7519);
   U8044 : OAI21_X1 port map( B1 => n9250, B2 => n11862, A => n9257, ZN => 
                           n7520);
   U8045 : XNOR2_X1 port map( A => n7520, B => n7519, ZN => n7521);
   U8046 : AOI22_X1 port map( A1 => n7517, A2 => n10094, B1 => n7521, B2 => 
                           n10426, ZN => n7522);
   U8047 : NOR2_X1 port map( A1 => n9252, A2 => n9254, ZN => n7523);
   U8048 : AOI21_X1 port map( B1 => n7519, B2 => n7523, A => n9993, ZN => n7524
                           );
   U8049 : OAI21_X1 port map( B1 => n7519, B2 => n7523, A => n7524, ZN => n7525
                           );
   U8050 : NAND3_X1 port map( A1 => n7898, A2 => DP_OP_751_130_6421_n1527, A3 
                           => n10035, ZN => n7526);
   U8051 : NAND4_X1 port map( A1 => n7515, A2 => n7522, A3 => n7525, A4 => 
                           n7526, ZN => n7527);
   U8052 : AOI22_X1 port map( A1 => DRAM_ADDRESS_7_port, A2 => n7791, B1 => 
                           n10429, B2 => n7527, ZN => n1998);
   U8053 : AOI22_X1 port map( A1 => IRAM_ADDRESS_1_port, A2 => n10417, B1 => 
                           n10418, B2 => i_RD1_1_port, ZN => n7528);
   U8054 : INV_X1 port map( A => intadd_0_n19, ZN => n7529);
   U8055 : NOR2_X1 port map( A1 => intadd_0_n18, A2 => n7529, ZN => n7530);
   U8056 : XOR2_X1 port map( A => n7594, B => n7530, Z => n7531);
   U8057 : OAI21_X1 port map( B1 => n7757, B2 => n7531, A => n7528, ZN => n7060
                           );
   U8058 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_30_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N34);
   U8059 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_28_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N32);
   U8060 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_27_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N31);
   U8061 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_26_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N30);
   U8062 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_25_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N29);
   U8063 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_24_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N28);
   U8064 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_23_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N27);
   U8065 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_22_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N26);
   U8066 : AND2_X1 port map( A1 => n8573, A2 => 
                           DataPath_RF_internal_out2_21_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N25);
   U8067 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_20_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N24);
   U8068 : AND2_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_internal_out2_11_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N15);
   U8069 : AND2_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_internal_out2_10_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N14);
   U8070 : AND2_X1 port map( A1 => n8579, A2 => 
                           DataPath_RF_internal_out2_9_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N13);
   U8071 : AND2_X1 port map( A1 => n8578, A2 => 
                           DataPath_RF_internal_out2_8_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N12);
   U8072 : AND2_X1 port map( A1 => n8572, A2 => 
                           DataPath_RF_internal_out2_7_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N11);
   U8073 : AND2_X1 port map( A1 => n8574, A2 => 
                           DataPath_RF_internal_out2_6_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N10);
   U8074 : AND2_X1 port map( A1 => n8580, A2 => 
                           DataPath_RF_internal_out2_5_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N9);
   U8075 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_4_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N8);
   U8076 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_3_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N7);
   U8077 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_2_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N6);
   U8078 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_1_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N5);
   U8079 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_0_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N4);
   U8080 : NOR2_X1 port map( A1 => n10390, A2 => n143, ZN => n7532);
   U8081 : NAND2_X1 port map( A1 => n10421, A2 => n7532, ZN => 
                           CU_I_CW_RF_RD2_EN_port);
   U8082 : AND2_X1 port map( A1 => n8570, A2 => 
                           DataPath_RF_internal_out1_12_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N16);
   U8083 : AND2_X1 port map( A1 => n8576, A2 => 
                           DataPath_RF_internal_out1_31_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N35);
   U8084 : OAI22_X1 port map( A1 => n7616, A2 => n9495, B1 => n8450, B2 => 
                           n7776, ZN => n7533);
   U8085 : XOR2_X1 port map( A => n7797, B => n7533, Z => 
                           DP_OP_751_130_6421_n1507);
   U8086 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1549, B2 => 
                           DP_OP_751_130_6421_n1505, A => 
                           DP_OP_751_130_6421_n1548, ZN => n7992);
   U8087 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1657, B2 => 
                           DP_OP_751_130_6421_n1610, A => n7954, ZN => n7953);
   U8088 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1667, B2 => 
                           DP_OP_751_130_6421_n1615, A => 
                           DP_OP_751_130_6421_n1666, ZN => n8058);
   U8089 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1347, B2 => 
                           DP_OP_751_130_6421_n1302, A => 
                           DP_OP_751_130_6421_n1346, ZN => n7878);
   U8090 : INV_X1 port map( A => DP_OP_751_130_6421_n1053, ZN => n7534);
   U8091 : INV_X1 port map( A => DP_OP_751_130_6421_n1002, ZN => n7535);
   U8092 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1002, B2 => 
                           DP_OP_751_130_6421_n1053, A => 
                           DP_OP_751_130_6421_n1052, ZN => n7536);
   U8093 : OAI21_X1 port map( B1 => n7534, B2 => n7535, A => n7536, ZN => 
                           DP_OP_751_130_6421_n953);
   U8094 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n857, B2 => 
                           DP_OP_751_130_6421_n802, A => 
                           DP_OP_751_130_6421_n856, ZN => n7537);
   U8095 : OAI21_X1 port map( B1 => n7538, B2 => n7539, A => n7537, ZN => 
                           DP_OP_751_130_6421_n757);
   U8096 : INV_X1 port map( A => DP_OP_751_130_6421_n857, ZN => n7538);
   U8097 : INV_X1 port map( A => DP_OP_751_130_6421_n802, ZN => n7539);
   U8098 : INV_X1 port map( A => n10477, ZN => n7540);
   U8099 : AOI221_X1 port map( B1 => n10475, B2 => n7540, C1 => n10478, C2 => 
                           n7540, A => n10476, ZN => n7541);
   U8100 : AOI221_X1 port map( B1 => n7541, B2 => n10450, C1 => n10451, C2 => 
                           n10450, A => n10447, ZN => n7542);
   U8101 : NOR2_X1 port map( A1 => n7542, A2 => n10452, ZN => n10496);
   U8102 : AOI22_X1 port map( A1 => n8242, A2 => DataPath_RF_c_win_3_port, B1 
                           => n826, B2 => DataPath_RF_c_win_1_port, ZN => n7543
                           );
   U8103 : OAI21_X1 port map( B1 => n826, B2 => DataPath_RF_c_win_1_port, A => 
                           n7543, ZN => n8377);
   U8104 : AOI211_X1 port map( C1 => n11868, C2 => n7875, A => n11850, B => 
                           n8969, ZN => n9214);
   U8105 : NOR3_X1 port map( A1 => n10267, A2 => n10279, A3 => 
                           IRAM_ADDRESS_29_port, ZN => n8070);
   U8106 : OAI21_X1 port map( B1 => DataPath_WRF_CUhw_curr_addr_28_port, B2 => 
                           DP_OP_1091J1_126_6973_n31, A => 
                           DataPath_WRF_CUhw_curr_addr_29_port, ZN => n7544);
   U8107 : INV_X1 port map( A => n7544, ZN => n8120);
   U8108 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n366, A2 => 
                           DP_OP_751_130_6421_n268, ZN => n8078);
   U8109 : NOR2_X1 port map( A1 => n9095, A2 => n9130, ZN => n7545);
   U8110 : XOR2_X1 port map( A => DP_OP_751_130_6421_n979, B => n7545, Z => 
                           DP_OP_751_130_6421_n880);
   U8111 : NOR2_X1 port map( A1 => n9095, A2 => n9130, ZN => n7546);
   U8112 : MUX2_X1 port map( A => n8149, B => DP_OP_751_130_6421_n979, S => 
                           n7546, Z => DP_OP_751_130_6421_n879);
   U8113 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1697, B => 
                           DP_OP_751_130_6421_n1760, Z => 
                           DP_OP_751_130_6421_n1692);
   U8114 : AOI22_X1 port map( A1 => DataPath_i_PIPLIN_A_2_port, A2 => n7618, B1
                           => DataPath_i_PIPLIN_IN1_2_port, B2 => n8225, ZN => 
                           n7547);
   U8115 : INV_X1 port map( A => n7547, ZN => n9156);
   U8116 : OAI21_X1 port map( B1 => n7821, B2 => DP_OP_751_130_6421_n404, A => 
                           DP_OP_751_130_6421_n469, ZN => n7548);
   U8117 : OAI21_X1 port map( B1 => n7549, B2 => n9914, A => n7548, ZN => 
                           DP_OP_751_130_6421_n369);
   U8118 : INV_X1 port map( A => DP_OP_751_130_6421_n404, ZN => n7549);
   U8119 : NOR2_X1 port map( A1 => n9317, A2 => n9936, ZN => n9319);
   U8120 : OAI21_X1 port map( B1 => n9333, B2 => n11869, A => n9334, ZN => 
                           n9365);
   U8121 : INV_X1 port map( A => n9011, ZN => n7550);
   U8122 : AOI21_X1 port map( B1 => n9137, B2 => n11861, A => n7550, ZN => 
                           n9533);
   U8123 : AOI22_X1 port map( A1 => n10081, A2 => n9547, B1 => n9585, B2 => 
                           n9657, ZN => n7551);
   U8124 : AOI22_X1 port map( A1 => n9602, A2 => n9542, B1 => n9583, B2 => 
                           n9762, ZN => n7552);
   U8125 : AOI22_X1 port map( A1 => n10100, A2 => n9704, B1 => n9582, B2 => 
                           n9469, ZN => n7553);
   U8126 : NAND3_X1 port map( A1 => n7788, A2 => n8229, A3 => n9584, ZN => 
                           n7554);
   U8127 : AND4_X1 port map( A1 => n7551, A2 => n7552, A3 => n7553, A4 => n7554
                           , ZN => n10105);
   U8128 : OAI21_X1 port map( B1 => n9303, B2 => n8406, A => n10047, ZN => 
                           n9741);
   U8129 : NOR2_X1 port map( A1 => n9298, A2 => n7727, ZN => n9777);
   U8130 : NAND2_X1 port map( A1 => n8160, A2 => DP_OP_751_130_6421_n138, ZN =>
                           n7555);
   U8131 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n137, A2 => n7555, ZN =>
                           DP_OP_751_130_6421_n132);
   U8132 : OAI22_X1 port map( A1 => n7750, A2 => n9130, B1 => n9133, B2 => 
                           n7726, ZN => n7556);
   U8133 : XNOR2_X1 port map( A => n8147, B => n7556, ZN => 
                           DP_OP_751_130_6421_n170);
   U8134 : INV_X1 port map( A => n9822, ZN => n7557);
   U8135 : NOR2_X1 port map( A1 => n9295, A2 => n7557, ZN => n10029);
   U8136 : NOR2_X1 port map( A1 => n9302, A2 => n8438, ZN => n10051);
   U8137 : XOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_0_port, B => 
                           n7998, Z => DP_OP_751_130_6421_n1765);
   U8138 : INV_X1 port map( A => n11775, ZN => n7558);
   U8139 : NAND4_X1 port map( A1 => n8224, A2 => n10160, A3 => IR_3_port, A4 =>
                           n7558, ZN => n10155);
   U8140 : OAI21_X1 port map( B1 => n10261, B2 => n172, A => n10263, ZN => 
                           n10319);
   U8141 : AOI21_X1 port map( B1 => IRAM_ADDRESS_8_port, B2 => n7846, A => 
                           n7610, ZN => n7559);
   U8142 : NOR2_X1 port map( A1 => n7846, A2 => n7609, ZN => n7560);
   U8143 : OAI21_X1 port map( B1 => n10348, B2 => n7560, A => n7559, ZN => 
                           n8934);
   U8144 : AOI21_X1 port map( B1 => n8131, B2 => n7601, A => n8130, ZN => n7561
                           );
   U8145 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_3_port, ZN => n7562);
   U8146 : OAI21_X1 port map( B1 => n7561, B2 => n7562, A => n10443, ZN => 
                           n7563);
   U8147 : AOI21_X1 port map( B1 => n7561, B2 => n7562, A => n7563, ZN => 
                           DRAMRF_ADDRESS_3_port);
   U8148 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_9_port, ZN => n7564);
   U8149 : OAI21_X1 port map( B1 => n7744, B2 => n7564, A => n10443, ZN => 
                           n7565);
   U8150 : AOI21_X1 port map( B1 => n7744, B2 => n7564, A => n7565, ZN => 
                           DRAMRF_ADDRESS_9_port);
   U8151 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_10_port, Z => n7566);
   U8152 : OAI21_X1 port map( B1 => n7599, B2 => n7566, A => n10443, ZN => 
                           n7567);
   U8153 : AOI21_X1 port map( B1 => n7599, B2 => n7566, A => n7567, ZN => 
                           DRAMRF_ADDRESS_10_port);
   U8154 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_11_port, Z => n7568);
   U8155 : OAI21_X1 port map( B1 => n7598, B2 => n7568, A => n10443, ZN => 
                           n7569);
   U8156 : AOI21_X1 port map( B1 => n7598, B2 => n7568, A => n7569, ZN => 
                           DRAMRF_ADDRESS_11_port);
   U8157 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_13_port, Z => n7570);
   U8158 : OAI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n20, B2 => n7570, A 
                           => n10443, ZN => n7571);
   U8159 : AOI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n20, B2 => n7570, A 
                           => n7571, ZN => DRAMRF_ADDRESS_13_port);
   U8160 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_19_port, Z => n7572);
   U8161 : OAI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n14, B2 => n7572, A 
                           => n10443, ZN => n7573);
   U8162 : AOI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n14, B2 => n7572, A 
                           => n7573, ZN => DRAMRF_ADDRESS_19_port);
   U8163 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_20_port, Z => n7574);
   U8164 : OAI21_X1 port map( B1 => n7600, B2 => n7574, A => n10443, ZN => 
                           n7575);
   U8165 : AOI21_X1 port map( B1 => n7600, B2 => n7574, A => n7575, ZN => 
                           DRAMRF_ADDRESS_20_port);
   U8166 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_22_port, Z => n7576);
   U8167 : OAI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n11, B2 => n7576, A 
                           => n10443, ZN => n7577);
   U8168 : AOI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n11, B2 => n7576, A 
                           => n7577, ZN => DRAMRF_ADDRESS_22_port);
   U8169 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_24_port, ZN => n7578);
   U8170 : OAI21_X1 port map( B1 => n7725, B2 => n7578, A => n10443, ZN => 
                           n7579);
   U8171 : AOI21_X1 port map( B1 => n7725, B2 => n7578, A => n7579, ZN => 
                           DRAMRF_ADDRESS_24_port);
   U8172 : INV_X1 port map( A => n7868, ZN => n7580);
   U8173 : AOI21_X1 port map( B1 => n7869, B2 => n7872, A => n7580, ZN => n7581
                           );
   U8174 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_26_port, Z => n7582);
   U8175 : OAI21_X1 port map( B1 => n7581, B2 => n7582, A => n10443, ZN => 
                           n7583);
   U8176 : AOI21_X1 port map( B1 => n7581, B2 => n7582, A => n7583, ZN => 
                           DRAMRF_ADDRESS_26_port);
   U8177 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_27_port, Z => n7584);
   U8178 : OAI21_X1 port map( B1 => n7602, B2 => n7584, A => n10443, ZN => 
                           n7585);
   U8179 : AOI21_X1 port map( B1 => n7602, B2 => n7584, A => n7585, ZN => 
                           DRAMRF_ADDRESS_27_port);
   U8180 : NOR2_X1 port map( A1 => n8246, A2 => n8069, ZN => n7586);
   U8181 : AOI21_X1 port map( B1 => DataPath_i_PIPLIN_IN2_9_port, B2 => n7929, 
                           A => n7586, ZN => n7798);
   U8182 : NOR2_X1 port map( A1 => n159, A2 => n8418, ZN => n7587);
   U8183 : AOI21_X1 port map( B1 => IRAM_DATA(31), B2 => n8426, A => n7587, ZN 
                           => n8391);
   U8184 : INV_X1 port map( A => i_RD1_13_port, ZN => n7588);
   U8185 : NAND2_X1 port map( A1 => n10344, A2 => n10345, ZN => n7589);
   U8186 : AOI21_X1 port map( B1 => intadd_1_n23, B2 => n8267, A => intadd_1_n6
                           , ZN => n7590);
   U8187 : XNOR2_X1 port map( A => n7590, B => n7589, ZN => n7591);
   U8188 : OAI222_X1 port map( A1 => n7588, A2 => n11845, B1 => n8290, B2 => 
                           n10367, C1 => n7757, C2 => n7591, ZN => n7048);
   U8189 : NOR3_X1 port map( A1 => n10389, A2 => n10401, A3 => n10390, ZN => 
                           n7592);
   U8190 : OAI221_X1 port map( B1 => IR_26_port, B2 => n10372, C1 => n8223, C2 
                           => n10383, A => n7592, ZN => CU_I_CW_SEL_CMPB_port);
   U8191 : AND2_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_internal_out2_12_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N16);
   U8192 : AND2_X1 port map( A1 => n8570, A2 => 
                           DataPath_RF_internal_out1_30_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N34);
   U8193 : AND2_X1 port map( A1 => n8579, A2 => 
                           DataPath_RF_internal_out1_28_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N32);
   U8194 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out1_27_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N31);
   U8195 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out1_26_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N30);
   U8196 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out1_25_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N29);
   U8197 : AND2_X1 port map( A1 => n8580, A2 => 
                           DataPath_RF_internal_out1_24_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N28);
   U8198 : AND2_X1 port map( A1 => n8573, A2 => 
                           DataPath_RF_internal_out1_23_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N27);
   U8199 : AND2_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_internal_out1_22_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N26);
   U8200 : AND2_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_internal_out1_21_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N25);
   U8201 : AND2_X1 port map( A1 => n8579, A2 => 
                           DataPath_RF_internal_out1_20_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N24);
   U8202 : AND2_X1 port map( A1 => n8574, A2 => 
                           DataPath_RF_internal_out1_11_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N15);
   U8203 : AND2_X1 port map( A1 => n8571, A2 => 
                           DataPath_RF_internal_out1_10_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N14);
   U8204 : AND2_X1 port map( A1 => n8578, A2 => 
                           DataPath_RF_internal_out1_9_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N13);
   U8205 : AND2_X1 port map( A1 => n8577, A2 => 
                           DataPath_RF_internal_out1_8_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N12);
   U8206 : AND2_X1 port map( A1 => n8576, A2 => 
                           DataPath_RF_internal_out1_7_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N11);
   U8207 : AND2_X1 port map( A1 => n8580, A2 => 
                           DataPath_RF_internal_out1_6_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N10);
   U8208 : AND2_X1 port map( A1 => n8582, A2 => 
                           DataPath_RF_internal_out1_5_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N9);
   U8209 : AND2_X1 port map( A1 => n8574, A2 => 
                           DataPath_RF_internal_out1_4_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N8);
   U8210 : AND2_X1 port map( A1 => n8581, A2 => 
                           DataPath_RF_internal_out1_3_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N7);
   U8211 : AND2_X1 port map( A1 => n8570, A2 => 
                           DataPath_RF_internal_out1_2_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N6);
   U8212 : AND2_X1 port map( A1 => n8574, A2 => 
                           DataPath_RF_internal_out1_1_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N5);
   U8213 : AND2_X1 port map( A1 => n8578, A2 => 
                           DataPath_RF_internal_out1_0_port, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N4);
   U8214 : NOR2_X1 port map( A1 => n10231, A2 => n10395, ZN => n7593);
   U8215 : AOI21_X1 port map( B1 => n7593, B2 => n10221, A => n11753, ZN => 
                           CU_I_CW_IF_MEM_EN_port);
   U8216 : AND2_X1 port map( A1 => n8575, A2 => 
                           DataPath_RF_internal_out2_31_port, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N35);
   U8217 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_27_port, A2 => n8555, 
                           ZN => n9473);
   U8218 : NOR2_X1 port map( A1 => n7652, A2 => n7653, ZN => 
                           DP_OP_751_130_6421_n1663);
   U8219 : OR2_X2 port map( A1 => n10369, A2 => n211, ZN => n7594);
   U8220 : BUF_X1 port map( A => n9165, Z => n8004);
   U8221 : BUF_X1 port map( A => DP_OP_751_130_6421_n470, Z => n7595);
   U8222 : INV_X1 port map( A => n8359, ZN => n7596);
   U8223 : OR2_X1 port map( A1 => IRAM_ADDRESS_29_port, A2 => n10278, ZN => 
                           n7597);
   U8224 : BUF_X1 port map( A => DP_OP_1091J1_126_6973_n22, Z => n7598);
   U8225 : BUF_X1 port map( A => DP_OP_1091J1_126_6973_n23, Z => n7599);
   U8226 : BUF_X1 port map( A => DP_OP_1091J1_126_6973_n13, Z => n7600);
   U8227 : BUF_X1 port map( A => n8143, Z => n7601);
   U8228 : BUF_X1 port map( A => DP_OP_1091J1_126_6973_n6, Z => n7602);
   U8229 : OAI211_X1 port map( C1 => n8202, C2 => n8389, A => n7855, B => n7607
                           , ZN => n7603);
   U8230 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1724, B => 
                           DP_OP_751_130_6421_n1754, Z => 
                           DP_OP_751_130_6421_n1680);
   U8231 : BUF_X1 port map( A => DP_OP_751_130_6421_n96, Z => n7605);
   U8232 : AND2_X1 port map( A1 => IR_29_port, A2 => n10149, ZN => n8354);
   U8233 : NAND2_X1 port map( A1 => n8103, A2 => n8101, ZN => n10282);
   U8234 : AND2_X1 port map( A1 => n8103, A2 => n8100, ZN => n10289);
   U8235 : OAI21_X1 port map( B1 => n8139, B2 => n10236, A => n10235, ZN => 
                           n10340);
   U8236 : OR2_X1 port map( A1 => n7749, A2 => n10239, ZN => n10261);
   U8237 : INV_X2 port map( A => n9253, ZN => n9248);
   U8238 : BUF_X2 port map( A => n9074, Z => n8453);
   U8239 : AND2_X2 port map( A1 => DataPath_i_PIPLIN_A_22_port, A2 => n8557, ZN
                           => n7606);
   U8240 : NAND2_X2 port map( A1 => DataPath_i_PIPLIN_A_21_port, A2 => n7617, 
                           ZN => n9961);
   U8241 : BUF_X2 port map( A => n161, Z => n8396);
   U8242 : INV_X2 port map( A => n7755, ZN => n7774);
   U8243 : INV_X2 port map( A => n8433, ZN => n7799);
   U8244 : INV_X2 port map( A => n9602, ZN => n9600);
   U8245 : INV_X4 port map( A => n9985, ZN => n9986);
   U8246 : INV_X4 port map( A => n9903, ZN => n9188);
   U8247 : CLKBUF_X3 port map( A => i_ALU_OP_2_port, Z => n8566);
   U8248 : BUF_X2 port map( A => n10017, Z => n8403);
   U8249 : CLKBUF_X3 port map( A => n10017, Z => n8404);
   U8250 : INV_X2 port map( A => n10016, ZN => n10017);
   U8251 : INV_X2 port map( A => n9785, ZN => n7727);
   U8252 : OAI21_X2 port map( B1 => n8320, B2 => n8069, A => n9066, ZN => n9241
                           );
   U8253 : NAND2_X2 port map( A1 => n10188, A2 => n10421, ZN => n8420);
   U8254 : CLKBUF_X3 port map( A => n8420, Z => n8421);
   U8255 : INV_X1 port map( A => n8448, ZN => n8449);
   U8256 : OR3_X1 port map( A1 => n7926, A2 => n8396, A3 => n8223, ZN => n10421
                           );
   U8257 : BUF_X1 port map( A => n9059, Z => n7751);
   U8258 : OR2_X1 port map( A1 => n7859, A2 => n8389, ZN => n7607);
   U8259 : OR2_X1 port map( A1 => n10199, A2 => n10400, ZN => n7608);
   U8260 : BUF_X4 port map( A => n8419, Z => n7621);
   U8261 : NOR2_X1 port map( A1 => n7850, A2 => n7848, ZN => n7609);
   U8262 : BUF_X1 port map( A => n10373, Z => n7926);
   U8263 : INV_X1 port map( A => n10429, ZN => n11885);
   U8264 : NAND2_X2 port map( A1 => DataPath_i_PIPLIN_A_24_port, A2 => n7618, 
                           ZN => n9528);
   U8265 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_31_port, ZN => n7612);
   U8266 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_28_port, ZN => n7613);
   U8267 : NOR2_X1 port map( A1 => n11884, A2 => n514, ZN => n7614);
   U8268 : BUF_X1 port map( A => DataPath_RF_c_win_4_port, Z => n8564);
   U8269 : BUF_X2 port map( A => n9069, Z => n7615);
   U8270 : INV_X4 port map( A => n9137, ZN => n9133);
   U8271 : NAND2_X2 port map( A1 => n9004, A2 => n9003, ZN => n9137);
   U8272 : BUF_X2 port map( A => n8556, Z => n7618);
   U8273 : INV_X1 port map( A => n8558, ZN => n8556);
   U8274 : NOR2_X1 port map( A1 => n7654, A2 => n7655, ZN => 
                           DP_OP_751_130_6421_n1667);
   U8275 : INV_X1 port map( A => DP_OP_751_130_6421_n1748, ZN => n7654);
   U8276 : INV_X1 port map( A => DP_OP_751_130_6421_n1746, ZN => n7652);
   U8277 : OAI211_X1 port map( C1 => n9165, C2 => DP_OP_751_130_6421_I2, A => 
                           n7844, B => n7845, ZN => n7619);
   U8278 : BUF_X1 port map( A => n8441, Z => n7620);
   U8279 : INV_X1 port map( A => n10348, ZN => n8920);
   U8280 : NAND2_X1 port map( A1 => n10348, A2 => n206, ZN => n8921);
   U8281 : BUF_X2 port map( A => n8140, Z => n7622);
   DRAMRF_ADDRESS_1_port <= '0';
   DRAMRF_ADDRESS_0_port <= '0';
   U8284 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_26_port, A2 => n8576, ZN => 
                           n7623);
   U8285 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_27_port, A2 => n8575, ZN => 
                           n7624);
   U8286 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_25_port, A2 => n8577, ZN => 
                           n7625);
   U8287 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_28_port, A2 => n8571, ZN => 
                           n7626);
   U8288 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_24_port, A2 => n8574, ZN => 
                           n7627);
   U8289 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_23_port, A2 => n8573, ZN => 
                           n7628);
   U8290 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_22_port, A2 => n8578, ZN => 
                           n7629);
   U8291 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_21_port, A2 => n8575, ZN => 
                           n7630);
   U8292 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_20_port, A2 => n8572, ZN => 
                           n7631);
   U8293 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_19_port, A2 => n8571, ZN => 
                           n7632);
   U8294 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_18_port, A2 => n8574, ZN => 
                           n7633);
   U8295 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_17_port, A2 => n8573, ZN => 
                           n7634);
   U8296 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_16_port, A2 => n8578, ZN => 
                           n7635);
   U8297 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_15_port, A2 => n8580, ZN => 
                           n7636);
   U8298 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_14_port, A2 => n8574, ZN => 
                           n7637);
   U8299 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_13_port, A2 => n8570, ZN => 
                           n7638);
   U8300 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_12_port, A2 => n8581, ZN => 
                           n7639);
   U8301 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_11_port, A2 => n8582, ZN => 
                           n7640);
   U8302 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_9_port, A2 => n8576, ZN => 
                           n7641);
   U8303 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_10_port, A2 => n8572, ZN => 
                           n7642);
   U8304 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_8_port, A2 => n8576, ZN => 
                           n7643);
   U8305 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_7_port, A2 => n8580, ZN => 
                           n7644);
   U8306 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_6_port, A2 => n8570, ZN => 
                           n7645);
   U8307 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_5_port, A2 => n8578, ZN => 
                           n7646);
   U8308 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_4_port, A2 => n8582, ZN => 
                           n7647);
   U8309 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_3_port, A2 => n8573, ZN => 
                           n7648);
   U8310 : AND2_X1 port map( A1 => DRAMRF_ADDRESS_2_port, A2 => n8576, ZN => 
                           n7649);
   U8311 : NAND2_X1 port map( A1 => n7947, A2 => n7650, ZN => 
                           DP_OP_751_130_6421_n1453);
   U8312 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1507, B2 => 
                           DP_OP_751_130_6421_n1553, A => n7948, ZN => n7650);
   U8313 : XNOR2_X1 port map( A => n7651, B => n7958, ZN => n7948);
   U8314 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1607, B => 
                           DP_OP_751_130_6421_n1651, ZN => n7651);
   U8315 : XNOR2_X1 port map( A => n7653, B => DP_OP_751_130_6421_n1746, ZN => 
                           DP_OP_751_130_6421_n1664);
   U8316 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_18_port, B => 
                           n8146, ZN => n7653);
   U8317 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1748, B => n7655, ZN => 
                           DP_OP_751_130_6421_n1668);
   U8318 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_16_port, B => 
                           n8146, ZN => n7655);
   U8319 : OAI21_X1 port map( B1 => n7656, B2 => n7874, A => n7873, ZN => n6992
                           );
   U8320 : XNOR2_X1 port map( A => n7659, B => n7657, ZN => n7656);
   U8321 : XNOR2_X1 port map( A => n7658, B => n7937, ZN => n7657);
   U8322 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n267, B => 
                           DP_OP_751_130_6421_n365, ZN => n7658);
   U8323 : AOI21_X1 port map( B1 => DP_OP_751_130_6421_n64, B2 => n8078, A => 
                           n8077, ZN => n7659);
   U8324 : AND2_X1 port map( A1 => n7668, A2 => n7669, ZN => 
                           DP_OP_751_130_6421_n64);
   U8325 : NAND2_X1 port map( A1 => n7661, A2 => n7660, ZN => n6993);
   U8326 : AOI21_X1 port map( B1 => n9412, B2 => n10429, A => n7614, ZN => 
                           n7660);
   U8327 : NAND2_X1 port map( A1 => n7664, A2 => n7662, ZN => n7661);
   U8328 : NOR2_X1 port map( A1 => n11885, A2 => n7663, ZN => n7662);
   U8329 : INV_X1 port map( A => n10094, ZN => n7663);
   U8330 : XNOR2_X1 port map( A => n7665, B => DP_OP_751_130_6421_n64, ZN => 
                           n7664);
   U8331 : NAND2_X1 port map( A1 => n8078, A2 => DP_OP_751_130_6421_n63, ZN => 
                           n7665);
   U8332 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n466, B => n7666, ZN => 
                           DP_OP_751_130_6421_n368);
   U8333 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n467, B => 
                           DP_OP_751_130_6421_n403, ZN => n7666);
   U8334 : INV_X1 port map( A => n7667, ZN => n8369);
   U8335 : OAI21_X1 port map( B1 => n8371, B2 => n8370, A => n8373, ZN => n7667
                           );
   U8336 : OAI21_X1 port map( B1 => n8385, B2 => n8387, A => n8271, ZN => n8370
                           );
   U8337 : NAND3_X1 port map( A1 => n7832, A2 => n7973, A3 => n8050, ZN => 
                           n7668);
   U8338 : NAND2_X1 port map( A1 => n7973, A2 => n7670, ZN => n7669);
   U8339 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n368, A2 => 
                           DP_OP_751_130_6421_n369, ZN => n7670);
   U8340 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n66, A2 => n8042, ZN => 
                           n7832);
   U8341 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1359, B => 
                           DP_OP_751_130_6421_n1308, Z => n7671);
   U8342 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1358, B => n7671, Z => 
                           DP_OP_751_130_6421_n1260);
   U8343 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1457, A2 => 
                           DP_OP_751_130_6421_n1408, ZN => n7672);
   U8344 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1457, A2 => 
                           DP_OP_751_130_6421_n1456, ZN => n7673);
   U8345 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1408, A2 => 
                           DP_OP_751_130_6421_n1456, ZN => n7674);
   U8346 : NAND3_X1 port map( A1 => n7672, A2 => n7673, A3 => n7674, ZN => 
                           DP_OP_751_130_6421_n1357);
   U8347 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1359, A2 => 
                           DP_OP_751_130_6421_n1308, ZN => n7675);
   U8348 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1359, A2 => 
                           DP_OP_751_130_6421_n1358, ZN => n7676);
   U8349 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1308, A2 => 
                           DP_OP_751_130_6421_n1358, ZN => n7677);
   U8350 : NAND3_X1 port map( A1 => n7675, A2 => n7676, A3 => n7677, ZN => 
                           DP_OP_751_130_6421_n1259);
   U8351 : INV_X1 port map( A => n7606, ZN => n7714);
   U8352 : AND2_X2 port map( A1 => n8556, A2 => DataPath_i_PIPLIN_A_23_port, ZN
                           => n9602);
   U8353 : OR2_X1 port map( A1 => n8567, A2 => n8268, ZN => n7678);
   U8354 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1453, A2 => 
                           DP_OP_751_130_6421_n1406, ZN => n7909);
   U8355 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1460, B => n7679, ZN => 
                           DP_OP_751_130_6421_n1362);
   U8356 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1461, B => 
                           DP_OP_751_130_6421_n1410, ZN => n7679);
   U8357 : XNOR2_X1 port map( A => n7680, B => DP_OP_751_130_6421_n1064, ZN => 
                           DP_OP_751_130_6421_n966);
   U8358 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1065, B => 
                           DP_OP_751_130_6421_n1008, ZN => n7680);
   U8359 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n768, B => n7681, ZN => 
                           DP_OP_751_130_6421_n670);
   U8360 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n769, B => 
                           DP_OP_751_130_6421_n707, ZN => n7681);
   U8361 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1553, A2 => 
                           DP_OP_751_130_6421_n1507, ZN => n7947);
   U8362 : XOR2_X1 port map( A => DP_OP_751_130_6421_n955, B => 
                           DP_OP_751_130_6421_n902, Z => n7682);
   U8363 : XOR2_X1 port map( A => n7682, B => DP_OP_751_130_6421_n954, Z => 
                           DP_OP_751_130_6421_n856);
   U8364 : XOR2_X1 port map( A => DP_OP_751_130_6421_n857, B => 
                           DP_OP_751_130_6421_n802, Z => n7683);
   U8365 : XOR2_X1 port map( A => n7683, B => DP_OP_751_130_6421_n856, Z => 
                           DP_OP_751_130_6421_n758);
   U8366 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n955, A2 => 
                           DP_OP_751_130_6421_n902, ZN => n7684);
   U8367 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n955, A2 => 
                           DP_OP_751_130_6421_n954, ZN => n7685);
   U8368 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n902, A2 => 
                           DP_OP_751_130_6421_n954, ZN => n7686);
   U8369 : NAND3_X1 port map( A1 => n7684, A2 => n7685, A3 => n7686, ZN => 
                           DP_OP_751_130_6421_n855);
   U8370 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1281, B => 
                           DP_OP_751_130_6421_n1218, Z => n7687);
   U8371 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1280, B => n7687, Z => 
                           DP_OP_751_130_6421_n1182);
   U8372 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1280, A2 => 
                           DP_OP_751_130_6421_n1281, ZN => n7688);
   U8373 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1280, A2 => 
                           DP_OP_751_130_6421_n1218, ZN => n7689);
   U8374 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1281, A2 => 
                           DP_OP_751_130_6421_n1218, ZN => n7690);
   U8375 : NAND3_X1 port map( A1 => n7688, A2 => n7689, A3 => n7690, ZN => 
                           DP_OP_751_130_6421_n1181);
   U8376 : INV_X1 port map( A => n9961, ZN => n9962);
   U8377 : AND2_X1 port map( A1 => DP_OP_751_130_6421_n878, A2 => 
                           DP_OP_751_130_6421_n879, ZN => n7691);
   U8378 : OR2_X1 port map( A1 => n7692, A2 => n8225, ZN => n8964);
   U8379 : BUF_X4 port map( A => DP_OP_751_130_6421_n1527, Z => n7797);
   U8380 : CLKBUF_X3 port map( A => n8568, Z => n8069);
   U8381 : AND2_X1 port map( A1 => DP_OP_751_130_6421_n776, A2 => 
                           DP_OP_751_130_6421_n777, ZN => n7693);
   U8382 : XNOR2_X1 port map( A => n7694, B => DP_OP_751_130_6421_n870, ZN => 
                           DP_OP_751_130_6421_n772);
   U8383 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n871, B => 
                           DP_OP_751_130_6421_n809, ZN => n7694);
   U8384 : XOR2_X1 port map( A => DP_OP_751_130_6421_n565, B => 
                           DP_OP_751_130_6421_n503, Z => n7695);
   U8385 : XOR2_X1 port map( A => n7695, B => DP_OP_751_130_6421_n564, Z => 
                           DP_OP_751_130_6421_n466);
   U8386 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n565, A2 => 
                           DP_OP_751_130_6421_n503, ZN => n7696);
   U8387 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n565, A2 => 
                           DP_OP_751_130_6421_n564, ZN => n7697);
   U8388 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n503, A2 => 
                           DP_OP_751_130_6421_n564, ZN => n7698);
   U8389 : NAND3_X1 port map( A1 => n7696, A2 => n7697, A3 => n7698, ZN => 
                           DP_OP_751_130_6421_n465);
   U8390 : BUF_X2 port map( A => n9063, Z => n8444);
   U8391 : INV_X1 port map( A => n9727, ZN => n9504);
   U8392 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n119, B2 => 
                           DP_OP_751_130_6421_n117, A => 
                           DP_OP_751_130_6421_n118, ZN => n7699);
   U8393 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n119, B2 => 
                           DP_OP_751_130_6421_n117, A => 
                           DP_OP_751_130_6421_n118, ZN => 
                           DP_OP_751_130_6421_n116);
   U8394 : INV_X2 port map( A => n8438, ZN => n8439);
   U8395 : XOR2_X1 port map( A => DP_OP_751_130_6421_n969, B => 
                           DP_OP_751_130_6421_n909, Z => n7700);
   U8396 : XOR2_X1 port map( A => n7700, B => DP_OP_751_130_6421_n968, Z => 
                           DP_OP_751_130_6421_n870);
   U8397 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n969, A2 => 
                           DP_OP_751_130_6421_n909, ZN => n7701);
   U8398 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n969, A2 => 
                           DP_OP_751_130_6421_n968, ZN => n7702);
   U8399 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n909, A2 => 
                           DP_OP_751_130_6421_n968, ZN => n7703);
   U8400 : NAND3_X1 port map( A1 => n7701, A2 => n7702, A3 => n7703, ZN => 
                           DP_OP_751_130_6421_n869);
   U8401 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n871, A2 => 
                           DP_OP_751_130_6421_n809, ZN => n7704);
   U8402 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n871, A2 => 
                           DP_OP_751_130_6421_n870, ZN => n7705);
   U8403 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n809, A2 => 
                           DP_OP_751_130_6421_n870, ZN => n7706);
   U8404 : NAND3_X1 port map( A1 => n7704, A2 => n7705, A3 => n7706, ZN => 
                           DP_OP_751_130_6421_n771);
   U8405 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1460, A2 => 
                           DP_OP_751_130_6421_n1461, ZN => n7707);
   U8406 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1460, A2 => 
                           DP_OP_751_130_6421_n1410, ZN => n7708);
   U8407 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1461, A2 => 
                           DP_OP_751_130_6421_n1410, ZN => n7709);
   U8408 : NAND3_X1 port map( A1 => n7707, A2 => n7708, A3 => n7709, ZN => 
                           DP_OP_751_130_6421_n1361);
   U8409 : NAND2_X1 port map( A1 => n8103, A2 => n7712, ZN => n7710);
   U8410 : AND2_X1 port map( A1 => n7710, A2 => n7711, ZN => n8002);
   U8411 : OR2_X1 port map( A1 => IRAM_ADDRESS_30_port, A2 => n8070, ZN => 
                           n7711);
   U8412 : AND2_X1 port map( A1 => n8098, A2 => n8003, ZN => n7712);
   U8413 : AND2_X1 port map( A1 => n8103, A2 => n7713, ZN => n10273);
   U8414 : AND2_X1 port map( A1 => n8098, A2 => n10271, ZN => n7713);
   U8415 : BUF_X2 port map( A => n10054, Z => n8405);
   U8416 : MUX2_X2 port map( A => n10096, B => n9370, S => n8560, Z => n9063);
   U8417 : XNOR2_X1 port map( A => n7715, B => DP_OP_751_130_6421_n1166, ZN => 
                           DP_OP_751_130_6421_n1068);
   U8418 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1167, B => 
                           DP_OP_751_130_6421_n1110, ZN => n7715);
   U8419 : OR2_X2 port map( A1 => n8889, A2 => n10150, ZN => n8419);
   U8420 : INV_X2 port map( A => n8434, ZN => n7776);
   U8421 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1265, B => 
                           DP_OP_751_130_6421_n1210, Z => n7716);
   U8422 : XOR2_X1 port map( A => n7716, B => DP_OP_751_130_6421_n1264, Z => 
                           DP_OP_751_130_6421_n1166);
   U8423 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1265, A2 => 
                           DP_OP_751_130_6421_n1210, ZN => n7717);
   U8424 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1265, A2 => 
                           DP_OP_751_130_6421_n1264, ZN => n7718);
   U8425 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1210, A2 => 
                           DP_OP_751_130_6421_n1264, ZN => n7719);
   U8426 : NAND3_X1 port map( A1 => n7717, A2 => n7718, A3 => n7719, ZN => 
                           DP_OP_751_130_6421_n1165);
   U8427 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1167, A2 => 
                           DP_OP_751_130_6421_n1110, ZN => n7720);
   U8428 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1167, A2 => 
                           DP_OP_751_130_6421_n1166, ZN => n7721);
   U8429 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1110, A2 => 
                           DP_OP_751_130_6421_n1166, ZN => n7722);
   U8430 : NAND3_X1 port map( A1 => n7720, A2 => n7721, A3 => n7722, ZN => 
                           DP_OP_751_130_6421_n1067);
   U8431 : INV_X1 port map( A => n7840, ZN => n7723);
   U8432 : AND2_X1 port map( A1 => DP_OP_751_130_6421_n1713, A2 => 
                           DP_OP_751_130_6421_n1743, ZN => 
                           DP_OP_751_130_6421_n1657);
   U8433 : NAND2_X1 port map( A1 => n10263, A2 => n10262, ZN => n10293);
   U8434 : BUF_X1 port map( A => n11998, Z => n7724);
   U8435 : AOI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n10, B2 => n8027, A 
                           => n8026, ZN => n7725);
   U8436 : AOI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n10, B2 => n8027, A 
                           => n8026, ZN => n8009);
   U8437 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1742, B => 
                           DP_OP_751_130_6421_n1712, Z => n7954);
   U8438 : BUF_X4 port map( A => n8359, Z => n7726);
   U8439 : INV_X1 port map( A => n9785, ZN => n9784);
   U8440 : BUF_X2 port map( A => n9063, Z => n8445);
   U8441 : CLKBUF_X1 port map( A => n7596, Z => n8020);
   U8442 : NOR2_X1 port map( A1 => n8397, A2 => n10238, ZN => n10422);
   U8443 : NOR2_X1 port map( A1 => n10191, A2 => n10149, ZN => n10402);
   U8444 : XNOR2_X1 port map( A => n7595, B => DP_OP_751_130_6421_n471, ZN => 
                           n8041);
   U8445 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n768, A2 => 
                           DP_OP_751_130_6421_n769, ZN => n7729);
   U8446 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n768, A2 => 
                           DP_OP_751_130_6421_n707, ZN => n7730);
   U8447 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n769, A2 => 
                           DP_OP_751_130_6421_n707, ZN => n7731);
   U8448 : NAND3_X1 port map( A1 => n7729, A2 => n7730, A3 => n7731, ZN => 
                           DP_OP_751_130_6421_n669);
   U8449 : OR2_X1 port map( A1 => n9883, A2 => n7755, ZN => n10096);
   U8450 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1569, A2 => 
                           DP_OP_751_130_6421_n1515, ZN => n8059);
   U8451 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1569, B2 => 
                           DP_OP_751_130_6421_n1515, A => n8061, ZN => n8060);
   U8452 : NAND2_X1 port map( A1 => n8358, A2 => n11800, ZN => n11998);
   U8453 : NOR2_X1 port map( A1 => CU_I_CW_MUXA_SEL_port, A2 => n10402, ZN => 
                           n8603);
   U8454 : BUF_X1 port map( A => n8221, Z => n7732);
   U8455 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1261, B => 
                           DP_OP_751_130_6421_n1208, Z => n7733);
   U8456 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1260, B => n7733, Z => 
                           DP_OP_751_130_6421_n1162);
   U8457 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1260, A2 => 
                           DP_OP_751_130_6421_n1261, ZN => n7734);
   U8458 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1260, A2 => 
                           DP_OP_751_130_6421_n1208, ZN => n7735);
   U8459 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1261, A2 => 
                           DP_OP_751_130_6421_n1208, ZN => n7736);
   U8460 : NAND3_X1 port map( A1 => n7734, A2 => n7735, A3 => n7736, ZN => 
                           DP_OP_751_130_6421_n1161);
   U8461 : AND2_X2 port map( A1 => DP_OP_751_130_6421_n1710, A2 => n7188, ZN =>
                           DP_OP_751_130_6421_n1651);
   U8462 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1657, A2 => 
                           DP_OP_751_130_6421_n1610, ZN => n7952);
   U8463 : XNOR2_X1 port map( A => n7841, B => n8148, ZN => n7746);
   U8464 : XOR2_X1 port map( A => DP_OP_751_130_6421_n1163, B => 
                           DP_OP_751_130_6421_n1108, Z => n7737);
   U8465 : XOR2_X1 port map( A => n7737, B => DP_OP_751_130_6421_n1162, Z => 
                           DP_OP_751_130_6421_n1064);
   U8466 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1163, A2 => 
                           DP_OP_751_130_6421_n1108, ZN => n7738);
   U8467 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1163, A2 => 
                           DP_OP_751_130_6421_n1162, ZN => n7739);
   U8468 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1108, A2 => 
                           DP_OP_751_130_6421_n1162, ZN => n7740);
   U8469 : NAND3_X1 port map( A1 => n7738, A2 => n7739, A3 => n7740, ZN => 
                           DP_OP_751_130_6421_n1063);
   U8470 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1065, A2 => 
                           DP_OP_751_130_6421_n1008, ZN => n7741);
   U8471 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1065, A2 => 
                           DP_OP_751_130_6421_n1064, ZN => n7742);
   U8472 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1008, A2 => 
                           DP_OP_751_130_6421_n1064, ZN => n7743);
   U8473 : NAND3_X1 port map( A1 => n7741, A2 => n7742, A3 => n7743, ZN => 
                           DP_OP_751_130_6421_n965);
   U8474 : AND3_X2 port map( A1 => n8181, A2 => n8180, A3 => n8179, ZN => n7744
                           );
   U8475 : BUF_X1 port map( A => DP_OP_751_130_6421_n66, Z => n7745);
   U8476 : NAND2_X1 port map( A1 => n7832, A2 => n8050, ZN => n7747);
   U8477 : AND2_X1 port map( A1 => n8193, A2 => DataPath_i_PIPLIN_IN2_5_port, 
                           ZN => n7839);
   U8478 : BUF_X1 port map( A => DP_OP_751_130_6421_n88, Z => n7918);
   U8479 : BUF_X1 port map( A => DP_OP_751_130_6421_n83, Z => n7922);
   U8480 : NAND2_X1 port map( A1 => n8939, A2 => n8940, ZN => 
                           DP_OP_751_130_6421_n1731);
   U8481 : CLKBUF_X3 port map( A => n9064, Z => n8446);
   U8482 : OAI21_X2 port map( B1 => n9743, B2 => DP_OP_751_130_6421_n915, A => 
                           n9093, ZN => n9094);
   U8483 : XNOR2_X2 port map( A => DP_OP_751_130_6421_n1017, B => n9743, ZN => 
                           n9095);
   U8484 : BUF_X1 port map( A => DP_OP_751_130_6421_n67, Z => n7999);
   U8485 : XNOR2_X1 port map( A => n7745, B => n8049, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_60_port);
   U8486 : BUF_X1 port map( A => n10240, Z => n7748);
   U8487 : BUF_X2 port map( A => n10240, Z => n7749);
   U8488 : NAND2_X1 port map( A1 => n8912, A2 => n8911, ZN => n10240);
   U8489 : XNOR2_X1 port map( A => n7747, B => n8052, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_61_port);
   U8490 : INV_X1 port map( A => n9041, ZN => n9059);
   U8491 : AND2_X2 port map( A1 => n8557, A2 => DataPath_i_PIPLIN_A_25_port, ZN
                           => n9936);
   U8492 : INV_X2 port map( A => n8559, ZN => n8557);
   U8493 : OAI21_X1 port map( B1 => n7754, B2 => n8004, A => n8988, ZN => n7753
                           );
   U8494 : INV_X2 port map( A => n9843, ZN => n9844);
   U8495 : BUF_X4 port map( A => n9844, Z => n8401);
   U8496 : BUF_X1 port map( A => n9843, Z => n7828);
   U8497 : NAND2_X1 port map( A1 => n7678, A2 => n8938, ZN => n7754);
   U8498 : BUF_X4 port map( A => DP_OP_751_130_6421_I2, Z => n8148);
   U8499 : NAND2_X1 port map( A1 => n8939, A2 => n8940, ZN => n7755);
   U8500 : BUF_X4 port map( A => DP_OP_751_130_6421_n1731, Z => n8146);
   U8501 : BUF_X1 port map( A => DP_OP_751_130_6421_n91, Z => n7876);
   U8502 : INV_X2 port map( A => n9041, ZN => n7756);
   U8503 : INV_X2 port map( A => n8194, ZN => n7757);
   U8504 : BUF_X2 port map( A => n8425, Z => n8426);
   U8505 : AOI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n6, B2 => n8106, A =>
                           n7807, ZN => n8115);
   U8506 : INV_X4 port map( A => n11846, ZN => n7758);
   U8507 : AND2_X1 port map( A1 => n8808, A2 => n8834, ZN => n8691);
   U8508 : NOR2_X2 port map( A1 => n10498, A2 => n10485, ZN => n8465);
   U8509 : NOR2_X2 port map( A1 => n10499, A2 => n10502, ZN => n8471);
   U8510 : NOR2_X2 port map( A1 => n10500, A2 => n10486, ZN => n8467);
   U8511 : NOR2_X2 port map( A1 => n10501, A2 => n10485, ZN => n8462);
   U8512 : NOR2_X2 port map( A1 => n10502, A2 => n10486, ZN => n8468);
   U8513 : NOR2_X2 port map( A1 => n10503, A2 => n10502, ZN => n8477);
   U8514 : NOR2_X2 port map( A1 => n10503, A2 => n10502, ZN => n8478);
   U8515 : NOR2_X2 port map( A1 => n10500, A2 => n10499, ZN => n8474);
   U8516 : NOR2_X2 port map( A1 => n10500, A2 => n10486, ZN => n8466);
   U8517 : NOR2_X2 port map( A1 => n10500, A2 => n10499, ZN => n8475);
   U8518 : NOR2_X2 port map( A1 => n10501, A2 => n10485, ZN => n8461);
   U8519 : NOR2_X2 port map( A1 => n10502, A2 => n10486, ZN => n8469);
   U8520 : NOR2_X2 port map( A1 => n10499, A2 => n10501, ZN => n8473);
   U8521 : NOR2_X2 port map( A1 => n10498, A2 => n10486, ZN => n8460);
   U8522 : OAI22_X1 port map( A1 => n10127, A2 => n11881, B1 => n11884, B2 => 
                           n515, ZN => n7978);
   U8523 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1255, A2 => 
                           DP_OP_751_130_6421_n1205, ZN => n7884);
   U8524 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1353, A2 => 
                           DP_OP_751_130_6421_n1305, ZN => n7882);
   U8525 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1353, B2 => 
                           DP_OP_751_130_6421_n1305, A => 
                           DP_OP_751_130_6421_n1352, ZN => n7883);
   U8526 : INV_X2 port map( A => n11554, ZN => n11553);
   U8527 : INV_X2 port map( A => n11148, ZN => n11147);
   U8528 : INV_X2 port map( A => n8410, ZN => n7759);
   U8529 : INV_X2 port map( A => n11101, ZN => n11100);
   U8530 : INV_X2 port map( A => n11145, ZN => n11144);
   U8531 : INV_X2 port map( A => n11368, ZN => n11367);
   U8532 : INV_X2 port map( A => n8408, ZN => n7760);
   U8533 : INV_X2 port map( A => n8409, ZN => n7761);
   U8534 : INV_X2 port map( A => n11142, ZN => n11141);
   U8535 : INV_X2 port map( A => n11566, ZN => n11565);
   U8536 : INV_X2 port map( A => n8411, ZN => n7762);
   U8537 : INV_X2 port map( A => n11560, ZN => n11559);
   U8538 : INV_X2 port map( A => n11152, ZN => n11151);
   U8539 : AND2_X2 port map( A1 => n8581, A2 => n11069, ZN => n11073);
   U8540 : INV_X1 port map( A => n8286, ZN => n7781);
   U8541 : INV_X2 port map( A => n11362, ZN => n11361);
   U8542 : INV_X2 port map( A => n11448, ZN => n11446);
   U8543 : INV_X2 port map( A => n11365, ZN => n11364);
   U8544 : INV_X2 port map( A => n8407, ZN => n7763);
   U8545 : AND2_X2 port map( A1 => n8577, A2 => n11334, ZN => n11335);
   U8546 : INV_X2 port map( A => n8528, ZN => n7764);
   U8547 : BUF_X2 port map( A => n11750, Z => n7765);
   U8548 : AND2_X2 port map( A1 => n8580, A2 => n11212, ZN => n11213);
   U8549 : INV_X2 port map( A => n11153, ZN => n11150);
   U8550 : INV_X2 port map( A => n11041, ZN => n11923);
   U8551 : INV_X2 port map( A => n8296, ZN => n7766);
   U8552 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1561, A2 => 
                           DP_OP_751_130_6421_n1511, ZN => n7833);
   U8553 : NOR2_X1 port map( A1 => n7863, A2 => n7807, ZN => n7862);
   U8554 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1615, A2 => 
                           DP_OP_751_130_6421_n1667, ZN => n8057);
   U8555 : BUF_X2 port map( A => n9088, Z => n7767);
   U8556 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1649, B2 => 
                           DP_OP_751_130_6421_n1606, A => n7934, ZN => n7933);
   U8557 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1649, A2 => 
                           DP_OP_751_130_6421_n1606, ZN => n7932);
   U8558 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1659, A2 => 
                           DP_OP_751_130_6421_n1611, ZN => n7890);
   U8559 : AND2_X1 port map( A1 => DP_OP_751_130_6421_n1709, A2 => 
                           DP_OP_751_130_6421_n1739, ZN => 
                           DP_OP_751_130_6421_n1649);
   U8560 : BUF_X1 port map( A => n9085, Z => n7785);
   U8561 : BUF_X1 port map( A => n9078, Z => n7787);
   U8562 : INV_X2 port map( A => n8569, ZN => n7768);
   U8563 : BUF_X1 port map( A => n9089, Z => n7790);
   U8564 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_2_17_port, B => 
                           n7772, ZN => DP_OP_751_130_6421_n1615);
   U8565 : INV_X2 port map( A => n10432, ZN => n11884);
   U8566 : INV_X1 port map( A => n9755, ZN => n7789);
   U8567 : BUF_X2 port map( A => n9078, Z => n7769);
   U8568 : BUF_X2 port map( A => n9080, Z => n7770);
   U8569 : BUF_X1 port map( A => DP_OP_751_130_6421_n1425, Z => n7792);
   U8570 : BUF_X2 port map( A => n9075, Z => n7771);
   U8571 : AOI21_X1 port map( B1 => n8187, B2 => n7802, A => n8129, ZN => n8128
                           );
   U8572 : INV_X1 port map( A => n8145, ZN => n7772);
   U8573 : NAND2_X1 port map( A1 => n8107, A2 => n7807, ZN => n8104);
   U8574 : NOR2_X1 port map( A1 => n8114, A2 => n7808, ZN => n8121);
   U8575 : INV_X2 port map( A => n7803, ZN => DP_OP_751_130_6421_n1323);
   U8576 : NOR3_X1 port map( A1 => n8176, A2 => n8170, A3 => n7484, ZN => n8133
                           );
   U8577 : BUF_X1 port map( A => n9370, Z => n7985);
   U8578 : BUF_X1 port map( A => n10096, Z => n7982);
   U8579 : INV_X1 port map( A => n7606, ZN => n7773);
   U8580 : BUF_X2 port map( A => DP_OP_751_130_6421_n1629, Z => n7775);
   U8581 : AOI21_X1 port map( B1 => n8111, B2 => n8177, A => n7808, ZN => n8107
                           );
   U8582 : AND2_X2 port map( A1 => n8978, A2 => n8977, ZN => n9122);
   U8583 : INV_X1 port map( A => n9495, ZN => n7777);
   U8584 : INV_X1 port map( A => n10443, ZN => n7778);
   U8585 : BUF_X4 port map( A => DP_OP_1091J1_126_6973_n72, Z => 
                           DP_OP_1091J1_126_6973_n31);
   U8586 : NOR2_X4 port map( A1 => n8292, A2 => i_ALU_OP_1_port, ZN => n10094);
   U8587 : CLKBUF_X1 port map( A => DP_OP_1091J1_126_6973_n72, Z => n7779);
   U8588 : AOI22_X1 port map( A1 => n8921, A2 => n10346, B1 => n8920, B2 => 
                           IRAM_ADDRESS_8_port, ZN => n8928);
   U8589 : AND2_X1 port map( A1 => n7860, A2 => n7859, ZN => n8390);
   U8590 : INV_X1 port map( A => n8098, ZN => n8097);
   U8591 : AOI21_X1 port map( B1 => n8098, B2 => n8096, A => n10267, ZN => 
                           n8095);
   U8592 : NOR2_X1 port map( A1 => n8099, A2 => n10284, ZN => n8098);
   U8593 : INV_X1 port map( A => n8101, ZN => n8099);
   U8594 : INV_X1 port map( A => n7851, ZN => n7850);
   U8595 : NOR2_X1 port map( A1 => n7857, A2 => n8389, ZN => n7856);
   U8596 : INV_X1 port map( A => n10265, ZN => n8096);
   U8597 : NAND2_X1 port map( A1 => n10287, A2 => n10266, ZN => n10267);
   U8598 : AND2_X1 port map( A1 => n8267, A2 => n10345, ZN => n7851);
   U8599 : INV_X1 port map( A => n10264, ZN => n8100);
   U8600 : INV_X1 port map( A => n10251, ZN => n7857);
   U8601 : INV_X1 port map( A => n7852, ZN => n7848);
   U8602 : NOR2_X1 port map( A1 => n8927, A2 => n8926, ZN => n7849);
   U8603 : INV_X1 port map( A => n11845, ZN => n10418);
   U8604 : INV_X1 port map( A => n10367, ZN => n10417);
   U8605 : AND2_X1 port map( A1 => n10367, A2 => n11834, ZN => n8194);
   U8606 : NAND2_X1 port map( A1 => n10367, A2 => i_NPC_SEL, ZN => n11845);
   U8607 : NAND2_X1 port map( A1 => n7880, A2 => n8913, ZN => n10367);
   U8608 : INV_X1 port map( A => n10355, ZN => n7780);
   U8609 : XNOR2_X1 port map( A => n7999, B => n8041, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_59_port);
   U8610 : XNOR2_X1 port map( A => n7895, B => n8019, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_58_port);
   U8611 : XNOR2_X1 port map( A => n8039, B => n7990, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_57_port);
   U8612 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n10, B => n8025, ZN =>
                           C620_DATA2_23);
   U8613 : AND2_X1 port map( A1 => n10200, A2 => n8887, ZN => n7972);
   U8614 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n12, B => n7986, ZN =>
                           C620_DATA2_21);
   U8615 : OAI21_X1 port map( B1 => n7979, B2 => n7989, A => n7988, ZN => 
                           DP_OP_1091J1_126_6973_n11);
   U8616 : INV_X1 port map( A => n7979, ZN => DP_OP_1091J1_126_6973_n12);
   U8617 : OR2_X1 port map( A1 => n8795, A2 => n8022, ZN => n8874);
   U8618 : INV_X1 port map( A => DP_OP_751_130_6421_n63, ZN => n8077);
   U8619 : NAND2_X1 port map( A1 => n7995, A2 => n7994, ZN => 
                           DP_OP_751_130_6421_n267);
   U8620 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n367, A2 => n7996, ZN =>
                           n7995);
   U8621 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n368, B => 
                           DP_OP_751_130_6421_n369, ZN => n8052);
   U8622 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n369, A2 => 
                           DP_OP_751_130_6421_n368, ZN => n7973);
   U8623 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n18, B => n8076, ZN =>
                           C620_DATA2_15);
   U8624 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n19, B => n8071, ZN =>
                           C620_DATA2_14);
   U8625 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n370, A2 => 
                           DP_OP_751_130_6421_n468, ZN => n8042);
   U8626 : NAND2_X1 port map( A1 => n8088, A2 => n8727, ZN => n8086);
   U8627 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n370, B => 
                           DP_OP_751_130_6421_n468, ZN => n8049);
   U8628 : NAND2_X1 port map( A1 => n8091, A2 => n8727, ZN => n8087);
   U8629 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n572, B => 
                           DP_OP_751_130_6421_n573, ZN => n8039);
   U8630 : NAND2_X1 port map( A1 => n8024, A2 => n8023, ZN => n8022);
   U8631 : INV_X1 port map( A => n8065, ZN => DP_OP_1091J1_126_6973_n19);
   U8632 : OAI21_X1 port map( B1 => n8092, B2 => n8090, A => n8089, ZN => n8088
                           );
   U8633 : AND2_X1 port map( A1 => n8094, A2 => n8801, ZN => n8091);
   U8634 : AOI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n20, B2 => n8066, A 
                           => n7970, ZN => n8065);
   U8635 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n469, B => n7969, ZN => 
                           DP_OP_751_130_6421_n370);
   U8636 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n472, B => 
                           DP_OP_751_130_6421_n570, ZN => n8019);
   U8637 : INV_X1 port map( A => n8792, ZN => n8023);
   U8638 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n472, A2 => 
                           DP_OP_751_130_6421_n570, ZN => n8016);
   U8639 : NOR2_X1 port map( A1 => n8794, A2 => n8793, ZN => n8024);
   U8640 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n472, A2 => 
                           DP_OP_751_130_6421_n570, ZN => n8018);
   U8641 : INV_X1 port map( A => n8801, ZN => n8090);
   U8642 : INV_X1 port map( A => n8698, ZN => n8089);
   U8643 : OAI21_X1 port map( B1 => n8030, B2 => n8029, A => n8028, ZN => 
                           DP_OP_751_130_6421_n573);
   U8644 : AND2_X1 port map( A1 => n8846, A2 => n8800, ZN => n8727);
   U8645 : OAI21_X1 port map( B1 => n8055, B2 => n8054, A => n8053, ZN => 
                           DP_OP_751_130_6421_n675);
   U8646 : INV_X1 port map( A => DP_OP_751_130_6421_n673, ZN => n8030);
   U8647 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n775, B => n8056, ZN => 
                           DP_OP_751_130_6421_n676);
   U8648 : INV_X1 port map( A => DP_OP_751_130_6421_n775, ZN => n8055);
   U8649 : XNOR2_X1 port map( A => n7894, B => DP_OP_751_130_6421_n1154, ZN => 
                           DP_OP_751_130_6421_n1056);
   U8650 : INV_X1 port map( A => n11753, ZN => n8911);
   U8651 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n877, B => n7899, ZN => 
                           DP_OP_751_130_6421_n778);
   U8652 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1155, B => 
                           DP_OP_751_130_6421_n1104, ZN => n7894);
   U8653 : OR2_X1 port map( A1 => i_HAZARD_SIG_CU, A2 => n8585, ZN => n11753);
   U8654 : NAND2_X1 port map( A1 => n7885, A2 => n7884, ZN => 
                           DP_OP_751_130_6421_n1155);
   U8655 : INV_X1 port map( A => i_RD1_2_port, ZN => n7896);
   U8656 : NAND2_X1 port map( A1 => n7831, A2 => n7830, ZN => 
                           DP_OP_751_130_6421_n1251);
   U8657 : NAND2_X1 port map( A1 => n7878, A2 => n7877, ZN => 
                           DP_OP_751_130_6421_n1247);
   U8658 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1255, B2 => 
                           DP_OP_751_130_6421_n1205, A => n7886, ZN => n7885);
   U8659 : BUF_X1 port map( A => n11055, Z => n8485);
   U8660 : NAND2_X1 port map( A1 => n7883, A2 => n7882, ZN => 
                           DP_OP_751_130_6421_n1253);
   U8661 : BUF_X1 port map( A => n11498, Z => n8516);
   U8662 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1351, A2 => 
                           DP_OP_751_130_6421_n1304, ZN => n7830);
   U8663 : BUF_X1 port map( A => n11501, Z => n8518);
   U8664 : BUF_X1 port map( A => n11752, Z => n8540);
   U8665 : BUF_X1 port map( A => n11522, Z => n8525);
   U8666 : BUF_X1 port map( A => n11516, Z => n8523);
   U8667 : BUF_X1 port map( A => n11097, Z => n8494);
   U8668 : BUF_X1 port map( A => n11975, Z => n8551);
   U8669 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1346, B => n7879, ZN => 
                           DP_OP_751_130_6421_n1248);
   U8670 : BUF_X1 port map( A => n11058, Z => n8487);
   U8671 : BUF_X1 port map( A => n11023, Z => n8481);
   U8672 : AND2_X2 port map( A1 => n8576, A2 => n11888, ZN => n11889);
   U8673 : INV_X2 port map( A => n11038, ZN => n11037);
   U8674 : BUF_X1 port map( A => n11571, Z => n8527);
   U8675 : INV_X2 port map( A => n11577, ZN => n11576);
   U8676 : BUF_X1 port map( A => n11542, Z => n8526);
   U8677 : NAND2_X1 port map( A1 => n7910, A2 => n7909, ZN => 
                           DP_OP_751_130_6421_n1353);
   U8678 : NAND2_X1 port map( A1 => n7964, A2 => n7963, ZN => 
                           DP_OP_751_130_6421_n1351);
   U8679 : AND2_X2 port map( A1 => n8581, A2 => n11188, ZN => n11190);
   U8680 : BUF_X1 port map( A => n11957, Z => n8549);
   U8681 : BUF_X1 port map( A => n11505, Z => n8519);
   U8682 : INV_X2 port map( A => n11511, ZN => n11510);
   U8683 : AND2_X2 port map( A1 => n8580, A2 => n11318, ZN => n11322);
   U8684 : INV_X2 port map( A => n11353, ZN => n11352);
   U8685 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1347, B => 
                           DP_OP_751_130_6421_n1302, ZN => n7879);
   U8686 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1347, A2 => 
                           DP_OP_751_130_6421_n1302, ZN => n7877);
   U8687 : AND2_X2 port map( A1 => n8578, A2 => n11398, ZN => n11406);
   U8688 : BUF_X1 port map( A => n11514, Z => n8522);
   U8689 : AND2_X2 port map( A1 => n8576, A2 => n11904, ZN => n11905);
   U8690 : AND2_X2 port map( A1 => n8576, A2 => n11893, ZN => n11894);
   U8691 : AND2_X2 port map( A1 => n8576, A2 => n11944, ZN => n11956);
   U8692 : AND2_X2 port map( A1 => n8576, A2 => n11263, ZN => n11273);
   U8693 : BUF_X1 port map( A => n11499, Z => n8517);
   U8694 : AND2_X2 port map( A1 => n8577, A2 => n11337, ZN => n11338);
   U8695 : AND2_X2 port map( A1 => n8581, A2 => n11198, ZN => n11200);
   U8696 : AND2_X2 port map( A1 => n8578, A2 => n11370, ZN => n11371);
   U8697 : AND2_X2 port map( A1 => n8581, A2 => n11093, ZN => n11095);
   U8698 : INV_X2 port map( A => n11317, ZN => n11315);
   U8699 : AND2_X2 port map( A1 => n8580, A2 => n11219, ZN => n11220);
   U8700 : AND2_X2 port map( A1 => n8578, A2 => n11354, ZN => n11355);
   U8701 : AND2_X2 port map( A1 => n8581, A2 => n11136, ZN => n11134);
   U8702 : AND2_X2 port map( A1 => n8576, A2 => n10987, ZN => n11002);
   U8703 : AND2_X2 port map( A1 => n8576, A2 => n11006, ZN => n11007);
   U8704 : NAND2_X1 port map( A1 => n7905, A2 => n7904, ZN => 
                           DP_OP_751_130_6421_n1347);
   U8705 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1451, A2 => 
                           DP_OP_751_130_6421_n1405, ZN => n7963);
   U8706 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1405, B2 => 
                           DP_OP_751_130_6421_n1451, A => n7965, ZN => n7964);
   U8707 : INV_X2 port map( A => n11359, ZN => n11358);
   U8708 : INV_X2 port map( A => n11548, ZN => n11547);
   U8709 : BUF_X1 port map( A => n11251, Z => n7813);
   U8710 : AND2_X2 port map( A1 => n8577, A2 => n11340, ZN => n11341);
   U8711 : BUF_X1 port map( A => n11287, Z => n7819);
   U8712 : AND2_X2 port map( A1 => n8577, A2 => n11323, ZN => n11324);
   U8713 : AND2_X2 port map( A1 => n8581, A2 => n11081, ZN => n11079);
   U8714 : BUF_X1 port map( A => n11249, Z => n7814);
   U8715 : INV_X2 port map( A => n11043, ZN => n11042);
   U8716 : INV_X2 port map( A => n11411, ZN => n11410);
   U8717 : BUF_X1 port map( A => n11301, Z => n7811);
   U8718 : AND2_X2 port map( A1 => n8581, A2 => n11196, ZN => n11193);
   U8719 : INV_X2 port map( A => n11016, ZN => n11015);
   U8720 : BUF_X1 port map( A => n11284, Z => n7820);
   U8721 : AND2_X2 port map( A1 => n8581, A2 => n11090, ZN => n11091);
   U8722 : AND2_X2 port map( A1 => n8581, A2 => n11202, ZN => n11203);
   U8723 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n401, B => 
                           DP_OP_751_130_6421_n301, ZN => n7939);
   U8724 : BUF_X1 port map( A => n11283, Z => n7818);
   U8725 : BUF_X1 port map( A => n11257, Z => n7812);
   U8726 : NAND2_X1 port map( A1 => n7834, A2 => n7833, ZN => 
                           DP_OP_751_130_6421_n1461);
   U8727 : NAND2_X1 port map( A1 => n8060, A2 => n8059, ZN => 
                           DP_OP_751_130_6421_n1469);
   U8728 : BUF_X1 port map( A => n11258, Z => n7815);
   U8729 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1447, A2 => 
                           DP_OP_751_130_6421_n1403, ZN => n7904);
   U8730 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1447, B2 => 
                           DP_OP_751_130_6421_n1403, A => n7906, ZN => n7905);
   U8731 : OR4_X1 port map( A1 => n9482, A2 => n9481, A3 => n9480, A4 => n9479,
                           ZN => n9970);
   U8732 : NAND2_X1 port map( A1 => n7943, A2 => n7942, ZN => 
                           DP_OP_751_130_6421_n1445);
   U8733 : NAND2_X1 port map( A1 => n7953, A2 => n7952, ZN => 
                           DP_OP_751_130_6421_n1557);
   U8734 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1545, B2 => 
                           DP_OP_751_130_6421_n1503, A => n7944, ZN => n7943);
   U8735 : BUF_X1 port map( A => n11153, Z => n8483);
   U8736 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1511, B2 => 
                           DP_OP_751_130_6421_n1561, A => n7835, ZN => n7834);
   U8737 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1549, A2 => 
                           DP_OP_751_130_6421_n1505, ZN => n7991);
   U8738 : NAND2_X1 port map( A1 => n7957, A2 => n7956, ZN => 
                           DP_OP_751_130_6421_n1551);
   U8739 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1016, B => 
                           DP_OP_751_130_6421_n1017, ZN => n8006);
   U8740 : AND2_X1 port map( A1 => DP_OP_751_130_6421_n1697, A2 => 
                           DP_OP_751_130_6421_n1760, ZN => 
                           DP_OP_751_130_6421_n1691);
   U8741 : NAND2_X1 port map( A1 => n7933, A2 => n7932, ZN => 
                           DP_OP_751_130_6421_n1549);
   U8742 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n506, B => 
                           DP_OP_751_130_6421_n507, ZN => n8008);
   U8743 : NAND2_X1 port map( A1 => n7941, A2 => n7940, ZN => 
                           DP_OP_751_130_6421_n1543);
   U8744 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1545, A2 => 
                           DP_OP_751_130_6421_n1503, ZN => n7942);
   U8745 : AND2_X1 port map( A1 => DataPath_RF_c_swin_1_port, A2 => n11449, ZN 
                           => n8296);
   U8746 : NAND2_X1 port map( A1 => n7891, A2 => n7890, ZN => 
                           DP_OP_751_130_6421_n1559);
   U8747 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n710, A2 => 
                           DP_OP_751_130_6421_n711, ZN => n8054);
   U8748 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n812, B => 
                           DP_OP_751_130_6421_n813, ZN => n7899);
   U8749 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n710, B => 
                           DP_OP_751_130_6421_n711, ZN => n8056);
   U8750 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n710, A2 => 
                           DP_OP_751_130_6421_n711, ZN => n8053);
   U8751 : INV_X1 port map( A => n10437, ZN => n11084);
   U8752 : AND2_X1 port map( A1 => DP_OP_751_130_6421_n1734, A2 => n7959, ZN =>
                           DP_OP_751_130_6421_n1639);
   U8753 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1603, B2 => 
                           DP_OP_751_130_6421_n1643, A => 
                           DP_OP_751_130_6421_n1642, ZN => n7941);
   U8754 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1643, A2 => 
                           DP_OP_751_130_6421_n1603, ZN => n7940);
   U8755 : BUF_X2 port map( A => n11041, Z => n7782);
   U8756 : INV_X1 port map( A => n10197, ZN => i_ADD_WS1_2_port);
   U8757 : BUF_X2 port map( A => n11276, Z => n7783);
   U8758 : BUF_X2 port map( A => n11409, Z => n7784);
   U8759 : INV_X1 port map( A => n8412, ZN => n11449);
   U8760 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n1696, A2 => 
                           DP_OP_751_130_6421_n1762, ZN => 
                           DP_OP_751_130_6421_n166);
   U8761 : NOR2_X2 port map( A1 => n10423, A2 => n176, ZN => i_ADD_RS2_0_port);
   U8762 : OR2_X1 port map( A1 => n11885, A2 => n7663, ZN => n7874);
   U8763 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n302, A2 => n7816, ZN => 
                           n7996);
   U8764 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n302, A2 => n7816, ZN =>
                           n7994);
   U8765 : AND2_X1 port map( A1 => DP_OP_751_130_6421_n1707, A2 => 
                           DP_OP_751_130_6421_n1737, ZN => 
                           DP_OP_751_130_6421_n1645);
   U8766 : AND2_X1 port map( A1 => DP_OP_751_130_6421_n1706, A2 => 
                           DP_OP_751_130_6421_n1736, ZN => 
                           DP_OP_751_130_6421_n1643);
   U8767 : INV_X1 port map( A => n7960, ZN => n7959);
   U8768 : NOR2_X1 port map( A1 => n7865, A2 => n8082, ZN => n7863);
   U8769 : AOI21_X1 port map( B1 => n8127, B2 => n8130, A => n8125, ZN => n8124
                           );
   U8770 : OR2_X1 port map( A1 => n7866, A2 => n8082, ZN => n7864);
   U8771 : AND2_X1 port map( A1 => n7724, A2 => n8583, ZN => n10437);
   U8772 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n302, B => n7816, ZN => 
                           n7997);
   U8773 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n608, A2 => n7817, ZN =>
                           n8028);
   U8774 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n608, A2 => n7817, ZN => 
                           n8029);
   U8775 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n608, B => n7817, ZN => 
                           n8031);
   U8776 : AND2_X1 port map( A1 => DP_OP_751_130_6421_n1712, A2 => 
                           DP_OP_751_130_6421_n1742, ZN => 
                           DP_OP_751_130_6421_n1655);
   U8777 : AND2_X1 port map( A1 => DP_OP_751_130_6421_n1708, A2 => 
                           DP_OP_751_130_6421_n1738, ZN => 
                           DP_OP_751_130_6421_n1647);
   U8778 : INV_X2 port map( A => i_SEL_CMPB, ZN => n8569);
   U8779 : INV_X1 port map( A => n7867, ZN => n7866);
   U8780 : NAND2_X1 port map( A1 => n8126, A2 => n8186, ZN => n8125);
   U8781 : NOR2_X1 port map( A1 => n8121, A2 => n8120, ZN => n8116);
   U8782 : BUF_X2 port map( A => n11988, Z => n7786);
   U8783 : INV_X2 port map( A => n8563, ZN => DP_OP_751_130_6421_n1017);
   U8784 : NOR2_X1 port map( A1 => n8360, A2 => n8240, ZN => n8594);
   U8785 : BUF_X2 port map( A => n10099, Z => n7788);
   U8786 : OR2_X1 port map( A1 => n8127, A2 => n8128, ZN => n8123);
   U8787 : NAND2_X1 port map( A1 => n8128, A2 => n8130, ZN => n8126);
   U8788 : INV_X2 port map( A => n8227, ZN => DP_OP_751_130_6421_n1221);
   U8789 : BUF_X2 port map( A => n10432, Z => n7791);
   U8790 : BUF_X1 port map( A => n10402, Z => n7949);
   U8791 : NAND2_X1 port map( A1 => n8113, A2 => n8132, ZN => n8112);
   U8792 : AND4_X1 port map( A1 => n8239, A2 => n8192, A3 => n8355, A4 => n8376
                           , ZN => n11800);
   U8793 : INV_X1 port map( A => n8187, ZN => n8130);
   U8794 : BUF_X2 port map( A => DP_OP_751_130_6421_n1119, Z => n7793);
   U8795 : NAND2_X1 port map( A1 => n8133, A2 => n8114, ZN => n8113);
   U8796 : BUF_X1 port map( A => n9156, Z => n7913);
   U8797 : BUF_X1 port map( A => n9064, Z => n8447);
   U8798 : INV_X1 port map( A => DP_OP_751_130_6421_n813, ZN => n7794);
   U8799 : AND2_X2 port map( A1 => CU_I_CW_MEM_MEM_EN_port, A2 => n10439, ZN =>
                           n11987);
   U8800 : AND3_X1 port map( A1 => n8119, A2 => n8118, A3 => n8175, ZN => n8117
                           );
   U8801 : NOR2_X1 port map( A1 => n10384, A2 => n10389, ZN => n8007);
   U8802 : OR2_X1 port map( A1 => n8602, A2 => IR_29_port, ZN => n10191);
   U8803 : NOR2_X1 port map( A1 => n7871, A2 => n7870, ZN => n7869);
   U8804 : NAND2_X1 port map( A1 => n8176, A2 => 
                           DataPath_WRF_CUhw_curr_addr_29_port, ZN => n8118);
   U8805 : NAND2_X1 port map( A1 => n8176, A2 => DP_OP_1091J1_126_6973_n31, ZN 
                           => n8119);
   U8806 : BUF_X1 port map( A => n9785, Z => n7983);
   U8807 : NOR2_X1 port map( A1 => n8176, A2 => n8108, ZN => n8105);
   U8808 : INV_X2 port map( A => n9821, ZN => n9822);
   U8809 : BUF_X1 port map( A => n9903, Z => n7875);
   U8810 : BUF_X1 port map( A => n9985, Z => n7827);
   U8811 : BUF_X1 port map( A => DP_OP_751_130_6421_n609, Z => n7817);
   U8812 : BUF_X1 port map( A => n10016, Z => n7824);
   U8813 : BUF_X1 port map( A => n9253, Z => n7898);
   U8814 : BUF_X2 port map( A => n10433, Z => n7796);
   U8815 : BUF_X1 port map( A => DP_OP_751_130_6421_n303, Z => n7816);
   U8816 : INV_X1 port map( A => n11790, ZN => n10439);
   U8817 : BUF_X1 port map( A => n9934, Z => n8402);
   U8818 : BUF_X1 port map( A => n10053, Z => n7924);
   U8819 : OR2_X1 port map( A1 => n8415, A2 => n8414, ZN => n8379);
   U8820 : NOR2_X1 port map( A1 => n8111, A2 => n8110, ZN => n8109);
   U8821 : INV_X1 port map( A => n8032, ZN => n7870);
   U8822 : INV_X1 port map( A => n8111, ZN => n8106);
   U8823 : INV_X1 port map( A => n8136, ZN => n8137);
   U8824 : BUF_X1 port map( A => n9122, Z => n7800);
   U8825 : AND2_X2 port map( A1 => n8945, A2 => n8944, ZN => n10032);
   U8826 : BUF_X1 port map( A => n8435, Z => n7801);
   U8827 : CLKBUF_X1 port map( A => n10376, Z => n7903);
   U8828 : NOR2_X1 port map( A1 => n8177, A2 => n8110, ZN => n8108);
   U8829 : NAND2_X2 port map( A1 => n8574, A2 => n11639, ZN => n11640);
   U8830 : INV_X1 port map( A => n8131, ZN => n7802);
   U8831 : INV_X1 port map( A => n8596, ZN => n10376);
   U8832 : AND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_13_port, ZN => n7970);
   U8833 : OR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_10_port, ZN => n8068);
   U8834 : NAND2_X2 port map( A1 => n8573, A2 => n11626, ZN => n11627);
   U8835 : NAND2_X2 port map( A1 => n8573, A2 => n11644, ZN => n11676);
   U8836 : NOR2_X1 port map( A1 => n10393, A2 => n10229, ZN => n8888);
   U8837 : NAND2_X2 port map( A1 => n8574, A2 => n11618, ZN => n11619);
   U8838 : INV_X1 port map( A => n9473, ZN => n7804);
   U8839 : NOR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_27_port, ZN => n8111);
   U8840 : NOR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_19_port, ZN => n7961);
   U8841 : OR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_23_port, ZN => n8027);
   U8842 : INV_X1 port map( A => n9883, ZN => n8021);
   U8843 : OR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_15_port, ZN => n8075);
   U8844 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_21_port, ZN => n7986);
   U8845 : OR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_22_port, ZN => n8011);
   U8846 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_14_port, ZN => n8071);
   U8847 : INV_X1 port map( A => n9528, ZN => n7805);
   U8848 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_15_port, ZN => n8076);
   U8849 : INV_X1 port map( A => n11879, ZN => n7806);
   U8850 : NOR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_27_port, ZN => n8082);
   U8851 : AND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_20_port, ZN => n7900);
   U8852 : AND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_22_port, ZN => n8010);
   U8853 : NAND2_X1 port map( A1 => n8938, A2 => n8200, ZN => 
                           DP_OP_751_130_6421_n1764);
   U8854 : AND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_25_port, ZN => n7871);
   U8855 : AND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_23_port, ZN => n8026);
   U8856 : INV_X1 port map( A => n8177, ZN => n7807);
   U8857 : AND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_28_port, ZN => n8176);
   U8858 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_23_port, ZN => n8025);
   U8859 : OR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_13_port, ZN => n8066);
   U8860 : OR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_20_port, ZN => n7980);
   U8861 : NOR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_28_port, ZN => n8114);
   U8862 : INV_X1 port map( A => DP_OP_1091J1_126_6973_n31, ZN => n7808);
   U8863 : NAND2_X2 port map( A1 => n466, A2 => n465, ZN => n10443);
   U8864 : NAND2_X1 port map( A1 => n8941, A2 => n8942, ZN => n9883);
   U8865 : INV_X1 port map( A => n8601, ZN => n8889);
   U8866 : BUF_X1 port map( A => n10387, Z => n8051);
   U8867 : BUF_X1 port map( A => n10128, Z => n7962);
   U8868 : AND2_X1 port map( A1 => n10128, A2 => n8356, ZN => n8587);
   U8869 : BUF_X1 port map( A => n10226, Z => n8005);
   U8870 : NOR2_X1 port map( A1 => n11976, A2 => DRAM_READY, ZN => n2867);
   U8871 : INV_X2 port map( A => n8566, ZN => n7809);
   U8872 : INV_X1 port map( A => n576, ZN => n11814);
   U8873 : NOR2_X1 port map( A1 => IR_29_port, A2 => n8586, ZN => n10387);
   U8874 : INV_X2 port map( A => DRAMRF_READY, ZN => n11993);
   U8875 : BUF_X1 port map( A => n11973, Z => n8550);
   U8876 : BUF_X1 port map( A => n11054, Z => n8484);
   U8877 : INV_X1 port map( A => n9970, ZN => n7810);
   U8878 : AND2_X2 port map( A1 => n8021, A2 => n8146, ZN => n10103);
   U8879 : NOR2_X2 port map( A1 => n10499, A2 => n10501, ZN => n8217);
   U8880 : OAI211_X2 port map( C1 => n176, C2 => n10405, A => n10404, B => 
                           n10403, ZN => i_ADD_WS1_0_port);
   U8881 : NOR2_X2 port map( A1 => n10498, A2 => n10485, ZN => n8216);
   U8882 : NOR3_X2 port map( A1 => i_ADD_WB_3_port, A2 => n8209, A3 => n8306, 
                           ZN => n11082);
   U8883 : OAI22_X2 port map( A1 => n576, A2 => n11924, B1 => n11922, B2 => 
                           n11153, ZN => n11087);
   U8884 : NOR2_X2 port map( A1 => n10503, A2 => n10500, ZN => n8215);
   U8885 : AOI211_X2 port map( C1 => n7789, C2 => n9557, A => n9556, B => n9555
                           , ZN => n10057);
   U8886 : OAI21_X1 port map( B1 => n8201, B2 => n7929, A => n9106, ZN => 
                           DP_OP_751_130_6421_n609);
   U8887 : INV_X1 port map( A => n11508, ZN => n11507);
   U8888 : BUF_X1 port map( A => n11521, Z => n8524);
   U8889 : AOI211_X2 port map( C1 => n7789, C2 => n9424, A => n9423, B => n9422
                           , ZN => n9922);
   U8890 : NOR2_X2 port map( A1 => RST, A2 => n11078, ZN => n11178);
   U8891 : NOR2_X2 port map( A1 => RST, A2 => n11072, ZN => n11186);
   U8892 : NOR2_X2 port map( A1 => RST, A2 => n11077, ZN => n11174);
   U8893 : NOR2_X2 port map( A1 => RST, A2 => n11086, ZN => n11182);
   U8894 : NOR2_X2 port map( A1 => n10499, A2 => n10502, ZN => n8213);
   U8895 : NOR2_X2 port map( A1 => n10503, A2 => n10500, ZN => n8214);
   U8896 : NOR2_X2 port map( A1 => n10498, A2 => n10486, ZN => n8212);
   U8897 : OAI22_X2 port map( A1 => n8529, A2 => n11891, B1 => n11892, B2 => 
                           n8191, ZN => n11499);
   U8898 : INV_X1 port map( A => n8296, ZN => n8529);
   U8899 : OAI22_X2 port map( A1 => n575, A2 => n11924, B1 => n11922, B2 => 
                           n11281, ZN => n11211);
   U8900 : AOI211_X2 port map( C1 => n9704, C2 => n9541, A => n9540, B => n9539
                           , ZN => n10061);
   U8901 : BUF_X1 port map( A => n11491, Z => n8515);
   U8902 : OAI22_X2 port map( A1 => n7766, A2 => n11886, B1 => n11887, B2 => 
                           n8191, ZN => n11491);
   U8903 : OAI22_X2 port map( A1 => n7766, A2 => n11513, B1 => n11512, B2 => 
                           n8191, ZN => n11514);
   U8904 : NOR2_X2 port map( A1 => n8541, A2 => n11816, ZN => n10961);
   U8905 : NOR2_X2 port map( A1 => n9627, A2 => n11879, ZN => n9586);
   U8906 : NOR2_X2 port map( A1 => n9052, A2 => n9128, ZN => n10117);
   U8907 : AOI22_X2 port map( A1 => n7783, A2 => n11466, B1 => n11659, B2 => 
                           n11281, ZN => n11297);
   U8908 : AOI22_X2 port map( A1 => n7783, A2 => n11319, B1 => n11665, B2 => 
                           n11281, ZN => n11303);
   U8909 : OAI21_X4 port map( B1 => n9102, B2 => n8137, A => n9101, ZN => 
                           DP_OP_751_130_6421_n711);
   U8910 : OAI21_X4 port map( B1 => n9097, B2 => n7929, A => n9096, ZN => 
                           DP_OP_751_130_6421_n813);
   U8911 : OAI21_X4 port map( B1 => n7766, B2 => n11569, A => n8338, ZN => 
                           n11570);
   U8912 : NOR3_X2 port map( A1 => i_ADD_WB_4_port, A2 => i_ADD_WB_3_port, A3 
                           => n8306, ZN => n11642);
   U8913 : INV_X1 port map( A => n9914, ZN => n7821);
   U8914 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n404, B => 
                           DP_OP_751_130_6421_n405, ZN => n7969);
   U8915 : XNOR2_X1 port map( A => n7822, B => n8148, ZN => 
                           DP_OP_751_130_6421_n1746);
   U8916 : OAI22_X1 port map( A1 => n7751, A2 => n8405, B1 => n7726, B2 => 
                           n9495, ZN => n7822);
   U8917 : BUF_X2 port map( A => DP_OP_751_130_6421_n1629, Z => n8145);
   U8918 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1611, B2 => 
                           DP_OP_751_130_6421_n1659, A => 
                           DP_OP_751_130_6421_n1658, ZN => n7891);
   U8919 : INV_X1 port map( A => DP_OP_751_130_6421_n1764, ZN => 
                           DP_OP_751_130_6421_I2);
   U8920 : OR2_X1 port map( A1 => n8621, A2 => n7896, ZN => n8802);
   U8921 : NAND2_X1 port map( A1 => n8618, A2 => n8617, ZN => n8621);
   U8922 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1052, B => n7825, ZN => 
                           DP_OP_751_130_6421_n954);
   U8923 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1053, B => 
                           DP_OP_751_130_6421_n1002, ZN => n7825);
   U8924 : XNOR2_X1 port map( A => n7826, B => DP_OP_751_130_6421_n1350, ZN => 
                           DP_OP_751_130_6421_n1252);
   U8925 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1351, B => 
                           DP_OP_751_130_6421_n1304, ZN => n7826);
   U8926 : AND2_X1 port map( A1 => DP_OP_751_130_6421_n1711, A2 => n7746, ZN =>
                           DP_OP_751_130_6421_n1653);
   U8927 : XNOR2_X1 port map( A => n7841, B => n7837, ZN => n7914);
   U8928 : INV_X4 port map( A => n9156, ZN => n9168);
   U8929 : INV_X1 port map( A => n8874, ZN => n8856);
   U8930 : NAND2_X1 port map( A1 => n8856, A2 => n8855, ZN => n10199);
   U8931 : INV_X1 port map( A => n8193, ZN => n7840);
   U8932 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n1764, A2 => n7755, ZN => 
                           n7844);
   U8933 : XNOR2_X1 port map( A => n7829, B => n8148, ZN => 
                           DP_OP_751_130_6421_n1745);
   U8934 : OAI22_X1 port map( A1 => n7756, A2 => n9495, B1 => n7726, B2 => 
                           n9692, ZN => n7829);
   U8935 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n673, B => n8031, ZN => 
                           DP_OP_751_130_6421_n574);
   U8936 : NAND2_X1 port map( A1 => n8015, A2 => n8043, ZN => 
                           DP_OP_751_130_6421_n66);
   U8937 : XNOR2_X1 port map( A => n7836, B => n7835, ZN => 
                           DP_OP_751_130_6421_n1462);
   U8938 : XNOR2_X1 port map( A => n7892, B => DP_OP_751_130_6421_n1658, ZN => 
                           n7835);
   U8939 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1561, B => 
                           DP_OP_751_130_6421_n1511, ZN => n7836);
   U8940 : NOR2_X2 port map( A1 => DP_OP_751_130_6421_n980, A2 => 
                           DP_OP_751_130_6421_n981, ZN => n8155);
   U8941 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1453, B => 
                           DP_OP_751_130_6421_n1406, ZN => n7911);
   U8942 : XNOR2_X1 port map( A => n7912, B => n7837, ZN => n7916);
   U8943 : INV_X1 port map( A => n8148, ZN => n7837);
   U8944 : XNOR2_X1 port map( A => n7838, B => n7948, ZN => 
                           DP_OP_751_130_6421_n1454);
   U8945 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1553, B => 
                           DP_OP_751_130_6421_n1507, ZN => n7838);
   U8946 : INV_X4 port map( A => n9060, ZN => n9130);
   U8947 : AOI21_X2 port map( B1 => n7840, B2 => DataPath_i_PIPLIN_B_5_port, A 
                           => n7839, ZN => n8560);
   U8948 : OAI22_X1 port map( A1 => n8134, A2 => n7714, B1 => n7726, B2 => 
                           n9600, ZN => n7841);
   U8949 : XNOR2_X1 port map( A => n7843, B => n7842, ZN => n7908);
   U8950 : INV_X1 port map( A => n8147, ZN => n7842);
   U8951 : OAI22_X1 port map( A1 => n7750, A2 => n9692, B1 => n7726, B2 => 
                           n9312, ZN => n7843);
   U8952 : OAI211_X1 port map( C1 => n9165, C2 => DP_OP_751_130_6421_I2, A => 
                           n7844, B => n7845, ZN => n9061);
   U8953 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1731, A2 => n9165, ZN 
                           => n7845);
   U8954 : NOR2_X1 port map( A1 => n7850, A2 => n7847, ZN => n7846);
   U8955 : INV_X1 port map( A => n7853, ZN => n7847);
   U8956 : NOR2_X1 port map( A1 => n8926, A2 => n206, ZN => n7852);
   U8957 : NOR2_X1 port map( A1 => n8926, A2 => n7854, ZN => n7853);
   U8958 : INV_X1 port map( A => n10346, ZN => n7854);
   U8959 : OAI211_X1 port map( C1 => n8202, C2 => n8389, A => n7855, B => n7607
                           , ZN => n8388);
   U8960 : NAND2_X1 port map( A1 => n10324, A2 => n7856, ZN => n7855);
   U8961 : NAND2_X1 port map( A1 => n10324, A2 => n10251, ZN => n7860);
   U8962 : OAI21_X1 port map( B1 => n8388, B2 => n8386, A => n8273, ZN => n8385
                           );
   U8963 : AND2_X1 port map( A1 => n7860, A2 => n7858, ZN => n10252);
   U8964 : INV_X1 port map( A => n7936, ZN => n7858);
   U8965 : OAI21_X1 port map( B1 => n8009, B2 => n7866, A => n7865, ZN => 
                           DP_OP_1091J1_126_6973_n6);
   U8966 : AND2_X1 port map( A1 => n7861, A2 => n7862, ZN => n8084);
   U8967 : OR2_X1 port map( A1 => n7725, A2 => n7864, ZN => n7861);
   U8968 : OR2_X1 port map( A1 => n8009, A2 => n8033, ZN => n7872);
   U8969 : AOI21_X1 port map( B1 => n10093, B2 => n10429, A => n7978, ZN => 
                           n7873);
   U8970 : AOI21_X1 port map( B1 => n8187, B2 => n7802, A => n7808, ZN => n8127
                           );
   U8971 : NAND2_X1 port map( A1 => n7881, A2 => DP_OP_751_130_6421_n79, ZN => 
                           DP_OP_751_130_6421_n74);
   U8972 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n80, A2 => n8159, ZN => 
                           n7881);
   U8973 : XNOR2_X1 port map( A => n7888, B => n7886, ZN => 
                           DP_OP_751_130_6421_n1156);
   U8974 : XNOR2_X1 port map( A => n7887, B => DP_OP_751_130_6421_n1352, ZN => 
                           n7886);
   U8975 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1353, B => 
                           DP_OP_751_130_6421_n1305, ZN => n7887);
   U8976 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1255, B => 
                           DP_OP_751_130_6421_n1205, ZN => n7888);
   U8977 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1651, B2 => 
                           DP_OP_751_130_6421_n1607, A => n7958, ZN => n7957);
   U8978 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n571, B => n8008, ZN => 
                           DP_OP_751_130_6421_n472);
   U8979 : NAND2_X1 port map( A1 => n10387, A2 => n8598, ZN => n10373);
   U8980 : NOR2_X1 port map( A1 => n167, A2 => n8195, ZN => n8598);
   U8981 : XNOR2_X1 port map( A => n7889, B => DP_OP_751_130_6421_n1054, ZN => 
                           DP_OP_751_130_6421_n956);
   U8982 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1055, B => 
                           DP_OP_751_130_6421_n1003, ZN => n7889);
   U8983 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1659, B => 
                           DP_OP_751_130_6421_n1611, ZN => n7892);
   U8984 : BUF_X1 port map( A => DP_OP_751_130_6421_n68, Z => n7895);
   U8985 : AOI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n13, B2 => n7980, A 
                           => n7900, ZN => n7979);
   U8986 : OAI21_X1 port map( B1 => n7902, B2 => n7961, A => n7901, ZN => 
                           DP_OP_1091J1_126_6973_n13);
   U8987 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_19_port, ZN => n7901);
   U8988 : INV_X1 port map( A => DP_OP_1091J1_126_6973_n14, ZN => n7902);
   U8989 : XNOR2_X1 port map( A => n7907, B => n7906, ZN => 
                           DP_OP_751_130_6421_n1348);
   U8990 : XNOR2_X1 port map( A => n7946, B => n7944, ZN => n7906);
   U8991 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1447, B => 
                           DP_OP_751_130_6421_n1403, ZN => n7907);
   U8992 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1406, B2 => 
                           DP_OP_751_130_6421_n1453, A => 
                           DP_OP_751_130_6421_n1452, ZN => n7910);
   U8993 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1714, B => n7908, ZN => 
                           DP_OP_751_130_6421_n1660);
   U8994 : XNOR2_X1 port map( A => n7911, B => DP_OP_751_130_6421_n1452, ZN => 
                           DP_OP_751_130_6421_n1354);
   U8995 : OAI22_X1 port map( A1 => n7756, A2 => n9600, B1 => n7726, B2 => 
                           n9528, ZN => n7912);
   U8996 : OR2_X1 port map( A1 => n8567, A2 => n8268, ZN => n8200);
   U8997 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1711, B => n7914, ZN => 
                           DP_OP_751_130_6421_n1654);
   U8998 : NAND2_X1 port map( A1 => n8058, A2 => n8057, ZN => 
                           DP_OP_751_130_6421_n1567);
   U8999 : XNOR2_X1 port map( A => n7915, B => n8148, ZN => 
                           DP_OP_751_130_6421_n1736);
   U9000 : OAI22_X1 port map( A1 => n7756, A2 => n9473, B1 => n7726, B2 => 
                           n9660, ZN => n7915);
   U9001 : INV_X1 port map( A => DP_OP_751_130_6421_n1737, ZN => n7921);
   U9002 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1707, B => n7921, ZN => 
                           DP_OP_751_130_6421_n1646);
   U9003 : XNOR2_X1 port map( A => n7916, B => DP_OP_751_130_6421_n1710, ZN => 
                           DP_OP_751_130_6421_n1652);
   U9004 : NAND2_X1 port map( A1 => n10128, A2 => n10226, ZN => n10150);
   U9005 : NOR2_X1 port map( A1 => IR_26_port, A2 => n10149, ZN => n10226);
   U9006 : XNOR2_X1 port map( A => n7917, B => n8148, ZN => 
                           DP_OP_751_130_6421_n1743);
   U9007 : OAI22_X1 port map( A1 => n7750, A2 => n9312, B1 => n7726, B2 => 
                           n9961, ZN => n7917);
   U9008 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_20_port, B => 
                           n7774, ZN => DP_OP_751_130_6421_n1714);
   U9009 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n982, A2 => 
                           DP_OP_751_130_6421_n1080, ZN => 
                           DP_OP_751_130_6421_n105);
   U9010 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1081, B => n8006, ZN => 
                           DP_OP_751_130_6421_n982);
   U9011 : NOR2_X1 port map( A1 => n7919, A2 => n8918, ZN => n10348);
   U9012 : AOI21_X1 port map( B1 => n10356, B2 => n10358, A => n7920, ZN => 
                           n7919);
   U9013 : NAND2_X1 port map( A1 => n7780, A2 => n8919, ZN => n7920);
   U9014 : BUF_X2 port map( A => n9063, Z => n8443);
   U9015 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_25_port, B => 
                           n7774, ZN => DP_OP_751_130_6421_n1709);
   U9016 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n463, B => n7939, ZN => 
                           n7938);
   U9017 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n462, B => n7938, ZN => 
                           n7937);
   U9018 : AND2_X2 port map( A1 => n8359, A2 => DP_OP_751_130_6421_n1764, ZN =>
                           n9041);
   U9019 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1706, B => n7923, ZN => 
                           DP_OP_751_130_6421_n1644);
   U9020 : INV_X1 port map( A => DP_OP_751_130_6421_n1736, ZN => n7923);
   U9021 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_19_port, B => 
                           n7774, ZN => DP_OP_751_130_6421_n1715);
   U9022 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_24_port, B => 
                           n7774, ZN => DP_OP_751_130_6421_n1710);
   U9023 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_23_port, B => 
                           n7774, ZN => DP_OP_751_130_6421_n1711);
   U9024 : BUF_X1 port map( A => DP_OP_751_130_6421_n74, Z => n7925);
   U9025 : AOI21_X1 port map( B1 => n7927, B2 => n8815, A => n8774, ZN => n8795
                           );
   U9026 : NAND2_X1 port map( A1 => n8854, A2 => n7928, ZN => n7927);
   U9027 : AND2_X1 port map( A1 => n8737, A2 => n8738, ZN => n7928);
   U9028 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_28_port, B => 
                           n7774, ZN => DP_OP_751_130_6421_n1706);
   U9029 : XNOR2_X1 port map( A => n7930, B => n8148, ZN => 
                           DP_OP_751_130_6421_n1738);
   U9030 : OAI22_X1 port map( A1 => n7751, A2 => n9934, B1 => n7726, B2 => 
                           n9504, ZN => n7930);
   U9031 : NAND2_X1 port map( A1 => n10280, A2 => n7931, ZN => n10415);
   U9032 : AND2_X1 port map( A1 => n10271, A2 => IRAM_ADDRESS_29_port, ZN => 
                           n7931);
   U9033 : XNOR2_X1 port map( A => n7935, B => n7934, ZN => 
                           DP_OP_751_130_6421_n1550);
   U9034 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1649, B => 
                           DP_OP_751_130_6421_n1606, ZN => n7935);
   U9035 : AND2_X1 port map( A1 => n10250, A2 => IRAM_ADDRESS_19_port, ZN => 
                           n7936);
   U9036 : NAND2_X1 port map( A1 => n7992, A2 => n7991, ZN => 
                           DP_OP_751_130_6421_n1449);
   U9037 : XNOR2_X1 port map( A => n7945, B => DP_OP_751_130_6421_n1642, ZN => 
                           n7944);
   U9038 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1603, B => 
                           DP_OP_751_130_6421_n1643, ZN => n7945);
   U9039 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1545, B => 
                           DP_OP_751_130_6421_n1503, ZN => n7946);
   U9040 : BUF_X1 port map( A => DP_OP_751_130_6421_n80, Z => n7950);
   U9041 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n67, A2 => n7951, ZN => 
                           n8015);
   U9042 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n470, A2 => 
                           DP_OP_751_130_6421_n471, ZN => n7951);
   U9043 : NAND2_X1 port map( A1 => n8017, A2 => n8016, ZN => 
                           DP_OP_751_130_6421_n67);
   U9044 : XNOR2_X1 port map( A => n7955, B => n7954, ZN => 
                           DP_OP_751_130_6421_n1558);
   U9045 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1657, B => 
                           DP_OP_751_130_6421_n1610, ZN => n7955);
   U9046 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1734, B => n7960, ZN => 
                           DP_OP_751_130_6421_n1640);
   U9047 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_30_port, B => 
                           n8146, ZN => n7960);
   U9048 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n367, B => n7997, ZN => 
                           DP_OP_751_130_6421_n268);
   U9049 : XNOR2_X1 port map( A => n7966, B => n7965, ZN => 
                           DP_OP_751_130_6421_n1352);
   U9050 : XNOR2_X1 port map( A => n7993, B => DP_OP_751_130_6421_n1548, ZN => 
                           n7965);
   U9051 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1451, B => 
                           DP_OP_751_130_6421_n1405, ZN => n7966);
   U9052 : NOR2_X1 port map( A1 => n7967, A2 => n8156, ZN => 
                           DP_OP_751_130_6421_n99);
   U9053 : NOR2_X1 port map( A1 => n8155, A2 => n7968, ZN => n7967);
   U9054 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n111, A2 => n8152, ZN => 
                           n7968);
   U9055 : OAI21_X1 port map( B1 => n7972, B2 => n7971, A => n10385, ZN => 
                           n7977);
   U9056 : OAI21_X1 port map( B1 => n10200, B2 => n8888, A => n7608, ZN => 
                           n7971);
   U9057 : INV_X1 port map( A => n10373, ZN => n10389);
   U9058 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n74, A2 => n8158, ZN => 
                           n8038);
   U9059 : INV_X1 port map( A => n8419, ZN => n8397);
   U9060 : AOI21_X1 port map( B1 => n10329, B2 => n10327, A => n10326, ZN => 
                           n10324);
   U9061 : AOI21_X1 port map( B1 => n7728, B2 => n10248, A => n7975, ZN => 
                           n10329);
   U9062 : AND2_X1 port map( A1 => n10247, A2 => IRAM_ADDRESS_17_port, ZN => 
                           n7975);
   U9063 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_26_port, B => 
                           n7774, ZN => DP_OP_751_130_6421_n1708);
   U9064 : NAND2_X1 port map( A1 => n7977, A2 => n7976, ZN => n8912);
   U9065 : AND2_X1 port map( A1 => n8893, A2 => n8007, ZN => n7976);
   U9066 : OAI21_X1 port map( B1 => n8568, B2 => n8235, A => n7984, ZN => n9191
                           );
   U9067 : NAND2_X1 port map( A1 => n8193, A2 => DataPath_i_PIPLIN_IN2_0_port, 
                           ZN => n7984);
   U9068 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_2_26_port, B => 
                           n7772, ZN => DP_OP_751_130_6421_n1606);
   U9069 : INV_X1 port map( A => n7987, ZN => DP_OP_1091J1_126_6973_n10);
   U9070 : AOI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n11, B2 => n8011, A 
                           => n8010, ZN => n7987);
   U9071 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_21_port, ZN => n7988);
   U9072 : NOR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_21_port, ZN => n7989);
   U9073 : BUF_X1 port map( A => n8037, Z => n7990);
   U9074 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_2_25_port, B => 
                           n7772, ZN => DP_OP_751_130_6421_n1607);
   U9075 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1549, B => 
                           DP_OP_751_130_6421_n1505, ZN => n7993);
   U9076 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_2_16_port, B => 
                           n7772, ZN => DP_OP_751_130_6421_n1616);
   U9077 : BUF_X2 port map( A => n7842, Z => n7998);
   U9078 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_2_27_port, B => 
                           n7772, ZN => DP_OP_751_130_6421_n1605);
   U9079 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_2_22_port, B => 
                           n7772, ZN => DP_OP_751_130_6421_n1610);
   U9080 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_2_21_port, B => 
                           n7772, ZN => DP_OP_751_130_6421_n1611);
   U9081 : XNOR2_X1 port map( A => n8000, B => n8048, ZN => n8047);
   U9082 : NAND2_X1 port map( A1 => n8002, A2 => n8001, ZN => n8000);
   U9083 : NAND2_X1 port map( A1 => n10415, A2 => IRAM_ADDRESS_30_port, ZN => 
                           n8001);
   U9084 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_27_port, B => 
                           n7774, ZN => DP_OP_751_130_6421_n1707);
   U9085 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_21_port, B => 
                           n7774, ZN => DP_OP_751_130_6421_n1713);
   U9086 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_29_port, B => 
                           n7774, ZN => DP_OP_751_130_6421_n1705);
   U9087 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_22_port, B => 
                           n7774, ZN => DP_OP_751_130_6421_n1712);
   U9088 : XNOR2_X1 port map( A => DataPath_ALUhw_MULT_mux_out_1_14_port, B => 
                           n7774, ZN => DP_OP_751_130_6421_n1720);
   U9089 : AOI21_X1 port map( B1 => n8012, B2 => n8883, A => n8882, ZN => n8884
                           );
   U9090 : NAND2_X1 port map( A1 => n8874, A2 => n8013, ZN => n8012);
   U9091 : AND2_X1 port map( A1 => n8871, A2 => n8014, ZN => n8013);
   U9092 : AND2_X1 port map( A1 => n8872, A2 => n8873, ZN => n8014);
   U9093 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n68, A2 => n8018, ZN => 
                           n8017);
   U9094 : INV_X1 port map( A => n8221, ZN => n8567);
   U9095 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_24_port, ZN => n8032);
   U9096 : NOR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_24_port, ZN => n8033);
   U9097 : NAND2_X1 port map( A1 => n8035, A2 => n8034, ZN => 
                           DP_OP_751_130_6421_n68);
   U9098 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n572, A2 => 
                           DP_OP_751_130_6421_n573, ZN => n8034);
   U9099 : NAND2_X1 port map( A1 => n8037, A2 => n8036, ZN => n8035);
   U9100 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n572, A2 => 
                           DP_OP_751_130_6421_n573, ZN => n8036);
   U9101 : NAND2_X1 port map( A1 => n8038, A2 => DP_OP_751_130_6421_n73, ZN => 
                           n8037);
   U9102 : NAND2_X1 port map( A1 => n8040, A2 => n8074, ZN => 
                           DP_OP_1091J1_126_6973_n17);
   U9103 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n18, A2 => n8075, ZN 
                           => n8040);
   U9104 : OAI21_X1 port map( B1 => n8065, B2 => n8073, A => n8072, ZN => 
                           DP_OP_1091J1_126_6973_n18);
   U9105 : NAND2_X1 port map( A1 => n10272, A2 => n8070, ZN => n10416);
   U9106 : NAND2_X1 port map( A1 => n8103, A2 => n8098, ZN => n10272);
   U9107 : NAND2_X1 port map( A1 => n7595, A2 => DP_OP_751_130_6421_n471, ZN =>
                           n8043);
   U9108 : NAND2_X1 port map( A1 => n8044, A2 => n8067, ZN => 
                           DP_OP_1091J1_126_6973_n22);
   U9109 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n23, A2 => n8068, ZN 
                           => n8044);
   U9110 : OAI21_X1 port map( B1 => n7744, B2 => n8046, A => n8045, ZN => 
                           DP_OP_1091J1_126_6973_n23);
   U9111 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_9_port, ZN => n8045);
   U9112 : NOR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_9_port, ZN => n8046);
   U9113 : OAI21_X1 port map( B1 => n8047, B2 => n7757, A => n10419, ZN => 
                           n7030);
   U9114 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n370, A2 => 
                           DP_OP_751_130_6421_n468, ZN => n8050);
   U9115 : XNOR2_X1 port map( A => n8063, B => n8061, ZN => 
                           DP_OP_751_130_6421_n1470);
   U9116 : XNOR2_X1 port map( A => n8062, B => DP_OP_751_130_6421_n1666, ZN => 
                           n8061);
   U9117 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1615, B => 
                           DP_OP_751_130_6421_n1667, ZN => n8062);
   U9118 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1569, B => 
                           DP_OP_751_130_6421_n1515, ZN => n8063);
   U9119 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1458, B => n8064, ZN => 
                           DP_OP_751_130_6421_n1360);
   U9120 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1459, B => 
                           DP_OP_751_130_6421_n1409, ZN => n8064);
   U9121 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n22, A2 => 
                           DP_OP_1091J1_126_6973_n31, ZN => n8185);
   U9122 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_10_port, ZN => n8067);
   U9123 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_14_port, ZN => n8072);
   U9124 : NOR2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_14_port, ZN => n8073);
   U9125 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n17, A2 => 
                           DP_OP_1091J1_126_6973_n31, ZN => n8173);
   U9126 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_15_port, ZN => n8074);
   U9127 : NAND2_X1 port map( A1 => n8123, A2 => n8143, ZN => n8122);
   U9128 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n75, B => n7808, ZN =>
                           n8143);
   U9129 : XNOR2_X1 port map( A => n8079, B => n7612, ZN => C620_DATA2_31);
   U9130 : AOI21_X1 port map( B1 => n8080, B2 => n8178, A => n8112, ZN => n8079
                           );
   U9131 : AOI21_X1 port map( B1 => DP_OP_1091J1_126_6973_n6, B2 => 
                           DP_OP_1091J1_126_6973_n31, A => n8081, ZN => n8080);
   U9132 : NAND2_X1 port map( A1 => n8133, A2 => n8177, ZN => n8081);
   U9133 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n6, A2 => 
                           DataPath_WRF_CUhw_curr_addr_27_port, ZN => n8178);
   U9134 : NOR2_X1 port map( A1 => n8083, A2 => n7778, ZN => 
                           DRAMRF_ADDRESS_28_port);
   U9135 : XNOR2_X1 port map( A => n8084, B => n7613, ZN => n8083);
   U9136 : OAI211_X1 port map( C1 => n8085, C2 => n8087, A => n8086, B => n8269
                           , ZN => n8854);
   U9137 : INV_X1 port map( A => n8682, ZN => n8085);
   U9138 : AOI21_X1 port map( B1 => n8691, B2 => n8805, A => n8093, ZN => n8092
                           );
   U9139 : INV_X1 port map( A => n8845, ZN => n8093);
   U9140 : AND2_X1 port map( A1 => n8691, A2 => n8842, ZN => n8094);
   U9141 : NAND2_X1 port map( A1 => n10295, A2 => n10265, ZN => n8103);
   U9142 : OAI21_X2 port map( B1 => n10295, B2 => n8097, A => n8095, ZN => 
                           n10280);
   U9143 : NOR2_X1 port map( A1 => n10264, A2 => n8102, ZN => n8101);
   U9144 : INV_X1 port map( A => n10288, ZN => n8102);
   U9145 : OAI21_X1 port map( B1 => n8115, B2 => n8116, A => n8117, ZN => n8142
                           );
   U9146 : NAND2_X1 port map( A1 => n8124, A2 => n8122, ZN => 
                           DP_OP_1091J1_126_6973_n29);
   U9147 : OR2_X1 port map( A1 => n7748, A2 => n177, ZN => n10237);
   U9148 : INV_X2 port map( A => n9041, ZN => n8134);
   U9149 : OAI21_X1 port map( B1 => intadd_0_n8, B2 => intadd_0_n6, A => 
                           intadd_0_n7, ZN => n8135);
   U9150 : OAI21_X1 port map( B1 => intadd_0_n8, B2 => intadd_0_n6, A => 
                           intadd_0_n7, ZN => intadd_0_CO);
   U9151 : AOI21_X1 port map( B1 => n10358, B2 => n10356, A => n10355, ZN => 
                           n8138);
   U9152 : AOI21_X1 port map( B1 => n8934, B2 => n8933, A => n8932, ZN => n8139
                           );
   U9153 : NAND2_X1 port map( A1 => n10422, A2 => n8603, ZN => n8140);
   U9154 : NAND2_X1 port map( A1 => n10422, A2 => n8603, ZN => n8703);
   U9155 : OR3_X2 port map( A1 => n8703, A2 => n177, A3 => 
                           CU_I_CW_ID_UNSIGNED_ID_port, ZN => n8829);
   U9156 : AND2_X1 port map( A1 => C620_DATA2_29, A2 => n8277, ZN => n8395);
   U9157 : AND2_X1 port map( A1 => C620_DATA2_29, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_29_port);
   U9158 : AOI21_X1 port map( B1 => n8928, B2 => n8927, A => n8926, ZN => n8141
                           );
   U9159 : AND2_X1 port map( A1 => C620_DATA2_30, A2 => n8277, ZN => n8394);
   U9160 : AND2_X1 port map( A1 => C620_DATA2_30, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_30_port);
   U9161 : NOR2_X1 port map( A1 => n10442, A2 => n8379, ZN => n11803);
   U9162 : AOI21_X1 port map( B1 => n11803, B2 => n8594, A => n8593, ZN => 
                           n8412);
   U9163 : INV_X1 port map( A => DP_OP_751_130_6421_n115, ZN => 
                           DP_OP_751_130_6421_n113);
   U9164 : INV_X1 port map( A => DP_OP_751_130_6421_n131, ZN => 
                           DP_OP_751_130_6421_n129);
   U9165 : INV_X1 port map( A => DP_OP_751_130_6421_n145, ZN => 
                           DP_OP_751_130_6421_n143);
   U9166 : INV_X1 port map( A => DP_OP_751_130_6421_n153, ZN => 
                           DP_OP_751_130_6421_n151);
   U9167 : INV_X1 port map( A => DP_OP_751_130_6421_n167, ZN => 
                           DP_OP_751_130_6421_n165);
   U9168 : INV_X1 port map( A => DP_OP_751_130_6421_n174, ZN => 
                           DP_OP_751_130_6421_n172);
   U9169 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_31_port, ZN => 
                           DP_OP_751_130_6421_n1768);
   U9170 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_29_port, ZN => 
                           DP_OP_751_130_6421_n1770);
   U9171 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_27_port, ZN => 
                           DP_OP_751_130_6421_n1772);
   U9172 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_25_port, ZN => 
                           DP_OP_751_130_6421_n1774);
   U9173 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_22_port, ZN => 
                           DP_OP_751_130_6421_n1777);
   U9174 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_17_port, ZN => 
                           DP_OP_751_130_6421_n1782);
   U9175 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_16_port, ZN => 
                           DP_OP_751_130_6421_n1783);
   U9176 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_14_port, ZN => 
                           DP_OP_751_130_6421_n1785);
   U9177 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_12_port, ZN => 
                           DP_OP_751_130_6421_n1787);
   U9178 : INV_X1 port map( A => DP_OP_751_130_6421_n81, ZN => 
                           DP_OP_751_130_6421_n179);
   U9179 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_9_port, ZN => 
                           DP_OP_751_130_6421_n1790);
   U9180 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_8_port, ZN => 
                           DP_OP_751_130_6421_n1791);
   U9181 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_5_port, ZN => 
                           DP_OP_751_130_6421_n1794);
   U9182 : INV_X1 port map( A => DataPath_ALUhw_MULT_mux_out_0_4_port, ZN => 
                           DP_OP_751_130_6421_n1795);
   U9183 : INV_X1 port map( A => DP_OP_751_130_6421_n89, ZN => 
                           DP_OP_751_130_6421_n181);
   U9184 : INV_X1 port map( A => DP_OP_751_130_6421_n97, ZN => 
                           DP_OP_751_130_6421_n183);
   U9185 : INV_X1 port map( A => DP_OP_751_130_6421_n125, ZN => 
                           DP_OP_751_130_6421_n190);
   U9186 : INV_X1 port map( A => DP_OP_751_130_6421_n139, ZN => 
                           DP_OP_751_130_6421_n193);
   U9187 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n147, B2 => 
                           DP_OP_751_130_6421_n149, A => 
                           DP_OP_751_130_6421_n148, ZN => 
                           DP_OP_751_130_6421_n146);
   U9188 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n97, B2 => 
                           DP_OP_751_130_6421_n99, A => DP_OP_751_130_6421_n98,
                           ZN => DP_OP_751_130_6421_n96);
   U9189 : AOI21_X1 port map( B1 => n8161, B2 => DP_OP_751_130_6421_n146, A => 
                           DP_OP_751_130_6421_n143, ZN => 
                           DP_OP_751_130_6421_n141);
   U9190 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n139, B2 => 
                           DP_OP_751_130_6421_n141, A => 
                           DP_OP_751_130_6421_n140, ZN => 
                           DP_OP_751_130_6421_n138);
   U9191 : NAND2_X1 port map( A1 => n8157, A2 => DP_OP_751_130_6421_n153, ZN =>
                           DP_OP_751_130_6421_n23);
   U9192 : XOR2_X1 port map( A => DP_OP_751_130_6421_n8, B => n7876, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_52_port);
   U9193 : XNOR2_X1 port map( A => n7605, B => DP_OP_751_130_6421_n9, ZN => 
                           DataPath_ALUhw_i_Q_EXTENDED_51_port);
   U9194 : XOR2_X1 port map( A => DP_OP_751_130_6421_n20, B => 
                           DP_OP_751_130_6421_n141, Z => 
                           DataPath_ALUhw_i_Q_EXTENDED_40_port);
   U9195 : OAI21_X1 port map( B1 => n8154, B2 => n8155, A => 
                           DP_OP_751_130_6421_n103, ZN => n8156);
   U9196 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1186, A2 => 
                           DP_OP_751_130_6421_n1284, ZN => 
                           DP_OP_751_130_6421_n123);
   U9197 : INV_X1 port map( A => DP_OP_751_130_6421_n109, ZN => n8150);
   U9198 : INV_X1 port map( A => DP_OP_751_130_6421_n105, ZN => n8151);
   U9199 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n980, A2 => 
                           DP_OP_751_130_6421_n981, ZN => 
                           DP_OP_751_130_6421_n103);
   U9200 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n1592, A2 => 
                           DP_OP_751_130_6421_n1593, ZN => n8157);
   U9201 : NOR2_X1 port map( A1 => DP_OP_751_130_6421_n1082, A2 => 
                           DP_OP_751_130_6421_n1083, ZN => 
                           DP_OP_751_130_6421_n109);
   U9202 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n574, A2 => 
                           DP_OP_751_130_6421_n672, ZN => n8158);
   U9203 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n674, A2 => 
                           DP_OP_751_130_6421_n675, ZN => n8159);
   U9204 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n1084, A2 => 
                           DP_OP_751_130_6421_n1182, ZN => n8168);
   U9205 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n1186, A2 => 
                           DP_OP_751_130_6421_n1284, ZN => n8163);
   U9206 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n1388, A2 => 
                           DP_OP_751_130_6421_n1389, ZN => n8160);
   U9207 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n1490, A2 => 
                           DP_OP_751_130_6421_n1491, ZN => n8161);
   U9208 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n1594, A2 => 
                           DP_OP_751_130_6421_n1692, ZN => n8162);
   U9209 : AND2_X1 port map( A1 => DP_OP_751_130_6421_n170, A2 => 
                           DP_OP_751_130_6421_n172, ZN => n8167);
   U9210 : AOI21_X1 port map( B1 => n8157, B2 => DP_OP_751_130_6421_n154, A => 
                           DP_OP_751_130_6421_n151, ZN => 
                           DP_OP_751_130_6421_n149);
   U9211 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n1288, A2 => 
                           DP_OP_751_130_6421_n1386, ZN => n8166);
   U9212 : AOI21_X1 port map( B1 => DP_OP_751_130_6421_n132, B2 => n8166, A => 
                           DP_OP_751_130_6421_n129, ZN => 
                           DP_OP_751_130_6421_n127);
   U9213 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n127, B2 => 
                           DP_OP_751_130_6421_n125, A => 
                           DP_OP_751_130_6421_n126, ZN => 
                           DP_OP_751_130_6421_n124);
   U9214 : NAND2_X1 port map( A1 => n8151, A2 => n8150, ZN => n8152);
   U9215 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n105, B2 => 
                           DP_OP_751_130_6421_n110, A => 
                           DP_OP_751_130_6421_n106, ZN => n8153);
   U9216 : INV_X1 port map( A => n8153, ZN => n8154);
   U9217 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n878, A2 => 
                           DP_OP_751_130_6421_n879, ZN => n8165);
   U9218 : AOI21_X1 port map( B1 => DP_OP_751_130_6421_n96, B2 => n8165, A => 
                           n7691, ZN => DP_OP_751_130_6421_n91);
   U9219 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n91, B2 => 
                           DP_OP_751_130_6421_n89, A => DP_OP_751_130_6421_n90,
                           ZN => DP_OP_751_130_6421_n88);
   U9220 : OR2_X1 port map( A1 => DP_OP_751_130_6421_n777, A2 => 
                           DP_OP_751_130_6421_n776, ZN => n8164);
   U9221 : AOI21_X1 port map( B1 => DP_OP_751_130_6421_n88, B2 => n8164, A => 
                           n7693, ZN => DP_OP_751_130_6421_n83);
   U9222 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n83, B2 => 
                           DP_OP_751_130_6421_n81, A => DP_OP_751_130_6421_n82,
                           ZN => DP_OP_751_130_6421_n80);
   U9223 : BUF_X1 port map( A => DP_OP_751_130_6421_n1425, Z => n8144);
   U9224 : BUF_X1 port map( A => DP_OP_751_130_6421_n915, Z => n8149);
   U9225 : BUF_X1 port map( A => DP_OP_751_130_6421_I2, Z => n8147);
   U9226 : AND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_30_port, ZN => n8170);
   U9227 : XNOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_30_port, ZN => n8169);
   U9228 : XNOR2_X1 port map( A => n8142, B => n8169, ZN => C620_DATA2_30);
   U9229 : NAND3_X1 port map( A1 => n8173, A2 => n8172, A3 => n8171, ZN => 
                           DP_OP_1091J1_126_6973_n16);
   U9230 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_16_port, ZN => n8171);
   U9231 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n17, A2 => 
                           DataPath_WRF_CUhw_curr_addr_16_port, ZN => n8172);
   U9232 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n17, B => n8174, Z => 
                           C620_DATA2_16);
   U9233 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_16_port, Z => n8174);
   U9234 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_29_port, ZN => n8175);
   U9235 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_27_port, ZN => n8177);
   U9236 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_8_port, ZN => n8179);
   U9237 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n25, A2 => 
                           DataPath_WRF_CUhw_curr_addr_8_port, ZN => n8180);
   U9238 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n25, A2 => 
                           DP_OP_1091J1_126_6973_n31, ZN => n8181);
   U9239 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n25, B => n8182, Z => 
                           C620_DATA2_8);
   U9240 : XOR2_X1 port map( A => DP_OP_1091J1_126_6973_n31, B => 
                           DataPath_WRF_CUhw_curr_addr_8_port, Z => n8182);
   U9241 : NAND3_X1 port map( A1 => n8185, A2 => n8184, A3 => n8183, ZN => 
                           DP_OP_1091J1_126_6973_n21);
   U9242 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n31, A2 => 
                           DataPath_WRF_CUhw_curr_addr_11_port, ZN => n8183);
   U9243 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n22, A2 => 
                           DataPath_WRF_CUhw_curr_addr_11_port, ZN => n8184);
   U9244 : NAND2_X1 port map( A1 => n7779, A2 => 
                           DataPath_WRF_CUhw_curr_addr_3_port, ZN => n8186);
   U9245 : NAND2_X1 port map( A1 => n7779, A2 => 
                           DataPath_WRF_CUhw_curr_addr_2_port, ZN => n8187);
   U9246 : AND2_X1 port map( A1 => C620_DATA2_31, A2 => n8277, ZN => n8393);
   U9247 : INV_X1 port map( A => n11228, ZN => n11227);
   U9248 : INV_X1 port map( A => n11280, ZN => n11279);
   U9249 : INV_X1 port map( A => n11241, ZN => n11240);
   U9250 : INV_X1 port map( A => n11233, ZN => n11232);
   U9251 : INV_X1 port map( A => n11237, ZN => n11236);
   U9252 : INV_X1 port map( A => n11247, ZN => n11246);
   U9253 : BUF_X1 port map( A => n11356, Z => n8512);
   U9254 : BUF_X1 port map( A => n11372, Z => n8513);
   U9255 : BUF_X1 port map( A => n11336, Z => n8508);
   U9256 : BUF_X1 port map( A => n11214, Z => n8501);
   U9257 : AND2_X1 port map( A1 => n8580, A2 => n11217, ZN => n11215);
   U9258 : AOI22_X1 port map( A1 => n7783, A2 => n11450, B1 => n11645, B2 => 
                           n11281, ZN => n11283);
   U9259 : AOI22_X1 port map( A1 => n7783, A2 => n11454, B1 => n11649, B2 => 
                           n11281, ZN => n11287);
   U9260 : AND2_X1 port map( A1 => n8577, A2 => n11330, ZN => n11331);
   U9261 : BUF_X1 port map( A => n11332, Z => n8507);
   U9262 : BUF_X1 port map( A => n11050, Z => n8482);
   U9263 : BUF_X1 port map( A => n11216, Z => n8502);
   U9264 : BUF_X1 port map( A => n11221, Z => n8503);
   U9265 : BUF_X1 port map( A => n11197, Z => n8497);
   U9266 : AOI22_X1 port map( A1 => n7783, A2 => n11451, B1 => n11646, B2 => 
                           n11281, ZN => n11284);
   U9267 : BUF_X1 port map( A => n11210, Z => n8500);
   U9268 : BUF_X1 port map( A => n11089, Z => n8490);
   U9269 : BUF_X1 port map( A => n11508, Z => n8520);
   U9270 : BUF_X1 port map( A => n11906, Z => n8547);
   U9271 : BUF_X1 port map( A => n11008, Z => n8480);
   U9272 : BUF_X1 port map( A => n11895, Z => n8546);
   U9273 : BUF_X1 port map( A => n11135, Z => n8495);
   U9274 : BUF_X1 port map( A => n11074, Z => n8488);
   U9275 : NAND2_X1 port map( A1 => n8573, A2 => n8529, ZN => n11496);
   U9276 : OR2_X1 port map( A1 => n11993, A2 => n10946, ZN => n11832);
   U9277 : INV_X1 port map( A => n8420, ZN => n10404);
   U9278 : INV_X1 port map( A => n8357, ZN => n8360);
   U9279 : NOR2_X1 port map( A1 => n10423, A2 => n174, ZN => i_ADD_RS2_2_port);
   U9280 : BUF_X1 port map( A => n8420, Z => n8422);
   U9281 : BUF_X1 port map( A => n11321, Z => n8505);
   U9282 : BUF_X1 port map( A => n11189, Z => n8496);
   U9283 : BUF_X1 port map( A => n11890, Z => n8545);
   U9284 : BUF_X1 port map( A => n11407, Z => n8514);
   U9285 : BUF_X1 port map( A => n11274, Z => n8504);
   U9286 : BUF_X1 port map( A => n11342, Z => n8510);
   U9287 : BUF_X1 port map( A => n11096, Z => n8492);
   U9288 : BUF_X1 port map( A => n11204, Z => n8499);
   U9289 : BUF_X1 port map( A => n11003, Z => n8479);
   U9290 : BUF_X1 port map( A => n11325, Z => n8506);
   U9291 : BUF_X1 port map( A => n11339, Z => n8509);
   U9292 : BUF_X1 port map( A => n11092, Z => n8491);
   U9293 : BUF_X1 port map( A => n11201, Z => n8498);
   U9294 : BUF_X1 port map( A => n11988, Z => n8553);
   U9295 : NOR2_X1 port map( A1 => RST, A2 => n11987, ZN => n11988);
   U9296 : BUF_X1 port map( A => n11080, Z => n8489);
   U9297 : INV_X2 port map( A => n11409, ZN => n11412);
   U9298 : AND2_X1 port map( A1 => n8581, A2 => n11087, ZN => n11088);
   U9299 : AND2_X1 port map( A1 => n8580, A2 => n11211, ZN => n11209);
   U9300 : INV_X2 port map( A => n11276, ZN => n11281);
   U9301 : AND2_X1 port map( A1 => n8580, A2 => n11504, ZN => n11503);
   U9302 : AND2_X1 port map( A1 => n8581, A2 => n11541, ZN => n11540);
   U9303 : NOR2_X1 port map( A1 => RST, A2 => n8517, ZN => n11501);
   U9304 : AND2_X1 port map( A1 => n8580, A2 => n8524, ZN => n11520);
   U9305 : NOR2_X1 port map( A1 => RST, A2 => n8515, ZN => n11498);
   U9306 : NOR2_X1 port map( A1 => RST, A2 => n8522, ZN => n11516);
   U9307 : NOR2_X1 port map( A1 => RST, A2 => n8486, ZN => n11058);
   U9308 : NOR2_X1 port map( A1 => RST, A2 => n8493, ZN => n11097);
   U9309 : NOR2_X1 port map( A1 => RST, A2 => n8550, ZN => n11975);
   U9310 : NOR2_X1 port map( A1 => RST, A2 => n8484, ZN => n11055);
   U9311 : BUF_X1 port map( A => n10434, Z => n8418);
   U9312 : INV_X1 port map( A => n8561, ZN => DP_OP_751_130_6421_n1527);
   U9313 : INV_X1 port map( A => n8560, ZN => DP_OP_751_130_6421_n1629);
   U9314 : NOR2_X1 port map( A1 => RST, A2 => n11506, ZN => n11508);
   U9315 : NOR2_X1 port map( A1 => RST, A2 => n11541, ZN => n11542);
   U9316 : NOR2_X1 port map( A1 => RST, A2 => n11024, ZN => n11023);
   U9317 : NOR2_X1 port map( A1 => RST, A2 => n11570, ZN => n11571);
   U9318 : AND2_X1 port map( A1 => n8579, A2 => n11533, ZN => n11596);
   U9319 : AND2_X1 port map( A1 => n8580, A2 => n11502, ZN => n11608);
   U9320 : NOR2_X1 port map( A1 => RST, A2 => n8524, ZN => n11522);
   U9321 : AND2_X1 port map( A1 => n8579, A2 => n11535, ZN => n11598);
   U9322 : AND2_X1 port map( A1 => n8579, A2 => n11537, ZN => n11600);
   U9323 : AND2_X1 port map( A1 => n8579, A2 => n11534, ZN => n11597);
   U9324 : AND2_X1 port map( A1 => n8579, A2 => n11529, ZN => n11590);
   U9325 : AND2_X1 port map( A1 => n8579, A2 => n11536, ZN => n11599);
   U9326 : AND2_X1 port map( A1 => n8580, A2 => n11519, ZN => n11612);
   U9327 : AND2_X1 port map( A1 => n8580, A2 => n11539, ZN => n11607);
   U9328 : AND2_X1 port map( A1 => n8579, A2 => n11538, ZN => n11604);
   U9329 : AND2_X1 port map( A1 => n8582, A2 => n11117, ZN => n11169);
   U9330 : AND2_X1 port map( A1 => n8582, A2 => n11115, ZN => n11167);
   U9331 : INV_X1 port map( A => n11846, ZN => n11848);
   U9332 : AND2_X1 port map( A1 => n8582, A2 => n11111, ZN => n11163);
   U9333 : AND2_X1 port map( A1 => n8581, A2 => n11125, ZN => n11177);
   U9334 : AND2_X1 port map( A1 => n8582, A2 => n11114, ZN => n11166);
   U9335 : AND2_X1 port map( A1 => n8582, A2 => n11121, ZN => n11173);
   U9336 : AND2_X1 port map( A1 => n8582, A2 => n11113, ZN => n11165);
   U9337 : AND2_X1 port map( A1 => n8582, A2 => n11103, ZN => n11155);
   U9338 : NAND2_X2 port map( A1 => n11449, A2 => DataPath_RF_c_swin_4_port, ZN
                           => n11153);
   U9339 : INV_X1 port map( A => n7806, ZN => n9531);
   U9340 : INV_X1 port map( A => n7798, ZN => DP_OP_751_130_6421_n1425);
   U9341 : INV_X1 port map( A => n403, ZN => n8561);
   U9342 : AND2_X1 port map( A1 => n7724, A2 => n8583, ZN => n8417);
   U9343 : NOR2_X1 port map( A1 => n10423, A2 => n172, ZN => i_ADD_RS2_4_port);
   U9344 : NOR2_X1 port map( A1 => n10423, A2 => n175, ZN => i_ADD_RS2_1_port);
   U9345 : NAND3_X1 port map( A1 => n10422, A2 => i_RF2, A3 => n10421, ZN => 
                           n10423);
   U9346 : AND2_X1 port map( A1 => n8595, A2 => n8903, ZN => n8604);
   U9347 : OAI21_X1 port map( B1 => i_DATAMEM_WM, B2 => i_DATAMEM_RM, A => 
                           CU_I_CW_MEM_MEM_EN_port, ZN => n11976);
   U9348 : INV_X1 port map( A => n8286, ZN => n8548);
   U9349 : BUF_X1 port map( A => n11987, Z => n8552);
   U9350 : NOR2_X1 port map( A1 => RST, A2 => n11330, ZN => n11332);
   U9351 : AND2_X1 port map( A1 => n8581, A2 => n11264, ZN => n11306);
   U9352 : NOR2_X1 port map( A1 => n825, A2 => n8412, ZN => n11409);
   U9353 : NOR2_X1 port map( A1 => RST, A2 => n11211, ZN => n11210);
   U9354 : NOR2_X1 port map( A1 => n826, A2 => n8412, ZN => n11276);
   U9355 : NOR2_X1 port map( A1 => RST, A2 => n11087, ZN => n11089);
   U9356 : NOR2_X1 port map( A1 => RST, A2 => n7765, ZN => n11752);
   U9357 : NOR2_X1 port map( A1 => RST, A2 => n11504, ZN => n11505);
   U9358 : NOR2_X1 port map( A1 => RST, A2 => n11944, ZN => n11957);
   U9359 : AND2_X1 port map( A1 => n8582, A2 => n11106, ZN => n11158);
   U9360 : AND2_X1 port map( A1 => n8582, A2 => n11110, ZN => n11162);
   U9361 : AND2_X1 port map( A1 => n8579, A2 => n11530, ZN => n11592);
   U9362 : AND2_X1 port map( A1 => n8578, A2 => n11528, ZN => n11589);
   U9363 : AND2_X1 port map( A1 => n8578, A2 => n11525, ZN => n11586);
   U9364 : AND2_X1 port map( A1 => n8578, A2 => n11526, ZN => n11587);
   U9365 : AND2_X1 port map( A1 => n8578, A2 => n11527, ZN => n11588);
   U9366 : AND2_X1 port map( A1 => n8579, A2 => n11532, ZN => n11594);
   U9367 : AND2_X1 port map( A1 => n8579, A2 => n11531, ZN => n11593);
   U9368 : AND2_X1 port map( A1 => n8582, A2 => n11124, ZN => n11176);
   U9369 : AND2_X1 port map( A1 => n8581, A2 => n11132, ZN => n11184);
   U9370 : AND2_X1 port map( A1 => n8582, A2 => n11107, ZN => n11159);
   U9371 : AND2_X1 port map( A1 => n8582, A2 => n11116, ZN => n11168);
   U9372 : AND2_X1 port map( A1 => n8582, A2 => n11109, ZN => n11161);
   U9373 : AND2_X1 port map( A1 => n8582, A2 => n11105, ZN => n11157);
   U9374 : AND2_X1 port map( A1 => n8581, A2 => n11129, ZN => n11181);
   U9375 : AND2_X1 port map( A1 => n8582, A2 => n11104, ZN => n11156);
   U9376 : AND2_X1 port map( A1 => n8582, A2 => n11123, ZN => n11175);
   U9377 : NOR2_X2 port map( A1 => n11831, A2 => n11830, ZN => n10947);
   U9378 : INV_X1 port map( A => n11051, ZN => n11830);
   U9379 : AND2_X1 port map( A1 => n8576, A2 => n11953, ZN => n11919);
   U9380 : NOR2_X1 port map( A1 => n8242, A2 => n8412, ZN => n11041);
   U9381 : NOR2_X2 port map( A1 => n11832, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_15_port, ZN => 
                           n11831);
   U9382 : INV_X1 port map( A => n10428, ZN => n11881);
   U9383 : BUF_X1 port map( A => n9086, Z => n8456);
   U9384 : BUF_X1 port map( A => n9081, Z => n8455);
   U9385 : BUF_X1 port map( A => n9079, Z => n8454);
   U9386 : INV_X1 port map( A => n8221, ZN => n8568);
   U9387 : NAND2_X1 port map( A1 => n10440, A2 => n8582, ZN => n11790);
   U9388 : INV_X1 port map( A => n2867, ZN => n10440);
   U9389 : INV_X1 port map( A => n8604, ZN => n8605);
   U9390 : NAND2_X1 port map( A1 => i_BUSY_WINDOW, A2 => n159, ZN => n8357);
   U9391 : BUF_X1 port map( A => n11623, Z => n8531);
   U9392 : BUF_X1 port map( A => n11636, Z => n8536);
   U9393 : BUF_X1 port map( A => n11631, Z => n8534);
   U9394 : NOR2_X1 port map( A1 => RST, A2 => n11188, ZN => n11189);
   U9395 : NOR2_X1 port map( A1 => RST, A2 => n11398, ZN => n11407);
   U9396 : NOR2_X1 port map( A1 => RST, A2 => n11263, ZN => n11274);
   U9397 : NOR2_X1 port map( A1 => RST, A2 => n11340, ZN => n11342);
   U9398 : NOR2_X1 port map( A1 => RST, A2 => n11093, ZN => n11096);
   U9399 : NOR2_X1 port map( A1 => RST, A2 => n11202, ZN => n11204);
   U9400 : NOR2_X1 port map( A1 => RST, A2 => n10987, ZN => n11003);
   U9401 : NOR2_X1 port map( A1 => RST, A2 => n11323, ZN => n11325);
   U9402 : NOR2_X1 port map( A1 => RST, A2 => n11337, ZN => n11339);
   U9403 : NOR2_X1 port map( A1 => RST, A2 => n11090, ZN => n11092);
   U9404 : NOR2_X1 port map( A1 => RST, A2 => n11198, ZN => n11201);
   U9405 : AND2_X1 port map( A1 => n8577, A2 => n11375, ZN => n11416);
   U9406 : NOR2_X1 port map( A1 => RST, A2 => n11354, ZN => n11356);
   U9407 : NOR2_X1 port map( A1 => RST, A2 => n11081, ZN => n11080);
   U9408 : NOR2_X1 port map( A1 => RST, A2 => n11370, ZN => n11372);
   U9409 : NOR2_X1 port map( A1 => RST, A2 => n11334, ZN => n11336);
   U9410 : AND2_X1 port map( A1 => n8577, A2 => n11396, ZN => n11437);
   U9411 : NOR2_X1 port map( A1 => RST, A2 => n11212, ZN => n11214);
   U9412 : AND2_X1 port map( A1 => n8579, A2 => n11255, ZN => n11293);
   U9413 : AND2_X1 port map( A1 => n8577, A2 => n11376, ZN => n11417);
   U9414 : AND2_X1 port map( A1 => n8577, A2 => n11400, ZN => n11441);
   U9415 : AND2_X1 port map( A1 => n8577, A2 => n11382, ZN => n11423);
   U9416 : NOR2_X1 port map( A1 => RST, A2 => n11048, ZN => n11050);
   U9417 : NOR2_X1 port map( A1 => RST, A2 => n11217, ZN => n11216);
   U9418 : NOR2_X1 port map( A1 => RST, A2 => n11219, ZN => n11221);
   U9419 : NOR2_X1 port map( A1 => RST, A2 => n11196, ZN => n11197);
   U9420 : AND2_X1 port map( A1 => n8577, A2 => n11403, ZN => n11444);
   U9421 : AND2_X1 port map( A1 => n8580, A2 => n11270, ZN => n11313);
   U9422 : INV_X1 port map( A => n11226, ZN => n11277);
   U9423 : AND2_X1 port map( A1 => n8581, A2 => n11256, ZN => n11294);
   U9424 : NOR2_X1 port map( A1 => RST, A2 => n11904, ZN => n11906);
   U9425 : NOR2_X1 port map( A1 => RST, A2 => n11006, ZN => n11008);
   U9426 : NOR2_X1 port map( A1 => RST, A2 => n11893, ZN => n11895);
   U9427 : NOR2_X1 port map( A1 => RST, A2 => n11136, ZN => n11135);
   U9428 : NOR2_X1 port map( A1 => RST, A2 => n11069, ZN => n11074);
   U9429 : AOI22_X1 port map( A1 => n8417, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_4_port, B1 => 
                           n11085, B2 => n11084, ZN => n11922);
   U9430 : AND2_X1 port map( A1 => n8579, A2 => n11932, ZN => n11965);
   U9431 : AND2_X1 port map( A1 => n8572, A2 => n11899, ZN => n11972);
   U9432 : AND2_X1 port map( A1 => n8578, A2 => n11935, ZN => n11969);
   U9433 : AND2_X1 port map( A1 => n8576, A2 => n11934, ZN => n11968);
   U9434 : AOI22_X1 port map( A1 => n8417, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_12_port, B1 => 
                           n11031, B2 => n11084, ZN => n11569);
   U9435 : AOI22_X1 port map( A1 => n8417, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_6_port, B1 => 
                           n10977, B2 => n11084, ZN => n11518);
   U9436 : AOI22_X1 port map( A1 => n10437, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_1_port, B1 => 
                           n11057, B2 => n11084, ZN => n11891);
   U9437 : AOI22_X1 port map( A1 => n8417, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_7_port, B1 => 
                           n11005, B2 => n11084, ZN => n11523);
   U9438 : AND2_X1 port map( A1 => n8580, A2 => n11931, ZN => n11964);
   U9439 : AND2_X1 port map( A1 => n8571, A2 => n11929, ZN => n11962);
   U9440 : AND2_X1 port map( A1 => n8579, A2 => n11898, ZN => n11966);
   U9441 : AND2_X1 port map( A1 => n8579, A2 => n11936, ZN => n11970);
   U9442 : AND2_X1 port map( A1 => n8574, A2 => n11937, ZN => n11971);
   U9443 : AND2_X1 port map( A1 => n8582, A2 => n11927, ZN => n11960);
   U9444 : AND2_X1 port map( A1 => n8576, A2 => n11941, ZN => n11911);
   U9445 : AND2_X1 port map( A1 => n8576, A2 => n11946, ZN => n11912);
   U9446 : AND2_X1 port map( A1 => n8576, A2 => n11903, ZN => n11945);
   U9447 : AND2_X1 port map( A1 => n8576, A2 => n11902, ZN => n11943);
   U9448 : AND2_X1 port map( A1 => n8579, A2 => n11925, ZN => n11958);
   U9449 : AND2_X1 port map( A1 => n8577, A2 => n11928, ZN => n11961);
   U9450 : AND2_X1 port map( A1 => n8579, A2 => n11926, ZN => n11959);
   U9451 : AND2_X1 port map( A1 => n8576, A2 => n11950, ZN => n11916);
   U9452 : OAI22_X1 port map( A1 => n11513, A2 => n11923, B1 => n8219, B2 => 
                           n11512, ZN => n11973);
   U9453 : AOI22_X1 port map( A1 => n10437, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_5_port, B1 => 
                           n10969, B2 => n11084, ZN => n11513);
   U9454 : OAI22_X1 port map( A1 => n576, A2 => n11887, B1 => n11886, B2 => 
                           n8483, ZN => n11054);
   U9455 : NOR2_X1 port map( A1 => n7796, A2 => RST, ZN => n10432);
   U9456 : AND2_X1 port map( A1 => n10429, A2 => n9897, ZN => n10428);
   U9457 : INV_X1 port map( A => n10036, ZN => n10088);
   U9458 : AND2_X1 port map( A1 => n7796, A2 => n217, ZN => n10429);
   U9459 : NOR2_X1 port map( A1 => n11790, A2 => n8301, ZN => n10433);
   U9460 : NAND2_X1 port map( A1 => n10238, A2 => n8605, ZN => n10188);
   U9461 : NOR2_X1 port map( A1 => IR_29_port, A2 => n159, ZN => n8601);
   U9462 : AND2_X1 port map( A1 => n8219, A2 => DataPath_RF_c_swin_4_port, ZN 
                           => n8415);
   U9463 : NOR2_X2 port map( A1 => n163, A2 => n161, ZN => n10128);
   U9464 : BUF_X1 port map( A => n11677, Z => n8539);
   U9465 : BUF_X1 port map( A => n11628, Z => n8533);
   U9466 : BUF_X1 port map( A => n11641, Z => n8538);
   U9467 : BUF_X1 port map( A => n11620, Z => n8530);
   U9468 : BUF_X1 port map( A => n11817, Z => n8541);
   U9469 : BUF_X1 port map( A => n11632, Z => n8535);
   U9470 : BUF_X1 port map( A => n11624, Z => n8532);
   U9471 : BUF_X1 port map( A => n11637, Z => n8537);
   U9472 : INV_X1 port map( A => n11791, ZN => n11981);
   U9473 : NOR2_X1 port map( A1 => RST, A2 => n11241, ZN => n11239);
   U9474 : NOR2_X1 port map( A1 => RST, A2 => n11318, ZN => n11321);
   U9475 : AND2_X1 port map( A1 => n8577, A2 => n11377, ZN => n11418);
   U9476 : AND2_X1 port map( A1 => n8578, A2 => n11381, ZN => n11422);
   U9477 : AND2_X1 port map( A1 => n8577, A2 => n11380, ZN => n11421);
   U9478 : AND2_X1 port map( A1 => n8577, A2 => n11378, ZN => n11419);
   U9479 : AND2_X1 port map( A1 => n8577, A2 => n11374, ZN => n11415);
   U9480 : AND2_X1 port map( A1 => n8578, A2 => n11384, ZN => n11425);
   U9481 : NOR2_X1 port map( A1 => RST, A2 => n11888, ZN => n11890);
   U9482 : AND2_X1 port map( A1 => n8579, A2 => n11248, ZN => n11285);
   U9483 : AND2_X1 port map( A1 => n8579, A2 => n11253, ZN => n11291);
   U9484 : AND2_X1 port map( A1 => n8580, A2 => n11252, ZN => n11290);
   U9485 : INV_X1 port map( A => n10846, ZN => n10945);
   U9486 : INV_X1 port map( A => n11350, ZN => n11397);
   U9487 : INV_X1 port map( A => n11344, ZN => n11379);
   U9488 : AND2_X1 port map( A1 => n8579, A2 => n11230, ZN => n11305);
   U9489 : INV_X1 port map( A => n11205, ZN => n11259);
   U9490 : INV_X1 port map( A => n11207, ZN => n11262);
   U9491 : INV_X1 port map( A => n11224, ZN => n11261);
   U9492 : INV_X1 port map( A => n11349, ZN => n11393);
   U9493 : INV_X1 port map( A => n11346, ZN => n11389);
   U9494 : INV_X1 port map( A => n11351, ZN => n11405);
   U9495 : INV_X1 port map( A => n11345, ZN => n11383);
   U9496 : INV_X1 port map( A => n11348, ZN => n11391);
   U9497 : AND2_X1 port map( A1 => n8580, A2 => n11267, ZN => n11310);
   U9498 : OAI22_X1 port map( A1 => n575, A2 => n11517, B1 => n11518, B2 => 
                           n11281, ZN => n11217);
   U9499 : OAI22_X1 port map( A1 => n575, A2 => n11524, B1 => n11523, B2 => 
                           n11281, ZN => n11219);
   U9500 : OAI22_X1 port map( A1 => n575, A2 => n11892, B1 => n11891, B2 => 
                           n11281, ZN => n11196);
   U9501 : AND2_X1 port map( A1 => n8578, A2 => n11392, ZN => n11433);
   U9502 : AND2_X1 port map( A1 => n8578, A2 => n11395, ZN => n11436);
   U9503 : AND2_X1 port map( A1 => n8578, A2 => n11385, ZN => n11426);
   U9504 : AND2_X1 port map( A1 => n8578, A2 => n11394, ZN => n11435);
   U9505 : AND2_X1 port map( A1 => n8578, A2 => n11387, ZN => n11428);
   U9506 : AND2_X1 port map( A1 => n8578, A2 => n11386, ZN => n11427);
   U9507 : AND2_X1 port map( A1 => n8578, A2 => n11388, ZN => n11429);
   U9508 : AOI22_X1 port map( A1 => n7783, A2 => n11465, B1 => n11658, B2 => 
                           n11281, ZN => n11258);
   U9509 : INV_X1 port map( A => n11223, ZN => n11254);
   U9510 : OAI22_X1 port map( A1 => n8529, A2 => n11907, B1 => n11908, B2 => 
                           n8191, ZN => n11506);
   U9511 : AOI22_X1 port map( A1 => n10437, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_3_port, B1 => 
                           n11076, B2 => n11084, ZN => n11907);
   U9512 : AOI22_X1 port map( A1 => n8417, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_2_port, B1 => 
                           n11061, B2 => n11084, ZN => n11896);
   U9513 : INV_X1 port map( A => n11102, ZN => n11552);
   U9514 : INV_X1 port map( A => n11567, ZN => n11243);
   U9515 : AOI22_X1 port map( A1 => n8417, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_11_port, B1 => 
                           n11027, B2 => n11084, ZN => n11561);
   U9516 : NOR2_X1 port map( A1 => n11025, A2 => n11630, ZN => n11564);
   U9517 : INV_X1 port map( A => n11137, ZN => n11558);
   U9518 : INV_X1 port map( A => n11584, ZN => n11414);
   U9519 : OAI22_X1 port map( A1 => n7766, A2 => n11518, B1 => n11517, B2 => 
                           n8191, ZN => n11521);
   U9520 : INV_X1 port map( A => n10984, ZN => n11652);
   U9521 : NOR2_X1 port map( A1 => i_ADD_WB_4_port, A2 => n11010, ZN => n11044)
                           ;
   U9522 : NOR2_X1 port map( A1 => n8209, A2 => n11010, ZN => n11045);
   U9523 : INV_X1 port map( A => n10991, ZN => n11659);
   U9524 : NOR2_X1 port map( A1 => RST, A2 => n11062, ZN => n11160);
   U9525 : BUF_X2 port map( A => n11059, Z => n8486);
   U9526 : OAI22_X1 port map( A1 => n576, A2 => n11892, B1 => n11891, B2 => 
                           n8483, ZN => n11059);
   U9527 : BUF_X2 port map( A => n11098, Z => n8493);
   U9528 : OAI22_X1 port map( A1 => n576, A2 => n11524, B1 => n11523, B2 => 
                           n8483, ZN => n11098);
   U9529 : NAND2_X1 port map( A1 => n8573, A2 => n11679, ZN => n11847);
   U9530 : INV_X1 port map( A => n10989, ZN => n11657);
   U9531 : INV_X1 port map( A => n10972, ZN => n11666);
   U9532 : INV_X1 port map( A => n10981, ZN => n11648);
   U9533 : INV_X1 port map( A => n10985, ZN => n11653);
   U9534 : INV_X1 port map( A => n10982, ZN => n11649);
   U9535 : INV_X1 port map( A => n10990, ZN => n11658);
   U9536 : INV_X1 port map( A => n10973, ZN => n11667);
   U9537 : INV_X1 port map( A => n10983, ZN => n11651);
   U9538 : INV_X1 port map( A => n10980, ZN => n11647);
   U9539 : INV_X1 port map( A => n10988, ZN => n11656);
   U9540 : INV_X1 port map( A => n10979, ZN => n11646);
   U9541 : INV_X1 port map( A => n10970, ZN => n11663);
   U9542 : INV_X1 port map( A => n10971, ZN => n11665);
   U9543 : NOR2_X1 port map( A1 => RST, A2 => n11071, ZN => n11185);
   U9544 : INV_X1 port map( A => n10986, ZN => n11655);
   U9545 : INV_X1 port map( A => n10974, ZN => n11671);
   U9546 : INV_X1 port map( A => n10975, ZN => n11674);
   U9547 : NOR2_X1 port map( A1 => RST, A2 => n11068, ZN => n11180);
   U9548 : NOR2_X1 port map( A1 => RST, A2 => n11063, ZN => n11164);
   U9549 : NOR2_X1 port map( A1 => RST, A2 => n11070, ZN => n11183);
   U9550 : BUF_X1 port map( A => i_S3, Z => n8565);
   U9551 : OAI22_X1 port map( A1 => n11053, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_0_port, B1 => 
                           n8417, B2 => n11052, ZN => n11886);
   U9552 : INV_X1 port map( A => n10978, ZN => n11645);
   U9553 : NOR2_X1 port map( A1 => n556, A2 => n11726, ZN => n11727);
   U9554 : NOR2_X1 port map( A1 => n554, A2 => n11723, ZN => n11724);
   U9555 : NOR2_X1 port map( A1 => n552, A2 => n11720, ZN => n11721);
   U9556 : NOR2_X1 port map( A1 => n550, A2 => n11717, ZN => n11718);
   U9557 : NOR2_X1 port map( A1 => n548, A2 => n11714, ZN => n11715);
   U9558 : NOR2_X1 port map( A1 => n546, A2 => n11711, ZN => n11712);
   U9559 : OAI211_X1 port map( C1 => n172, C2 => n10405, A => n10404, B => 
                           n10192, ZN => i_ADD_WS1_4_port);
   U9560 : OAI211_X1 port map( C1 => n175, C2 => n10405, A => n10404, B => 
                           n10198, ZN => i_ADD_WS1_1_port);
   U9561 : NAND2_X1 port map( A1 => n7621, A2 => n10191, ZN => n10405);
   U9562 : INV_X1 port map( A => n10116, ZN => n10046);
   U9563 : INV_X1 port map( A => n10117, ZN => n10056);
   U9564 : BUF_X1 port map( A => n9202, Z => n8398);
   U9565 : BUF_X1 port map( A => n9100, Z => n8457);
   U9566 : NAND2_X1 port map( A1 => n10434, A2 => IRAM_READY, ZN => n8913);
   U9567 : NOR2_X1 port map( A1 => n10423, A2 => n173, ZN => i_ADD_RS2_3_port);
   U9568 : INV_X2 port map( A => n8419, ZN => n10401);
   U9569 : AND2_X1 port map( A1 => DataPath_RF_c_win_4_port, A2 => n8334, ZN =>
                           n8414);
   U9570 : OAI211_X1 port map( C1 => DataPath_RF_c_swin_2_port, C2 => n575, A 
                           => n8349, B => n8347, ZN => n10442);
   U9571 : OR2_X1 port map( A1 => DataPath_RF_c_win_3_port, A2 => n8242, ZN => 
                           n8376);
   U9572 : INV_X2 port map( A => n11847, ZN => n8543);
   U9573 : INV_X2 port map( A => n11847, ZN => n8544);
   U9574 : NOR2_X1 port map( A1 => RST, A2 => n11233, ZN => n11231);
   U9575 : NOR2_X1 port map( A1 => RST, A2 => n11247, ZN => n11245);
   U9576 : NOR2_X1 port map( A1 => RST, A2 => n11343, ZN => n11353);
   U9577 : AND2_X1 port map( A1 => n8579, A2 => n7813, ZN => n11289);
   U9578 : AND2_X1 port map( A1 => n8579, A2 => n7814, ZN => n11286);
   U9579 : AND2_X1 port map( A1 => n8577, A2 => n7811, ZN => n11244);
   U9580 : AND2_X1 port map( A1 => n8580, A2 => n7815, ZN => n11296);
   U9581 : INV_X1 port map( A => n11329, ZN => n11402);
   U9582 : OR2_X2 port map( A1 => RST, A2 => n11909, ZN => n8286);
   U9583 : INV_X1 port map( A => n10835, ZN => n10902);
   U9584 : INV_X1 port map( A => n11333, ZN => n11404);
   U9585 : INV_X1 port map( A => n11347, ZN => n11390);
   U9586 : INV_X1 port map( A => n11327, ZN => n11399);
   U9587 : OAI21_X1 port map( B1 => n11412, B2 => n11569, A => n8341, ZN => 
                           n11370);
   U9588 : OAI22_X1 port map( A1 => n575, A2 => n11512, B1 => n11513, B2 => 
                           n11281, ZN => n11212);
   U9589 : INV_X1 port map( A => n11191, ZN => n11250);
   U9590 : INV_X1 port map( A => n11208, ZN => n11265);
   U9591 : OAI22_X1 port map( A1 => n8333, A2 => n11897, B1 => n11412, B2 => 
                           n11896, ZN => n11330);
   U9592 : NOR2_X1 port map( A1 => RST, A2 => n11199, ZN => n11311);
   U9593 : NOR2_X1 port map( A1 => RST, A2 => n11509, ZN => n11511);
   U9594 : AND2_X1 port map( A1 => n8580, A2 => n7812, ZN => n11295);
   U9595 : INV_X1 port map( A => n11218, ZN => n11269);
   U9596 : NOR2_X1 port map( A1 => RST, A2 => n11195, ZN => n11316);
   U9597 : OAI22_X1 port map( A1 => n8219, A2 => n11924, B1 => n11923, B2 => 
                           n11922, ZN => n11944);
   U9598 : INV_X2 port map( A => n11033, ZN => n8409);
   U9599 : INV_X2 port map( A => n11020, ZN => n8407);
   U9600 : AOI22_X1 port map( A1 => n10437, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_9_port, B1 => 
                           n11018, B2 => n11084, ZN => n11549);
   U9601 : INV_X2 port map( A => n11029, ZN => n8408);
   U9602 : AOI22_X1 port map( A1 => n10437, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_10_port, B1 => 
                           n11022, B2 => n11084, ZN => n11555);
   U9603 : INV_X1 port map( A => n11501, ZN => n11500);
   U9604 : INV_X1 port map( A => n11498, ZN => n11497);
   U9605 : INV_X1 port map( A => n11494, ZN => n11678);
   U9606 : INV_X1 port map( A => n11474, ZN => n11664);
   U9607 : INV_X1 port map( A => n11488, ZN => n11673);
   U9608 : INV_X1 port map( A => n11486, ZN => n11672);
   U9609 : INV_X1 port map( A => n11471, ZN => n11662);
   U9610 : INV_X1 port map( A => n11492, ZN => n11675);
   U9611 : INV_X1 port map( A => n11516, ZN => n11515);
   U9612 : INV_X1 port map( A => n11469, ZN => n11661);
   U9613 : INV_X1 port map( A => n11455, ZN => n11650);
   U9614 : INV_X1 port map( A => n11467, ZN => n11660);
   U9615 : INV_X1 port map( A => n11460, ZN => n11654);
   U9616 : INV_X1 port map( A => n11483, ZN => n11670);
   U9617 : INV_X1 port map( A => n11481, ZN => n11669);
   U9618 : INV_X1 port map( A => n11479, ZN => n11668);
   U9619 : INV_X1 port map( A => n11373, ZN => n11575);
   U9620 : OAI22_X1 port map( A1 => n11084, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_13_port, B1 => 
                           n11035, B2 => n8417, ZN => n11373);
   U9621 : AOI22_X1 port map( A1 => n10437, A2 => n8211, B1 => n11039, B2 => 
                           n11084, ZN => n11581);
   U9622 : NAND2_X1 port map( A1 => i_ADD_WB_3_port, A2 => i_WF, ZN => n11010);
   U9623 : INV_X1 port map( A => n575, ZN => n8554);
   U9624 : AOI22_X1 port map( A1 => n10437, A2 => n8308, B1 => n11009, B2 => 
                           n11084, ZN => n11546);
   U9625 : NOR2_X1 port map( A1 => RST, A2 => n11065, ZN => n11171);
   U9626 : NOR2_X1 port map( A1 => RST, A2 => n11000, ZN => n11920);
   U9627 : NOR2_X1 port map( A1 => RST, A2 => n10999, ZN => n11918);
   U9628 : NOR2_X1 port map( A1 => RST, A2 => n10994, ZN => n11942);
   U9629 : NOR2_X1 port map( A1 => RST, A2 => n11066, ZN => n11172);
   U9630 : NOR2_X1 port map( A1 => RST, A2 => n11064, ZN => n11170);
   U9631 : NOR2_X1 port map( A1 => RST, A2 => n11067, ZN => n11179);
   U9632 : NOR2_X1 port map( A1 => n564, A2 => n11738, ZN => n11739);
   U9633 : NOR2_X1 port map( A1 => n562, A2 => n11735, ZN => n11736);
   U9634 : NOR2_X1 port map( A1 => n560, A2 => n11732, ZN => n11733);
   U9635 : NOR2_X1 port map( A1 => n558, A2 => n11729, ZN => n11730);
   U9636 : NOR2_X1 port map( A1 => n544, A2 => n11708, ZN => n11709);
   U9637 : INV_X1 port map( A => n10120, ZN => n10059);
   U9638 : INV_X1 port map( A => n10110, ZN => n9977);
   U9639 : INV_X1 port map( A => n10121, ZN => n10002);
   U9640 : INV_X1 port map( A => n10066, ZN => n10113);
   U9641 : INV_X1 port map( A => n10045, ZN => n10104);
   U9642 : INV_X1 port map( A => n10430, ZN => n10106);
   U9643 : NAND2_X1 port map( A1 => n8188, A2 => n11852, ZN => n11879);
   U9644 : AND2_X1 port map( A1 => n9041, A2 => n9146, ZN => n10110);
   U9645 : AND2_X1 port map( A1 => n9127, A2 => n9126, ZN => n10035);
   U9646 : AND2_X1 port map( A1 => DataPath_RF_POP_ADDRGEN_curr_state_1_port, 
                           A2 => n866, ZN => n8593);
   U9647 : OR2_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_state_0_port, 
                           A2 => n838, ZN => n8583);
   U9648 : NOR2_X1 port map( A1 => n466, A2 => n465, ZN => 
                           DP_OP_1091J1_126_6973_n72);
   U9649 : NOR2_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_addr_15_port, 
                           A2 => n11818, ZN => n11817);
   U9650 : OAI21_X1 port map( B1 => n11622, B2 => n11634, A => n8571, ZN => 
                           n11623);
   U9651 : OAI21_X1 port map( B1 => n11635, B2 => n11634, A => n8580, ZN => 
                           n11636);
   U9652 : OAI21_X1 port map( B1 => n11630, B2 => n11634, A => n8580, ZN => 
                           n11631);
   U9653 : INV_X1 port map( A => n11807, ZN => n11811);
   U9654 : INV_X2 port map( A => n11847, ZN => n8542);
   U9655 : NOR2_X1 port map( A1 => RST, A2 => n11228, ZN => n11225);
   U9656 : NOR2_X1 port map( A1 => RST, A2 => n11237, ZN => n11235);
   U9657 : BUF_X2 port map( A => n11353, Z => n8511);
   U9658 : OR2_X1 port map( A1 => n10941, A2 => n10919, ZN => n10893);
   U9659 : OAI22_X1 port map( A1 => n8333, A2 => n11908, B1 => n11412, B2 => 
                           n11907, ZN => n11334);
   U9660 : NOR2_X1 port map( A1 => RST, A2 => n11194, ZN => n11314);
   U9661 : AOI22_X1 port map( A1 => n7783, A2 => n11473, B1 => n11663, B2 => 
                           n11281, ZN => n11301);
   U9662 : NOR2_X1 port map( A1 => RST, A2 => n11326, ZN => n11439);
   U9663 : NOR2_X1 port map( A1 => RST, A2 => n11328, ZN => n11442);
   U9664 : NOR2_X1 port map( A1 => RST, A2 => n11192, ZN => n11308);
   U9665 : INV_X2 port map( A => n11582, ZN => n8528);
   U9666 : NOR2_X1 port map( A1 => RST, A2 => n11333, ZN => n11445);
   U9667 : NOR2_X1 port map( A1 => RST, A2 => n11329, ZN => n11443);
   U9668 : BUF_X2 port map( A => n11511, Z => n8521);
   U9669 : NOR2_X1 port map( A1 => RST, A2 => n11208, ZN => n11307);
   U9670 : AOI22_X1 port map( A1 => n7783, A2 => n11464, B1 => n11657, B2 => 
                           n11281, ZN => n11257);
   U9671 : NOR2_X1 port map( A1 => RST, A2 => n11206, ZN => n11299);
   U9672 : AOI22_X1 port map( A1 => n7783, A2 => n11457, B1 => n11651, B2 => 
                           n11281, ZN => n11251);
   U9673 : AOI22_X1 port map( A1 => n7783, A2 => n11453, B1 => n11648, B2 => 
                           n11281, ZN => n11249);
   U9674 : OAI22_X1 port map( A1 => n8219, A2 => n11892, B1 => n11923, B2 => 
                           n11891, ZN => n11893);
   U9675 : OAI22_X1 port map( A1 => n576, A2 => n11897, B1 => n11896, B2 => 
                           n8483, ZN => n11069);
   U9676 : NOR2_X1 port map( A1 => RST, A2 => n11014, ZN => n11974);
   U9677 : AOI211_X1 port map( C1 => n11243, C2 => n11814, A => RST, B => 
                           n11032, ZN => n11033);
   U9678 : AOI211_X1 port map( C1 => n11552, C2 => n11814, A => RST, B => 
                           n11019, ZN => n11020);
   U9679 : AOI211_X1 port map( C1 => n11564, C2 => n11814, A => RST, B => 
                           n11028, ZN => n11029);
   U9680 : INV_X1 port map( A => n11629, ZN => n11630);
   U9681 : NOR3_X1 port map( A1 => i_ADD_WB_0_port, A2 => n525, A3 => 
                           i_ADD_WB_1_port, ZN => n11629);
   U9682 : INV_X2 port map( A => n11139, ZN => n8410);
   U9683 : AOI211_X1 port map( C1 => n11558, C2 => n11814, A => RST, B => 
                           n11138, ZN => n11139);
   U9684 : INV_X2 port map( A => n11187, ZN => n8411);
   U9685 : AOI211_X1 port map( C1 => n11414, C2 => n11814, A => RST, B => 
                           n11154, ZN => n11187);
   U9686 : AOI22_X1 port map( A1 => n10437, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_15_port, B1 => 
                           n11047, B2 => n11084, ZN => n11585);
   U9687 : NOR2_X1 port map( A1 => RST, A2 => n10998, ZN => n11917);
   U9688 : NOR2_X1 port map( A1 => RST, A2 => n10992, ZN => n11910);
   U9689 : NOR2_X1 port map( A1 => RST, A2 => n11001, ZN => n11921);
   U9690 : NOR2_X1 port map( A1 => RST, A2 => n11013, ZN => n11967);
   U9691 : NOR2_X1 port map( A1 => RST, A2 => n10995, ZN => n11913);
   U9692 : NOR3_X1 port map( A1 => n525, A2 => n523, A3 => i_ADD_WB_1_port, ZN 
                           => n11625);
   U9693 : NOR3_X1 port map( A1 => i_ADD_WB_2_port, A2 => n8276, A3 => n523, ZN
                           => n11633);
   U9694 : INV_X1 port map( A => n11694, ZN => n11458);
   U9695 : NOR3_X1 port map( A1 => n523, A2 => i_ADD_WB_1_port, A3 => 
                           i_ADD_WB_2_port, ZN => n11643);
   U9696 : INV_X1 port map( A => n11700, ZN => n11466);
   U9697 : NOR3_X1 port map( A1 => i_ADD_WB_0_port, A2 => n8276, A3 => n525, ZN
                           => n11621);
   U9698 : NAND3_X1 port map( A1 => CU_I_CW_ID_ID_EN_port, A2 => n10440, A3 => 
                           n8582, ZN => n11846);
   U9699 : NOR2_X1 port map( A1 => RST, A2 => n10997, ZN => n11915);
   U9700 : NOR2_X1 port map( A1 => RST, A2 => n11012, ZN => n11963);
   U9701 : INV_X1 port map( A => n11698, ZN => n11464);
   U9702 : INV_X1 port map( A => n11702, ZN => n11477);
   U9703 : NOR2_X1 port map( A1 => RST, A2 => n10996, ZN => n11914);
   U9704 : NOR2_X1 port map( A1 => RST, A2 => n10993, ZN => n11940);
   U9705 : INV_X1 port map( A => n11691, ZN => n11453);
   U9706 : INV_X1 port map( A => n11695, ZN => n11459);
   U9707 : INV_X1 port map( A => n11692, ZN => n11454);
   U9708 : INV_X1 port map( A => n11699, ZN => n11465);
   U9709 : INV_X1 port map( A => n11703, ZN => n11478);
   U9710 : INV_X1 port map( A => n11693, ZN => n11457);
   U9711 : INV_X1 port map( A => n11690, ZN => n11452);
   U9712 : INV_X1 port map( A => n11697, ZN => n11463);
   U9713 : INV_X1 port map( A => n11689, ZN => n11451);
   U9714 : INV_X1 port map( A => n11701, ZN => n11473);
   U9715 : INV_X1 port map( A => n11476, ZN => n11319);
   U9716 : INV_X1 port map( A => n11696, ZN => n11462);
   U9717 : INV_X1 port map( A => n11704, ZN => n11485);
   U9718 : NOR3_X1 port map( A1 => i_ADD_WB_2_port, A2 => i_ADD_WB_0_port, A3 
                           => n8276, ZN => n11638);
   U9719 : INV_X1 port map( A => n11490, ZN => n11320);
   U9720 : INV_X1 port map( A => n11688, ZN => n11450);
   U9721 : NOR2_X1 port map( A1 => n461, A2 => n11679, ZN => DECODEhw_i_WR1);
   U9722 : NAND2_X1 port map( A1 => CU_I_CW_ID_ID_EN_port, A2 => n10440, ZN => 
                           n11679);
   U9723 : INV_X1 port map( A => n10434, ZN => n10413);
   U9724 : INV_X1 port map( A => n9897, ZN => n9748);
   U9725 : INV_X1 port map( A => n9704, ZN => n9755);
   U9726 : INV_X1 port map( A => n10038, ZN => n10112);
   U9727 : AND2_X1 port map( A1 => i_ALU_OP_0_port, A2 => i_ALU_OP_1_port, ZN 
                           => n9897);
   U9728 : INV_X1 port map( A => n10035, ZN => n10084);
   U9729 : INV_X1 port map( A => n11878, ZN => n9780);
   U9730 : OAI21_X1 port map( B1 => n8243, B2 => n8137, A => n9115, ZN => 
                           DP_OP_751_130_6421_n405);
   U9731 : BUF_X1 port map( A => n9202, Z => n8399);
   U9732 : INV_X1 port map( A => RST, ZN => n8571);
   U9733 : INV_X1 port map( A => RST, ZN => n8570);
   U9734 : OR2_X1 port map( A1 => RST, A2 => i_RF2, ZN => 
                           DataPath_RF_RDPORT1_OUTLATCH_N3);
   U9735 : OR2_X1 port map( A1 => RST, A2 => i_RF1, ZN => 
                           DataPath_RF_RDPORT0_OUTLATCH_N3);
   U9736 : OR3_X1 port map( A1 => n8592, A2 => n8901, A3 => n8590, ZN => n10231
                           );
   U9737 : INV_X1 port map( A => RST, ZN => n8575);
   U9738 : BUF_X1 port map( A => n10815, Z => n8463);
   U9739 : BUF_X1 port map( A => n10826, Z => n8472);
   U9740 : BUF_X1 port map( A => n10828, Z => n8476);
   U9741 : BUF_X1 port map( A => n10824, Z => n8470);
   U9742 : NOR2_X1 port map( A1 => n10499, A2 => n10498, ZN => n10824);
   U9743 : NOR2_X1 port map( A1 => n10503, A2 => n10501, ZN => n10828);
   U9744 : OR2_X1 port map( A1 => n10497, A2 => n10496, ZN => n10499);
   U9745 : BUF_X1 port map( A => n10817, Z => n8459);
   U9746 : NOR2_X1 port map( A1 => n10501, A2 => n10486, ZN => n10817);
   U9747 : NAND2_X1 port map( A1 => n10479, A2 => n10481, ZN => n10501);
   U9748 : BUF_X1 port map( A => n10813, Z => n8464);
   U9749 : NOR2_X1 port map( A1 => n10502, A2 => n10485, ZN => n10813);
   U9750 : OR2_X1 port map( A1 => n10495, A2 => n10494, ZN => n10485);
   U9751 : INV_X1 port map( A => n10448, ZN => n10449);
   U9752 : NAND3_X1 port map( A1 => n11638, A2 => n11642, A3 => n8581, ZN => 
                           n11641);
   U9753 : NAND3_X1 port map( A1 => n11617, A2 => n11642, A3 => n8570, ZN => 
                           n11620);
   U9754 : NAND3_X1 port map( A1 => n11643, A2 => n11642, A3 => n8579, ZN => 
                           n11677);
   U9755 : NAND3_X1 port map( A1 => n11625, A2 => n11642, A3 => n8576, ZN => 
                           n11628);
   U9756 : NAND3_X1 port map( A1 => n11621, A2 => n11642, A3 => n8575, ZN => 
                           n11624);
   U9757 : NAND3_X1 port map( A1 => n11633, A2 => n11642, A3 => n8576, ZN => 
                           n11637);
   U9758 : NAND3_X1 port map( A1 => n11629, A2 => n11642, A3 => n8571, ZN => 
                           n11632);
   U9759 : NAND2_X1 port map( A1 => n8572, A2 => n8458, ZN => n11791);
   U9760 : NOR2_X1 port map( A1 => DRAM_READY, A2 => n11976, ZN => n8458);
   U9761 : INV_X1 port map( A => RST, ZN => n8572);
   U9762 : NOR2_X1 port map( A1 => RST, A2 => n11280, ZN => n11278);
   U9763 : NOR2_X1 port map( A1 => RST, A2 => n11327, ZN => n11440);
   U9764 : NOR2_X1 port map( A1 => n10898, A2 => n10895, ZN => n10926);
   U9765 : NOR2_X1 port map( A1 => n8293, A2 => n10896, ZN => n10898);
   U9766 : NOR2_X1 port map( A1 => i_DATAMEM_RM, A2 => n10846, ZN => n10941);
   U9767 : INV_X1 port map( A => n10867, ZN => n10940);
   U9768 : INV_X1 port map( A => n11328, ZN => n11401);
   U9769 : NOR2_X1 port map( A1 => RST, A2 => n11218, ZN => n11312);
   U9770 : AND2_X2 port map( A1 => n8580, A2 => n11048, ZN => n11049);
   U9771 : INV_X1 port map( A => n11206, ZN => n11260);
   U9772 : INV_X1 port map( A => n11194, ZN => n11271);
   U9773 : NOR2_X1 port map( A1 => RST, A2 => n11191, ZN => n11288);
   U9774 : INV_X1 port map( A => RST, ZN => n8577);
   U9775 : INV_X1 port map( A => n11012, ZN => n11930);
   U9776 : INV_X1 port map( A => n11013, ZN => n11933);
   U9777 : INV_X1 port map( A => n10997, ZN => n11949);
   U9778 : INV_X1 port map( A => n10996, ZN => n11948);
   U9779 : INV_X1 port map( A => n11001, ZN => n11955);
   U9780 : INV_X1 port map( A => n10992, ZN => n11939);
   U9781 : INV_X1 port map( A => n10998, ZN => n11951);
   U9782 : INV_X1 port map( A => n10995, ZN => n11947);
   U9783 : INV_X1 port map( A => n11014, ZN => n11938);
   U9784 : INV_X1 port map( A => RST, ZN => n8578);
   U9785 : INV_X1 port map( A => RST, ZN => n8580);
   U9786 : INV_X1 port map( A => RST, ZN => n8579);
   U9787 : INV_X1 port map( A => RST, ZN => n8574);
   U9788 : INV_X1 port map( A => RST, ZN => n8573);
   U9789 : INV_X1 port map( A => RST, ZN => n8581);
   U9790 : INV_X1 port map( A => RST, ZN => n8576);
   U9791 : NOR3_X1 port map( A1 => n525, A2 => n523, A3 => n8276, ZN => n11617)
                           ;
   U9792 : INV_X1 port map( A => RST, ZN => n8582);
   U9793 : OR2_X1 port map( A1 => i_ALU_OP_1_port, A2 => i_ALU_OP_0_port, ZN =>
                           n11878);
   U9794 : BUF_X1 port map( A => n8435, Z => n8436);
   U9795 : AND2_X1 port map( A1 => n8557, A2 => DataPath_i_PIPLIN_A_31_port, ZN
                           => n10081);
   U9796 : INV_X1 port map( A => n10070, ZN => n9619);
   U9797 : AND2_X1 port map( A1 => n8557, A2 => DataPath_i_PIPLIN_A_30_port, ZN
                           => n10070);
   U9798 : INV_X1 port map( A => DP_OP_751_130_6421_n405, ZN => n9914);
   U9799 : INV_X1 port map( A => DP_OP_751_130_6421_n507, ZN => n9461);
   U9800 : INV_X1 port map( A => n9912, ZN => n9913);
   U9801 : AND2_X1 port map( A1 => n8557, A2 => DataPath_i_PIPLIN_A_29_port, ZN
                           => n9912);
   U9802 : INV_X1 port map( A => n9442, ZN => n9660);
   U9803 : AND2_X1 port map( A1 => n8557, A2 => DataPath_i_PIPLIN_A_28_port, ZN
                           => n9442);
   U9804 : AND2_X1 port map( A1 => n8557, A2 => DataPath_i_PIPLIN_A_26_port, ZN
                           => n9727);
   U9805 : INV_X1 port map( A => n9312, ZN => n8433);
   U9806 : XNOR2_X1 port map( A => n9651, B => DP_OP_751_130_6421_n915, ZN => 
                           n9100);
   U9807 : INV_X1 port map( A => n9936, ZN => n9934);
   U9808 : INV_X1 port map( A => DP_OP_751_130_6421_n915, ZN => n9693);
   U9809 : OAI21_X1 port map( B1 => n8252, B2 => n7929, A => n9090, ZN => 
                           DP_OP_751_130_6421_n915);
   U9810 : OAI21_X1 port map( B1 => n8249, B2 => n7929, A => n9082, ZN => 
                           DP_OP_751_130_6421_n1119);
   U9811 : BUF_X1 port map( A => n9074, Z => n8452);
   U9812 : BUF_X1 port map( A => n10054, Z => n8406);
   U9813 : AND2_X1 port map( A1 => n8557, A2 => DataPath_i_PIPLIN_A_17_port, ZN
                           => n10053);
   U9814 : INV_X1 port map( A => n460, ZN => n8558);
   U9815 : NOR2_X1 port map( A1 => n10420, A2 => n8232, ZN => i_ADD_RS1_0_port)
                           ;
   U9816 : NOR2_X1 port map( A1 => n10420, A2 => n8231, ZN => i_ADD_RS1_3_port)
                           ;
   U9817 : NOR2_X1 port map( A1 => n10420, A2 => n170, ZN => i_ADD_RS1_2_port);
   U9818 : NOR2_X1 port map( A1 => n10420, A2 => n171, ZN => i_ADD_RS1_1_port);
   U9819 : NOR2_X1 port map( A1 => n10420, A2 => n169, ZN => i_ADD_RS1_4_port);
   U9820 : INV_X1 port map( A => n10422, ZN => n10420);
   U9821 : AOI211_X4 port map( C1 => n7783, C2 => n11546, A => RST, B => n11222
                           , ZN => n11228);
   U9822 : AOI211_X4 port map( C1 => n7783, C2 => n11581, A => RST, B => n11275
                           , ZN => n11280);
   U9823 : OAI22_X1 port map( A1 => n575, A2 => n11887, B1 => n11281, B2 => 
                           n11886, ZN => n11188);
   U9824 : AOI211_X4 port map( C1 => DataPath_RF_c_win_1_port, C2 => n11564, A 
                           => RST, B => n11238, ZN => n11241);
   U9825 : OAI22_X1 port map( A1 => n8219, A2 => n11887, B1 => n11886, B2 => 
                           n11923, ZN => n11888);
   U9826 : AOI211_X4 port map( C1 => DataPath_RF_c_win_1_port, C2 => n11552, A 
                           => RST, B => n11229, ZN => n11233);
   U9827 : OAI21_X1 port map( B1 => n11412, B2 => n11373, A => n8344, ZN => 
                           n11398);
   U9828 : AOI211_X4 port map( C1 => n11558, C2 => n8554, A => RST, B => n11234
                           , ZN => n11237);
   U9829 : AOI211_X4 port map( C1 => DataPath_RF_c_win_1_port, C2 => n11243, A 
                           => RST, B => n11242, ZN => n11247);
   U9830 : AOI211_X4 port map( C1 => n7784, C2 => n11581, A => RST, B => n11408
                           , ZN => n11411);
   U9831 : AOI211_X4 port map( C1 => n7784, C2 => n11546, A => RST, B => n11357
                           , ZN => n11359);
   U9832 : AOI211_X4 port map( C1 => n7782, C2 => n11581, A => RST, B => n11040
                           , ZN => n11043);
   U9833 : AOI211_X4 port map( C1 => n7782, C2 => n11546, A => RST, B => n11011
                           , ZN => n11016);
   U9834 : AOI211_X4 port map( C1 => n7782, C2 => n11575, A => RST, B => n11036
                           , ZN => n11038);
   U9835 : NOR2_X2 port map( A1 => n10872, A2 => n10893, ZN => n10929);
   U9836 : OAI22_X1 port map( A1 => n8333, A2 => n11524, B1 => n11412, B2 => 
                           n11523, ZN => n11354);
   U9837 : OAI22_X1 port map( A1 => n576, A2 => n11908, B1 => n11907, B2 => 
                           n11153, ZN => n11081);
   U9838 : AOI211_X4 port map( C1 => n11414, C2 => n8554, A => RST, B => n11282
                           , ZN => n11317);
   U9839 : AOI211_X4 port map( C1 => DataPath_RF_c_win_0_port, C2 => n11552, A 
                           => RST, B => n11360, ZN => n11362);
   U9840 : AOI211_X4 port map( C1 => DataPath_RF_c_win_0_port, C2 => n11564, A 
                           => RST, B => n11366, ZN => n11368);
   U9841 : AOI211_X4 port map( C1 => n8296, C2 => n11546, A => RST, B => n11545
                           , ZN => n11548);
   U9842 : AOI211_X4 port map( C1 => n8296, C2 => n11575, A => RST, B => n11574
                           , ZN => n11577);
   U9843 : AOI211_X4 port map( C1 => DataPath_RF_c_win_1_port, C2 => n11558, A 
                           => RST, B => n11363, ZN => n11365);
   U9844 : AOI211_X4 port map( C1 => DataPath_RF_c_win_1_port, C2 => n11414, A 
                           => RST, B => n11413, ZN => n11448);
   U9845 : AOI211_X4 port map( C1 => DataPath_RF_c_win_4_port, C2 => n11564, A 
                           => RST, B => n11563, ZN => n11566);
   U9846 : AOI211_X4 port map( C1 => n8564, C2 => n11552, A => RST, B => n11551
                           , ZN => n11554);
   U9847 : AOI211_X4 port map( C1 => DataPath_RF_c_win_0_port, C2 => n11558, A 
                           => RST, B => n11557, ZN => n11560);
   U9848 : AOI211_X4 port map( C1 => n11243, C2 => n8554, A => RST, B => n11143
                           , ZN => n11145);
   U9849 : AOI211_X4 port map( C1 => n11564, C2 => n8554, A => RST, B => n11140
                           , ZN => n11142);
   U9850 : OAI222_X4 port map( A1 => n11137, A2 => n8219, B1 => n11556, B2 => 
                           n576, C1 => n11555, C2 => n11923, ZN => n11024);
   U9851 : OAI22_X2 port map( A1 => n11678, A2 => n11496, B1 => n3204, B2 => 
                           n7766, ZN => n11751);
   U9852 : OAI22_X2 port map( A1 => n11665, A2 => n11496, B1 => n3217, B2 => 
                           n7766, ZN => n11606);
   U9853 : OAI22_X2 port map( A1 => n11664, A2 => n11496, B1 => n3218, B2 => 
                           n7766, ZN => n11605);
   U9854 : OAI22_X2 port map( A1 => n11673, A2 => n11496, B1 => n3209, B2 => 
                           n7766, ZN => n11614);
   U9855 : OAI22_X2 port map( A1 => n11672, A2 => n11496, B1 => n3210, B2 => 
                           n7766, ZN => n11613);
   U9856 : OAI22_X2 port map( A1 => n11662, A2 => n11496, B1 => n3220, B2 => 
                           n7766, ZN => n11603);
   U9857 : OAI22_X2 port map( A1 => n11675, A2 => n11496, B1 => n3207, B2 => 
                           n7766, ZN => n11616);
   U9858 : OAI22_X2 port map( A1 => n11661, A2 => n11496, B1 => n3221, B2 => 
                           n7766, ZN => n11602);
   U9859 : AOI22_X2 port map( A1 => n11650, A2 => n7766, B1 => n11496, B2 => 
                           n3232, ZN => n11591);
   U9860 : AOI22_X2 port map( A1 => n11660, A2 => n7766, B1 => n11496, B2 => 
                           n3222, ZN => n11601);
   U9861 : AOI22_X2 port map( A1 => n11654, A2 => n7766, B1 => n11496, B2 => 
                           n3228, ZN => n11595);
   U9862 : AOI22_X2 port map( A1 => n11674, A2 => n7766, B1 => n11496, B2 => 
                           n3208, ZN => n11615);
   U9863 : AOI22_X2 port map( A1 => n11670, A2 => n7766, B1 => n11496, B2 => 
                           n3212, ZN => n11611);
   U9864 : AOI22_X2 port map( A1 => n11669, A2 => n7766, B1 => n11496, B2 => 
                           n3213, ZN => n11610);
   U9865 : AOI22_X2 port map( A1 => n11668, A2 => n7766, B1 => n11496, B2 => 
                           n3214, ZN => n11609);
   U9866 : AOI211_X4 port map( C1 => n11150, C2 => n11575, A => RST, B => 
                           n11146, ZN => n11148);
   U9867 : AOI211_X4 port map( C1 => n11150, C2 => n11581, A => RST, B => 
                           n11149, ZN => n11152);
   U9868 : AOI211_X4 port map( C1 => n11150, C2 => n11546, A => RST, B => 
                           n11099, ZN => n11101);
   U9869 : NOR3_X1 port map( A1 => i_ADD_WB_1_port, A2 => i_ADD_WB_0_port, A3 
                           => i_ADD_WB_2_port, ZN => n11046);
   U9870 : OAI21_X1 port map( B1 => DataPath_RF_POP_ADDRGEN_curr_state_1_port, 
                           B2 => n866, A => n10946, ZN => n11051);
   U9871 : NAND2_X1 port map( A1 => DataPath_RF_POP_ADDRGEN_curr_state_1_port, 
                           A2 => n866, ZN => n10946);
   U9872 : NOR2_X2 port map( A1 => n9058, A2 => n9169, ZN => n10120);
   U9873 : NOR2_X2 port map( A1 => n9146, A2 => n7756, ZN => n10121);
   U9874 : NOR2_X2 port map( A1 => n9052, A2 => n8432, ZN => n10116);
   U9875 : NOR2_X2 port map( A1 => n9025, A2 => n9024, ZN => n10045);
   U9876 : NOR2_X2 port map( A1 => n9058, A2 => n9053, ZN => n10430);
   U9877 : OAI21_X2 port map( B1 => n8288, B2 => n7929, A => n9111, ZN => 
                           DP_OP_751_130_6421_n507);
   U9878 : INV_X1 port map( A => n460, ZN => n8559);
   U9879 : OR2_X2 port map( A1 => n10237, A2 => n10238, ZN => n10263);
   U9880 : OR2_X1 port map( A1 => n825, A2 => DataPath_RF_c_win_0_port, ZN => 
                           n8239);
   U9881 : NOR2_X2 port map( A1 => n11846, A2 => n10187, ZN => n10190);
   U9882 : OAI21_X1 port map( B1 => n7752, B2 => n10434, A => n11767, ZN => 
                           n7122);
   U9883 : INV_X1 port map( A => i_NPC_SEL, ZN => n11834);
   U9884 : NOR2_X1 port map( A1 => n10392, A2 => n8890, ZN => n10374);
   U9885 : NAND2_X1 port map( A1 => n10397, A2 => n10396, ZN => 
                           CU_I_CW_RF_RD1_EN_port);
   U9886 : OAI21_X1 port map( B1 => n10393, B2 => n10392, A => n10391, ZN => 
                           n10394);
   U9887 : NOR2_X1 port map( A1 => n10228, A2 => n10225, ZN => 
                           CU_I_CW_DATA_SIZE_0_port);
   U9888 : NOR2_X1 port map( A1 => n10228, A2 => n10227, ZN => 
                           CU_I_CW_DATA_SIZE_1_port);
   U9889 : NOR2_X1 port map( A1 => n10230, A2 => n10224, ZN => n10228);
   U9890 : INV_X1 port map( A => n10223, ZN => n10224);
   U9891 : NOR2_X1 port map( A1 => n10397, A2 => n10223, ZN => 
                           CU_I_CW_WB_MUX_SEL_port);
   U9892 : INV_X1 port map( A => n10222, ZN => n10397);
   U9893 : OAI22_X1 port map( A1 => n8592, A2 => n8591, B1 => n10395, B2 => 
                           n10231, ZN => n6692);
   U9894 : INV_X1 port map( A => n8901, ZN => n8588);
   U9895 : NAND2_X1 port map( A1 => n10234, A2 => n10233, ZN => 
                           CU_I_CW_MUXB_SEL_port);
   U9896 : INV_X1 port map( A => n10231, ZN => n10234);
   U9897 : OAI211_X1 port map( C1 => n8596, C2 => n10400, A => n8589, B => 
                           n10150, ZN => n8590);
   U9898 : INV_X1 port map( A => n8587, ZN => n8589);
   U9899 : OAI211_X1 port map( C1 => n10382, C2 => n10383, A => n10381, B => 
                           n10380, ZN => CU_I_CW_UNSIGNED_ID_port);
   U9900 : AOI21_X1 port map( B1 => n10379, B2 => n8195, A => n10378, ZN => 
                           n10380);
   U9901 : INV_X1 port map( A => n10377, ZN => n10379);
   U9902 : OR2_X1 port map( A1 => n10223, A2 => n10149, ZN => n10377);
   U9903 : NAND2_X1 port map( A1 => n8601, A2 => n8396, ZN => n10223);
   U9904 : AOI22_X1 port map( A1 => n7903, A2 => n10375, B1 => n10374, B2 => 
                           n10400, ZN => n10381);
   U9905 : OAI22_X1 port map( A1 => n8396, A2 => n7926, B1 => n8223, B2 => 
                           n10372, ZN => CU_I_CW_NPC_SEL_port);
   U9906 : NAND2_X1 port map( A1 => n10391, A2 => n10388, ZN => n10390);
   U9907 : OAI211_X1 port map( C1 => n8223, C2 => n8195, A => n8051, B => 
                           n10386, ZN => n10388);
   U9908 : INV_X1 port map( A => n10385, ZN => n10391);
   U9909 : NOR2_X1 port map( A1 => n8383, A2 => n7778, ZN => 
                           DRAMRF_ADDRESS_31_port);
   U9910 : INV_X1 port map( A => n7724, ZN => n10445);
   U9911 : OAI21_X1 port map( B1 => n8909, B2 => n8908, A => n10439, ZN => 
                           n11787);
   U9912 : OAI211_X1 port map( C1 => n8907, C2 => n10392, A => n8906, B => 
                           n8905, ZN => n8908);
   U9913 : INV_X1 port map( A => n10378, ZN => n8906);
   U9914 : INV_X1 port map( A => n8902, ZN => n8909);
   U9915 : OAI222_X1 port map( A1 => n11784, A2 => n10163, B1 => n11791, B2 => 
                           n219, C1 => n8223, C2 => n11783, ZN => n7088);
   U9916 : NAND2_X1 port map( A1 => n10439, A2 => n8901, ZN => n11783);
   U9917 : NAND2_X1 port map( A1 => n8904, A2 => n8905, ZN => n8901);
   U9918 : OR2_X1 port map( A1 => n8903, A2 => n10149, ZN => n8905);
   U9919 : NAND2_X1 port map( A1 => n8896, A2 => n8354, ZN => n8904);
   U9920 : OR2_X1 port map( A1 => n11781, A2 => n8900, ZN => n11784);
   U9921 : OAI22_X1 port map( A1 => n10210, A2 => n11846, B1 => n486, B2 => 
                           n11847, ZN => n7026);
   U9922 : INV_X1 port map( A => n10209, ZN => n10210);
   U9923 : OAI22_X1 port map( A1 => n10216, A2 => n11846, B1 => n11847, B2 => 
                           n8316, ZN => n7023);
   U9924 : INV_X1 port map( A => n10215, ZN => n10216);
   U9925 : OAI22_X1 port map( A1 => n10212, A2 => n11846, B1 => n11847, B2 => 
                           n8315, ZN => n7025);
   U9926 : INV_X1 port map( A => n10211, ZN => n10212);
   U9927 : OAI22_X1 port map( A1 => n10214, A2 => n11846, B1 => n11847, B2 => 
                           n8326, ZN => n7024);
   U9928 : INV_X1 port map( A => n10213, ZN => n10214);
   U9929 : INV_X1 port map( A => n8899, ZN => n8910);
   U9930 : INV_X1 port map( A => n8898, ZN => n11779);
   U9931 : OAI22_X1 port map( A1 => n11790, A2 => n8897, B1 => n8332, B2 => 
                           n11791, ZN => n8898);
   U9932 : OAI21_X1 port map( B1 => n10375, B2 => n8354, A => n8896, ZN => 
                           n8897);
   U9933 : INV_X1 port map( A => n8907, ZN => n8896);
   U9934 : NOR2_X1 port map( A1 => n10392, A2 => n8223, ZN => n10375);
   U9935 : AND2_X1 port map( A1 => n8899, A2 => n8895, ZN => n11781);
   U9936 : NAND2_X1 port map( A1 => n10156, A2 => IR_3_port, ZN => n8899);
   U9937 : AOI22_X1 port map( A1 => n10184, A2 => n11848, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_5_port, ZN => n2380);
   U9938 : AOI22_X1 port map( A1 => n10179, A2 => n11848, B1 => n8544, B2 => 
                           DataPath_i_PIPLIN_IN2_15_port, ZN => n2365);
   U9939 : AOI22_X1 port map( A1 => n10190, A2 => n8282, B1 => 
                           DataPath_i_PIPLIN_IN1_14_port, B2 => n8542, ZN => 
                           n2842);
   U9940 : AOI22_X1 port map( A1 => n10190, A2 => IR_1_port, B1 => 
                           DataPath_i_PIPLIN_IN1_1_port, B2 => n8542, ZN => 
                           n2858);
   U9941 : AOI22_X1 port map( A1 => n10190, A2 => n8280, B1 => 
                           DataPath_i_PIPLIN_IN1_11_port, B2 => n8542, ZN => 
                           n2845);
   U9942 : AOI22_X1 port map( A1 => n10190, A2 => IR_13_port, B1 => 
                           DataPath_i_PIPLIN_IN1_13_port, B2 => n8542, ZN => 
                           n2843);
   U9943 : AOI22_X1 port map( A1 => n10190, A2 => IR_3_port, B1 => 
                           DataPath_i_PIPLIN_IN1_3_port, B2 => n8542, ZN => 
                           n2853);
   U9944 : AOI22_X1 port map( A1 => n10190, A2 => IR_7_port, B1 => 
                           DataPath_i_PIPLIN_IN1_7_port, B2 => n8542, ZN => 
                           n2849);
   U9945 : AOI22_X1 port map( A1 => n10190, A2 => IR_10_port, B1 => 
                           DataPath_i_PIPLIN_IN1_10_port, B2 => n8542, ZN => 
                           n2846);
   U9946 : AOI22_X1 port map( A1 => n10190, A2 => IR_9_port, B1 => 
                           DataPath_i_PIPLIN_IN1_9_port, B2 => n8542, ZN => 
                           n2847);
   U9947 : AOI22_X1 port map( A1 => n10190, A2 => IR_5_port, B1 => 
                           DataPath_i_PIPLIN_IN1_5_port, B2 => n8542, ZN => 
                           n2851);
   U9948 : AOI22_X1 port map( A1 => n10190, A2 => n8196, B1 => 
                           DataPath_i_PIPLIN_IN1_12_port, B2 => n8542, ZN => 
                           n2844);
   U9949 : AOI22_X1 port map( A1 => n10190, A2 => IR_4_port, B1 => 
                           DataPath_i_PIPLIN_IN1_4_port, B2 => n8542, ZN => 
                           n2852);
   U9950 : AOI22_X1 port map( A1 => n10190, A2 => n8309, B1 => 
                           DataPath_i_PIPLIN_IN1_0_port, B2 => n8542, ZN => 
                           n2859);
   U9951 : AOI22_X1 port map( A1 => n10190, A2 => IR_8_port, B1 => 
                           DataPath_i_PIPLIN_IN1_8_port, B2 => n8542, ZN => 
                           n2848);
   U9952 : AOI22_X1 port map( A1 => n10190, A2 => IR_6_port, B1 => 
                           DataPath_i_PIPLIN_IN1_6_port, B2 => n8544, ZN => 
                           n2850);
   U9953 : OAI211_X1 port map( C1 => n10399, C2 => n10225, A => n10141, B => 
                           n10140, ZN => n7092);
   U9954 : AOI22_X1 port map( A1 => n10139, A2 => n10393, B1 => n11981, B2 => 
                           i_ALU_OP_3_port, ZN => n10140);
   U9955 : NAND2_X1 port map( A1 => n10138, A2 => n10137, ZN => n10141);
   U9956 : OAI21_X1 port map( B1 => n10142, B2 => IR_1_port, A => n10136, ZN =>
                           n10137);
   U9957 : INV_X1 port map( A => n10163, ZN => n10138);
   U9958 : AOI22_X1 port map( A1 => n10190, A2 => n8210, B1 => n8543, B2 => 
                           DataPath_i_PIPLIN_IN1_15_port, ZN => n2840);
   U9959 : AOI222_X1 port map( A1 => n11814, A2 => n11813, B1 => 
                           DataPath_RF_c_win_4_port, B2 => n11812, C1 => 
                           DataPath_RF_c_win_0_port, C2 => n11811, ZN => n11815
                           );
   U9960 : INV_X1 port map( A => n8594, ZN => n11802);
   U9961 : AOI21_X1 port map( B1 => n11801, B2 => n8358, A => n11996, ZN => 
                           n11805);
   U9962 : OAI211_X1 port map( C1 => n10399, C2 => n10232, A => n10148, B => 
                           n10147, ZN => n7091);
   U9963 : AOI22_X1 port map( A1 => n10146, A2 => n10145, B1 => i_ALU_OP_4_port
                           , B2 => n11981, ZN => n10147);
   U9964 : INV_X1 port map( A => n10155, ZN => n10145);
   U9965 : INV_X1 port map( A => n10142, ZN => n10143);
   U9966 : INV_X1 port map( A => n10229, ZN => n10232);
   U9967 : OAI211_X1 port map( C1 => n10135, C2 => n10142, A => n10398, B => 
                           n10134, ZN => n7094);
   U9968 : AOI21_X1 port map( B1 => i_ALU_OP_1_port, B2 => n11981, A => n10133,
                           ZN => n10134);
   U9969 : INV_X1 port map( A => n10399, ZN => n10133);
   U9970 : NAND2_X1 port map( A1 => n10156, A2 => n10129, ZN => n10142);
   U9971 : AOI21_X1 port map( B1 => n10146, B2 => n10160, A => n10144, ZN => 
                           n10135);
   U9972 : INV_X1 port map( A => n11782, ZN => n10144);
   U9973 : OAI211_X1 port map( C1 => n10400, C2 => n10399, A => n10398, B => 
                           n11777, ZN => n7095);
   U9974 : AOI211_X1 port map( C1 => n10139, C2 => n10225, A => n10132, B => 
                           n10161, ZN => n10398);
   U9975 : AOI21_X1 port map( B1 => n10155, B2 => n10136, A => n10130, ZN => 
                           n10132);
   U9976 : INV_X1 port map( A => n10146, ZN => n10130);
   U9977 : INV_X1 port map( A => n10131, ZN => n10129);
   U9978 : NOR2_X1 port map( A1 => n11790, A2 => n10383, ZN => n10139);
   U9979 : NAND2_X1 port map( A1 => n8051, A2 => n7962, ZN => n10383);
   U9980 : NAND2_X1 port map( A1 => n10439, A2 => n10374, ZN => n10399);
   U9981 : INV_X1 port map( A => n10162, ZN => n7093);
   U9982 : AOI211_X1 port map( C1 => n10161, C2 => n10160, A => n10159, B => 
                           n10158, ZN => n10162);
   U9983 : NOR3_X1 port map( A1 => n11780, A2 => IR_3_port, A3 => n10157, ZN =>
                           n10158);
   U9984 : INV_X1 port map( A => n10156, ZN => n10157);
   U9985 : AND2_X1 port map( A1 => n8894, A2 => n8190, ZN => n10156);
   U9986 : OAI21_X1 port map( B1 => n10163, B2 => n10155, A => n10154, ZN => 
                           n10159);
   U9987 : AOI22_X1 port map( A1 => n10439, A2 => n10153, B1 => n11981, B2 => 
                           i_ALU_OP_2_port, ZN => n10154);
   U9988 : OAI22_X1 port map( A1 => n10152, A2 => n10392, B1 => n10151, B2 => 
                           n10150, ZN => n10153);
   U9989 : INV_X1 port map( A => n8051, ZN => n10151);
   U9990 : AOI22_X1 port map( A1 => n10393, A2 => n8396, B1 => n7903, B2 => 
                           n10149, ZN => n10152);
   U9991 : NAND2_X1 port map( A1 => n10146, A2 => n8309, ZN => n10163);
   U9992 : NOR3_X1 port map( A1 => n11782, A2 => n11775, A3 => n10131, ZN => 
                           n10161);
   U9993 : NAND2_X1 port map( A1 => n8226, A2 => IR_2_port, ZN => n10131);
   U9994 : NAND4_X1 port map( A1 => n8190, A2 => n8228, A3 => n8198, A4 => 
                           n11754, ZN => n11775);
   U9995 : NAND2_X1 port map( A1 => n10146, A2 => n193, ZN => n11782);
   U9996 : NOR2_X1 port map( A1 => n11790, A2 => n10194, ZN => n10146);
   U9997 : AOI22_X1 port map( A1 => n10177, A2 => n7758, B1 => n8544, B2 => 
                           DataPath_i_PIPLIN_IN2_17_port, ZN => n2361);
   U9998 : AOI22_X1 port map( A1 => n10180, A2 => n7758, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_11_port, ZN => n2370);
   U9999 : AOI22_X1 port map( A1 => n10176, A2 => n7758, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_18_port, ZN => n2359);
   U10000 : AOI22_X1 port map( A1 => n10178, A2 => n7758, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_16_port, ZN => n2363);
   U10001 : AOI22_X1 port map( A1 => i_ADD_WS1_0_port, A2 => n7758, B1 => n8543
                           , B2 => DataPath_i_PIPLIN_WRB1_0_port, ZN => n2865);
   U10002 : AOI22_X1 port map( A1 => i_ADD_WS1_2_port, A2 => n7758, B1 => n8543
                           , B2 => DataPath_i_PIPLIN_WRB1_2_port, ZN => n2863);
   U10003 : AOI22_X1 port map( A1 => i_ADD_WS1_1_port, A2 => n7758, B1 => n8543
                           , B2 => DataPath_i_PIPLIN_WRB1_1_port, ZN => n2864);
   U10004 : AOI22_X1 port map( A1 => n10181, A2 => n7758, B1 => n8543, B2 => 
                           DataPath_i_PIPLIN_IN2_9_port, ZN => n2373);
   U10005 : AOI22_X1 port map( A1 => i_ADD_WS1_4_port, A2 => n7758, B1 => n8543
                           , B2 => DataPath_i_PIPLIN_WRB1_4_port, ZN => n2861);
   U10006 : AOI22_X1 port map( A1 => i_ADD_WS1_3_port, A2 => n7758, B1 => n8543
                           , B2 => DataPath_i_PIPLIN_WRB1_3_port, ZN => n2862);
   U10007 : INV_X1 port map( A => n10204, ZN => n7029);
   U10008 : AOI222_X1 port map( A1 => n10190, A2 => IR_2_port, B1 => n10189, B2
                           => n7758, C1 => DataPath_i_PIPLIN_IN1_2_port, C2 => 
                           n8542, ZN => n2854);
   U10009 : INV_X1 port map( A => n10188, ZN => n10189);
   U10010 : AOI22_X1 port map( A1 => n10172, A2 => n7758, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_23_port, ZN => n2348);
   U10011 : AOI22_X1 port map( A1 => n10168, A2 => n7758, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_27_port, ZN => n2340);
   U10012 : AOI22_X1 port map( A1 => n10174, A2 => n7758, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_21_port, ZN => n2352);
   U10013 : AOI22_X1 port map( A1 => n10170, A2 => n7758, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_25_port, ZN => n2344);
   U10014 : AOI22_X1 port map( A1 => n10164, A2 => n7758, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_31_port, ZN => n2332);
   U10015 : AOI22_X1 port map( A1 => n10165, A2 => n7758, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_30_port, ZN => n2334);
   U10016 : AOI22_X1 port map( A1 => n10173, A2 => n7758, B1 => n8543, B2 => 
                           DataPath_i_PIPLIN_IN2_22_port, ZN => n2350);
   U10017 : AOI22_X1 port map( A1 => n10169, A2 => n7758, B1 => n8543, B2 => 
                           DataPath_i_PIPLIN_IN2_26_port, ZN => n2342);
   U10018 : AOI22_X1 port map( A1 => n10183, A2 => n7758, B1 => n8543, B2 => 
                           DataPath_i_PIPLIN_IN2_7_port, ZN => n2377);
   U10019 : AOI22_X1 port map( A1 => n10175, A2 => n7758, B1 => n8543, B2 => 
                           DataPath_i_PIPLIN_IN2_19_port, ZN => n2357);
   U10020 : AOI22_X1 port map( A1 => n10166, A2 => n7758, B1 => n8543, B2 => 
                           DataPath_i_PIPLIN_IN2_29_port, ZN => n2336);
   U10021 : AOI22_X1 port map( A1 => n10167, A2 => n7758, B1 => n8543, B2 => 
                           DataPath_i_PIPLIN_IN2_28_port, ZN => n2338);
   U10022 : AOI22_X1 port map( A1 => n10171, A2 => n7758, B1 => n8543, B2 => 
                           DataPath_i_PIPLIN_IN2_24_port, ZN => n2346);
   U10023 : AOI22_X1 port map( A1 => n10182, A2 => n7758, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_8_port, ZN => n2375);
   U10024 : INV_X1 port map( A => n10206, ZN => n7028);
   U10025 : AOI22_X1 port map( A1 => n10205, A2 => n7758, B1 => n8544, B2 => 
                           DataPath_i_PIPLIN_IN2_3_port, ZN => n10206);
   U10026 : INV_X1 port map( A => n10218, ZN => n7022);
   U10027 : AOI22_X1 port map( A1 => n10217, A2 => n7758, B1 => n8544, B2 => 
                           DataPath_i_PIPLIN_IN2_14_port, ZN => n10218);
   U10028 : INV_X1 port map( A => n10220, ZN => n7021);
   U10029 : AOI22_X1 port map( A1 => n10219, A2 => n7758, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_20_port, ZN => n10220);
   U10030 : INV_X1 port map( A => n10208, ZN => n7027);
   U10031 : AOI22_X1 port map( A1 => n10207, A2 => n7758, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_4_port, ZN => n10208);
   U10032 : AND2_X1 port map( A1 => C620_DATA2_4, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_4_port);
   U10033 : AND2_X1 port map( A1 => C620_DATA2_5, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_5_port);
   U10034 : AND2_X1 port map( A1 => C620_DATA2_6, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_6_port);
   U10035 : NOR2_X1 port map( A1 => n8346, A2 => n8345, ZN => n8344);
   U10036 : NOR2_X1 port map( A1 => n11572, A2 => n8191, ZN => n8345);
   U10037 : NOR2_X1 port map( A1 => n11573, A2 => n8333, ZN => n8346);
   U10038 : AND2_X1 port map( A1 => C620_DATA2_7, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_7_port);
   U10039 : OAI22_X1 port map( A1 => n11578, A2 => n8191, B1 => n11579, B2 => 
                           n8333, ZN => n11408);
   U10040 : OAI22_X1 port map( A1 => n11543, A2 => n8191, B1 => n11544, B2 => 
                           n8333, ZN => n11357);
   U10041 : NOR2_X1 port map( A1 => n8343, A2 => n8342, ZN => n8341);
   U10042 : NOR2_X1 port map( A1 => n11568, A2 => n8333, ZN => n8342);
   U10043 : NOR2_X1 port map( A1 => n11567, A2 => n8191, ZN => n8343);
   U10044 : OAI22_X1 port map( A1 => n11544, A2 => n8191, B1 => n11543, B2 => 
                           n8219, ZN => n11545);
   U10045 : OAI22_X1 port map( A1 => n11572, A2 => n8219, B1 => n11573, B2 => 
                           n8191, ZN => n11574);
   U10046 : OAI22_X1 port map( A1 => n11578, A2 => n8219, B1 => n11579, B2 => 
                           n8191, ZN => n11580);
   U10047 : OAI21_X1 port map( B1 => n11412, B2 => n11555, A => n8294, ZN => 
                           n11363);
   U10048 : AND2_X1 port map( A1 => C620_DATA2_8, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_8_port);
   U10049 : OAI21_X1 port map( B1 => n11412, B2 => n11585, A => n8295, ZN => 
                           n11413);
   U10050 : OAI22_X1 port map( A1 => n8529, A2 => n11922, B1 => n11924, B2 => 
                           n8191, ZN => n11509);
   U10051 : OAI21_X1 port map( B1 => n7766, B2 => n11585, A => n8335, ZN => 
                           n11750);
   U10052 : NOR2_X1 port map( A1 => n8337, A2 => n8336, ZN => n8335);
   U10053 : NOR2_X1 port map( A1 => n11584, A2 => n8191, ZN => n8336);
   U10054 : NOR2_X1 port map( A1 => n11583, A2 => n8219, ZN => n8337);
   U10055 : OAI22_X1 port map( A1 => n8529, A2 => n11561, B1 => n11562, B2 => 
                           n8191, ZN => n11563);
   U10056 : OAI22_X1 port map( A1 => n8529, A2 => n11549, B1 => n11550, B2 => 
                           n8191, ZN => n11551);
   U10057 : NOR2_X1 port map( A1 => n8340, A2 => n8339, ZN => n8338);
   U10058 : NOR2_X1 port map( A1 => n11568, A2 => n8191, ZN => n8339);
   U10059 : NOR2_X1 port map( A1 => n11567, A2 => n8219, ZN => n8340);
   U10060 : OAI21_X1 port map( B1 => n11847, B2 => n492, A => n10201, ZN => 
                           n7117);
   U10061 : OAI22_X1 port map( A1 => n10202, A2 => n10201, B1 => n493, B2 => 
                           n11847, ZN => n7116);
   U10062 : INV_X1 port map( A => n10200, ZN => n10202);
   U10063 : OAI211_X1 port map( C1 => n9175, C2 => n9748, A => n9174, B => 
                           n9173, ZN => n11855);
   U10064 : AOI211_X1 port map( C1 => n9172, C2 => n10088, A => n9171, B => 
                           n9170, ZN => n9173);
   U10065 : NOR3_X1 port map( A1 => n10084, A2 => n9169, A3 => n9168, ZN => 
                           n9170);
   U10066 : OAI211_X1 port map( C1 => n11859, C2 => n8304, A => n9167, B => 
                           n9166, ZN => n9171);
   U10067 : XNOR2_X1 port map( A => n9168, B => n7974, ZN => n9172);
   U10068 : NAND2_X1 port map( A1 => DataPath_ALUhw_i_Q_EXTENDED_34_port, A2 =>
                           n10094, ZN => n9174);
   U10069 : NOR3_X1 port map( A1 => n9164, A2 => n9163, A3 => n9162, ZN => 
                           n9175);
   U10070 : OAI22_X1 port map( A1 => n10004, A2 => n10106, B1 => n10001, B2 => 
                           n10056, ZN => n9162);
   U10071 : OAI22_X1 port map( A1 => n9975, A2 => n10038, B1 => n9885, B2 => 
                           n10059, ZN => n9163);
   U10072 : OAI211_X1 port map( C1 => n9153, C2 => n10104, A => n9152, B => 
                           n9151, ZN => n9164);
   U10073 : AOI22_X1 port map( A1 => n9247, A2 => n10116, B1 => n10110, B2 => 
                           n9972, ZN => n9151);
   U10074 : AOI22_X1 port map( A1 => n9150, A2 => n10113, B1 => n10121, B2 => 
                           n9888, ZN => n9152);
   U10075 : INV_X1 port map( A => n9150, ZN => n9185);
   U10076 : OAI21_X1 port map( B1 => n9148, B2 => n9147, A => n9193, ZN => 
                           n11857);
   U10077 : NOR2_X1 port map( A1 => n9131, A2 => n9130, ZN => n9147);
   U10078 : INV_X1 port map( A => n9132, ZN => n9148);
   U10079 : NOR2_X1 port map( A1 => n9129, A2 => n9196, ZN => n9132);
   U10080 : INV_X1 port map( A => n9193, ZN => n9129);
   U10081 : OAI21_X1 port map( B1 => n9196, B2 => n9149, A => n9193, ZN => 
                           n11856);
   U10082 : AND2_X1 port map( A1 => n9194, A2 => n9198, ZN => n10427);
   U10083 : AND2_X1 port map( A1 => C620_DATA2_12, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_12_port);
   U10084 : NAND2_X1 port map( A1 => n9131, A2 => n9130, ZN => n9149);
   U10085 : XNOR2_X1 port map( A => n8020, B => n8566, ZN => n9131);
   U10086 : NAND2_X1 port map( A1 => n9780, A2 => n8566, ZN => n11859);
   U10087 : NOR2_X1 port map( A1 => n9017, A2 => n9016, ZN => n9134);
   U10088 : OAI21_X1 port map( B1 => n9015, B2 => n9757, A => n9014, ZN => 
                           n9016);
   U10089 : AOI22_X1 port map( A1 => n9586, A2 => n9139, B1 => n9140, B2 => 
                           n7789, ZN => n9014);
   U10090 : OAI211_X1 port map( C1 => n9009, C2 => n8402, A => n9008, B => 
                           n9007, ZN => n9017);
   U10091 : AOI22_X1 port map( A1 => n9047, A2 => n9348, B1 => n9542, B2 => 
                           n9532, ZN => n9007);
   U10092 : NAND2_X1 port map( A1 => n9005, A2 => n9137, ZN => n9008);
   U10093 : OAI21_X1 port map( B1 => n8398, B2 => n9002, A => n9001, ZN => 
                           n9150);
   U10094 : AOI211_X1 port map( C1 => n9586, C2 => n9176, A => n9000, B => 
                           n8999, ZN => n9001);
   U10095 : OAI21_X1 port map( B1 => n9015, B2 => n9472, A => n8998, ZN => 
                           n8999);
   U10096 : AOI22_X1 port map( A1 => n9047, A2 => n9707, B1 => n9542, B2 => 
                           n9470, ZN => n8998);
   U10097 : OAI22_X1 port map( A1 => n9658, A2 => n8992, B1 => n11865, B2 => 
                           n7985, ZN => n9000);
   U10098 : INV_X1 port map( A => n10431, ZN => n8992);
   U10099 : INV_X1 port map( A => n9005, ZN => n9002);
   U10100 : AOI211_X1 port map( C1 => n7913, C2 => n9005, A => n8987, B => 
                           n8986, ZN => n9153);
   U10101 : OAI211_X1 port map( C1 => n9015, C2 => n9499, A => n8985, B => 
                           n8984, ZN => n8986);
   U10102 : NAND2_X1 port map( A1 => n9542, A2 => n9501, ZN => n8984);
   U10103 : AOI22_X1 port map( A1 => n9047, A2 => n8981, B1 => n9586, B2 => 
                           n9158, ZN => n8985);
   U10104 : INV_X1 port map( A => n9384, ZN => n8981);
   U10105 : AOI21_X1 port map( B1 => n9009, B2 => n9755, A => n9504, ZN => 
                           n8987);
   U10106 : INV_X1 port map( A => n9030, ZN => n9009);
   U10107 : INV_X1 port map( A => n9888, ZN => n9135);
   U10108 : OAI222_X1 port map( A1 => n11881, A2 => n9996, B1 => n11880, B2 => 
                           n9995, C1 => n11884, C2 => n8317, ZN => n7017);
   U10109 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_37_port, B2 =>
                           n10094, A => n9994, ZN => n9995);
   U10110 : OAI211_X1 port map( C1 => n9993, C2 => n9992, A => n9991, B => 
                           n9990, ZN => n9994);
   U10111 : AOI211_X1 port map( C1 => n9989, C2 => n10088, A => n9988, B => 
                           n9987, ZN => n9990);
   U10112 : NOR3_X1 port map( A1 => n10084, A2 => n9986, A3 => n8560, ZN => 
                           n9987);
   U10113 : NOR3_X1 port map( A1 => n10082, A2 => n7827, A3 => n7775, ZN => 
                           n9988);
   U10114 : XNOR2_X1 port map( A => n9986, B => n7775, ZN => n9989);
   U10115 : NAND2_X1 port map( A1 => n10426, A2 => n9984, ZN => n9991);
   U10116 : XNOR2_X1 port map( A => n9983, B => n9982, ZN => n9984);
   U10117 : XNOR2_X1 port map( A => n9983, B => n9981, ZN => n9992);
   U10118 : NOR3_X1 port map( A1 => n9980, A2 => n9979, A3 => n9978, ZN => 
                           n9996);
   U10119 : OAI22_X1 port map( A1 => n10004, A2 => n10046, B1 => n10003, B2 => 
                           n9977, ZN => n9978);
   U10120 : OAI22_X1 port map( A1 => n9976, A2 => n10002, B1 => n10001, B2 => 
                           n10059, ZN => n9979);
   U10121 : OAI211_X1 port map( C1 => n9975, C2 => n10104, A => n9974, B => 
                           n9973, ZN => n9980);
   U10122 : AOI22_X1 port map( A1 => n10044, A2 => n10430, B1 => n9972, B2 => 
                           n10112, ZN => n9973);
   U10123 : AOI22_X1 port map( A1 => n9971, A2 => n10113, B1 => n9997, B2 => 
                           n10117, ZN => n9974);
   U10124 : OAI222_X1 port map( A1 => n11881, A2 => n10025, B1 => n11880, B2 =>
                           n10024, C1 => n11884, C2 => n8318, ZN => n7014);
   U10125 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_41_port, B2 =>
                           n10094, A => n10023, ZN => n10024);
   U10126 : OAI21_X1 port map( B1 => n10022, B2 => n11878, A => n10021, ZN => 
                           n10023);
   U10127 : AOI211_X1 port map( C1 => n10020, C2 => n10088, A => n10019, B => 
                           n10018, ZN => n10021);
   U10128 : NOR3_X1 port map( A1 => n10084, A2 => n10017, A3 => n7798, ZN => 
                           n10018);
   U10129 : NOR3_X1 port map( A1 => n10082, A2 => n7824, A3 => 
                           DP_OP_751_130_6421_n1425, ZN => n10019);
   U10130 : XNOR2_X1 port map( A => n10017, B => DP_OP_751_130_6421_n1425, ZN 
                           => n10020);
   U10131 : XNOR2_X1 port map( A => n10015, B => n10014, ZN => n10022);
   U10132 : NOR2_X1 port map( A1 => n10013, A2 => n10012, ZN => n10014);
   U10133 : INV_X1 port map( A => n10011, ZN => n10013);
   U10134 : AOI21_X1 port map( B1 => n10010, B2 => n10009, A => n10008, ZN => 
                           n10015);
   U10135 : NOR3_X1 port map( A1 => n10007, A2 => n10006, A3 => n10005, ZN => 
                           n10025);
   U10136 : OAI22_X1 port map( A1 => n10004, A2 => n10066, B1 => n10040, B2 => 
                           n10046, ZN => n10005);
   U10137 : OAI22_X1 port map( A1 => n10003, A2 => n10002, B1 => n10001, B2 => 
                           n10104, ZN => n10006);
   U10138 : OAI211_X1 port map( C1 => n10039, C2 => n10056, A => n10000, B => 
                           n9999, ZN => n10007);
   U10139 : AOI22_X1 port map( A1 => n10120, A2 => n10044, B1 => n10043, B2 => 
                           n10110, ZN => n9999);
   U10140 : AOI22_X1 port map( A1 => n9998, A2 => n10430, B1 => n10112, B2 => 
                           n9997, ZN => n10000);
   U10141 : OAI22_X1 port map( A1 => n9879, A2 => n11885, B1 => n499, B2 => 
                           n11884, ZN => n7013);
   U10142 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_42_port, B2 =>
                           n10094, A => n9878, ZN => n9879);
   U10143 : OAI211_X1 port map( C1 => n9877, C2 => n11878, A => n9876, B => 
                           n9875, ZN => n9878);
   U10144 : OAI21_X1 port map( B1 => n9870, B2 => n9869, A => n9897, ZN => 
                           n9876);
   U10145 : OAI211_X1 port map( C1 => n9868, C2 => n10002, A => n9867, B => 
                           n9866, ZN => n9869);
   U10146 : NAND2_X1 port map( A1 => n9865, A2 => n10120, ZN => n9866);
   U10147 : AOI22_X1 port map( A1 => n9890, A2 => n10045, B1 => n10113, B2 => 
                           n11866, ZN => n9867);
   U10148 : OAI211_X1 port map( C1 => n10067, C2 => n10106, A => n9864, B => 
                           n9863, ZN => n9870);
   U10149 : AOI22_X1 port map( A1 => n10112, A2 => n10044, B1 => n10043, B2 => 
                           n10116, ZN => n9863);
   U10150 : AOI22_X1 port map( A1 => n9998, A2 => n10117, B1 => n10110, B2 => 
                           n9862, ZN => n9864);
   U10151 : XNOR2_X1 port map( A => n9861, B => n9860, ZN => n9877);
   U10152 : XNOR2_X1 port map( A => n9859, B => n9871, ZN => n9860);
   U10153 : OAI22_X1 port map( A1 => n9858, A2 => n11885, B1 => n500, B2 => 
                           n11884, ZN => n7012);
   U10154 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_43_port, B2 =>
                           n10094, A => n9857, ZN => n9858);
   U10155 : OAI211_X1 port map( C1 => n9856, C2 => n11878, A => n9855, B => 
                           n9854, ZN => n9857);
   U10156 : OAI21_X1 port map( B1 => n9853, B2 => n9852, A => n9897, ZN => 
                           n9854);
   U10157 : OAI211_X1 port map( C1 => n10067, C2 => n10056, A => n9851, B => 
                           n9850, ZN => n9852);
   U10158 : AOI22_X1 port map( A1 => n10121, A2 => n10044, B1 => n10043, B2 => 
                           n10120, ZN => n9850);
   U10159 : AOI22_X1 port map( A1 => n9862, A2 => n10116, B1 => n10430, B2 => 
                           n10064, ZN => n9851);
   U10160 : INV_X1 port map( A => n10039, ZN => n9862);
   U10161 : OAI211_X1 port map( C1 => n9868, C2 => n10066, A => n9849, B => 
                           n9848, ZN => n9853);
   U10162 : AOI22_X1 port map( A1 => n11866, A2 => n10045, B1 => n9865, B2 => 
                           n10112, ZN => n9848);
   U10163 : NAND2_X1 port map( A1 => n9998, A2 => n10110, ZN => n9849);
   U10164 : AOI211_X1 port map( C1 => n9847, C2 => n10088, A => n9846, B => 
                           n9845, ZN => n9855);
   U10165 : NOR3_X1 port map( A1 => n10084, A2 => n8401, A3 => n7803, ZN => 
                           n9845);
   U10166 : NOR3_X1 port map( A1 => n10082, A2 => n7828, A3 => 
                           DP_OP_751_130_6421_n1323, ZN => n9846);
   U10167 : XNOR2_X1 port map( A => n8401, B => DP_OP_751_130_6421_n1323, ZN =>
                           n9847);
   U10168 : XNOR2_X1 port map( A => n9842, B => n9841, ZN => n9856);
   U10169 : NOR2_X1 port map( A1 => n9840, A2 => n9839, ZN => n9841);
   U10170 : INV_X1 port map( A => n9838, ZN => n9840);
   U10171 : OAI22_X1 port map( A1 => n9906, A2 => n11885, B1 => n496, B2 => 
                           n11884, ZN => n7018);
   U10172 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_36_port, B2 =>
                           n10094, A => n9905, ZN => n9906);
   U10173 : OAI211_X1 port map( C1 => n9904, C2 => n7875, A => n9902, B => 
                           n9901, ZN => n9905);
   U10174 : OAI21_X1 port map( B1 => n9900, B2 => n9899, A => n10426, ZN => 
                           n9901);
   U10175 : INV_X1 port map( A => n9981, ZN => n9899);
   U10176 : INV_X1 port map( A => n9982, ZN => n9900);
   U10177 : AOI22_X1 port map( A1 => n9898, A2 => n9897, B1 => n7875, B2 => 
                           n9896, ZN => n9902);
   U10178 : OAI21_X1 port map( B1 => n9993, B2 => n9895, A => n9894, ZN => 
                           n9896);
   U10179 : AOI22_X1 port map( A1 => n9997, A2 => n10430, B1 => n9890, B2 => 
                           n10110, ZN => n9891);
   U10180 : AOI22_X1 port map( A1 => n11866, A2 => n10117, B1 => n9889, B2 => 
                           n10116, ZN => n9892);
   U10181 : AOI211_X1 port map( C1 => n10045, C2 => n9888, A => n9887, B => 
                           n9886, ZN => n9893);
   U10182 : OAI22_X1 port map( A1 => n9975, A2 => n10066, B1 => n9885, B2 => 
                           n10002, ZN => n9886);
   U10183 : INV_X1 port map( A => n9971, ZN => n9885);
   U10184 : AOI211_X1 port map( C1 => n9030, C2 => n9912, A => n8959, B => 
                           n8958, ZN => n9975);
   U10185 : OAI211_X1 port map( C1 => n9986, C2 => n9505, A => n8957, B => 
                           n8956, ZN => n8958);
   U10186 : AOI22_X1 port map( A1 => n9047, A2 => n9228, B1 => n9586, B2 => 
                           n9227, ZN => n8956);
   U10187 : AOI21_X1 port map( B1 => n9037, B2 => n7827, A => n8950, ZN => 
                           n8957);
   U10188 : OAI22_X1 port map( A1 => n8949, A2 => n9496, B1 => n9755, B2 => 
                           n9913, ZN => n8950);
   U10189 : INV_X1 port map( A => n9419, ZN => n8949);
   U10190 : NOR2_X1 port map( A1 => n9015, A2 => n9674, ZN => n8959);
   U10191 : INV_X1 port map( A => n9045, ZN => n9015);
   U10192 : OAI22_X1 port map( A1 => n9976, A2 => n10038, B1 => n9884, B2 => 
                           n10059, ZN => n9887);
   U10193 : INV_X1 port map( A => n9247, ZN => n9976);
   U10194 : NAND4_X1 port map( A1 => n8976, A2 => n8975, A3 => n8974, A4 => 
                           n8973, ZN => n9888);
   U10195 : AOI22_X1 port map( A1 => n9586, A2 => n9209, B1 => n7789, B2 => 
                           n9427, ZN => n8973);
   U10196 : AOI22_X1 port map( A1 => n9047, A2 => n8968, B1 => n9542, B2 => 
                           n9430, ZN => n8974);
   U10197 : INV_X1 port map( A => n9659, ZN => n8968);
   U10198 : AOI22_X1 port map( A1 => n9045, A2 => n9208, B1 => n9442, B2 => 
                           n9030, ZN => n8975);
   U10199 : NAND2_X1 port map( A1 => n9005, A2 => n7875, ZN => n8976);
   U10200 : NAND2_X1 port map( A1 => n8962, A2 => n9505, ZN => n9005);
   U10201 : INV_X1 port map( A => n9037, ZN => n8962);
   U10202 : AOI211_X1 port map( C1 => n10088, C2 => n9883, A => n9882, B => 
                           n9881, ZN => n9904);
   U10203 : NOR2_X1 port map( A1 => n9993, A2 => n9880, ZN => n9881);
   U10204 : NOR2_X1 port map( A1 => n9883, A2 => n10082, ZN => n9882);
   U10205 : OAI222_X1 port map( A1 => n11885, A2 => n9837, B1 => n11881, B2 => 
                           n9836, C1 => n11884, C2 => n501, ZN => n7011);
   U10206 : NOR4_X1 port map( A1 => n9835, A2 => n9834, A3 => n9833, A4 => 
                           n9832, ZN => n9836);
   U10207 : OAI21_X1 port map( B1 => n10067, B2 => n9977, A => n9831, ZN => 
                           n9832);
   U10208 : AOI22_X1 port map( A1 => n10113, A2 => n10044, B1 => n10043, B2 => 
                           n10112, ZN => n9831);
   U10209 : OAI22_X1 port map( A1 => n10039, A2 => n10059, B1 => n9830, B2 => 
                           n10056, ZN => n9833);
   U10210 : OAI22_X1 port map( A1 => n9868, A2 => n10104, B1 => n10040, B2 => 
                           n10002, ZN => n9834);
   U10211 : OAI22_X1 port map( A1 => n10058, A2 => n10046, B1 => n10041, B2 => 
                           n10106, ZN => n9835);
   U10212 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_44_port, B2 =>
                           n10094, A => n9829, ZN => n9837);
   U10213 : OAI21_X1 port map( B1 => n10037, B2 => n9828, A => n9827, ZN => 
                           n9829);
   U10214 : AOI21_X1 port map( B1 => n10031, B2 => n9828, A => n9826, ZN => 
                           n9827);
   U10215 : OR2_X1 port map( A1 => n10029, A2 => n10027, ZN => n9828);
   U10216 : INV_X1 port map( A => n9972, ZN => n9884);
   U10217 : AOI21_X1 port map( B1 => n9037, B2 => n9240, A => n9036, ZN => 
                           n9038);
   U10218 : OAI22_X1 port map( A1 => n9496, A2 => n9035, B1 => n9327, B2 => 
                           n9034, ZN => n9036);
   U10219 : INV_X1 port map( A => n9366, ZN => n9035);
   U10220 : NOR2_X1 port map( A1 => n9658, A2 => n7809, ZN => n9037);
   U10221 : AOI22_X1 port map( A1 => n9045, A2 => n9620, B1 => n10070, B2 => 
                           n9030, ZN => n9039);
   U10222 : NOR2_X1 port map( A1 => n9658, A2 => i_ALU_OP_2_port, ZN => n9030);
   U10223 : AOI21_X1 port map( B1 => n9586, B2 => n9221, A => n9028, ZN => 
                           n9040);
   U10224 : OAI22_X1 port map( A1 => n8400, A2 => n9505, B1 => n9755, B2 => 
                           n9619, ZN => n9028);
   U10225 : AND2_X1 port map( A1 => C620_DATA2_14, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_14_port);
   U10226 : INV_X1 port map( A => n9034, ZN => n9047);
   U10227 : NAND2_X1 port map( A1 => n10103, A2 => n8951, ZN => n9034);
   U10228 : NAND2_X1 port map( A1 => n8189, A2 => i_ALU_OP_2_port, ZN => n8951)
                           ;
   U10229 : NOR2_X1 port map( A1 => n9246, A2 => n8189, ZN => n9045);
   U10230 : NAND2_X1 port map( A1 => n9255, A2 => n9207, ZN => n11862);
   U10231 : NOR2_X1 port map( A1 => n9256, A2 => n11878, ZN => n10426);
   U10232 : NAND2_X1 port map( A1 => n9256, A2 => n9780, ZN => n9993);
   U10233 : INV_X1 port map( A => n9257, ZN => n9252);
   U10234 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_40_port, B2 =>
                           n10094, A => n9281, ZN => n11863);
   U10235 : OAI211_X1 port map( C1 => n9280, C2 => n9279, A => n9278, B => 
                           n9277, ZN => n9281);
   U10236 : OAI211_X1 port map( C1 => n9276, C2 => n10010, A => n9275, B => 
                           n9780, ZN => n9277);
   U10237 : OAI21_X1 port map( B1 => n8437, B2 => n9274, A => n10010, ZN => 
                           n9275);
   U10238 : INV_X1 port map( A => n10009, ZN => n9276);
   U10239 : AOI22_X1 port map( A1 => n9273, A2 => n9897, B1 => n9279, B2 => 
                           n9272, ZN => n9278);
   U10240 : OR3_X1 port map( A1 => n9270, A2 => n9269, A3 => n9268, ZN => n9273
                           );
   U10241 : OAI22_X1 port map( A1 => n10004, A2 => n10002, B1 => n10003, B2 => 
                           n10038, ZN => n9268);
   U10242 : INV_X1 port map( A => n11866, ZN => n10003);
   U10243 : NAND4_X1 port map( A1 => n9184, A2 => n9183, A3 => n9182, A4 => 
                           n9181, ZN => n11866);
   U10244 : NAND2_X1 port map( A1 => n9703, A2 => n7789, ZN => n9181);
   U10245 : NAND2_X1 port map( A1 => n9245, A2 => n9706, ZN => n9182);
   U10246 : AOI22_X1 port map( A1 => n9586, A2 => n7804, B1 => n9730, B2 => 
                           n9702, ZN => n9183);
   U10247 : INV_X1 port map( A => n9178, ZN => n9184);
   U10248 : OAI21_X1 port map( B1 => n9246, B2 => n9355, A => n9177, ZN => 
                           n9178);
   U10249 : NAND2_X1 port map( A1 => n9176, A2 => n10103, ZN => n9177);
   U10250 : NAND2_X1 port map( A1 => n9477, A2 => n8991, ZN => n9176);
   U10251 : NAND2_X1 port map( A1 => n9013, A2 => n8434, ZN => n8991);
   U10252 : INV_X1 port map( A => n9890, ZN => n10004);
   U10253 : OAI211_X1 port map( C1 => n9161, C2 => n9755, A => n9160, B => 
                           n9159, ZN => n9890);
   U10254 : AOI22_X1 port map( A1 => n9730, A2 => n9507, B1 => n9158, B2 => 
                           n10103, ZN => n9159);
   U10255 : NAND2_X1 port map( A1 => n9494, A2 => n8980, ZN => n9158);
   U10256 : NAND2_X1 port map( A1 => n9013, A2 => n7777, ZN => n8980);
   U10257 : AOI22_X1 port map( A1 => n9155, A2 => n9725, B1 => n9729, B2 => 
                           n9245, ZN => n9160);
   U10258 : AOI21_X1 port map( B1 => n7806, B2 => n9504, A => n9627, ZN => 
                           n9155);
   U10259 : INV_X1 port map( A => n9731, ZN => n9161);
   U10260 : OAI22_X1 port map( A1 => n9267, A2 => n10046, B1 => n10001, B2 => 
                           n10066, ZN => n9269);
   U10261 : INV_X1 port map( A => n9889, ZN => n10001);
   U10262 : NAND4_X1 port map( A1 => n9144, A2 => n9143, A3 => n9142, A4 => 
                           n9141, ZN => n9889);
   U10263 : NAND2_X1 port map( A1 => n9768, A2 => n7789, ZN => n9141);
   U10264 : NAND2_X1 port map( A1 => n9140, A2 => n7788, ZN => n9142);
   U10265 : AOI22_X1 port map( A1 => n10103, A2 => n9139, B1 => n9730, B2 => 
                           n9138, ZN => n9143);
   U10266 : INV_X1 port map( A => n9764, ZN => n9138);
   U10267 : NAND2_X1 port map( A1 => n9533, A2 => n9012, ZN => n9139);
   U10268 : NAND2_X1 port map( A1 => n7924, A2 => n7806, ZN => n9012);
   U10269 : NAND2_X1 port map( A1 => n9245, A2 => n9136, ZN => n9144);
   U10270 : INV_X1 port map( A => n9757, ZN => n9136);
   U10271 : INV_X1 port map( A => n10044, ZN => n9267);
   U10272 : OAI211_X1 port map( C1 => n10039, C2 => n10106, A => n9266, B => 
                           n9265, ZN => n9270);
   U10273 : AOI22_X1 port map( A1 => n10117, A2 => n10043, B1 => n9972, B2 => 
                           n10045, ZN => n9265);
   U10274 : AOI22_X1 port map( A1 => n9997, A2 => n10120, B1 => n10110, B2 => 
                           n9865, ZN => n9266);
   U10275 : INV_X1 port map( A => n9868, ZN => n9997);
   U10276 : NOR2_X1 port map( A1 => n9218, A2 => n9217, ZN => n9868);
   U10277 : OAI211_X1 port map( C1 => n9246, C2 => n9659, A => n9216, B => 
                           n9215, ZN => n9217);
   U10278 : NAND2_X1 port map( A1 => n9542, A2 => n7875, ZN => n9215);
   U10279 : NAND2_X1 port map( A1 => n9664, A2 => n7789, ZN => n9216);
   U10280 : NAND2_X1 port map( A1 => n9586, A2 => n9442, ZN => n9210);
   U10281 : AOI22_X1 port map( A1 => n9547, A2 => n9821, B1 => n10103, B2 => 
                           n9209, ZN => n9211);
   U10282 : OAI211_X1 port map( C1 => n7799, C2 => n9531, A => n8971, B => 
                           n8970, ZN => n9209);
   U10283 : NAND2_X1 port map( A1 => n7875, A2 => n11861, ZN => n8970);
   U10284 : INV_X1 port map( A => n8969, ZN => n8971);
   U10285 : NAND2_X1 port map( A1 => n9245, A2 => n9208, ZN => n9212);
   U10286 : INV_X1 port map( A => n9656, ZN => n9208);
   U10287 : AOI21_X1 port map( B1 => n9263, B2 => n9780, A => n9262, ZN => 
                           n9280);
   U10288 : XNOR2_X1 port map( A => n10010, B => n9274, ZN => n9263);
   U10289 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(19), ZN => n11761);
   U10290 : AOI22_X1 port map( A1 => n8426, A2 => IRAM_DATA(13), B1 => 
                           IR_13_port, B2 => n10413, ZN => n2883);
   U10291 : AOI22_X1 port map( A1 => n8426, A2 => IRAM_DATA(21), B1 => 
                           IR_21_port, B2 => n10413, ZN => n2878);
   U10292 : AOI22_X1 port map( A1 => n8426, A2 => IRAM_DATA(24), B1 => 
                           IR_24_port, B2 => n10413, ZN => n2875);
   U10293 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(20), ZN => n11762);
   U10294 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(18), ZN => n11760);
   U10295 : AOI22_X1 port map( A1 => n8426, A2 => n11769, B1 => n8396, B2 => 
                           n10413, ZN => n7119);
   U10296 : AOI22_X1 port map( A1 => n8426, A2 => IRAM_DATA(10), B1 => 
                           IR_10_port, B2 => n10413, ZN => n2886);
   U10297 : AOI22_X1 port map( A1 => n8426, A2 => n11768, B1 => n163, B2 => 
                           n10413, ZN => n7121);
   U10298 : OAI211_X1 port map( C1 => n173, C2 => n10405, A => n10404, B => 
                           n10193, ZN => i_ADD_WS1_3_port);
   U10299 : AOI211_X1 port map( C1 => n8287, C2 => n10196, A => n8424, B => 
                           n10195, ZN => n10197);
   U10300 : OAI22_X1 port map( A1 => n10194, A2 => n8199, B1 => n170, B2 => 
                           n7621, ZN => n10195);
   U10301 : INV_X1 port map( A => n10405, ZN => n10196);
   U10302 : AOI22_X1 port map( A1 => n8426, A2 => n11766, B1 => n8223, B2 => 
                           n10413, ZN => n7123);
   U10303 : NAND4_X1 port map( A1 => n9238, A2 => n9237, A3 => n9236, A4 => 
                           n9235, ZN => n10044);
   U10304 : NAND2_X1 port map( A1 => n9704, A2 => n9669, ZN => n9235);
   U10305 : NAND2_X1 port map( A1 => n9245, A2 => n9233, ZN => n9236);
   U10306 : INV_X1 port map( A => n9674, ZN => n9233);
   U10307 : AND2_X1 port map( A1 => n9232, A2 => n9231, ZN => n9237);
   U10308 : NAND2_X1 port map( A1 => n9230, A2 => n9730, ZN => n9231);
   U10309 : INV_X1 port map( A => n9670, ZN => n9230);
   U10310 : INV_X1 port map( A => n9668, ZN => n9228);
   U10311 : AOI22_X1 port map( A1 => n9586, A2 => n9912, B1 => n10103, B2 => 
                           n9227, ZN => n9238);
   U10312 : NAND2_X1 port map( A1 => n9416, A2 => n8955, ZN => n9227);
   U10313 : NAND2_X1 port map( A1 => n9013, A2 => n9962, ZN => n8955);
   U10314 : INV_X1 port map( A => n9865, ZN => n10040);
   U10315 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(15), ZN => n11757);
   U10316 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(17), ZN => n11759);
   U10317 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(16), ZN => n11758);
   U10318 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(12), ZN => n11999);
   U10319 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(11), ZN => n12000);
   U10320 : OAI21_X1 port map( B1 => n8418, B2 => n8234, A => n10406, ZN => n41
                           );
   U10321 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(7), ZN => n10406);
   U10322 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(8), ZN => n11755);
   U10323 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(2), ZN => n12001);
   U10324 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(25), ZN => n11765);
   U10325 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(22), ZN => n11763);
   U10326 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(0), ZN => n12002);
   U10327 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(14), ZN => n11756);
   U10328 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(23), ZN => n11764);
   U10329 : AND2_X1 port map( A1 => C620_DATA2_15, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_15_port);
   U10330 : AOI22_X1 port map( A1 => n8426, A2 => IRAM_DATA(29), B1 => 
                           IR_29_port, B2 => n10413, ZN => n10414);
   U10331 : INV_X1 port map( A => n10409, ZN => n38);
   U10332 : AOI22_X1 port map( A1 => n8426, A2 => IRAM_DATA(4), B1 => IR_4_port
                           , B2 => n10413, ZN => n10409);
   U10333 : INV_X1 port map( A => n10412, ZN => n7134);
   U10334 : AOI22_X1 port map( A1 => n8426, A2 => IRAM_DATA(9), B1 => IR_9_port
                           , B2 => n10413, ZN => n10412);
   U10335 : INV_X1 port map( A => n10410, ZN => n37);
   U10336 : AOI22_X1 port map( A1 => n8426, A2 => IRAM_DATA(3), B1 => IR_3_port
                           , B2 => n10413, ZN => n10410);
   U10337 : AOI22_X1 port map( A1 => n8426, A2 => IRAM_DATA(1), B1 => IR_1_port
                           , B2 => n10413, ZN => n10411);
   U10338 : OAI21_X1 port map( B1 => n8418, B2 => n8228, A => n10407, ZN => n40
                           );
   U10339 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(6), ZN => n10407);
   U10340 : OAI21_X1 port map( B1 => n8418, B2 => n8198, A => n10408, ZN => n39
                           );
   U10341 : NAND2_X1 port map( A1 => n8426, A2 => IRAM_DATA(5), ZN => n10408);
   U10342 : OAI222_X1 port map( A1 => n11885, A2 => n9820, B1 => n11881, B2 => 
                           n9819, C1 => n11884, C2 => n502, ZN => n7009);
   U10343 : NOR3_X1 port map( A1 => n9818, A2 => n9817, A3 => n9816, ZN => 
                           n9819);
   U10344 : OAI211_X1 port map( C1 => n10067, C2 => n10059, A => n9815, B => 
                           n9814, ZN => n9816);
   U10345 : AOI22_X1 port map( A1 => n10113, A2 => n10043, B1 => n9865, B2 => 
                           n10045, ZN => n9814);
   U10346 : NAND4_X1 port map( A1 => n9226, A2 => n9225, A3 => n9224, A4 => 
                           n9223, ZN => n9865);
   U10347 : OAI211_X1 port map( C1 => n10070, C2 => n9531, A => n9623, B => 
                           n7788, ZN => n9223);
   U10348 : AOI22_X1 port map( A1 => n9222, A2 => n9730, B1 => n10103, B2 => 
                           n9221, ZN => n9224);
   U10349 : INV_X1 port map( A => n9362, ZN => n9222);
   U10350 : NAND2_X1 port map( A1 => n9219, A2 => n7789, ZN => n9225);
   U10351 : INV_X1 port map( A => n9628, ZN => n9219);
   U10352 : NAND2_X1 port map( A1 => n9245, A2 => n9620, ZN => n9226);
   U10353 : AOI22_X1 port map( A1 => n10065, A2 => n10430, B1 => n10116, B2 => 
                           n10064, ZN => n9815);
   U10354 : OAI22_X1 port map( A1 => n10039, A2 => n10002, B1 => n10060, B2 => 
                           n10056, ZN => n9817);
   U10355 : OAI22_X1 port map( A1 => n10058, A2 => n10038, B1 => n10041, B2 => 
                           n9977, ZN => n9818);
   U10356 : INV_X1 port map( A => n10063, ZN => n10041);
   U10357 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_46_port, B2 =>
                           n10094, A => n9813, ZN => n9820);
   U10358 : OAI211_X1 port map( C1 => n10037, C2 => n9812, A => n9811, B => 
                           n9810, ZN => n9813);
   U10359 : NAND2_X1 port map( A1 => n10031, A2 => n9805, ZN => n9811);
   U10360 : AND2_X1 port map( A1 => C620_DATA2_16, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_16_port);
   U10361 : OAI222_X1 port map( A1 => n11885, A2 => n9801, B1 => n11881, B2 => 
                           n9800, C1 => n11884, C2 => n503, ZN => n7008);
   U10362 : NOR3_X1 port map( A1 => n9799, A2 => n9798, A3 => n9797, ZN => 
                           n9800);
   U10363 : OAI22_X1 port map( A1 => n9796, A2 => n10056, B1 => n10067, B2 => 
                           n10038, ZN => n9797);
   U10364 : INV_X1 port map( A => n10065, ZN => n9796);
   U10365 : OAI22_X1 port map( A1 => n9830, A2 => n10059, B1 => n10060, B2 => 
                           n9977, ZN => n9798);
   U10366 : OAI211_X1 port map( C1 => n10039, C2 => n10066, A => n9795, B => 
                           n9794, ZN => n9799);
   U10367 : AOI22_X1 port map( A1 => n10045, A2 => n10043, B1 => n10062, B2 => 
                           n10430, ZN => n9794);
   U10368 : NAND2_X1 port map( A1 => n7788, A2 => n11853, ZN => n9246);
   U10369 : NOR2_X1 port map( A1 => n10098, A2 => n8189, ZN => n9245);
   U10370 : OR2_X1 port map( A1 => n9583, A2 => n8303, ZN => n9244);
   U10371 : AND2_X1 port map( A1 => n10081, A2 => n7806, ZN => n9243);
   U10372 : AOI22_X1 port map( A1 => n9998, A2 => n10121, B1 => n10116, B2 => 
                           n10063, ZN => n9795);
   U10373 : INV_X1 port map( A => n10058, ZN => n9998);
   U10374 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_47_port, B2 =>
                           n10094, A => n9793, ZN => n9801);
   U10375 : OAI21_X1 port map( B1 => n9792, B2 => n10037, A => n9791, ZN => 
                           n9793);
   U10376 : AOI21_X1 port map( B1 => n10031, B2 => n9790, A => n9789, ZN => 
                           n9791);
   U10377 : OAI211_X1 port map( C1 => n9788, C2 => n10036, A => n9787, B => 
                           n9786, ZN => n9789);
   U10378 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1119, B => n7983, ZN =>
                           n9788);
   U10379 : XNOR2_X1 port map( A => n9783, B => n9782, ZN => n9790);
   U10380 : NOR2_X1 port map( A1 => n9781, A2 => n11878, ZN => n10031);
   U10381 : NAND2_X1 port map( A1 => n9781, A2 => n9780, ZN => n10037);
   U10382 : XNOR2_X1 port map( A => n9779, B => n9782, ZN => n9792);
   U10383 : NOR2_X1 port map( A1 => n9778, A2 => n9777, ZN => n9782);
   U10384 : INV_X1 port map( A => n9776, ZN => n9778);
   U10385 : NOR2_X1 port map( A1 => n9775, A2 => n9783, ZN => n9779);
   U10386 : AOI21_X1 port map( B1 => n9803, B2 => n9804, A => n9774, ZN => 
                           n9783);
   U10387 : INV_X1 port map( A => n9773, ZN => n9774);
   U10388 : AND2_X1 port map( A1 => n9773, A2 => n9772, ZN => n9804);
   U10389 : OAI21_X1 port map( B1 => n9771, B2 => n10029, A => n9770, ZN => 
                           n9803);
   U10390 : INV_X1 port map( A => n9769, ZN => n9771);
   U10391 : AND2_X1 port map( A1 => C620_DATA2_17, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_17_port);
   U10392 : AOI211_X1 port map( C1 => n7788, C2 => n9768, A => n9767, B => 
                           n9766, ZN => n10058);
   U10393 : OAI21_X1 port map( B1 => n9765, B2 => n9764, A => n9763, ZN => 
                           n9766);
   U10394 : AOI21_X1 port map( B1 => n9762, B2 => n9761, A => n9760, ZN => 
                           n9763);
   U10395 : OAI22_X1 port map( A1 => n9759, A2 => n9758, B1 => n9757, B2 => 
                           n7982, ZN => n9760);
   U10396 : NAND2_X1 port map( A1 => n9013, A2 => n9936, ZN => n9758);
   U10397 : NOR2_X1 port map( A1 => n8566, A2 => n11864, ZN => n9013);
   U10398 : AND2_X1 port map( A1 => n9348, A2 => n11853, ZN => n9761);
   U10399 : NOR2_X1 port map( A1 => n9756, A2 => n9755, ZN => n9767);
   U10400 : OAI21_X1 port map( B1 => n9347, B2 => n9531, A => n9533, ZN => 
                           n9768);
   U10401 : AND2_X1 port map( A1 => C620_DATA2_18, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_18_port);
   U10402 : OAI222_X1 port map( A1 => n11885, A2 => n9718, B1 => n11881, B2 => 
                           n9717, C1 => n11884, C2 => n506, ZN => n7004);
   U10403 : NOR3_X1 port map( A1 => n9716, A2 => n9715, A3 => n9714, ZN => 
                           n9717);
   U10404 : OAI22_X1 port map( A1 => n7810, A2 => n10106, B1 => n10057, B2 => 
                           n10046, ZN => n9714);
   U10405 : OAI211_X1 port map( C1 => n9968, C2 => n10056, A => n9713, B => 
                           n9712, ZN => n9715);
   U10406 : AOI22_X1 port map( A1 => n10042, A2 => n10121, B1 => n10112, B2 => 
                           n10065, ZN => n9712);
   U10407 : AOI22_X1 port map( A1 => n10063, A2 => n10113, B1 => n10120, B2 => 
                           n10062, ZN => n9713);
   U10408 : OAI22_X1 port map( A1 => n10061, A2 => n9977, B1 => n9830, B2 => 
                           n10104, ZN => n9716);
   U10409 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_51_port, B2 =>
                           n10094, A => n9700, ZN => n9718);
   U10410 : OAI211_X1 port map( C1 => n9699, C2 => n10055, A => n9698, B => 
                           n9697, ZN => n9700);
   U10411 : AOI211_X1 port map( C1 => n10088, C2 => n9696, A => n9695, B => 
                           n9694, ZN => n9697);
   U10412 : NOR3_X1 port map( A1 => n10084, A2 => n9693, A3 => n7776, ZN => 
                           n9694);
   U10413 : NOR3_X1 port map( A1 => n10082, A2 => n8434, A3 => 
                           DP_OP_751_130_6421_n915, ZN => n9695);
   U10414 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n915, B => n7776, ZN => 
                           n9696);
   U10415 : INV_X1 port map( A => n9687, ZN => n9691);
   U10416 : XNOR2_X1 port map( A => n9685, B => n9689, ZN => n9699);
   U10417 : OAI22_X1 port map( A1 => n9752, A2 => n11885, B1 => n505, B2 => 
                           n11884, ZN => n7005);
   U10418 : AOI211_X1 port map( C1 => DataPath_ALUhw_i_Q_EXTENDED_50_port, C2 
                           => n10094, A => n9751, B => n9750, ZN => n9752);
   U10419 : OAI211_X1 port map( C1 => n9749, C2 => n9748, A => n9747, B => 
                           n9746, ZN => n9750);
   U10420 : OAI211_X1 port map( C1 => n9742, C2 => n9741, A => n9740, B => 
                           n9739, ZN => n9747);
   U10421 : INV_X1 port map( A => n10055, ZN => n9740);
   U10422 : NAND2_X1 port map( A1 => n9686, A2 => n9780, ZN => n10055);
   U10423 : NOR3_X1 port map( A1 => n9738, A2 => n9737, A3 => n9736, ZN => 
                           n9749);
   U10424 : OAI22_X1 port map( A1 => n9830, A2 => n10066, B1 => n10060, B2 => 
                           n10038, ZN => n9736);
   U10425 : INV_X1 port map( A => n10064, ZN => n9830);
   U10426 : OAI211_X1 port map( C1 => n9711, C2 => n9759, A => n9710, B => 
                           n9709, ZN => n10064);
   U10427 : AOI22_X1 port map( A1 => n9708, A2 => n9707, B1 => n9730, B2 => 
                           n9706, ZN => n9709);
   U10428 : INV_X1 port map( A => n9472, ZN => n9706);
   U10429 : INV_X1 port map( A => n9355, ZN => n9707);
   U10430 : INV_X1 port map( A => n9658, ZN => n9708);
   U10431 : AOI22_X1 port map( A1 => n9705, A2 => n7789, B1 => n9703, B2 => 
                           n7788, ZN => n9710);
   U10432 : NAND2_X1 port map( A1 => n9180, A2 => n9477, ZN => n9703);
   U10433 : NAND2_X1 port map( A1 => n9470, A2 => n7806, ZN => n9180);
   U10434 : AOI21_X1 port map( B1 => n9702, B2 => n11879, A => n9701, ZN => 
                           n9711);
   U10435 : INV_X1 port map( A => n11865, ZN => n9701);
   U10436 : OAI211_X1 port map( C1 => n9968, C2 => n10106, A => n9735, B => 
                           n9734, ZN => n9737);
   U10437 : AOI22_X1 port map( A1 => n9733, A2 => n10045, B1 => n10120, B2 => 
                           n10065, ZN => n9734);
   U10438 : INV_X1 port map( A => n10067, ZN => n9733);
   U10439 : NAND2_X1 port map( A1 => n9154, A2 => n9494, ZN => n9731);
   U10440 : NAND2_X1 port map( A1 => n9501, A2 => n7806, ZN => n9154);
   U10441 : INV_X1 port map( A => n9499, ZN => n9729);
   U10442 : OAI21_X1 port map( B1 => n9384, B2 => n8189, A => n9531, ZN => 
                           n9725);
   U10443 : AOI22_X1 port map( A1 => n10063, A2 => n10121, B1 => n10116, B2 => 
                           n10062, ZN => n9735);
   U10444 : OAI22_X1 port map( A1 => n10061, A2 => n10056, B1 => n10057, B2 => 
                           n9977, ZN => n9738);
   U10445 : AOI211_X1 port map( C1 => n9723, C2 => n9722, A => n9721, B => 
                           n9720, ZN => n9751);
   U10446 : INV_X1 port map( A => n10052, ZN => n9720);
   U10447 : NOR2_X1 port map( A1 => n9686, A2 => n11878, ZN => n10052);
   U10448 : INV_X1 port map( A => n9719, ZN => n9721);
   U10449 : NAND2_X1 port map( A1 => n8425, A2 => IRAM_DATA(27), ZN => n11767);
   U10450 : OAI222_X1 port map( A1 => n8205, A2 => n7757, B1 => n11845, B2 => 
                           n11837, C1 => n8313, C2 => n10367, ZN => n7057);
   U10451 : OAI222_X1 port map( A1 => n8208, A2 => n7757, B1 => n11845, B2 => 
                           n11836, C1 => n8321, C2 => n10367, ZN => n7058);
   U10452 : OAI222_X1 port map( A1 => n10366, A2 => n7757, B1 => n10367, B2 => 
                           n207, C1 => n11845, C2 => n10365, ZN => n7056);
   U10453 : INV_X1 port map( A => i_RD1_5_port, ZN => n10365);
   U10454 : NOR2_X1 port map( A1 => n10363, A2 => n10362, ZN => n10364);
   U10455 : INV_X1 port map( A => n10361, ZN => n10363);
   U10456 : OAI211_X1 port map( C1 => n11835, C2 => n11845, A => n10371, B => 
                           n10370, ZN => n7061);
   U10457 : OR3_X1 port map( A1 => n10369, A2 => IRAM_ADDRESS_0_port, A3 => 
                           i_NPC_SEL, ZN => n10370);
   U10458 : OAI222_X1 port map( A1 => n11845, A2 => n10354, B1 => n10367, B2 =>
                           n8284, C1 => n7757, C2 => n10353, ZN => n7054);
   U10459 : XNOR2_X1 port map( A => n10351, B => IRAM_ADDRESS_7_port, ZN => 
                           n10352);
   U10460 : OAI222_X1 port map( A1 => n11885, A2 => n9684, B1 => n11881, B2 => 
                           n9683, C1 => n11884, C2 => n507, ZN => n7003);
   U10461 : NOR3_X1 port map( A1 => n9682, A2 => n9681, A3 => n9680, ZN => 
                           n9683);
   U10462 : OAI22_X1 port map( A1 => n7810, A2 => n10056, B1 => n9969, B2 => 
                           n10106, ZN => n9680);
   U10463 : OAI211_X1 port map( C1 => n9968, C2 => n9977, A => n9678, B => 
                           n9677, ZN => n9681);
   U10464 : AOI22_X1 port map( A1 => n10042, A2 => n10113, B1 => n10121, B2 => 
                           n10065, ZN => n9677);
   U10465 : AOI22_X1 port map( A1 => n10063, A2 => n10045, B1 => n10112, B2 => 
                           n10062, ZN => n9678);
   U10466 : OAI21_X1 port map( B1 => n9666, B2 => n9755, A => n9665, ZN => 
                           n10063);
   U10467 : AOI211_X1 port map( C1 => n7788, C2 => n9664, A => n9663, B => 
                           n9662, ZN => n9665);
   U10468 : OAI22_X1 port map( A1 => n9661, A2 => n9660, B1 => n9659, B2 => 
                           n9658, ZN => n9662);
   U10469 : INV_X1 port map( A => n9657, ZN => n9661);
   U10470 : OAI22_X1 port map( A1 => n7440, A2 => n9759, B1 => n7982, B2 => 
                           n9656, ZN => n9663);
   U10471 : OAI22_X1 port map( A1 => n10061, A2 => n10046, B1 => n10057, B2 => 
                           n10059, ZN => n9682);
   U10472 : AOI211_X1 port map( C1 => DataPath_ALUhw_i_Q_EXTENDED_52_port, C2 
                           => n10094, A => n9655, B => n9654, ZN => n9684);
   U10473 : OAI211_X1 port map( C1 => n9651, C2 => n10036, A => n9966, B => 
                           n9650, ZN => n9652);
   U10474 : NAND2_X1 port map( A1 => n10035, A2 => n9651, ZN => n9650);
   U10475 : OAI211_X1 port map( C1 => n9651, C2 => n10082, A => n9649, B => 
                           n9648, ZN => n9653);
   U10476 : NAND2_X1 port map( A1 => n10088, A2 => n9651, ZN => n9648);
   U10477 : NAND2_X1 port map( A1 => n9964, A2 => n9647, ZN => n9649);
   U10478 : OAI22_X1 port map( A1 => n9647, A2 => n9966, B1 => n9960, B2 => 
                           n9959, ZN => n9655);
   U10479 : INV_X1 port map( A => n10060, ZN => n10042);
   U10480 : AOI21_X1 port map( B1 => n9676, B2 => n9724, A => n9675, ZN => 
                           n10060);
   U10481 : OAI211_X1 port map( C1 => n9674, C2 => n7982, A => n9673, B => 
                           n9672, ZN => n9675);
   U10482 : OAI211_X1 port map( C1 => n11879, C2 => n9912, A => n9671, B => 
                           n10103, ZN => n9672);
   U10483 : NAND2_X1 port map( A1 => n9670, A2 => n11879, ZN => n9671);
   U10484 : NAND2_X1 port map( A1 => n9669, A2 => n7788, ZN => n9673);
   U10485 : NAND2_X1 port map( A1 => n9234, A2 => n9416, ZN => n9669);
   U10486 : NAND2_X1 port map( A1 => n9419, A2 => n7806, ZN => n9234);
   U10487 : OAI21_X1 port map( B1 => n8943, B2 => n9668, A => n9667, ZN => 
                           n9676);
   U10488 : INV_X1 port map( A => n9964, ZN => n9960);
   U10489 : NAND2_X1 port map( A1 => n9646, A2 => n9959, ZN => n9966);
   U10490 : OAI222_X1 port map( A1 => n10350, A2 => n7757, B1 => n10367, B2 => 
                           n206, C1 => n11845, C2 => n10349, ZN => n7053);
   U10491 : XNOR2_X1 port map( A => n10346, B => IRAM_ADDRESS_8_port, ZN => 
                           n10347);
   U10492 : AOI22_X1 port map( A1 => n10418, A2 => i_RD1_9_port, B1 => n10417, 
                           B2 => IRAM_ADDRESS_9_port, ZN => n11838);
   U10493 : NAND2_X1 port map( A1 => n8924, A2 => n8927, ZN => n8925);
   U10494 : INV_X1 port map( A => n8926, ZN => n8924);
   U10495 : OAI22_X1 port map( A1 => n9614, A2 => n11885, B1 => n509, B2 => 
                           n11884, ZN => n7000);
   U10496 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_55_port, B2 =>
                           n10094, A => n9613, ZN => n9614);
   U10497 : OAI21_X1 port map( B1 => n9612, B2 => n9611, A => n9610, ZN => 
                           n9613);
   U10498 : AOI211_X1 port map( C1 => n9897, C2 => n9609, A => n9608, B => 
                           n9607, ZN => n9610);
   U10499 : NOR3_X1 port map( A1 => n9958, A2 => n9606, A3 => n9618, ZN => 
                           n9607);
   U10500 : OAI211_X1 port map( C1 => n9605, C2 => n10036, A => n9604, B => 
                           n9603, ZN => n9608);
   U10501 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n711, B => n9602, ZN => 
                           n9605);
   U10502 : AOI22_X1 port map( A1 => n10121, A2 => n9596, B1 => n9970, B2 => 
                           n10120, ZN => n9597);
   U10503 : INV_X1 port map( A => n10061, ZN => n9596);
   U10504 : AOI22_X1 port map( A1 => n9967, A2 => n10110, B1 => n10116, B2 => 
                           n9679, ZN => n9598);
   U10505 : AOI211_X1 port map( C1 => n10113, C2 => n9595, A => n9594, B => 
                           n9593, ZN => n9599);
   U10506 : OAI22_X1 port map( A1 => n9968, A2 => n10038, B1 => n9592, B2 => 
                           n10056, ZN => n9593);
   U10507 : OAI22_X1 port map( A1 => n9591, A2 => n10104, B1 => n10105, B2 => 
                           n10106, ZN => n9594);
   U10508 : INV_X1 port map( A => n10062, ZN => n9591);
   U10509 : INV_X1 port map( A => n10057, ZN => n9595);
   U10510 : XNOR2_X1 port map( A => n9580, B => n9606, ZN => n9611);
   U10511 : XNOR2_X1 port map( A => n9579, B => n9602, ZN => n9606);
   U10512 : NOR2_X1 port map( A1 => n9578, A2 => n11872, ZN => n9580);
   U10513 : INV_X1 port map( A => n9634, ZN => n9578);
   U10514 : AOI21_X1 port map( B1 => n9646, B2 => n9618, A => n9964, ZN => 
                           n9612);
   U10515 : INV_X1 port map( A => n9958, ZN => n9646);
   U10516 : OAI21_X1 port map( B1 => n10360, B2 => n7757, A => n10359, ZN => 
                           n7055);
   U10517 : AOI22_X1 port map( A1 => n10418, A2 => i_RD1_6_port, B1 => 
                           IRAM_ADDRESS_6_port, B2 => n10417, ZN => n10359);
   U10518 : NAND2_X1 port map( A1 => n7780, A2 => n10356, ZN => n10357);
   U10519 : INV_X1 port map( A => n10368, ZN => n7059);
   U10520 : AOI222_X1 port map( A1 => IRAM_ADDRESS_2_port, A2 => n10417, B1 => 
                           n8194, B2 => intadd_0_SUM_1_port, C1 => n10418, C2 
                           => i_RD1_2_port, ZN => n10368);
   U10521 : AND2_X1 port map( A1 => C620_DATA2_21, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_21_port);
   U10522 : OAI22_X1 port map( A1 => n9645, A2 => n11885, B1 => n508, B2 => 
                           n11884, ZN => n7001);
   U10523 : AOI211_X1 port map( C1 => DataPath_ALUhw_i_Q_EXTENDED_54_port, C2 
                           => n10094, A => n9644, B => n9643, ZN => n9645);
   U10524 : OAI211_X1 port map( C1 => n9642, C2 => n9748, A => n9641, B => 
                           n9640, ZN => n9643);
   U10525 : OAI211_X1 port map( C1 => n9636, C2 => n9635, A => n9964, B => 
                           n9634, ZN => n9641);
   U10526 : NOR2_X1 port map( A1 => n9577, A2 => n11878, ZN => n9964);
   U10527 : NOR3_X1 port map( A1 => n9633, A2 => n9632, A3 => n9631, ZN => 
                           n9642);
   U10528 : OAI211_X1 port map( C1 => n9968, C2 => n10059, A => n9630, B => 
                           n9629, ZN => n9631);
   U10529 : AOI22_X1 port map( A1 => n9679, A2 => n10110, B1 => n10062, B2 => 
                           n10113, ZN => n9629);
   U10530 : NAND4_X1 port map( A1 => n9590, A2 => n9589, A3 => n9588, A4 => 
                           n9587, ZN => n10062);
   U10531 : NAND2_X1 port map( A1 => n9586, A2 => n9585, ZN => n9587);
   U10532 : OAI211_X1 port map( C1 => n11879, C2 => n10081, A => n9584, B => 
                           n10103, ZN => n9588);
   U10533 : AOI22_X1 port map( A1 => n7788, A2 => n9583, B1 => n9730, B2 => 
                           n9582, ZN => n9589);
   U10534 : OAI21_X1 port map( B1 => n9581, B2 => n7789, A => n8229, ZN => 
                           n9590);
   U10535 : NOR2_X1 port map( A1 => n9658, A2 => n7353, ZN => n9581);
   U10536 : OR2_X1 port map( A1 => n7985, A2 => n8943, ZN => n9658);
   U10537 : AOI22_X1 port map( A1 => n10065, A2 => n10045, B1 => n9948, B2 => 
                           n10430, ZN => n9630);
   U10538 : OAI211_X1 port map( C1 => n9628, C2 => n9627, A => n9626, B => 
                           n9625, ZN => n10065);
   U10539 : OAI21_X1 port map( B1 => n9327, B2 => n8189, A => n9531, ZN => 
                           n9623);
   U10540 : INV_X1 port map( A => n7985, ZN => n9724);
   U10541 : AOI22_X1 port map( A1 => n9622, A2 => n9621, B1 => n9730, B2 => 
                           n9620, ZN => n9626);
   U10542 : INV_X1 port map( A => n9333, ZN => n9620);
   U10543 : OAI21_X1 port map( B1 => n9759, B2 => n9619, A => n9728, ZN => 
                           n9622);
   U10544 : AOI21_X1 port map( B1 => n9366, B2 => n7806, A => n9332, ZN => 
                           n9628);
   U10545 : OAI22_X1 port map( A1 => n7810, A2 => n10046, B1 => n9922, B2 => 
                           n10056, ZN => n9632);
   U10546 : OAI22_X1 port map( A1 => n10061, A2 => n10038, B1 => n10057, B2 => 
                           n10002, ZN => n9633);
   U10547 : AOI21_X1 port map( B1 => n9618, B2 => n9617, A => n9958, ZN => 
                           n9644);
   U10548 : NAND2_X1 port map( A1 => n9577, A2 => n9780, ZN => n9958);
   U10549 : NAND2_X1 port map( A1 => n9616, A2 => n9615, ZN => n9617);
   U10550 : INV_X1 port map( A => n9635, ZN => n9615);
   U10551 : NAND2_X1 port map( A1 => n9576, A2 => n9635, ZN => n9618);
   U10552 : INV_X1 port map( A => n9616, ZN => n9576);
   U10553 : NOR2_X1 port map( A1 => n9575, A2 => n9574, ZN => n9616);
   U10554 : OAI22_X1 port map( A1 => n9573, A2 => n11885, B1 => n510, B2 => 
                           n11884, ZN => n6999);
   U10555 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_56_port, B2 =>
                           n10094, A => n9572, ZN => n9573);
   U10556 : OAI211_X1 port map( C1 => n9571, C2 => n9570, A => n9569, B => 
                           n9568, ZN => n9572);
   U10557 : AOI211_X1 port map( C1 => n9567, C2 => n9566, A => n9565, B => 
                           n9564, ZN => n9568);
   U10558 : NOR2_X1 port map( A1 => n9563, A2 => n9748, ZN => n9564);
   U10559 : NOR3_X1 port map( A1 => n9562, A2 => n9561, A3 => n9560, ZN => 
                           n9563);
   U10560 : OAI211_X1 port map( C1 => n9968, C2 => n10002, A => n9559, B => 
                           n9558, ZN => n9560);
   U10561 : AOI22_X1 port map( A1 => n9947, A2 => n10117, B1 => n10120, B2 => 
                           n9679, ZN => n9558);
   U10562 : AOI22_X1 port map( A1 => n10114, A2 => n10430, B1 => n10110, B2 => 
                           n9948, ZN => n9559);
   U10563 : OAI22_X1 port map( A1 => n7810, A2 => n10038, B1 => n9922, B2 => 
                           n10046, ZN => n9561);
   U10564 : OAI22_X1 port map( A1 => n10061, A2 => n10066, B1 => n10057, B2 => 
                           n10104, ZN => n9562);
   U10565 : OAI211_X1 port map( C1 => n9554, C2 => n9553, A => n9552, B => 
                           n9551, ZN => n9555);
   U10566 : OAI211_X1 port map( C1 => n9550, C2 => n7806, A => n10103, B => 
                           n9549, ZN => n9551);
   U10567 : OR2_X1 port map( A1 => n9380, A2 => n11879, ZN => n9549);
   U10568 : INV_X1 port map( A => n9379, ZN => n9550);
   U10569 : AOI22_X1 port map( A1 => n9762, A2 => n9548, B1 => n9547, B2 => 
                           n7805, ZN => n9552);
   U10570 : NAND2_X1 port map( A1 => n9022, A2 => n9021, ZN => n9548);
   U10571 : NAND2_X1 port map( A1 => n7805, A2 => n11851, ZN => n9021);
   U10572 : NAND2_X1 port map( A1 => n9060, A2 => n11861, ZN => n9022);
   U10573 : INV_X1 port map( A => n9546, ZN => n9553);
   U10574 : OAI21_X1 port map( B1 => n9545, B2 => n9544, A => n9543, ZN => 
                           n9556);
   U10575 : NAND2_X1 port map( A1 => n9542, A2 => n8438, ZN => n9543);
   U10576 : NOR2_X1 port map( A1 => n9529, A2 => n9567, ZN => n9565);
   U10577 : NAND2_X1 port map( A1 => n9527, A2 => n9571, ZN => n9569);
   U10578 : NOR2_X1 port map( A1 => n10425, A2 => n9933, ZN => n9571);
   U10579 : OAI222_X1 port map( A1 => n8204, A2 => n7757, B1 => n11845, B2 => 
                           n8679, C1 => n8314, C2 => n10367, ZN => n7051);
   U10580 : OAI222_X1 port map( A1 => n8207, A2 => n7757, B1 => n11845, B2 => 
                           n11840, C1 => n8312, C2 => n10367, ZN => n7050);
   U10581 : OAI222_X1 port map( A1 => n8206, A2 => n7757, B1 => n11845, B2 => 
                           n8686, C1 => n8311, C2 => n10367, ZN => n7049);
   U10582 : OAI222_X1 port map( A1 => n8328, A2 => n11884, B1 => n11880, B2 => 
                           n9956, C1 => n11881, C2 => n9955, ZN => n6998);
   U10583 : NOR3_X1 port map( A1 => n9954, A2 => n9953, A3 => n9952, ZN => 
                           n9955);
   U10584 : OAI22_X1 port map( A1 => n7810, A2 => n10002, B1 => n9969, B2 => 
                           n10038, ZN => n9952);
   U10585 : INV_X1 port map( A => n9679, ZN => n9969);
   U10586 : OAI22_X1 port map( A1 => n10061, A2 => n10104, B1 => n9951, B2 => 
                           n10106, ZN => n9953);
   U10587 : OAI211_X1 port map( C1 => n9545, C2 => n9764, A => n9538, B => 
                           n9537, ZN => n9539);
   U10588 : AOI22_X1 port map( A1 => n9762, A2 => n9536, B1 => n9535, B2 => 
                           n9730, ZN => n9537);
   U10589 : INV_X1 port map( A => n9534, ZN => n9535);
   U10590 : INV_X1 port map( A => n9533, ZN => n9536);
   U10591 : OAI21_X1 port map( B1 => n9532, B2 => n9531, A => n9530, ZN => 
                           n9538);
   U10592 : AOI21_X1 port map( B1 => n9757, B2 => n11879, A => n9759, ZN => 
                           n9530);
   U10593 : NOR2_X1 port map( A1 => n9756, A2 => n9554, ZN => n9540);
   U10594 : OAI211_X1 port map( C1 => n9968, C2 => n10066, A => n9950, B => 
                           n9949, ZN => n9954);
   U10595 : AOI22_X1 port map( A1 => n10114, A2 => n10117, B1 => n10116, B2 => 
                           n9948, ZN => n9949);
   U10596 : AOI22_X1 port map( A1 => n9967, A2 => n10120, B1 => n10110, B2 => 
                           n9947, ZN => n9950);
   U10597 : INV_X1 port map( A => n9922, ZN => n9967);
   U10598 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_57_port, B2 =>
                           n10094, A => n9946, ZN => n9956);
   U10599 : OAI21_X1 port map( B1 => n9945, B2 => n9944, A => n9943, ZN => 
                           n9946);
   U10600 : AOI21_X1 port map( B1 => n9942, B2 => n9941, A => n9940, ZN => 
                           n9943);
   U10601 : OAI211_X1 port map( C1 => n9939, C2 => n10036, A => n9938, B => 
                           n9937, ZN => n9940);
   U10602 : INV_X1 port map( A => n10082, ZN => n10033);
   U10603 : XNOR2_X1 port map( A => n7817, B => n9936, ZN => n9939);
   U10604 : OAI21_X1 port map( B1 => n9933, B2 => n9932, A => n9931, ZN => 
                           n9941);
   U10605 : XNOR2_X1 port map( A => n9932, B => n10425, ZN => n9944);
   U10606 : AND2_X1 port map( A1 => C620_DATA2_23, A2 => n10443, ZN => 
                           DRAMRF_ADDRESS_23_port);
   U10607 : AOI22_X1 port map( A1 => n8930, A2 => n8194, B1 => 
                           IRAM_ADDRESS_14_port, B2 => n10417, ZN => n11841);
   U10608 : XNOR2_X1 port map( A => n8931, B => n8279, ZN => n8929);
   U10609 : AOI22_X1 port map( A1 => n10418, A2 => i_RD1_15_port, B1 => 
                           IRAM_ADDRESS_15_port, B2 => n10417, ZN => n11843);
   U10610 : NAND2_X1 port map( A1 => n8936, A2 => n10235, ZN => n8937);
   U10611 : INV_X1 port map( A => n10236, ZN => n8936);
   U10612 : OAI22_X1 port map( A1 => n9526, A2 => n11885, B1 => n511, B2 => 
                           n11884, ZN => n6997);
   U10613 : AOI211_X1 port map( C1 => DataPath_ALUhw_i_Q_EXTENDED_58_port, C2 
                           => n10094, A => n9525, B => n9524, ZN => n9526);
   U10614 : OAI211_X1 port map( C1 => n9523, C2 => n9748, A => n9522, B => 
                           n9521, ZN => n9524);
   U10615 : OAI211_X1 port map( C1 => n9517, C2 => n9516, A => n9942, B => 
                           n9515, ZN => n9522);
   U10616 : INV_X1 port map( A => n9570, ZN => n9942);
   U10617 : NOR3_X1 port map( A1 => n9514, A2 => n9513, A3 => n9512, ZN => 
                           n9523);
   U10618 : OAI211_X1 port map( C1 => n9968, C2 => n10104, A => n9511, B => 
                           n9510, ZN => n9512);
   U10619 : AOI22_X1 port map( A1 => n9947, A2 => n10116, B1 => n10121, B2 => 
                           n9679, ZN => n9510);
   U10620 : AOI22_X1 port map( A1 => n10114, A2 => n10110, B1 => n10430, B2 => 
                           n10111, ZN => n9511);
   U10621 : NOR2_X1 port map( A1 => n9509, A2 => n9508, ZN => n9968);
   U10622 : NOR3_X1 port map( A1 => n9726, A2 => n9732, A3 => n9627, ZN => 
                           n9508);
   U10623 : NOR2_X1 port map( A1 => n9507, A2 => n7806, ZN => n9732);
   U10624 : NOR2_X1 port map( A1 => n9506, A2 => n9531, ZN => n9726);
   U10625 : OAI211_X1 port map( C1 => n9505, C2 => n9504, A => n9503, B => 
                           n9502, ZN => n9509);
   U10626 : OAI211_X1 port map( C1 => n11879, C2 => n9501, A => n10103, B => 
                           n9500, ZN => n9502);
   U10627 : NAND2_X1 port map( A1 => n9499, A2 => n9531, ZN => n9500);
   U10628 : AOI21_X1 port map( B1 => n9704, B2 => n9498, A => n9497, ZN => 
                           n9503);
   U10629 : OAI22_X1 port map( A1 => n9496, A2 => n9495, B1 => n9494, B2 => 
                           n10098, ZN => n9497);
   U10630 : OAI22_X1 port map( A1 => n9951, A2 => n10056, B1 => n9592, B2 => 
                           n10059, ZN => n9513);
   U10631 : OAI22_X1 port map( A1 => n7810, A2 => n10066, B1 => n9922, B2 => 
                           n10038, ZN => n9514);
   U10632 : NOR2_X1 port map( A1 => n9945, A2 => n9493, ZN => n9525);
   U10633 : XNOR2_X1 port map( A => n9492, B => n9491, ZN => n9493);
   U10634 : INV_X1 port map( A => n9527, ZN => n9945);
   U10635 : NAND2_X1 port map( A1 => n10343, A2 => n10342, ZN => n7045);
   U10636 : AOI22_X1 port map( A1 => n10418, A2 => i_RD1_16_port, B1 => 
                           IRAM_ADDRESS_16_port, B2 => n10417, ZN => n10342);
   U10637 : OAI222_X1 port map( A1 => n11885, A2 => n9490, B1 => n11881, B2 => 
                           n9489, C1 => n11884, C2 => n512, ZN => n6996);
   U10638 : NOR3_X1 port map( A1 => n9488, A2 => n9487, A3 => n9486, ZN => 
                           n9489);
   U10639 : OAI211_X1 port map( C1 => n9592, C2 => n10038, A => n9485, B => 
                           n9484, ZN => n9486);
   U10640 : AOI22_X1 port map( A1 => n9947, A2 => n10120, B1 => n10113, B2 => 
                           n9679, ZN => n9484);
   U10641 : INV_X1 port map( A => n10105, ZN => n9947);
   U10642 : AOI22_X1 port map( A1 => n10114, A2 => n10116, B1 => n10117, B2 => 
                           n10111, ZN => n9485);
   U10643 : INV_X1 port map( A => n9948, ZN => n9592);
   U10644 : OAI22_X1 port map( A1 => n9951, A2 => n9977, B1 => n9483, B2 => 
                           n10106, ZN => n9487);
   U10645 : INV_X1 port map( A => n10119, ZN => n9483);
   U10646 : INV_X1 port map( A => n10122, ZN => n9951);
   U10647 : OAI22_X1 port map( A1 => n7810, A2 => n10104, B1 => n9922, B2 => 
                           n10002, ZN => n9488);
   U10648 : OAI22_X1 port map( A1 => n9545, A2 => n9478, B1 => n9477, B2 => 
                           n10098, ZN => n9479);
   U10649 : INV_X1 port map( A => n9702, ZN => n9478);
   U10650 : OAI22_X1 port map( A1 => n9554, A2 => n9476, B1 => n9475, B2 => 
                           n9755, ZN => n9480);
   U10651 : INV_X1 port map( A => n9474, ZN => n9475);
   U10652 : INV_X1 port map( A => n9705, ZN => n9476);
   U10653 : INV_X1 port map( A => n9586, ZN => n9554);
   U10654 : OAI22_X1 port map( A1 => n9473, A2 => n9505, B1 => n9496, B2 => 
                           n7776, ZN => n9481);
   U10655 : AOI21_X1 port map( B1 => n9472, B2 => n11879, A => n9471, ZN => 
                           n9482);
   U10656 : AOI21_X1 port map( B1 => n10103, B2 => n9470, A => n9469, ZN => 
                           n9471);
   U10657 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_59_port, B2 =>
                           n10094, A => n9468, ZN => n9490);
   U10658 : OAI211_X1 port map( C1 => n9467, C2 => n9570, A => n9466, B => 
                           n9465, ZN => n9468);
   U10659 : AOI211_X1 port map( C1 => n10088, C2 => n9464, A => n9463, B => 
                           n9462, ZN => n9465);
   U10660 : NOR3_X1 port map( A1 => n10084, A2 => n9461, A3 => n9473, ZN => 
                           n9462);
   U10661 : NOR3_X1 port map( A1 => n10082, A2 => n7804, A3 => 
                           DP_OP_751_130_6421_n507, ZN => n9463);
   U10662 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n507, B => n9473, ZN => 
                           n9464);
   U10663 : NAND2_X1 port map( A1 => n9527, A2 => n9460, ZN => n9466);
   U10664 : XNOR2_X1 port map( A => n9459, B => n9458, ZN => n9460);
   U10665 : OAI21_X1 port map( B1 => n9492, B2 => n9491, A => n9457, ZN => 
                           n9459);
   U10666 : AOI21_X1 port map( B1 => n9932, B2 => n10425, A => n11876, ZN => 
                           n9492);
   U10667 : NOR2_X1 port map( A1 => n11875, A2 => n11878, ZN => n9527);
   U10668 : NAND2_X1 port map( A1 => n11875, A2 => n9780, ZN => n9570);
   U10669 : NAND2_X1 port map( A1 => n9515, A2 => n9457, ZN => n9456);
   U10670 : NAND2_X1 port map( A1 => n9517, A2 => n9516, ZN => n9515);
   U10671 : INV_X1 port map( A => n9491, ZN => n9516);
   U10672 : NAND2_X1 port map( A1 => n9457, A2 => n9455, ZN => n9491);
   U10673 : INV_X1 port map( A => n9454, ZN => n9517);
   U10674 : NAND2_X1 port map( A1 => n9453, A2 => n9452, ZN => n9458);
   U10675 : OAI222_X1 port map( A1 => n11845, A2 => n10302, B1 => n10367, B2 =>
                           n7611, C1 => n7757, C2 => n10301, ZN => n7037);
   U10676 : XNOR2_X1 port map( A => n10298, B => n7611, ZN => n10299);
   U10677 : OAI21_X1 port map( B1 => n10340, B2 => n8370, A => n8369, ZN => 
                           n10300);
   U10678 : INV_X1 port map( A => i_RD1_24_port, ZN => n10302);
   U10679 : OAI21_X1 port map( B1 => n10297, B2 => n7757, A => n10296, ZN => 
                           n7036);
   U10680 : AOI22_X1 port map( A1 => n10418, A2 => i_RD1_25_port, B1 => 
                           IRAM_ADDRESS_25_port, B2 => n10417, ZN => n10296);
   U10681 : XNOR2_X1 port map( A => n10295, B => n10294, ZN => n10297);
   U10682 : XNOR2_X1 port map( A => n10293, B => IRAM_ADDRESS_25_port, ZN => 
                           n10294);
   U10683 : OAI21_X1 port map( B1 => n10338, B2 => n7757, A => n10337, ZN => 
                           n7044);
   U10684 : AOI22_X1 port map( A1 => n10418, A2 => i_RD1_17_port, B1 => 
                           IRAM_ADDRESS_17_port, B2 => n10417, ZN => n10337);
   U10685 : OAI21_X1 port map( B1 => n10323, B2 => n7757, A => n10322, ZN => 
                           n7041);
   U10686 : AOI22_X1 port map( A1 => n10418, A2 => i_RD1_20_port, B1 => 
                           IRAM_ADDRESS_20_port, B2 => n10417, ZN => n10322);
   U10687 : OAI21_X1 port map( B1 => n10339, B2 => n8202, A => n10252, ZN => 
                           n10321);
   U10688 : OAI22_X1 port map( A1 => n9451, A2 => n11885, B1 => n513, B2 => 
                           n11884, ZN => n6995);
   U10689 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_60_port, B2 =>
                           n10094, A => n9450, ZN => n9451);
   U10690 : OAI21_X1 port map( B1 => n9449, B2 => n9660, A => n9448, ZN => 
                           n9450);
   U10691 : AOI211_X1 port map( C1 => n9897, C2 => n9447, A => n9446, B => 
                           n9445, ZN => n9448);
   U10692 : AOI21_X1 port map( B1 => n9444, B2 => n9443, A => n9442, ZN => 
                           n9445);
   U10693 : NAND2_X1 port map( A1 => n10078, A2 => n9440, ZN => n9444);
   U10694 : AOI21_X1 port map( B1 => n9908, B2 => n9910, A => n10091, ZN => 
                           n9446);
   U10695 : NAND4_X1 port map( A1 => n9439, A2 => n9438, A3 => n9437, A4 => 
                           n9436, ZN => n9447);
   U10696 : AOI22_X1 port map( A1 => n10111, A2 => n10110, B1 => n9948, B2 => 
                           n10121, ZN => n9436);
   U10697 : AOI22_X1 port map( A1 => n10115, A2 => n10430, B1 => n10117, B2 => 
                           n10119, ZN => n9437);
   U10698 : AOI22_X1 port map( A1 => n10122, A2 => n10116, B1 => n10045, B2 => 
                           n9679, ZN => n9438);
   U10699 : NAND4_X1 port map( A1 => n9435, A2 => n9434, A3 => n9433, A4 => 
                           n9432, ZN => n9679);
   U10700 : NAND2_X1 port map( A1 => n9586, A2 => n9431, ZN => n9432);
   U10701 : INV_X1 port map( A => n10099, ZN => n9627);
   U10702 : OAI211_X1 port map( C1 => n11879, C2 => n9430, A => n10103, B => 
                           n9429, ZN => n9433);
   U10703 : NAND2_X1 port map( A1 => n9656, A2 => n9531, ZN => n9429);
   U10704 : AOI22_X1 port map( A1 => n9428, A2 => n7788, B1 => n9730, B2 => 
                           n9427, ZN => n9434);
   U10705 : INV_X1 port map( A => n7982, ZN => n9730);
   U10706 : AOI22_X1 port map( A1 => n9664, A2 => n9762, B1 => n9426, B2 => 
                           n7789, ZN => n9435);
   U10707 : AOI21_X1 port map( B1 => n9214, B2 => n11860, A => n9213, ZN => 
                           n9664);
   U10708 : NOR2_X1 port map( A1 => n7875, A2 => n11860, ZN => n9213);
   U10709 : AOI21_X1 port map( B1 => n10120, B2 => n10114, A => n9425, ZN => 
                           n9439);
   U10710 : OAI22_X1 port map( A1 => n9922, A2 => n10066, B1 => n10105, B2 => 
                           n10038, ZN => n9425);
   U10711 : AOI21_X1 port map( B1 => n10078, B2 => n9414, A => n9413, ZN => 
                           n9449);
   U10712 : OAI222_X1 port map( A1 => n11845, A2 => n10333, B1 => n7757, B2 => 
                           n10332, C1 => n8322, C2 => n10367, ZN => n7043);
   U10713 : NAND2_X1 port map( A1 => n10328, A2 => n10327, ZN => n10331);
   U10714 : INV_X1 port map( A => n10326, ZN => n10328);
   U10715 : OAI222_X1 port map( A1 => n11845, A2 => n10292, B1 => n10367, B2 =>
                           n8323, C1 => n7757, C2 => n10291, ZN => n7035);
   U10716 : NAND2_X1 port map( A1 => n10288, A2 => n10287, ZN => n10290);
   U10717 : OAI21_X1 port map( B1 => n9930, B2 => n11880, A => n9929, ZN => 
                           n6994);
   U10718 : AOI22_X1 port map( A1 => n9928, A2 => n10428, B1 => n7791, B2 => 
                           DRAM_ADDRESS_29_port, ZN => n9929);
   U10719 : NAND4_X1 port map( A1 => n9927, A2 => n9926, A3 => n9925, A4 => 
                           n9924, ZN => n9928);
   U10720 : AOI22_X1 port map( A1 => n10111, A2 => n10116, B1 => n9948, B2 => 
                           n10113, ZN => n9924);
   U10721 : AOI22_X1 port map( A1 => n10115, A2 => n10117, B1 => n10110, B2 => 
                           n10119, ZN => n9925);
   U10722 : AOI22_X1 port map( A1 => n10120, A2 => n10122, B1 => n10109, B2 => 
                           n10430, ZN => n9926);
   U10723 : AOI21_X1 port map( B1 => n10112, B2 => n10114, A => n9923, ZN => 
                           n9927);
   U10724 : OAI22_X1 port map( A1 => n9922, A2 => n10104, B1 => n10105, B2 => 
                           n10002, ZN => n9923);
   U10725 : OAI211_X1 port map( C1 => n9670, C2 => n9545, A => n9421, B => 
                           n9420, ZN => n9422);
   U10726 : OAI211_X1 port map( C1 => n9531, C2 => n9419, A => n10103, B => 
                           n9418, ZN => n9420);
   U10727 : NAND2_X1 port map( A1 => n9674, A2 => n11879, ZN => n9418);
   U10728 : NAND2_X1 port map( A1 => n9417, A2 => n7788, ZN => n9421);
   U10729 : NAND2_X1 port map( A1 => n7788, A2 => n11879, ZN => n9545);
   U10730 : OAI22_X1 port map( A1 => n10098, A2 => n9416, B1 => n9415, B2 => 
                           n7982, ZN => n9423);
   U10731 : AOI21_X1 port map( B1 => n11861, B2 => n7827, A => n8954, ZN => 
                           n9416);
   U10732 : INV_X1 port map( A => n8953, ZN => n8954);
   U10733 : NAND2_X1 port map( A1 => n10429, A2 => n9748, ZN => n11880);
   U10734 : AOI21_X1 port map( B1 => DataPath_ALUhw_i_Q_EXTENDED_61_port, B2 =>
                           n10094, A => n9921, ZN => n9930);
   U10735 : OAI211_X1 port map( C1 => n9920, C2 => n10091, A => n9919, B => 
                           n9918, ZN => n9921);
   U10736 : AOI211_X1 port map( C1 => n10088, C2 => n9917, A => n9916, B => 
                           n9915, ZN => n9918);
   U10737 : NOR3_X1 port map( A1 => n10084, A2 => n9914, A3 => n9913, ZN => 
                           n9915);
   U10738 : NOR3_X1 port map( A1 => n10082, A2 => n9912, A3 => n7821, ZN => 
                           n9916);
   U10739 : XNOR2_X1 port map( A => n7821, B => n9913, ZN => n9917);
   U10740 : NAND2_X1 port map( A1 => n10078, A2 => n9911, ZN => n9919);
   U10741 : AOI21_X1 port map( B1 => n9909, B2 => n9908, A => n9907, ZN => 
                           n9920);
   U10742 : OAI21_X1 port map( B1 => n10286, B2 => n7757, A => n10285, ZN => 
                           n7034);
   U10743 : AOI22_X1 port map( A1 => n10418, A2 => i_RD1_27_port, B1 => 
                           IRAM_ADDRESS_27_port, B2 => n10417, ZN => n10285);
   U10744 : OAI211_X1 port map( C1 => n9411, C2 => n10091, A => n9410, B => 
                           n9409, ZN => n9412);
   U10745 : NAND2_X1 port map( A1 => n10078, A2 => n9408, ZN => n9409);
   U10746 : XNOR2_X1 port map( A => n10075, B => n10074, ZN => n9408);
   U10747 : AOI211_X1 port map( C1 => n9405, C2 => n9897, A => n9404, B => 
                           n9403, ZN => n9410);
   U10748 : OAI22_X1 port map( A1 => n10084, A2 => n9402, B1 => n10082, B2 => 
                           n9401, ZN => n9403);
   U10749 : INV_X1 port map( A => n9400, ZN => n9401);
   U10750 : INV_X1 port map( A => n9399, ZN => n9402);
   U10751 : NOR3_X1 port map( A1 => n9399, A2 => n10036, A3 => n9400, ZN => 
                           n9404);
   U10752 : NOR2_X1 port map( A1 => n9398, A2 => n10070, ZN => n9400);
   U10753 : NOR2_X1 port map( A1 => n9397, A2 => n9619, ZN => n9399);
   U10754 : INV_X1 port map( A => n9398, ZN => n9397);
   U10755 : NAND4_X1 port map( A1 => n9396, A2 => n9395, A3 => n9394, A4 => 
                           n9393, ZN => n9405);
   U10756 : AOI22_X1 port map( A1 => n10114, A2 => n10121, B1 => n10120, B2 => 
                           n10111, ZN => n9393);
   U10757 : AOI22_X1 port map( A1 => n10118, A2 => n10430, B1 => n10110, B2 => 
                           n10115, ZN => n9394);
   U10758 : AOI22_X1 port map( A1 => n10122, A2 => n10112, B1 => n10116, B2 => 
                           n10119, ZN => n9395);
   U10759 : AOI21_X1 port map( B1 => n10045, B2 => n9948, A => n9346, ZN => 
                           n9396);
   U10760 : OAI22_X1 port map( A1 => n9345, A2 => n10056, B1 => n10105, B2 => 
                           n10066, ZN => n9346);
   U10761 : INV_X1 port map( A => n10109, ZN => n9345);
   U10762 : NAND4_X1 port map( A1 => n9338, A2 => n9337, A3 => n9336, A4 => 
                           n9335, ZN => n9948);
   U10763 : NAND2_X1 port map( A1 => n9365, A2 => n7789, ZN => n9335);
   U10764 : AOI22_X1 port map( A1 => n9547, A2 => n10070, B1 => n9762, B2 => 
                           n9332, ZN => n9336);
   U10765 : NAND2_X1 port map( A1 => n9027, A2 => n9031, ZN => n9332);
   U10766 : NAND2_X1 port map( A1 => n9240, A2 => n11861, ZN => n9027);
   U10767 : NOR2_X1 port map( A1 => n9331, A2 => n9330, ZN => n9337);
   U10768 : NOR2_X1 port map( A1 => n9728, A2 => n9333, ZN => n9330);
   U10769 : OAI21_X1 port map( B1 => n9496, B2 => n7714, A => n9329, ZN => 
                           n9331);
   U10770 : NAND2_X1 port map( A1 => n9624, A2 => n9328, ZN => n9338);
   U10771 : AND2_X1 port map( A1 => n9621, A2 => n7788, ZN => n9328);
   U10772 : NAND2_X1 port map( A1 => n9362, A2 => n9531, ZN => n9621);
   U10773 : OR2_X1 port map( A1 => n9364, A2 => n9531, ZN => n9624);
   U10774 : XNOR2_X1 port map( A => n10072, B => n10071, ZN => n9411);
   U10775 : OAI21_X1 port map( B1 => n10309, B2 => n7757, A => n10308, ZN => 
                           n7038);
   U10776 : AOI22_X1 port map( A1 => n10418, A2 => i_RD1_23_port, B1 => 
                           IRAM_ADDRESS_23_port, B2 => n10417, ZN => n10308);
   U10777 : XNOR2_X1 port map( A => n10307, B => n10306, ZN => n10309);
   U10778 : XNOR2_X1 port map( A => n10305, B => IRAM_ADDRESS_23_port, ZN => 
                           n10306);
   U10779 : OAI21_X1 port map( B1 => n10313, B2 => n10312, A => n10311, ZN => 
                           n10307);
   U10780 : INV_X1 port map( A => n10304, ZN => n10312);
   U10781 : INV_X1 port map( A => n10303, ZN => n10315);
   U10782 : NAND2_X1 port map( A1 => n8384, A2 => n7603, ZN => n10317);
   U10783 : NAND2_X1 port map( A1 => n10339, A2 => n8390, ZN => n8384);
   U10784 : NAND2_X1 port map( A1 => n10340, A2 => n10341, ZN => n10339);
   U10785 : AND4_X1 port map( A1 => n10126, A2 => n10125, A3 => n10124, A4 => 
                           n10123, ZN => n10127);
   U10786 : AOI22_X1 port map( A1 => n10122, A2 => n10121, B1 => n10120, B2 => 
                           n10119, ZN => n10123);
   U10787 : NAND4_X1 port map( A1 => n9361, A2 => n9360, A3 => n9359, A4 => 
                           n9358, ZN => n10119);
   U10788 : NAND2_X1 port map( A1 => n9357, A2 => n8434, ZN => n9358);
   U10789 : INV_X1 port map( A => n9376, ZN => n9357);
   U10790 : AOI22_X1 port map( A1 => n9469, A2 => n10431, B1 => n9762, B2 => 
                           n9702, ZN => n9359);
   U10791 : NOR2_X1 port map( A1 => i_ALU_OP_2_port, A2 => n9473, ZN => n10431)
                           ;
   U10792 : AOI22_X1 port map( A1 => n10103, A2 => n9705, B1 => n9474, B2 => 
                           n7788, ZN => n9360);
   U10793 : OAI21_X1 port map( B1 => n11869, B2 => n9472, A => n9356, ZN => 
                           n9474);
   U10794 : AOI21_X1 port map( B1 => n8566, B2 => n7828, A => n8994, ZN => 
                           n9472);
   U10795 : NOR2_X1 port map( A1 => n8566, A2 => n7776, ZN => n8994);
   U10796 : OAI21_X1 port map( B1 => n11873, B2 => n9355, A => n9356, ZN => 
                           n9705);
   U10797 : NAND2_X1 port map( A1 => n9470, A2 => n11874, ZN => n9356);
   U10798 : NAND2_X1 port map( A1 => n9179, A2 => n8995, ZN => n9355);
   U10799 : NAND2_X1 port map( A1 => n8566, A2 => n7776, ZN => n8995);
   U10800 : OR2_X1 port map( A1 => n7828, A2 => i_ALU_OP_2_port, ZN => n9179);
   U10801 : AOI22_X1 port map( A1 => n9387, A2 => n7804, B1 => n9389, B2 => 
                           n9470, ZN => n9361);
   U10802 : NAND2_X1 port map( A1 => n7804, A2 => n11851, ZN => n8996);
   U10803 : NAND2_X1 port map( A1 => n7897, A2 => n11868, ZN => n8997);
   U10804 : INV_X1 port map( A => n7974, ZN => n9169);
   U10805 : OAI211_X1 port map( C1 => n9756, C2 => n9759, A => n9354, B => 
                           n9353, ZN => n10122);
   U10806 : AOI21_X1 port map( B1 => n9936, B2 => n9387, A => n9352, ZN => 
                           n9353);
   U10807 : OAI22_X1 port map( A1 => n9765, A2 => n9534, B1 => n10098, B2 => 
                           n9764, ZN => n9352);
   U10808 : AOI21_X1 port map( B1 => n9936, B2 => n7809, A => n9351, ZN => 
                           n9534);
   U10809 : AOI22_X1 port map( A1 => n9389, A2 => n9532, B1 => n9541, B2 => 
                           n7788, ZN => n9354);
   U10810 : OAI21_X1 port map( B1 => n11869, B2 => n9757, A => n9350, ZN => 
                           n9541);
   U10811 : INV_X1 port map( A => n9349, ZN => n9350);
   U10812 : AOI21_X1 port map( B1 => n8566, B2 => n7824, A => n9010, ZN => 
                           n9757);
   U10813 : NOR2_X1 port map( A1 => i_ALU_OP_2_port, A2 => n8405, ZN => n9010);
   U10814 : INV_X1 port map( A => n9347, ZN => n9532);
   U10815 : AOI21_X1 port map( B1 => n11868, B2 => n9348, A => n9349, ZN => 
                           n9756);
   U10816 : NOR2_X1 port map( A1 => n9347, A2 => n11867, ZN => n9349);
   U10817 : NAND2_X1 port map( A1 => n9936, A2 => n11851, ZN => n9011);
   U10818 : AND2_X1 port map( A1 => n7924, A2 => i_ALU_OP_2_port, ZN => n9351);
   U10819 : AOI22_X1 port map( A1 => n10118, A2 => n10117, B1 => n10116, B2 => 
                           n10115, ZN => n10124);
   U10820 : OAI211_X1 port map( C1 => n9666, C2 => n9759, A => n9375, B => 
                           n9374, ZN => n10115);
   U10821 : AOI22_X1 port map( A1 => n9387, A2 => n9442, B1 => n7788, B2 => 
                           n9426, ZN => n9374);
   U10822 : OAI21_X1 port map( B1 => n9821, B2 => n7809, A => n8966, ZN => 
                           n9656);
   U10823 : NAND2_X1 port map( A1 => n7809, A2 => n7799, ZN => n8966);
   U10824 : AOI21_X1 port map( B1 => n9389, B2 => n9430, A => n9372, ZN => 
                           n9375);
   U10825 : OAI22_X1 port map( A1 => n9765, A2 => n9371, B1 => n7985, B2 => 
                           n7440, ZN => n9372);
   U10826 : INV_X1 port map( A => n9427, ZN => n9371);
   U10827 : OAI21_X1 port map( B1 => n7809, B2 => n7799, A => n8972, ZN => 
                           n9427);
   U10828 : NAND2_X1 port map( A1 => n8188, A2 => n9442, ZN => n8972);
   U10829 : INV_X1 port map( A => n9431, ZN => n9666);
   U10830 : OAI21_X1 port map( B1 => n9659, B2 => n11873, A => n9373, ZN => 
                           n9431);
   U10831 : NAND2_X1 port map( A1 => n9430, A2 => n11874, ZN => n9373);
   U10832 : INV_X1 port map( A => n9214, ZN => n9430);
   U10833 : NOR2_X1 port map( A1 => n9660, A2 => n11849, ZN => n8969);
   U10834 : NAND2_X1 port map( A1 => n9369, A2 => n8967, ZN => n9659);
   U10835 : NAND2_X1 port map( A1 => n7799, A2 => i_ALU_OP_2_port, ZN => n8967)
                           ;
   U10836 : NAND2_X1 port map( A1 => n9822, A2 => n7809, ZN => n9369);
   U10837 : NAND2_X1 port map( A1 => n9146, A2 => n8020, ZN => n9052);
   U10838 : OAI211_X1 port map( C1 => n9383, C2 => n9619, A => n9368, B => 
                           n9367, ZN => n10118);
   U10839 : AOI22_X1 port map( A1 => n9389, A2 => n9366, B1 => n7788, B2 => 
                           n9365, ZN => n9367);
   U10840 : OAI21_X1 port map( B1 => n7893, B2 => n7809, A => n9029, ZN => 
                           n9333);
   U10841 : NAND2_X1 port map( A1 => n7809, A2 => n7714, ZN => n9029);
   U10842 : AOI21_X1 port map( B1 => n10103, B2 => n9364, A => n9363, ZN => 
                           n9368);
   U10843 : OAI22_X1 port map( A1 => n9376, A2 => n7714, B1 => n10098, B2 => 
                           n9362, ZN => n9363);
   U10844 : OAI21_X1 port map( B1 => n9327, B2 => n11873, A => n9334, ZN => 
                           n9364);
   U10845 : NAND2_X1 port map( A1 => n9366, A2 => n11874, ZN => n9334);
   U10846 : NAND2_X1 port map( A1 => n10070, A2 => n11851, ZN => n9031);
   U10847 : NAND2_X1 port map( A1 => n9240, A2 => n11868, ZN => n9032);
   U10848 : NAND2_X1 port map( A1 => n9220, A2 => n9033, ZN => n9327);
   U10849 : NAND2_X1 port map( A1 => n7773, A2 => n8566, ZN => n9033);
   U10850 : NAND2_X1 port map( A1 => n7981, A2 => n7809, ZN => n9220);
   U10851 : AOI22_X1 port map( A1 => n10114, A2 => n10113, B1 => n10112, B2 => 
                           n10111, ZN => n10125);
   U10852 : OAI211_X1 port map( C1 => n9392, C2 => n9759, A => n9391, B => 
                           n9390, ZN => n10111);
   U10853 : AOI22_X1 port map( A1 => n9389, A2 => n9501, B1 => n9498, B2 => 
                           n7788, ZN => n9390);
   U10854 : OAI21_X1 port map( B1 => n11869, B2 => n9499, A => n9388, ZN => 
                           n9498);
   U10855 : OAI21_X1 port map( B1 => n9871, B2 => n7809, A => n8979, ZN => 
                           n9499);
   U10856 : NAND2_X1 port map( A1 => n7809, A2 => n9495, ZN => n8979);
   U10857 : AOI22_X1 port map( A1 => n9387, A2 => n9727, B1 => n9762, B2 => 
                           n9507, ZN => n9391);
   U10858 : AOI21_X1 port map( B1 => n9386, B2 => n9385, A => n9506, ZN => 
                           n9392);
   U10859 : OAI21_X1 port map( B1 => n9384, B2 => n11873, A => n9388, ZN => 
                           n9506);
   U10860 : NAND2_X1 port map( A1 => n9501, A2 => n11874, ZN => n9388);
   U10861 : NAND2_X1 port map( A1 => n9727, A2 => n11851, ZN => n8982);
   U10862 : NAND2_X1 port map( A1 => n7913, A2 => n11868, ZN => n8983);
   U10863 : NAND2_X1 port map( A1 => n9157, A2 => n9385, ZN => n9384);
   U10864 : NAND2_X1 port map( A1 => n9122, A2 => n7809, ZN => n9157);
   U10865 : NAND2_X1 port map( A1 => n8566, A2 => n9495, ZN => n9385);
   U10866 : AOI21_X1 port map( B1 => n7809, B2 => n9504, A => n7806, ZN => 
                           n9386);
   U10867 : NAND4_X1 port map( A1 => n9025, A2 => n9053, A3 => n8988, A4 => 
                           n8020, ZN => n10038);
   U10868 : NAND2_X1 port map( A1 => n9019, A2 => n9128, ZN => n10066);
   U10869 : NOR2_X1 port map( A1 => n9146, A2 => n7726, ZN => n9019);
   U10870 : OAI211_X1 port map( C1 => n9383, C2 => n9528, A => n9382, B => 
                           n9381, ZN => n10114);
   U10871 : AOI22_X1 port map( A1 => n9389, A2 => n9380, B1 => n7788, B2 => 
                           n9557, ZN => n9381);
   U10872 : OAI21_X1 port map( B1 => n9379, B2 => n11869, A => n9378, ZN => 
                           n9557);
   U10873 : OAI21_X1 port map( B1 => n9279, B2 => n7809, A => n9020, ZN => 
                           n9379);
   U10874 : NAND2_X1 port map( A1 => n7809, A2 => n8439, ZN => n9020);
   U10875 : AOI21_X1 port map( B1 => n10103, B2 => n9546, A => n9377, ZN => 
                           n9382);
   U10876 : OAI22_X1 port map( A1 => n9376, A2 => n8439, B1 => n10098, B2 => 
                           n9544, ZN => n9377);
   U10877 : NAND2_X1 port map( A1 => n9055, A2 => n9054, ZN => n9544);
   U10878 : OR2_X1 port map( A1 => n9060, A2 => n8188, ZN => n9054);
   U10879 : NAND2_X1 port map( A1 => n9469, A2 => n8566, ZN => n9376);
   U10880 : OAI21_X1 port map( B1 => n9264, B2 => n11873, A => n9378, ZN => 
                           n9546);
   U10881 : NAND2_X1 port map( A1 => n9380, A2 => n11874, ZN => n9378);
   U10882 : NAND2_X1 port map( A1 => n9057, A2 => n9056, ZN => n9380);
   U10883 : NAND2_X1 port map( A1 => n9060, A2 => n11868, ZN => n9057);
   U10884 : NAND2_X1 port map( A1 => n9055, A2 => n9023, ZN => n9264);
   U10885 : NAND2_X1 port map( A1 => i_ALU_OP_2_port, A2 => n8439, ZN => n9023)
                           ;
   U10886 : NAND2_X1 port map( A1 => n8435, A2 => n7809, ZN => n9055);
   U10887 : AOI21_X1 port map( B1 => n9469, B2 => n7809, A => n9387, ZN => 
                           n9383);
   U10888 : INV_X1 port map( A => n9728, ZN => n9469);
   U10889 : AOI21_X1 port map( B1 => n10110, B2 => n10109, A => n10108, ZN => 
                           n10126);
   U10890 : OAI22_X1 port map( A1 => n10107, A2 => n10106, B1 => n10105, B2 => 
                           n10104, ZN => n10108);
   U10891 : OR2_X1 port map( A1 => n7974, A2 => n8020, ZN => n9024);
   U10892 : NAND2_X1 port map( A1 => n10097, A2 => n9531, ZN => n9584);
   U10893 : OR2_X1 port map( A1 => n9759, A2 => n7806, ZN => n9728);
   U10894 : NAND2_X1 port map( A1 => n9049, A2 => n9048, ZN => n9583);
   U10895 : NAND2_X1 port map( A1 => n10081, A2 => n11851, ZN => n9048);
   U10896 : NAND2_X1 port map( A1 => n7898, A2 => n11861, ZN => n9049);
   U10897 : INV_X1 port map( A => n10098, ZN => n9762);
   U10898 : NOR2_X1 port map( A1 => n9759, A2 => n11879, ZN => n9657);
   U10899 : OR2_X1 port map( A1 => n7998, A2 => n8020, ZN => n9058);
   U10900 : AOI211_X1 port map( C1 => n10103, C2 => n11882, A => n10102, B => 
                           n10101, ZN => n10107);
   U10901 : AND2_X1 port map( A1 => n10100, A2 => n7788, ZN => n10101);
   U10902 : NAND2_X1 port map( A1 => n9344, A2 => n9343, ZN => n10100);
   U10903 : NAND2_X1 port map( A1 => n9582, A2 => n11870, ZN => n9343);
   U10904 : NAND2_X1 port map( A1 => n9044, A2 => n9043, ZN => n9582);
   U10905 : NAND2_X1 port map( A1 => n7809, A2 => n9602, ZN => n9043);
   U10906 : NAND2_X1 port map( A1 => n7983, A2 => i_ALU_OP_2_port, ZN => n9044)
                           ;
   U10907 : OAI22_X1 port map( A1 => n10098, A2 => n10097, B1 => n7982, B2 => 
                           n10095, ZN => n10102);
   U10908 : OR2_X1 port map( A1 => n7898, A2 => n8188, ZN => n9242);
   U10909 : NAND2_X1 port map( A1 => n9284, A2 => n9344, ZN => n11882);
   U10910 : NAND2_X1 port map( A1 => n9585, A2 => n11874, ZN => n9344);
   U10911 : NAND2_X1 port map( A1 => n9051, A2 => n9050, ZN => n9585);
   U10912 : AOI21_X1 port map( B1 => n10081, B2 => n11851, A => n11850, ZN => 
                           n9050);
   U10913 : NAND2_X1 port map( A1 => n7898, A2 => n11868, ZN => n9051);
   U10914 : AOI22_X1 port map( A1 => n11868, A2 => n9283, B1 => n9282, B2 => 
                           n9531, ZN => n9284);
   U10915 : OAI21_X1 port map( B1 => n9600, B2 => n7809, A => n11883, ZN => 
                           n9282);
   U10916 : OAI211_X1 port map( C1 => n9667, C2 => n9759, A => n9342, B => 
                           n9341, ZN => n10109);
   U10917 : AOI22_X1 port map( A1 => n9387, A2 => n9912, B1 => n7788, B2 => 
                           n9424, ZN => n9341);
   U10918 : OAI21_X1 port map( B1 => n11869, B2 => n9674, A => n9340, ZN => 
                           n9424);
   U10919 : OAI21_X1 port map( B1 => n10034, B2 => n7809, A => n8946, ZN => 
                           n9674);
   U10920 : NAND2_X1 port map( A1 => n8188, A2 => n9961, ZN => n8946);
   U10921 : OAI21_X1 port map( B1 => n11873, B2 => n7985, A => n9496, ZN => 
                           n9387);
   U10922 : INV_X1 port map( A => n9542, ZN => n9496);
   U10923 : NOR2_X1 port map( A1 => n7982, A2 => n7809, ZN => n9542);
   U10924 : AOI21_X1 port map( B1 => n9389, B2 => n9419, A => n9339, ZN => 
                           n9342);
   U10925 : OAI22_X1 port map( A1 => n9765, A2 => n9415, B1 => n10098, B2 => 
                           n9670, ZN => n9339);
   U10926 : OR2_X1 port map( A1 => n7985, A2 => n7806, ZN => n10098);
   U10927 : NAND2_X1 port map( A1 => n10103, A2 => n11879, ZN => n9765);
   U10928 : NAND2_X1 port map( A1 => n9505, A2 => n11867, ZN => n9389);
   U10929 : INV_X1 port map( A => n9547, ZN => n9505);
   U10930 : NOR2_X1 port map( A1 => n7982, A2 => n8566, ZN => n9547);
   U10931 : INV_X1 port map( A => n10103, ZN => n9759);
   U10932 : INV_X1 port map( A => n9417, ZN => n9667);
   U10933 : OAI21_X1 port map( B1 => n9668, B2 => n11873, A => n9340, ZN => 
                           n9417);
   U10934 : NAND2_X1 port map( A1 => n9419, A2 => n11874, ZN => n9340);
   U10935 : NAND2_X1 port map( A1 => n9912, A2 => n11851, ZN => n8953);
   U10936 : INV_X1 port map( A => n11850, ZN => n9056);
   U10937 : NAND2_X1 port map( A1 => n7827, A2 => n11868, ZN => n8948);
   U10938 : NAND2_X1 port map( A1 => n9229, A2 => n8952, ZN => n9668);
   U10939 : NAND2_X1 port map( A1 => i_ALU_OP_2_port, A2 => n9961, ZN => n8952)
                           ;
   U10940 : NAND2_X1 port map( A1 => n8427, A2 => n7809, ZN => n9229);
   U10941 : OAI211_X1 port map( C1 => n10092, C2 => n10091, A => n10090, B => 
                           n10089, ZN => n10093);
   U10942 : AOI211_X1 port map( C1 => n10088, C2 => n10087, A => n10086, B => 
                           n10085, ZN => n10089);
   U10943 : NOR3_X1 port map( A1 => n10084, A2 => n10083, A3 => n10095, ZN => 
                           n10085);
   U10944 : NOR3_X1 port map( A1 => n10082, A2 => n10081, A3 => n7816, ZN => 
                           n10086);
   U10945 : NAND2_X1 port map( A1 => n9127, A2 => n8566, ZN => n10082);
   U10946 : NOR2_X1 port map( A1 => n9125, A2 => i_ALU_OP_0_port, ZN => n9127);
   U10947 : NAND2_X1 port map( A1 => i_ALU_OP_1_port, A2 => n11852, ZN => n9125
                           );
   U10948 : XNOR2_X1 port map( A => n8566, B => i_ALU_OP_4_port, ZN => n9126);
   U10949 : OAI211_X1 port map( C1 => n10080, C2 => n10079, A => n10078, B => 
                           n10077, ZN => n10090);
   U10950 : NAND2_X1 port map( A1 => n10079, A2 => n10076, ZN => n10077);
   U10951 : NOR2_X1 port map( A1 => n9406, A2 => n11878, ZN => n10078);
   U10952 : NOR2_X1 port map( A1 => n10075, A2 => n10074, ZN => n10079);
   U10953 : OAI22_X1 port map( A1 => n9909, A2 => n9910, B1 => n9407, B2 => 
                           n9913, ZN => n10075);
   U10954 : NAND2_X1 port map( A1 => n9440, A2 => n9442, ZN => n9910);
   U10955 : NAND2_X1 port map( A1 => n9406, A2 => n9780, ZN => n10091);
   U10956 : NAND2_X1 port map( A1 => n9326, A2 => n9453, ZN => n9406);
   U10957 : NAND2_X1 port map( A1 => n9325, A2 => n7804, ZN => n9453);
   U10958 : INV_X1 port map( A => n9324, ZN => n9325);
   U10959 : NAND2_X1 port map( A1 => n9324, A2 => n9473, ZN => n9452);
   U10960 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n507, B => n8566, ZN => 
                           n9324);
   U10961 : NAND2_X1 port map( A1 => n9322, A2 => n9504, ZN => n9455);
   U10962 : INV_X1 port map( A => n9321, ZN => n9322);
   U10963 : OAI21_X1 port map( B1 => n9454, B2 => n11877, A => n9457, ZN => 
                           n9323);
   U10964 : NAND2_X1 port map( A1 => n9321, A2 => n9727, ZN => n9457);
   U10965 : XNOR2_X1 port map( A => n9518, B => n8188, ZN => n9321);
   U10966 : OAI21_X1 port map( B1 => n9316, B2 => n9600, A => n9315, ZN => 
                           n11875);
   U10967 : OAI22_X1 port map( A1 => n9314, A2 => n11872, B1 => n9602, B2 => 
                           n9579, ZN => n9315);
   U10968 : AOI21_X1 port map( B1 => n9577, B2 => n9575, A => n9634, ZN => 
                           n9314);
   U10969 : NAND2_X1 port map( A1 => n9636, A2 => n9635, ZN => n9634);
   U10970 : XNOR2_X1 port map( A => n11871, B => n7606, ZN => n9635);
   U10971 : XNOR2_X1 port map( A => n9637, B => n8566, ZN => n11871);
   U10972 : NOR2_X1 port map( A1 => n9963, A2 => n9574, ZN => n9636);
   U10973 : INV_X1 port map( A => n9313, ZN => n9574);
   U10974 : NOR2_X1 port map( A1 => n9965, A2 => n9957, ZN => n9963);
   U10975 : NAND2_X1 port map( A1 => n9647, A2 => n7799, ZN => n9957);
   U10976 : NAND2_X1 port map( A1 => n9313, A2 => n9311, ZN => n9965);
   U10977 : NAND2_X1 port map( A1 => n9310, A2 => n9961, ZN => n9313);
   U10978 : AND2_X1 port map( A1 => n9959, A2 => n9311, ZN => n9575);
   U10979 : NAND2_X1 port map( A1 => n9309, A2 => n9962, ZN => n9311);
   U10980 : INV_X1 port map( A => n9310, ZN => n9309);
   U10981 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n813, B => 
                           i_ALU_OP_2_port, ZN => n9310);
   U10982 : NAND2_X1 port map( A1 => n9308, A2 => n8433, ZN => n9959);
   U10983 : INV_X1 port map( A => n9647, ZN => n9308);
   U10984 : XNOR2_X1 port map( A => n9651, B => i_ALU_OP_2_port, ZN => n9647);
   U10985 : AOI21_X1 port map( B1 => n9307, B2 => n9687, A => n9306, ZN => 
                           n9577);
   U10986 : NOR2_X1 port map( A1 => n9305, A2 => n7776, ZN => n9306);
   U10987 : AOI21_X1 port map( B1 => n9719, B2 => n9688, A => n9689, ZN => 
                           n9687);
   U10988 : XNOR2_X1 port map( A => n9305, B => n7776, ZN => n9689);
   U10989 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n915, B => n8566, ZN => 
                           n9305);
   U10990 : OR2_X1 port map( A1 => n9722, A2 => n9723, ZN => n9719);
   U10991 : INV_X1 port map( A => n9742, ZN => n9723);
   U10992 : NAND2_X1 port map( A1 => n10049, A2 => n9304, ZN => n9722);
   U10993 : NAND2_X1 port map( A1 => n9303, A2 => n8405, ZN => n9304);
   U10994 : NAND2_X1 port map( A1 => n10050, A2 => n10051, ZN => n10049);
   U10995 : NAND2_X1 port map( A1 => n9686, A2 => n9685, ZN => n9307);
   U10996 : AND2_X1 port map( A1 => n9739, A2 => n9688, ZN => n9685);
   U10997 : NAND2_X1 port map( A1 => n9301, A2 => n7777, ZN => n9688);
   U10998 : NAND2_X1 port map( A1 => n9741, A2 => n9742, ZN => n9739);
   U10999 : XNOR2_X1 port map( A => n9301, B => n9495, ZN => n9742);
   U11000 : XNOR2_X1 port map( A => n9743, B => n8188, ZN => n9301);
   U11001 : NAND2_X1 port map( A1 => n10050, A2 => n10048, ZN => n10047);
   U11002 : AND2_X1 port map( A1 => n9302, A2 => n8438, ZN => n10048);
   U11003 : XNOR2_X1 port map( A => n9754, B => n8188, ZN => n9302);
   U11004 : XNOR2_X1 port map( A => n9303, B => n7924, ZN => n10050);
   U11005 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1017, B => 
                           i_ALU_OP_2_port, ZN => n9303);
   U11006 : AOI21_X1 port map( B1 => n9300, B2 => n9299, A => n9777, ZN => 
                           n9686);
   U11007 : AND2_X1 port map( A1 => n9772, A2 => n9776, ZN => n9299);
   U11008 : NAND2_X1 port map( A1 => n9298, A2 => n7727, ZN => n9776);
   U11009 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1119, B => 
                           i_ALU_OP_2_port, ZN => n9298);
   U11010 : NAND2_X1 port map( A1 => n9297, A2 => n7981, ZN => n9772);
   U11011 : INV_X1 port map( A => n9296, ZN => n9297);
   U11012 : OAI21_X1 port map( B1 => n9781, B2 => n10030, A => n9775, ZN => 
                           n9300);
   U11013 : AND2_X1 port map( A1 => n9802, A2 => n9773, ZN => n9775);
   U11014 : NAND2_X1 port map( A1 => n9296, A2 => n7893, ZN => n9773);
   U11015 : XNOR2_X1 port map( A => n9807, B => n8188, ZN => n9296);
   U11016 : NAND2_X1 port map( A1 => n10026, A2 => n9769, ZN => n9802);
   U11017 : OR2_X1 port map( A1 => n10028, A2 => n10027, ZN => n10026);
   U11018 : AND2_X1 port map( A1 => n9295, A2 => n9821, ZN => n10027);
   U11019 : OR2_X1 port map( A1 => n10028, A2 => n10029, ZN => n10030);
   U11020 : XNOR2_X1 port map( A => n9823, B => n8188, ZN => n9295);
   U11021 : NAND2_X1 port map( A1 => n9769, A2 => n9770, ZN => n10028);
   U11022 : NAND2_X1 port map( A1 => n9294, A2 => n10034, ZN => n9770);
   U11023 : INV_X1 port map( A => n10032, ZN => n10034);
   U11024 : INV_X1 port map( A => n9293, ZN => n9294);
   U11025 : NAND2_X1 port map( A1 => n9293, A2 => n10032, ZN => n9769);
   U11026 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1221, B => 
                           i_ALU_OP_2_port, ZN => n9293);
   U11027 : AOI21_X1 port map( B1 => n9842, B2 => n9838, A => n9839, ZN => 
                           n9781);
   U11028 : AND2_X1 port map( A1 => n9292, A2 => n9843, ZN => n9839);
   U11029 : NAND2_X1 port map( A1 => n9291, A2 => n8401, ZN => n9838);
   U11030 : INV_X1 port map( A => n9292, ZN => n9291);
   U11031 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1323, B => n8188, ZN =>
                           n9292);
   U11032 : AOI21_X1 port map( B1 => n9861, B2 => n9290, A => n9289, ZN => 
                           n9842);
   U11033 : NOR2_X1 port map( A1 => n9859, A2 => n9871, ZN => n9289);
   U11034 : NAND2_X1 port map( A1 => n9859, A2 => n9871, ZN => n9290);
   U11035 : INV_X1 port map( A => n9122, ZN => n9871);
   U11036 : XNOR2_X1 port map( A => n9872, B => n8188, ZN => n9859);
   U11037 : AOI21_X1 port map( B1 => n9288, B2 => n10011, A => n10012, ZN => 
                           n9861);
   U11038 : AND2_X1 port map( A1 => n9287, A2 => n7824, ZN => n10012);
   U11039 : NAND2_X1 port map( A1 => n9286, A2 => n10017, ZN => n10011);
   U11040 : INV_X1 port map( A => n9287, ZN => n9286);
   U11041 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1425, B => n8188, ZN =>
                           n9287);
   U11042 : OAI21_X1 port map( B1 => n10010, B2 => n10008, A => n10009, ZN => 
                           n9288);
   U11043 : NAND2_X1 port map( A1 => n9274, A2 => n9279, ZN => n10009);
   U11044 : INV_X1 port map( A => n8435, ZN => n9279);
   U11045 : INV_X1 port map( A => n9285, ZN => n9274);
   U11046 : AND2_X1 port map( A1 => n9285, A2 => n8436, ZN => n10008);
   U11047 : XNOR2_X1 port map( A => n9271, B => i_ALU_OP_2_port, ZN => n9285);
   U11048 : AOI21_X1 port map( B1 => n9261, B2 => n9260, A => n9259, ZN => 
                           n10010);
   U11049 : AND2_X1 port map( A1 => n9258, A2 => n9257, ZN => n9260);
   U11050 : NAND2_X1 port map( A1 => n9186, A2 => n8400, ZN => n9257);
   U11051 : INV_X1 port map( A => n9187, ZN => n9186);
   U11052 : NAND2_X1 port map( A1 => n9249, A2 => n9248, ZN => n9258);
   U11053 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1527, B => 
                           i_ALU_OP_2_port, ZN => n9249);
   U11054 : OAI21_X1 port map( B1 => n9256, B2 => n9255, A => n9254, ZN => 
                           n9261);
   U11055 : NOR2_X1 port map( A1 => n9251, A2 => n9250, ZN => n9254);
   U11056 : AND2_X1 port map( A1 => n9187, A2 => n9240, ZN => n9250);
   U11057 : XNOR2_X1 port map( A => n9241, B => i_ALU_OP_2_port, ZN => n9187);
   U11058 : OAI21_X1 port map( B1 => n9983, B2 => n9981, A => n9207, ZN => 
                           n9251);
   U11059 : NAND2_X1 port map( A1 => n9895, A2 => n7875, ZN => n9981);
   U11060 : NAND2_X1 port map( A1 => n9207, A2 => n9206, ZN => n9983);
   U11061 : NAND2_X1 port map( A1 => n9190, A2 => n7827, ZN => n9207);
   U11062 : NAND2_X1 port map( A1 => n9982, A2 => n9206, ZN => n9255);
   U11063 : NAND2_X1 port map( A1 => n9189, A2 => n9986, ZN => n9206);
   U11064 : INV_X1 port map( A => n9190, ZN => n9189);
   U11065 : XNOR2_X1 port map( A => n7775, B => n7809, ZN => n9190);
   U11066 : NAND2_X1 port map( A1 => n9880, A2 => n9188, ZN => n9982);
   U11067 : INV_X1 port map( A => n9895, ZN => n9880);
   U11068 : XNOR2_X1 port map( A => n8021, B => i_ALU_OP_2_port, ZN => n9895);
   U11069 : NAND2_X1 port map( A1 => n9205, A2 => n9204, ZN => n9256);
   U11070 : NAND2_X1 port map( A1 => n9203, A2 => n8398, ZN => n9204);
   U11071 : INV_X1 port map( A => n9201, ZN => n9203);
   U11072 : NAND2_X1 port map( A1 => n9146, A2 => n7913, ZN => n9198);
   U11073 : NAND2_X1 port map( A1 => n9201, A2 => n7897, ZN => n9199);
   U11074 : XNOR2_X1 port map( A => n8146, B => n8188, ZN => n9201);
   U11075 : OAI211_X1 port map( C1 => n9196, C2 => n9195, A => n9194, B => 
                           n9193, ZN => n9200);
   U11076 : NAND2_X1 port map( A1 => n9128, A2 => n9133, ZN => n9193);
   U11077 : NAND2_X1 port map( A1 => n9145, A2 => n9168, ZN => n9194);
   U11078 : INV_X1 port map( A => n9146, ZN => n9145);
   U11079 : NAND2_X1 port map( A1 => n9053, A2 => n8961, ZN => n9146);
   U11080 : NAND2_X1 port map( A1 => n7974, A2 => n7809, ZN => n8961);
   U11081 : OR2_X1 port map( A1 => n7974, A2 => n8188, ZN => n9053);
   U11082 : OR2_X1 port map( A1 => DataPath_ALUhw_MULT_mux_out_0_0_port, A2 => 
                           n9192, ZN => n9195);
   U11083 : NOR2_X1 port map( A1 => n8020, A2 => n7809, ZN => n9192);
   U11084 : NOR2_X1 port map( A1 => n9128, A2 => n9133, ZN => n9196);
   U11085 : NAND2_X1 port map( A1 => n9025, A2 => n9018, ZN => n9128);
   U11086 : NAND2_X1 port map( A1 => n7998, A2 => i_ALU_OP_2_port, ZN => n9018)
                           ;
   U11087 : OR2_X1 port map( A1 => n7998, A2 => i_ALU_OP_2_port, ZN => n9025);
   U11088 : INV_X1 port map( A => n9579, ZN => n9316);
   U11089 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n711, B => n7809, ZN => 
                           n9579);
   U11090 : NOR2_X1 port map( A1 => n9318, A2 => n9528, ZN => n10425);
   U11091 : NAND2_X1 port map( A1 => n9931, A2 => n9320, ZN => n9454);
   U11092 : INV_X1 port map( A => n9319, ZN => n9320);
   U11093 : NAND2_X1 port map( A1 => n9932, A2 => n9933, ZN => n9931);
   U11094 : AND2_X1 port map( A1 => n9318, A2 => n9528, ZN => n9933);
   U11095 : XNOR2_X1 port map( A => n9567, B => n8566, ZN => n9318);
   U11096 : NOR2_X1 port map( A1 => n11876, A2 => n9319, ZN => n9932);
   U11097 : AND2_X1 port map( A1 => n9317, A2 => n9936, ZN => n11876);
   U11098 : XNOR2_X1 port map( A => n7817, B => n8188, ZN => n9317);
   U11099 : INV_X1 port map( A => n10080, ZN => n10092);
   U11100 : AOI22_X1 port map( A1 => n10072, A2 => n10071, B1 => n10070, B2 => 
                           n10069, ZN => n10073);
   U11101 : INV_X1 port map( A => n10074, ZN => n10071);
   U11102 : XNOR2_X1 port map( A => n10069, B => n10070, ZN => n10074);
   U11103 : XNOR2_X1 port map( A => n9398, B => n8188, ZN => n10069);
   U11104 : AOI21_X1 port map( B1 => n9407, B2 => n9913, A => n9907, ZN => 
                           n10072);
   U11105 : NOR2_X1 port map( A1 => n9909, A2 => n9908, ZN => n9907);
   U11106 : NAND2_X1 port map( A1 => n9414, A2 => n9660, ZN => n9908);
   U11107 : INV_X1 port map( A => n9440, ZN => n9414);
   U11108 : XNOR2_X1 port map( A => n9441, B => n8188, ZN => n9440);
   U11109 : XNOR2_X1 port map( A => n9407, B => n9913, ZN => n9909);
   U11110 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n405, B => n8566, ZN => 
                           n9407);
   U11111 : XNOR2_X1 port map( A => n10068, B => n7816, ZN => n10076);
   U11112 : OAI21_X1 port map( B1 => n10081, B2 => n7809, A => n11883, ZN => 
                           n10068);
   U11113 : NAND2_X1 port map( A1 => n8188, A2 => n10081, ZN => n11883);
   U11114 : NOR2_X1 port map( A1 => n8457, A2 => n9130, ZN => 
                           DataPath_ALUhw_MULT_mux_out_10_20_port);
   U11115 : OAI22_X1 port map( A1 => n9094, A2 => n9130, B1 => n9133, B2 => 
                           n9095, ZN => DataPath_ALUhw_MULT_mux_out_9_19_port);
   U11116 : OAI22_X1 port map( A1 => n7785, A2 => n9130, B1 => n9133, B2 => 
                           n9086, ZN => DataPath_ALUhw_MULT_mux_out_7_15_port);
   U11117 : NOR2_X1 port map( A1 => n7790, A2 => n9130, ZN => 
                           DataPath_ALUhw_MULT_mux_out_8_16_port);
   U11118 : AND2_X1 port map( A1 => n8020, A2 => n9060, ZN => 
                           DataPath_ALUhw_MULT_mux_out_0_0_port);
   U11119 : OAI22_X1 port map( A1 => n8442, A2 => n9130, B1 => n9133, B2 => 
                           n8430, ZN => DataPath_ALUhw_MULT_mux_out_1_3_port);
   U11120 : OAI22_X1 port map( A1 => n8445, A2 => n9130, B1 => n9133, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_5_port);
   U11121 : OAI22_X1 port map( A1 => n7756, A2 => n8398, B1 => n7726, B2 => 
                           n9188, ZN => DataPath_ALUhw_MULT_mux_out_0_4_port);
   U11122 : NOR2_X1 port map( A1 => n8450, A2 => n9130, ZN => 
                           DataPath_ALUhw_MULT_mux_out_3_6_port);
   U11123 : OAI22_X1 port map( A1 => n7615, A2 => n9130, B1 => n9133, B2 => 
                           n8449, ZN => DataPath_ALUhw_MULT_mux_out_3_7_port);
   U11124 : OAI22_X1 port map( A1 => n8444, A2 => n9133, B1 => n9168, B2 => 
                           n8447, ZN => DataPath_ALUhw_MULT_mux_out_2_6_port);
   U11125 : OAI22_X1 port map( A1 => n7750, A2 => n9188, B1 => n7726, B2 => 
                           n9986, ZN => DataPath_ALUhw_MULT_mux_out_0_5_port);
   U11126 : OAI22_X1 port map( A1 => n8442, A2 => n9168, B1 => n8399, B2 => 
                           n8429, ZN => DataPath_ALUhw_MULT_mux_out_1_5_port);
   U11127 : OAI22_X1 port map( A1 => n8453, A2 => n9130, B1 => n9133, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_9_port);
   U11128 : OAI22_X1 port map( A1 => n7616, A2 => n9133, B1 => n9168, B2 => 
                           n8449, ZN => DataPath_ALUhw_MULT_mux_out_3_8_port);
   U11129 : OAI22_X1 port map( A1 => n8444, A2 => n9168, B1 => n8399, B2 => 
                           n8447, ZN => DataPath_ALUhw_MULT_mux_out_2_7_port);
   U11130 : OAI22_X1 port map( A1 => n7769, A2 => n9130, B1 => n8454, B2 => 
                           n9133, ZN => DataPath_ALUhw_MULT_mux_out_5_11_port);
   U11131 : OAI22_X1 port map( A1 => n8452, A2 => n9133, B1 => n9168, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_10_port);
   U11132 : OAI22_X1 port map( A1 => n7616, A2 => n9168, B1 => n8399, B2 => 
                           n8450, ZN => DataPath_ALUhw_MULT_mux_out_3_9_port);
   U11133 : OAI22_X1 port map( A1 => n8443, A2 => n8398, B1 => n9188, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_8_port);
   U11134 : NOR2_X1 port map( A1 => n8455, A2 => n9130, ZN => 
                           DataPath_ALUhw_MULT_mux_out_6_12_port);
   U11135 : OAI22_X1 port map( A1 => n9080, A2 => n9133, B1 => n9081, B2 => 
                           n9168, ZN => DataPath_ALUhw_MULT_mux_out_6_14_port);
   U11136 : OAI22_X1 port map( A1 => n7787, A2 => n9168, B1 => n8454, B2 => 
                           n8399, ZN => DataPath_ALUhw_MULT_mux_out_5_13_port);
   U11137 : OAI22_X1 port map( A1 => n9080, A2 => n9130, B1 => n8455, B2 => 
                           n9133, ZN => DataPath_ALUhw_MULT_mux_out_6_13_port);
   U11138 : OAI22_X1 port map( A1 => n9074, A2 => n8398, B1 => n9188, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_12_port);
   U11139 : OAI22_X1 port map( A1 => n7787, A2 => n9133, B1 => n8454, B2 => 
                           n9168, ZN => DataPath_ALUhw_MULT_mux_out_5_12_port);
   U11140 : OAI22_X1 port map( A1 => n7615, A2 => n9188, B1 => n9986, B2 => 
                           n9070, ZN => DataPath_ALUhw_MULT_mux_out_3_11_port);
   U11141 : OAI22_X1 port map( A1 => n8453, A2 => n9168, B1 => n8399, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_11_port);
   U11142 : OAI22_X1 port map( A1 => n8443, A2 => n9986, B1 => n7795, B2 => 
                           n8447, ZN => DataPath_ALUhw_MULT_mux_out_2_10_port);
   U11143 : OAI22_X1 port map( A1 => n7615, A2 => n8398, B1 => n9188, B2 => 
                           n8449, ZN => DataPath_ALUhw_MULT_mux_out_3_10_port);
   U11144 : OAI22_X1 port map( A1 => n7756, A2 => n8435, B1 => n8403, B2 => 
                           n7726, ZN => DataPath_ALUhw_MULT_mux_out_0_9_port);
   U11145 : OAI22_X1 port map( A1 => n8445, A2 => n9188, B1 => n9986, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_9_port);
   U11146 : OAI22_X1 port map( A1 => n7756, A2 => n9248, B1 => n7726, B2 => 
                           n7801, ZN => DataPath_ALUhw_MULT_mux_out_0_8_port);
   U11147 : OAI22_X1 port map( A1 => n8441, A2 => n9986, B1 => n9239, B2 => 
                           n8430, ZN => DataPath_ALUhw_MULT_mux_out_1_8_port);
   U11148 : NOR2_X1 port map( A1 => n8456, A2 => n9130, ZN => 
                           DataPath_ALUhw_MULT_mux_out_7_14_port);
   U11149 : OAI22_X1 port map( A1 => n7767, A2 => n9133, B1 => n9168, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_18_port);
   U11150 : OAI22_X1 port map( A1 => n7785, A2 => n9168, B1 => n8399, B2 => 
                           n9086, ZN => DataPath_ALUhw_MULT_mux_out_7_17_port);
   U11151 : OAI22_X1 port map( A1 => n9088, A2 => n9130, B1 => n9133, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_17_port);
   U11152 : OAI22_X1 port map( A1 => n9080, A2 => n8398, B1 => n9081, B2 => 
                           n9188, ZN => DataPath_ALUhw_MULT_mux_out_6_16_port);
   U11153 : OAI22_X1 port map( A1 => n7785, A2 => n9133, B1 => n9168, B2 => 
                           n8456, ZN => DataPath_ALUhw_MULT_mux_out_7_16_port);
   U11154 : OAI22_X1 port map( A1 => n7787, A2 => n9188, B1 => n9079, B2 => 
                           n9986, ZN => DataPath_ALUhw_MULT_mux_out_5_15_port);
   U11155 : OAI22_X1 port map( A1 => n7770, A2 => n9168, B1 => n9081, B2 => 
                           n8399, ZN => DataPath_ALUhw_MULT_mux_out_6_15_port);
   U11156 : OAI22_X1 port map( A1 => n9074, A2 => n9986, B1 => n7823, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_14_port);
   U11157 : OAI22_X1 port map( A1 => n7769, A2 => n8398, B1 => n9079, B2 => 
                           n9188, ZN => DataPath_ALUhw_MULT_mux_out_5_14_port);
   U11158 : OAI22_X1 port map( A1 => n7616, A2 => n7823, B1 => n9248, B2 => 
                           n8449, ZN => DataPath_ALUhw_MULT_mux_out_3_13_port);
   U11159 : OAI22_X1 port map( A1 => n8453, A2 => n9188, B1 => n9986, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_13_port);
   U11160 : OAI22_X1 port map( A1 => n8443, A2 => n9248, B1 => n8436, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_12_port);
   U11161 : OAI22_X1 port map( A1 => n7616, A2 => n9986, B1 => n7823, B2 => 
                           n8449, ZN => DataPath_ALUhw_MULT_mux_out_3_12_port);
   U11162 : OAI22_X1 port map( A1 => n8440, A2 => n8435, B1 => n8403, B2 => 
                           n8431, ZN => DataPath_ALUhw_MULT_mux_out_1_11_port);
   U11163 : OAI22_X1 port map( A1 => n8444, A2 => n8400, B1 => n9248, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_11_port);
   U11164 : OAI22_X1 port map( A1 => n9248, A2 => n7620, B1 => n8437, B2 => 
                           n8429, ZN => DataPath_ALUhw_MULT_mux_out_1_10_port);
   U11165 : OAI22_X1 port map( A1 => n9099, A2 => n9130, B1 => n9133, B2 => 
                           n8457, ZN => DataPath_ALUhw_MULT_mux_out_10_21_port)
                           ;
   U11166 : OAI22_X1 port map( A1 => n9094, A2 => n9133, B1 => n9168, B2 => 
                           n9095, ZN => DataPath_ALUhw_MULT_mux_out_9_20_port);
   U11167 : OAI22_X1 port map( A1 => n9088, A2 => n9168, B1 => n8399, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_19_port);
   U11168 : OAI22_X1 port map( A1 => n7785, A2 => n8398, B1 => n9188, B2 => 
                           n8456, ZN => DataPath_ALUhw_MULT_mux_out_7_18_port);
   U11169 : OAI22_X1 port map( A1 => n7770, A2 => n9188, B1 => n8455, B2 => 
                           n9986, ZN => DataPath_ALUhw_MULT_mux_out_6_17_port);
   U11170 : OAI22_X1 port map( A1 => n7787, A2 => n9986, B1 => n8454, B2 => 
                           n7823, ZN => DataPath_ALUhw_MULT_mux_out_5_16_port);
   U11171 : OAI22_X1 port map( A1 => n8453, A2 => n7823, B1 => n9248, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_15_port);
   U11172 : OAI22_X1 port map( A1 => n7616, A2 => n9248, B1 => n8437, B2 => 
                           n8449, ZN => DataPath_ALUhw_MULT_mux_out_3_14_port);
   U11173 : BUF_X1 port map( A => n8435, Z => n8437);
   U11174 : OAI22_X1 port map( A1 => n8445, A2 => n8435, B1 => n8403, B2 => 
                           n8447, ZN => DataPath_ALUhw_MULT_mux_out_2_13_port);
   U11175 : OAI22_X1 port map( A1 => n8134, A2 => n9844, B1 => n7726, B2 => 
                           n9822, ZN => DataPath_ALUhw_MULT_mux_out_0_12_port);
   U11176 : OAI22_X1 port map( A1 => n8441, A2 => n8404, B1 => n9122, B2 => 
                           n8429, ZN => DataPath_ALUhw_MULT_mux_out_1_12_port);
   U11177 : NOR2_X1 port map( A1 => n9105, A2 => n9130, ZN => 
                           DataPath_ALUhw_MULT_mux_out_11_22_port);
   U11178 : OAI22_X1 port map( A1 => n9104, A2 => n9130, B1 => n9133, B2 => 
                           n9105, ZN => DataPath_ALUhw_MULT_mux_out_11_23_port)
                           ;
   U11179 : OAI22_X1 port map( A1 => n9099, A2 => n9133, B1 => n9168, B2 => 
                           n9100, ZN => DataPath_ALUhw_MULT_mux_out_10_22_port)
                           ;
   U11180 : OAI22_X1 port map( A1 => n9094, A2 => n9168, B1 => n8399, B2 => 
                           n9095, ZN => DataPath_ALUhw_MULT_mux_out_9_21_port);
   U11181 : OAI22_X1 port map( A1 => n7767, A2 => n8399, B1 => n9188, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_20_port);
   U11182 : OAI22_X1 port map( A1 => n7785, A2 => n9188, B1 => n9986, B2 => 
                           n9086, ZN => DataPath_ALUhw_MULT_mux_out_7_19_port);
   U11183 : OAI22_X1 port map( A1 => n9080, A2 => n9986, B1 => n8455, B2 => 
                           n7823, ZN => DataPath_ALUhw_MULT_mux_out_6_18_port);
   U11184 : OAI22_X1 port map( A1 => n7769, A2 => n7823, B1 => n8454, B2 => 
                           n9248, ZN => DataPath_ALUhw_MULT_mux_out_5_17_port);
   U11185 : OAI22_X1 port map( A1 => n8453, A2 => n9248, B1 => n8436, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_16_port);
   U11186 : OAI22_X1 port map( A1 => n7615, A2 => n7801, B1 => n8403, B2 => 
                           n8449, ZN => DataPath_ALUhw_MULT_mux_out_3_15_port);
   U11187 : OAI22_X1 port map( A1 => n8445, A2 => n8404, B1 => n9122, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_14_port);
   U11188 : OAI22_X1 port map( A1 => n8442, A2 => n9122, B1 => n9844, B2 => 
                           n8429, ZN => DataPath_ALUhw_MULT_mux_out_1_13_port);
   U11189 : NOR2_X1 port map( A1 => n9110, A2 => n9130, ZN => 
                           DataPath_ALUhw_MULT_mux_out_12_24_port);
   U11190 : OAI22_X1 port map( A1 => n9109, A2 => n9130, B1 => n9133, B2 => 
                           n9110, ZN => DataPath_ALUhw_MULT_mux_out_12_25_port)
                           ;
   U11191 : OAI22_X1 port map( A1 => n9104, A2 => n9133, B1 => n9168, B2 => 
                           n9105, ZN => DataPath_ALUhw_MULT_mux_out_11_24_port)
                           ;
   U11192 : OAI22_X1 port map( A1 => n9099, A2 => n9168, B1 => n8399, B2 => 
                           n8457, ZN => DataPath_ALUhw_MULT_mux_out_10_23_port)
                           ;
   U11193 : OAI22_X1 port map( A1 => n9094, A2 => n8398, B1 => n9188, B2 => 
                           n9095, ZN => DataPath_ALUhw_MULT_mux_out_9_22_port);
   U11194 : OAI22_X1 port map( A1 => n7767, A2 => n9188, B1 => n9986, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_21_port);
   U11195 : OAI22_X1 port map( A1 => n9085, A2 => n9986, B1 => n7823, B2 => 
                           n8456, ZN => DataPath_ALUhw_MULT_mux_out_7_20_port);
   U11196 : OAI22_X1 port map( A1 => n9080, A2 => n7823, B1 => n8455, B2 => 
                           n9248, ZN => DataPath_ALUhw_MULT_mux_out_6_19_port);
   U11197 : OAI22_X1 port map( A1 => n7787, A2 => n9248, B1 => n8454, B2 => 
                           n8435, ZN => DataPath_ALUhw_MULT_mux_out_5_18_port);
   U11198 : OAI22_X1 port map( A1 => n8453, A2 => n7801, B1 => n8403, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_17_port);
   U11199 : OAI22_X1 port map( A1 => n7615, A2 => n8404, B1 => n9122, B2 => 
                           n8451, ZN => DataPath_ALUhw_MULT_mux_out_3_16_port);
   U11200 : OAI22_X1 port map( A1 => n8443, A2 => n7800, B1 => n9844, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_15_port);
   U11201 : OAI22_X1 port map( A1 => n8134, A2 => n10032, B1 => n7726, B2 => 
                           n7309, ZN => DataPath_ALUhw_MULT_mux_out_0_14_port);
   U11202 : OAI22_X1 port map( A1 => n8440, A2 => n9844, B1 => n9822, B2 => 
                           n7753, ZN => DataPath_ALUhw_MULT_mux_out_1_14_port);
   U11203 : NOR2_X1 port map( A1 => n9114, A2 => n9130, ZN => 
                           DataPath_ALUhw_MULT_mux_out_13_26_port);
   U11204 : OAI22_X1 port map( A1 => n9113, A2 => n9130, B1 => n9133, B2 => 
                           n9114, ZN => DataPath_ALUhw_MULT_mux_out_13_27_port)
                           ;
   U11205 : OAI22_X1 port map( A1 => n9109, A2 => n9133, B1 => n9168, B2 => 
                           n9110, ZN => DataPath_ALUhw_MULT_mux_out_12_26_port)
                           ;
   U11206 : OAI22_X1 port map( A1 => n9099, A2 => n8398, B1 => n9188, B2 => 
                           n8457, ZN => DataPath_ALUhw_MULT_mux_out_10_24_port)
                           ;
   U11207 : OAI22_X1 port map( A1 => n9094, A2 => n9188, B1 => n9986, B2 => 
                           n9095, ZN => DataPath_ALUhw_MULT_mux_out_9_23_port);
   U11208 : OAI22_X1 port map( A1 => n9088, A2 => n9986, B1 => n7795, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_22_port);
   U11209 : OAI22_X1 port map( A1 => n9085, A2 => n7823, B1 => n9248, B2 => 
                           n8456, ZN => DataPath_ALUhw_MULT_mux_out_7_21_port);
   U11210 : OAI22_X1 port map( A1 => n7770, A2 => n9248, B1 => n8455, B2 => 
                           n8436, ZN => DataPath_ALUhw_MULT_mux_out_6_20_port);
   U11211 : OAI22_X1 port map( A1 => n7787, A2 => n8435, B1 => n9079, B2 => 
                           n8403, ZN => DataPath_ALUhw_MULT_mux_out_5_19_port);
   U11212 : OAI22_X1 port map( A1 => n8452, A2 => n8404, B1 => n9122, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_18_port);
   U11213 : OAI22_X1 port map( A1 => n7615, A2 => n9122, B1 => n8401, B2 => 
                           n8450, ZN => DataPath_ALUhw_MULT_mux_out_3_17_port);
   U11214 : OAI22_X1 port map( A1 => n8444, A2 => n9844, B1 => n9822, B2 => 
                           n8447, ZN => DataPath_ALUhw_MULT_mux_out_2_16_port);
   U11215 : OAI22_X1 port map( A1 => n7619, A2 => n9822, B1 => n10032, B2 => 
                           n7753, ZN => DataPath_ALUhw_MULT_mux_out_1_15_port);
   U11216 : NOR2_X1 port map( A1 => n9118, A2 => n9130, ZN => 
                           DataPath_ALUhw_MULT_mux_out_14_28_port);
   U11217 : OAI22_X1 port map( A1 => n9117, A2 => n9130, B1 => n9133, B2 => 
                           n9118, ZN => DataPath_ALUhw_MULT_mux_out_14_29_port)
                           ;
   U11218 : OAI22_X1 port map( A1 => n9113, A2 => n9133, B1 => n9168, B2 => 
                           n9114, ZN => DataPath_ALUhw_MULT_mux_out_13_28_port)
                           ;
   U11219 : OAI22_X1 port map( A1 => n9109, A2 => n9168, B1 => n8399, B2 => 
                           n9110, ZN => DataPath_ALUhw_MULT_mux_out_12_27_port)
                           ;
   U11220 : OAI22_X1 port map( A1 => n9104, A2 => n8398, B1 => n9188, B2 => 
                           n9105, ZN => DataPath_ALUhw_MULT_mux_out_11_26_port)
                           ;
   U11221 : OAI22_X1 port map( A1 => n9099, A2 => n9188, B1 => n9986, B2 => 
                           n9100, ZN => DataPath_ALUhw_MULT_mux_out_10_25_port)
                           ;
   U11222 : OAI22_X1 port map( A1 => n9094, A2 => n9986, B1 => n8400, B2 => 
                           n9095, ZN => DataPath_ALUhw_MULT_mux_out_9_24_port);
   U11223 : OAI22_X1 port map( A1 => n7767, A2 => n7823, B1 => n9248, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_23_port);
   U11224 : OAI22_X1 port map( A1 => n9085, A2 => n9248, B1 => n8436, B2 => 
                           n8456, ZN => DataPath_ALUhw_MULT_mux_out_7_22_port);
   U11225 : OAI22_X1 port map( A1 => n7770, A2 => n8436, B1 => n8455, B2 => 
                           n8403, ZN => DataPath_ALUhw_MULT_mux_out_6_21_port);
   U11226 : OAI22_X1 port map( A1 => n7769, A2 => n8404, B1 => n8454, B2 => 
                           n9122, ZN => DataPath_ALUhw_MULT_mux_out_5_20_port);
   U11227 : OAI22_X1 port map( A1 => n8453, A2 => n9122, B1 => n8401, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_19_port);
   U11228 : OAI22_X1 port map( A1 => n7616, A2 => n8401, B1 => n9822, B2 => 
                           n8451, ZN => DataPath_ALUhw_MULT_mux_out_3_18_port);
   U11229 : OAI22_X1 port map( A1 => n8443, A2 => n9822, B1 => n8427, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_17_port);
   U11230 : OAI22_X1 port map( A1 => n7756, A2 => n9784, B1 => n7726, B2 => 
                           n9753, ZN => DataPath_ALUhw_MULT_mux_out_0_16_port);
   U11231 : OAI22_X1 port map( A1 => n8441, A2 => n10032, B1 => n7309, B2 => 
                           n8430, ZN => DataPath_ALUhw_MULT_mux_out_1_16_port);
   U11232 : NOR2_X1 port map( A1 => n9124, A2 => n9130, ZN => 
                           DataPath_ALUhw_MULT_mux_out_15_30_port);
   U11233 : OAI22_X1 port map( A1 => n8134, A2 => n9619, B1 => n7726, B2 => 
                           n10095, ZN => DataPath_ALUhw_MULT_mux_out_0_31_port)
                           ;
   U11234 : OAI22_X1 port map( A1 => n7620, A2 => n9660, B1 => n8431, B2 => 
                           n9913, ZN => DataPath_ALUhw_MULT_mux_out_1_31_port);
   U11235 : OAI22_X1 port map( A1 => n8445, A2 => n9504, B1 => n9473, B2 => 
                           n8447, ZN => DataPath_ALUhw_MULT_mux_out_2_31_port);
   U11236 : OAI22_X1 port map( A1 => n7616, A2 => n9528, B1 => n8451, B2 => 
                           n8402, ZN => DataPath_ALUhw_MULT_mux_out_3_31_port);
   U11237 : OAI22_X1 port map( A1 => n9074, A2 => n7773, B1 => n9600, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_31_port);
   U11238 : OAI22_X1 port map( A1 => n7787, A2 => n7799, B1 => n8454, B2 => 
                           n9961, ZN => DataPath_ALUhw_MULT_mux_out_5_31_port);
   U11239 : OAI22_X1 port map( A1 => n7770, A2 => n9495, B1 => n8455, B2 => 
                           n7776, ZN => DataPath_ALUhw_MULT_mux_out_6_31_port);
   U11240 : OAI22_X1 port map( A1 => n7785, A2 => n8439, B1 => n8406, B2 => 
                           n8456, ZN => DataPath_ALUhw_MULT_mux_out_7_31_port);
   U11241 : OAI22_X1 port map( A1 => n9088, A2 => n7981, B1 => n7727, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_31_port);
   U11242 : OAI22_X1 port map( A1 => n9094, A2 => n9822, B1 => n8428, B2 => 
                           n9095, ZN => DataPath_ALUhw_MULT_mux_out_9_31_port);
   U11243 : OAI22_X1 port map( A1 => n9099, A2 => n7800, B1 => n8401, B2 => 
                           n9100, ZN => DataPath_ALUhw_MULT_mux_out_10_31_port)
                           ;
   U11244 : OAI22_X1 port map( A1 => n9104, A2 => n8435, B1 => n8404, B2 => 
                           n9105, ZN => DataPath_ALUhw_MULT_mux_out_11_31_port)
                           ;
   U11245 : OAI22_X1 port map( A1 => n9109, A2 => n7795, B1 => n9248, B2 => 
                           n9110, ZN => DataPath_ALUhw_MULT_mux_out_12_31_port)
                           ;
   U11246 : OAI22_X1 port map( A1 => n9113, A2 => n9188, B1 => n9986, B2 => 
                           n9114, ZN => DataPath_ALUhw_MULT_mux_out_13_31_port)
                           ;
   U11247 : OAI22_X1 port map( A1 => n9117, A2 => n9168, B1 => n8399, B2 => 
                           n9118, ZN => DataPath_ALUhw_MULT_mux_out_14_31_port)
                           ;
   U11248 : OAI22_X1 port map( A1 => n9123, A2 => n9130, B1 => n9133, B2 => 
                           n9124, ZN => DataPath_ALUhw_MULT_mux_out_15_31_port)
                           ;
   U11249 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n405, B => n9398, ZN => 
                           n9124);
   U11250 : OAI21_X1 port map( B1 => n8298, B2 => n8137, A => n9120, ZN => 
                           n9398);
   U11251 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_30_port
                           , ZN => n9120);
   U11252 : INV_X1 port map( A => n7816, ZN => n10083);
   U11253 : OAI21_X1 port map( B1 => n8297, B2 => n8137, A => n9119, ZN => 
                           DP_OP_751_130_6421_n303);
   U11254 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_31_port
                           , ZN => n9119);
   U11255 : OAI22_X1 port map( A1 => n7620, A2 => n9473, B1 => n9660, B2 => 
                           n8432, ZN => DataPath_ALUhw_MULT_mux_out_1_30_port);
   U11256 : OAI22_X1 port map( A1 => n8443, A2 => n8402, B1 => n9504, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_30_port);
   U11257 : OAI22_X1 port map( A1 => n7615, A2 => n9600, B1 => n9070, B2 => 
                           n9528, ZN => DataPath_ALUhw_MULT_mux_out_3_30_port);
   U11258 : OAI22_X1 port map( A1 => n9074, A2 => n9961, B1 => n7773, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_30_port);
   U11259 : OAI22_X1 port map( A1 => n7769, A2 => n7776, B1 => n8454, B2 => 
                           n7799, ZN => DataPath_ALUhw_MULT_mux_out_5_30_port);
   U11260 : OAI22_X1 port map( A1 => n9080, A2 => n8405, B1 => n8455, B2 => 
                           n9495, ZN => DataPath_ALUhw_MULT_mux_out_6_30_port);
   U11261 : OAI22_X1 port map( A1 => n7785, A2 => n7727, B1 => n8439, B2 => 
                           n8456, ZN => DataPath_ALUhw_MULT_mux_out_7_30_port);
   U11262 : OAI22_X1 port map( A1 => n7767, A2 => n8427, B1 => n7981, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_30_port);
   U11263 : OAI22_X1 port map( A1 => n9094, A2 => n8401, B1 => n9822, B2 => 
                           n9095, ZN => DataPath_ALUhw_MULT_mux_out_9_30_port);
   U11264 : OAI22_X1 port map( A1 => n9099, A2 => n10017, B1 => n9122, B2 => 
                           n9100, ZN => DataPath_ALUhw_MULT_mux_out_10_30_port)
                           ;
   U11265 : OAI22_X1 port map( A1 => n9104, A2 => n9248, B1 => n8435, B2 => 
                           n9105, ZN => DataPath_ALUhw_MULT_mux_out_11_30_port)
                           ;
   U11266 : OAI22_X1 port map( A1 => n9109, A2 => n9986, B1 => n8400, B2 => 
                           n9110, ZN => DataPath_ALUhw_MULT_mux_out_12_30_port)
                           ;
   U11267 : OAI22_X1 port map( A1 => n9113, A2 => n8398, B1 => n9188, B2 => 
                           n9114, ZN => DataPath_ALUhw_MULT_mux_out_13_30_port)
                           ;
   U11268 : OAI22_X1 port map( A1 => n9117, A2 => n9133, B1 => n9168, B2 => 
                           n9118, ZN => DataPath_ALUhw_MULT_mux_out_14_30_port)
                           ;
   U11269 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n507, B => n9441, ZN => 
                           n9118);
   U11270 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_1_port, A2 => n7618, 
                           ZN => n9003);
   U11271 : NAND2_X1 port map( A1 => n8225, A2 => DataPath_i_PIPLIN_IN1_1_port,
                           ZN => n9004);
   U11272 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_29_port
                           , ZN => n9115);
   U11273 : OAI21_X1 port map( B1 => n8299, B2 => n8137, A => n9116, ZN => 
                           n9441);
   U11274 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_28_port
                           , ZN => n9116);
   U11275 : OAI22_X1 port map( A1 => n8134, A2 => n9660, B1 => n7726, B2 => 
                           n9913, ZN => DataPath_ALUhw_MULT_mux_out_0_29_port);
   U11276 : OAI22_X1 port map( A1 => n8441, A2 => n9504, B1 => n9473, B2 => 
                           n8430, ZN => DataPath_ALUhw_MULT_mux_out_1_29_port);
   U11277 : OAI22_X1 port map( A1 => n8444, A2 => n9528, B1 => n8402, B2 => 
                           n8447, ZN => DataPath_ALUhw_MULT_mux_out_2_29_port);
   U11278 : OAI22_X1 port map( A1 => n7615, A2 => n7773, B1 => n8449, B2 => 
                           n9600, ZN => DataPath_ALUhw_MULT_mux_out_3_29_port);
   U11279 : OAI22_X1 port map( A1 => n8452, A2 => n7799, B1 => n9961, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_29_port);
   U11280 : OAI22_X1 port map( A1 => n7787, A2 => n9495, B1 => n8454, B2 => 
                           n7776, ZN => DataPath_ALUhw_MULT_mux_out_5_29_port);
   U11281 : OAI22_X1 port map( A1 => n9080, A2 => n8439, B1 => n8455, B2 => 
                           n8405, ZN => DataPath_ALUhw_MULT_mux_out_6_29_port);
   U11282 : OAI22_X1 port map( A1 => n7785, A2 => n7981, B1 => n9784, B2 => 
                           n8456, ZN => DataPath_ALUhw_MULT_mux_out_7_29_port);
   U11283 : OAI22_X1 port map( A1 => n7767, A2 => n9822, B1 => n8427, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_29_port);
   U11284 : OAI22_X1 port map( A1 => n9094, A2 => n9122, B1 => n8401, B2 => 
                           n9095, ZN => DataPath_ALUhw_MULT_mux_out_9_29_port);
   U11285 : OAI22_X1 port map( A1 => n9099, A2 => n8436, B1 => n10017, B2 => 
                           n9100, ZN => DataPath_ALUhw_MULT_mux_out_10_29_port)
                           ;
   U11286 : OAI22_X1 port map( A1 => n9104, A2 => n7795, B1 => n9248, B2 => 
                           n9105, ZN => DataPath_ALUhw_MULT_mux_out_11_29_port)
                           ;
   U11287 : OAI22_X1 port map( A1 => n9109, A2 => n9188, B1 => n9986, B2 => 
                           n9110, ZN => DataPath_ALUhw_MULT_mux_out_12_29_port)
                           ;
   U11288 : OAI22_X1 port map( A1 => n9113, A2 => n9168, B1 => n8399, B2 => 
                           n9114, ZN => DataPath_ALUhw_MULT_mux_out_13_29_port)
                           ;
   U11289 : XNOR2_X1 port map( A => n7817, B => n9518, ZN => n9114);
   U11290 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_27_port
                           , ZN => n9111);
   U11291 : OAI21_X1 port map( B1 => n8256, B2 => n7929, A => n9112, ZN => 
                           n9518);
   U11292 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_26_port
                           , ZN => n9112);
   U11293 : OAI22_X1 port map( A1 => n9934, A2 => n8442, B1 => n9504, B2 => 
                           n8432, ZN => DataPath_ALUhw_MULT_mux_out_1_28_port);
   U11294 : OAI22_X1 port map( A1 => n8443, A2 => n9600, B1 => n9528, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_28_port);
   U11295 : OAI22_X1 port map( A1 => n7615, A2 => n9961, B1 => n8450, B2 => 
                           n7773, ZN => DataPath_ALUhw_MULT_mux_out_3_28_port);
   U11296 : OAI22_X1 port map( A1 => n9074, A2 => n7776, B1 => n7799, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_28_port);
   U11297 : OAI22_X1 port map( A1 => n7787, A2 => n8405, B1 => n9079, B2 => 
                           n9495, ZN => DataPath_ALUhw_MULT_mux_out_5_28_port);
   U11298 : OAI22_X1 port map( A1 => n9080, A2 => n7727, B1 => n8455, B2 => 
                           n8439, ZN => DataPath_ALUhw_MULT_mux_out_6_28_port);
   U11299 : OAI22_X1 port map( A1 => n7785, A2 => n8427, B1 => n7981, B2 => 
                           n9086, ZN => DataPath_ALUhw_MULT_mux_out_7_28_port);
   U11300 : OAI22_X1 port map( A1 => n9088, A2 => n8401, B1 => n9822, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_28_port);
   U11301 : OAI22_X1 port map( A1 => n9094, A2 => n8404, B1 => n9122, B2 => 
                           n9095, ZN => DataPath_ALUhw_MULT_mux_out_9_28_port);
   U11302 : OAI22_X1 port map( A1 => n9099, A2 => n9248, B1 => n8437, B2 => 
                           n8457, ZN => DataPath_ALUhw_MULT_mux_out_10_28_port)
                           ;
   U11303 : OAI22_X1 port map( A1 => n9104, A2 => n9986, B1 => n8400, B2 => 
                           n9105, ZN => DataPath_ALUhw_MULT_mux_out_11_28_port)
                           ;
   U11304 : OAI22_X1 port map( A1 => n9109, A2 => n8398, B1 => n9188, B2 => 
                           n9110, ZN => DataPath_ALUhw_MULT_mux_out_12_28_port)
                           ;
   U11305 : NAND2_X1 port map( A1 => n8990, A2 => n8989, ZN => n9197);
   U11306 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_3_port, A2 => n8555, 
                           ZN => n8989);
   U11307 : NAND2_X1 port map( A1 => n8225, A2 => DataPath_i_PIPLIN_IN1_3_port,
                           ZN => n8990);
   U11308 : OAI21_X1 port map( B1 => n8255, B2 => n7929, A => n9107, ZN => 
                           n9567);
   U11309 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_24_port
                           , ZN => n9107);
   U11310 : INV_X1 port map( A => n7817, ZN => n9935);
   U11311 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_25_port
                           , ZN => n9106);
   U11312 : OAI22_X1 port map( A1 => n8134, A2 => n9504, B1 => n7726, B2 => 
                           n9473, ZN => DataPath_ALUhw_MULT_mux_out_0_27_port);
   U11313 : OAI22_X1 port map( A1 => n8442, A2 => n9528, B1 => n9934, B2 => 
                           n8430, ZN => DataPath_ALUhw_MULT_mux_out_1_27_port);
   U11314 : OAI22_X1 port map( A1 => n8445, A2 => n7773, B1 => n9600, B2 => 
                           n8447, ZN => DataPath_ALUhw_MULT_mux_out_2_27_port);
   U11315 : OAI22_X1 port map( A1 => n7615, A2 => n7799, B1 => n8451, B2 => 
                           n9961, ZN => DataPath_ALUhw_MULT_mux_out_3_27_port);
   U11316 : OAI22_X1 port map( A1 => n8453, A2 => n9495, B1 => n7776, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_27_port);
   U11317 : OAI22_X1 port map( A1 => n7769, A2 => n8439, B1 => n8454, B2 => 
                           n8405, ZN => DataPath_ALUhw_MULT_mux_out_5_27_port);
   U11318 : OAI22_X1 port map( A1 => n7770, A2 => n7981, B1 => n8455, B2 => 
                           n7727, ZN => DataPath_ALUhw_MULT_mux_out_6_27_port);
   U11319 : OAI22_X1 port map( A1 => n9085, A2 => n9822, B1 => n8428, B2 => 
                           n8456, ZN => DataPath_ALUhw_MULT_mux_out_7_27_port);
   U11320 : OAI22_X1 port map( A1 => n7767, A2 => n9122, B1 => n8401, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_27_port);
   U11321 : OAI22_X1 port map( A1 => n9094, A2 => n8435, B1 => n8404, B2 => 
                           n9095, ZN => DataPath_ALUhw_MULT_mux_out_9_27_port);
   U11322 : OAI22_X1 port map( A1 => n9099, A2 => n7795, B1 => n9248, B2 => 
                           n8457, ZN => DataPath_ALUhw_MULT_mux_out_10_27_port)
                           ;
   U11323 : OAI22_X1 port map( A1 => n9104, A2 => n9188, B1 => n9986, B2 => 
                           n9105, ZN => DataPath_ALUhw_MULT_mux_out_11_27_port)
                           ;
   U11324 : OAI21_X1 port map( B1 => n8259, B2 => n8557, A => n8963, ZN => 
                           n9903);
   U11325 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_4_port, A2 => n7617, 
                           ZN => n8963);
   U11326 : INV_X1 port map( A => DP_OP_751_130_6421_n711, ZN => n9601);
   U11327 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_23_port
                           , ZN => n9101);
   U11328 : OAI21_X1 port map( B1 => n8254, B2 => n7929, A => n9103, ZN => 
                           n9637);
   U11329 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_22_port
                           , ZN => n9103);
   U11330 : OAI22_X1 port map( A1 => n8440, A2 => n9600, B1 => n9528, B2 => 
                           n8432, ZN => DataPath_ALUhw_MULT_mux_out_1_26_port);
   U11331 : OAI22_X1 port map( A1 => n8443, A2 => n9961, B1 => n7773, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_26_port);
   U11332 : OAI22_X1 port map( A1 => n7616, A2 => n7776, B1 => n8451, B2 => 
                           n7799, ZN => DataPath_ALUhw_MULT_mux_out_3_26_port);
   U11333 : OAI22_X1 port map( A1 => n8452, A2 => n8405, B1 => n9495, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_26_port);
   U11334 : OAI22_X1 port map( A1 => n7787, A2 => n7727, B1 => n8454, B2 => 
                           n8439, ZN => DataPath_ALUhw_MULT_mux_out_5_26_port);
   U11335 : OAI22_X1 port map( A1 => n7770, A2 => n8428, B1 => n8455, B2 => 
                           n7981, ZN => DataPath_ALUhw_MULT_mux_out_6_26_port);
   U11336 : OAI22_X1 port map( A1 => n9085, A2 => n8401, B1 => n9822, B2 => 
                           n9086, ZN => DataPath_ALUhw_MULT_mux_out_7_26_port);
   U11337 : OAI22_X1 port map( A1 => n7767, A2 => n8403, B1 => n9122, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_26_port);
   U11338 : OAI22_X1 port map( A1 => n9094, A2 => n9248, B1 => n8436, B2 => 
                           n9095, ZN => DataPath_ALUhw_MULT_mux_out_9_26_port);
   U11339 : OAI22_X1 port map( A1 => n9099, A2 => n9986, B1 => n8400, B2 => 
                           n8457, ZN => DataPath_ALUhw_MULT_mux_out_10_26_port)
                           ;
   U11340 : OAI21_X1 port map( B1 => n8258, B2 => n8557, A => n8947, ZN => 
                           n9985);
   U11341 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_5_port, A2 => n8555, 
                           ZN => n8947);
   U11342 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_21_port
                           , ZN => n9096);
   U11343 : OAI22_X1 port map( A1 => n8134, A2 => n9528, B1 => n7726, B2 => 
                           n9934, ZN => DataPath_ALUhw_MULT_mux_out_0_25_port);
   U11344 : OAI22_X1 port map( A1 => n8440, A2 => n7714, B1 => n8431, B2 => 
                           n9600, ZN => DataPath_ALUhw_MULT_mux_out_1_25_port);
   U11345 : OAI22_X1 port map( A1 => n8444, A2 => n9312, B1 => n9961, B2 => 
                           n8447, ZN => DataPath_ALUhw_MULT_mux_out_2_25_port);
   U11346 : OAI22_X1 port map( A1 => n8453, A2 => n8439, B1 => n8406, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_25_port);
   U11347 : OAI22_X1 port map( A1 => n7769, A2 => n7981, B1 => n8454, B2 => 
                           n7727, ZN => DataPath_ALUhw_MULT_mux_out_5_25_port);
   U11348 : OAI22_X1 port map( A1 => n9080, A2 => n9822, B1 => n9081, B2 => 
                           n8427, ZN => DataPath_ALUhw_MULT_mux_out_6_25_port);
   U11349 : OAI22_X1 port map( A1 => n9085, A2 => n9122, B1 => n8401, B2 => 
                           n8456, ZN => DataPath_ALUhw_MULT_mux_out_7_25_port);
   U11350 : OAI22_X1 port map( A1 => n7767, A2 => n8437, B1 => n8404, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_25_port);
   U11351 : OAI22_X1 port map( A1 => n9094, A2 => n7795, B1 => n9248, B2 => 
                           n9095, ZN => DataPath_ALUhw_MULT_mux_out_9_25_port);
   U11352 : BUF_X1 port map( A => n9239, Z => n8400);
   U11353 : INV_X1 port map( A => n9240, ZN => n9239);
   U11354 : OAI21_X1 port map( B1 => n8263, B2 => n8557, A => n9026, ZN => 
                           n9240);
   U11355 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_6_port, A2 => n7617, 
                           ZN => n9026);
   U11356 : AOI21_X1 port map( B1 => n8563, B2 => n9743, A => n9092, ZN => 
                           n9093);
   U11357 : NOR2_X1 port map( A1 => n8563, A2 => n9693, ZN => n9092);
   U11358 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_19_port
                           , ZN => n9090);
   U11359 : OAI21_X1 port map( B1 => n8253, B2 => n7929, A => n9091, ZN => 
                           n9743);
   U11360 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_18_port
                           , ZN => n9091);
   U11361 : OAI22_X1 port map( A1 => n7619, A2 => n9961, B1 => n7753, B2 => 
                           n7714, ZN => DataPath_ALUhw_MULT_mux_out_1_24_port);
   U11362 : OAI22_X1 port map( A1 => n8444, A2 => n9692, B1 => n9312, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_24_port);
   U11363 : OAI22_X1 port map( A1 => n7616, A2 => n8405, B1 => n8449, B2 => 
                           n9495, ZN => DataPath_ALUhw_MULT_mux_out_3_24_port);
   U11364 : OAI22_X1 port map( A1 => n8453, A2 => n7727, B1 => n8439, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_24_port);
   U11365 : OAI22_X1 port map( A1 => n7769, A2 => n10032, B1 => n9079, B2 => 
                           n7981, ZN => DataPath_ALUhw_MULT_mux_out_5_24_port);
   U11366 : OAI22_X1 port map( A1 => n9085, A2 => n8403, B1 => n9122, B2 => 
                           n9086, ZN => DataPath_ALUhw_MULT_mux_out_7_24_port);
   U11367 : OAI22_X1 port map( A1 => n7767, A2 => n9248, B1 => n8436, B2 => 
                           n7790, ZN => DataPath_ALUhw_MULT_mux_out_8_24_port);
   U11368 : OAI21_X1 port map( B1 => n8264, B2 => n8557, A => n9046, ZN => 
                           n9253);
   U11369 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_7_port, A2 => n8555, 
                           ZN => n9046);
   U11370 : OAI21_X1 port map( B1 => n8251, B2 => n7929, A => n9087, ZN => 
                           n9754);
   U11371 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_16_port
                           , ZN => n9087);
   U11372 : OAI22_X1 port map( A1 => n7619, A2 => n9312, B1 => n7753, B2 => 
                           n9961, ZN => DataPath_ALUhw_MULT_mux_out_1_23_port);
   U11373 : OAI22_X1 port map( A1 => n8445, A2 => n9495, B1 => n9692, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_23_port);
   U11374 : OAI22_X1 port map( A1 => n7616, A2 => n8439, B1 => n8450, B2 => 
                           n8405, ZN => DataPath_ALUhw_MULT_mux_out_3_23_port);
   U11375 : OAI22_X1 port map( A1 => n8452, A2 => n7981, B1 => n7727, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_23_port);
   U11376 : OAI22_X1 port map( A1 => n7769, A2 => n9822, B1 => n9079, B2 => 
                           n8427, ZN => DataPath_ALUhw_MULT_mux_out_5_23_port);
   U11377 : OAI22_X1 port map( A1 => n7770, A2 => n9122, B1 => n9081, B2 => 
                           n8401, ZN => DataPath_ALUhw_MULT_mux_out_6_23_port);
   U11378 : OAI22_X1 port map( A1 => n7785, A2 => n8436, B1 => n8404, B2 => 
                           n8456, ZN => DataPath_ALUhw_MULT_mux_out_7_23_port);
   U11379 : OAI211_X1 port map( C1 => n9807, C2 => DP_OP_751_130_6421_n1119, A 
                           => n9084, B => n9083, ZN => n9085);
   U11380 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1221, A2 => 
                           DP_OP_751_130_6421_n1119, ZN => n9083);
   U11381 : NAND2_X1 port map( A1 => n8227, A2 => n9807, ZN => n9084);
   U11382 : NAND2_X1 port map( A1 => n8137, A2 => DataPath_i_PIPLIN_IN2_15_port
                           , ZN => n9082);
   U11383 : OAI22_X1 port map( A1 => n7751, A2 => n9961, B1 => n7726, B2 => 
                           n7714, ZN => DataPath_ALUhw_MULT_mux_out_0_22_port);
   U11384 : OAI22_X1 port map( A1 => n8440, A2 => n9692, B1 => n8429, B2 => 
                           n9312, ZN => DataPath_ALUhw_MULT_mux_out_1_22_port);
   U11385 : OAI22_X1 port map( A1 => n8445, A2 => n8405, B1 => n9495, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_22_port);
   U11386 : OAI22_X1 port map( A1 => n7615, A2 => n9784, B1 => n9070, B2 => 
                           n8439, ZN => DataPath_ALUhw_MULT_mux_out_3_22_port);
   U11387 : OAI22_X1 port map( A1 => n7769, A2 => n8401, B1 => n8454, B2 => 
                           n9822, ZN => DataPath_ALUhw_MULT_mux_out_5_22_port);
   U11388 : OAI22_X1 port map( A1 => n7770, A2 => n8404, B1 => n8455, B2 => 
                           n9122, ZN => DataPath_ALUhw_MULT_mux_out_6_22_port);
   U11389 : OAI21_X1 port map( B1 => n8261, B2 => n8557, A => n9006, ZN => 
                           n10016);
   U11390 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_9_port, A2 => n8555, 
                           ZN => n9006);
   U11391 : OAI22_X1 port map( A1 => n8441, A2 => n9495, B1 => n8429, B2 => 
                           n9692, ZN => DataPath_ALUhw_MULT_mux_out_1_21_port);
   U11392 : OAI22_X1 port map( A1 => n8443, A2 => n9753, B1 => n8406, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_21_port);
   U11393 : OAI22_X1 port map( A1 => n7615, A2 => n7309, B1 => n9784, B2 => 
                           n8451, ZN => DataPath_ALUhw_MULT_mux_out_3_21_port);
   U11394 : OAI22_X1 port map( A1 => n8452, A2 => n9822, B1 => n8428, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_21_port);
   U11395 : OAI22_X1 port map( A1 => n7787, A2 => n9122, B1 => n8454, B2 => 
                           n8401, ZN => DataPath_ALUhw_MULT_mux_out_5_21_port);
   U11396 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_10_port, A2 => n7618, 
                           ZN => n8977);
   U11397 : NAND2_X1 port map( A1 => n8225, A2 => DataPath_i_PIPLIN_IN1_10_port
                           , ZN => n8978);
   U11398 : OAI211_X1 port map( C1 => n9872, C2 => DP_OP_751_130_6421_n1323, A 
                           => n9077, B => n9076, ZN => n9078);
   U11399 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1323, A2 => 
                           DP_OP_751_130_6421_n1425, ZN => n9076);
   U11400 : NAND2_X1 port map( A1 => n7798, A2 => n9872, ZN => n9077);
   U11401 : OAI22_X1 port map( A1 => n8405, A2 => n7619, B1 => n7753, B2 => 
                           n9495, ZN => DataPath_ALUhw_MULT_mux_out_1_20_port);
   U11402 : OAI22_X1 port map( A1 => n8444, A2 => n9784, B1 => n9753, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_20_port);
   U11403 : OAI22_X1 port map( A1 => n7615, A2 => n8427, B1 => n7981, B2 => 
                           n8450, ZN => DataPath_ALUhw_MULT_mux_out_3_20_port);
   U11404 : OAI22_X1 port map( A1 => n8452, A2 => n8401, B1 => n9822, B2 => 
                           n7771, ZN => DataPath_ALUhw_MULT_mux_out_4_20_port);
   U11405 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1527, B => n9271, ZN =>
                           n9075);
   U11406 : OAI21_X1 port map( B1 => n8260, B2 => n8557, A => n8993, ZN => 
                           n9843);
   U11407 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_11_port, A2 => n7617, 
                           ZN => n8993);
   U11408 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1425, A2 => 
                           DP_OP_751_130_6421_n1527, ZN => n9072);
   U11409 : NAND2_X1 port map( A1 => n8561, A2 => n9271, ZN => n9073);
   U11410 : OAI21_X1 port map( B1 => n8247, B2 => n8069, A => n9071, ZN => 
                           n9271);
   U11411 : NAND2_X1 port map( A1 => n7723, A2 => DataPath_i_PIPLIN_IN2_8_port,
                           ZN => n9071);
   U11412 : OAI22_X1 port map( A1 => n7619, A2 => n9753, B1 => n8406, B2 => 
                           n7753, ZN => DataPath_ALUhw_MULT_mux_out_1_19_port);
   U11413 : BUF_X1 port map( A => n9062, Z => n8430);
   U11414 : OAI22_X1 port map( A1 => n8443, A2 => n7309, B1 => n7727, B2 => 
                           n8447, ZN => DataPath_ALUhw_MULT_mux_out_2_19_port);
   U11415 : OAI22_X1 port map( A1 => n7616, A2 => n9822, B1 => n8427, B2 => 
                           n8451, ZN => DataPath_ALUhw_MULT_mux_out_3_19_port);
   U11416 : NAND2_X1 port map( A1 => n8965, A2 => n8964, ZN => n9821);
   U11417 : NAND2_X1 port map( A1 => n8225, A2 => DataPath_i_PIPLIN_IN1_12_port
                           , ZN => n8965);
   U11418 : AOI21_X1 port map( B1 => n8561, B2 => n9241, A => n9067, ZN => 
                           n9068);
   U11419 : NOR2_X1 port map( A1 => n8561, A2 => n8560, ZN => n9067);
   U11420 : OAI21_X1 port map( B1 => n8245, B2 => n8069, A => n9065, ZN => n403
                           );
   U11421 : NAND2_X1 port map( A1 => n7723, A2 => DataPath_i_PIPLIN_IN2_7_port,
                           ZN => n9065);
   U11422 : NAND2_X1 port map( A1 => n7723, A2 => n486, ZN => n9066);
   U11423 : OAI22_X1 port map( A1 => n8442, A2 => n9784, B1 => n8432, B2 => 
                           n9753, ZN => DataPath_ALUhw_MULT_mux_out_1_18_port);
   U11424 : OAI22_X1 port map( A1 => n8443, A2 => n8428, B1 => n7309, B2 => 
                           n8446, ZN => DataPath_ALUhw_MULT_mux_out_2_18_port);
   U11425 : BUF_X1 port map( A => n10032, Z => n8428);
   U11426 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_13_port, A2 => n7617, 
                           ZN => n8944);
   U11427 : NAND2_X1 port map( A1 => n8558, A2 => DataPath_i_PIPLIN_IN1_13_port
                           , ZN => n8945);
   U11428 : NAND2_X1 port map( A1 => DP_OP_751_130_6421_n1731, A2 => n9883, ZN 
                           => n9370);
   U11429 : NAND2_X1 port map( A1 => n8193, A2 => DataPath_i_PIPLIN_IN2_4_port,
                           ZN => n8941);
   U11430 : NAND2_X1 port map( A1 => n7732, A2 => DataPath_i_PIPLIN_B_4_port, 
                           ZN => n8942);
   U11431 : OAI22_X1 port map( A1 => n7309, A2 => n8440, B1 => n7727, B2 => 
                           n8432, ZN => DataPath_ALUhw_MULT_mux_out_1_17_port);
   U11432 : BUF_X1 port map( A => n9062, Z => n8431);
   U11433 : OAI21_X1 port map( B1 => n7754, B2 => n8004, A => n8988, ZN => 
                           n9062);
   U11434 : NAND2_X1 port map( A1 => n7754, A2 => n9165, ZN => n8988);
   U11435 : OAI21_X1 port map( B1 => n8257, B2 => n8557, A => n9042, ZN => 
                           n9785);
   U11436 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_15_port, A2 => n8555, 
                           ZN => n9042);
   U11437 : OAI21_X1 port map( B1 => n8244, B2 => n8568, A => n8960, ZN => 
                           n9165);
   U11438 : NAND2_X1 port map( A1 => n8193, A2 => DataPath_i_PIPLIN_IN2_2_port,
                           ZN => n8960);
   U11439 : NAND2_X1 port map( A1 => n8568, A2 => DataPath_i_PIPLIN_IN2_1_port,
                           ZN => n8938);
   U11440 : NAND2_X1 port map( A1 => n8567, A2 => DataPath_i_PIPLIN_IN2_3_port,
                           ZN => n8939);
   U11441 : NAND2_X1 port map( A1 => n7732, A2 => DataPath_i_PIPLIN_B_3_port, 
                           ZN => n8940);
   U11442 : AOI22_X1 port map( A1 => n10278, A2 => n10276, B1 => i_RD1_29_port,
                           B2 => n10418, ZN => n10277);
   U11443 : NOR2_X1 port map( A1 => n10418, A2 => n10275, ZN => n10276);
   U11444 : OAI21_X1 port map( B1 => n10270, B2 => n7757, A => n10269, ZN => 
                           n7031);
   U11445 : AOI22_X1 port map( A1 => n10418, A2 => i_RD1_30_port, B1 => 
                           IRAM_ADDRESS_30_port, B2 => n10417, ZN => n10269);
   U11446 : XNOR2_X1 port map( A => n10268, B => IRAM_ADDRESS_30_port, ZN => 
                           n10270);
   U11447 : AOI22_X1 port map( A1 => n10418, A2 => i_RD1_31_port, B1 => 
                           IRAM_ADDRESS_31_port, B2 => n10417, ZN => n10419);
   U11448 : NOR2_X1 port map( A1 => n10293, A2 => n10281, ZN => n10271);
   U11449 : NAND2_X1 port map( A1 => n10293, A2 => n10281, ZN => n10279);
   U11450 : NAND2_X1 port map( A1 => n10293, A2 => IRAM_ADDRESS_27_port, ZN => 
                           n10266);
   U11451 : NAND2_X1 port map( A1 => n10293, A2 => IRAM_ADDRESS_26_port, ZN => 
                           n10287);
   U11452 : XNOR2_X1 port map( A => n10293, B => IRAM_ADDRESS_27_port, ZN => 
                           n10284);
   U11453 : OR2_X1 port map( A1 => n10293, A2 => IRAM_ADDRESS_26_port, ZN => 
                           n10288);
   U11454 : NOR2_X1 port map( A1 => n10293, A2 => IRAM_ADDRESS_25_port, ZN => 
                           n10264);
   U11455 : NAND2_X1 port map( A1 => n10293, A2 => IRAM_ADDRESS_25_port, ZN => 
                           n10265);
   U11456 : OR2_X1 port map( A1 => n7604, A2 => n169, ZN => n10262);
   U11457 : NAND2_X1 port map( A1 => n10260, A2 => n10259, ZN => n10295);
   U11458 : NAND2_X1 port map( A1 => n10298, A2 => n7611, ZN => n10259);
   U11459 : NAND2_X1 port map( A1 => n8935, A2 => IRAM_ADDRESS_15_port, ZN => 
                           n10235);
   U11460 : INV_X1 port map( A => n10237, ZN => n8935);
   U11461 : AND2_X1 port map( A1 => n10237, A2 => n8300, ZN => n10236);
   U11462 : NOR2_X1 port map( A1 => n8931, A2 => n8279, ZN => n8932);
   U11463 : NAND2_X1 port map( A1 => n8931, A2 => n8279, ZN => n8933);
   U11464 : OR2_X1 port map( A1 => intadd_1_B_2_port, A2 => 
                           IRAM_ADDRESS_12_port, ZN => n8222);
   U11465 : NOR2_X1 port map( A1 => n7749, A2 => n179, ZN => intadd_1_B_2_port)
                           ;
   U11466 : NOR2_X1 port map( A1 => n7749, A2 => n180, ZN => intadd_1_B_1_port)
                           ;
   U11467 : NOR2_X1 port map( A1 => n7749, A2 => n8233, ZN => intadd_1_B_0_port
                           );
   U11468 : AND2_X1 port map( A1 => n8922, A2 => n205, ZN => n8926);
   U11469 : NAND2_X1 port map( A1 => n8923, A2 => IRAM_ADDRESS_9_port, ZN => 
                           n8927);
   U11470 : INV_X1 port map( A => n8922, ZN => n8923);
   U11471 : OR2_X1 port map( A1 => n7880, A2 => n8241, ZN => n8922);
   U11472 : NOR2_X1 port map( A1 => n10351, A2 => n8284, ZN => n8918);
   U11473 : NAND2_X1 port map( A1 => n10351, A2 => n8284, ZN => n8919);
   U11474 : OR2_X1 port map( A1 => n7880, A2 => n8234, ZN => n10351);
   U11475 : AND2_X1 port map( A1 => n8917, A2 => n8307, ZN => n10355);
   U11476 : NAND2_X1 port map( A1 => n8916, A2 => IRAM_ADDRESS_6_port, ZN => 
                           n10356);
   U11477 : INV_X1 port map( A => n8917, ZN => n8916);
   U11478 : OR2_X1 port map( A1 => n7880, A2 => n8228, ZN => n8917);
   U11479 : NOR2_X1 port map( A1 => n8915, A2 => n207, ZN => n10362);
   U11480 : NAND2_X1 port map( A1 => n8915, A2 => n207, ZN => n10361);
   U11481 : OR2_X1 port map( A1 => n7880, A2 => n8198, ZN => n8915);
   U11482 : NOR2_X1 port map( A1 => n7880, A2 => n8190, ZN => intadd_0_B_3_port
                           );
   U11483 : AOI21_X1 port map( B1 => intadd_0_n9, B2 => intadd_0_n17, A => 
                           intadd_0_n10, ZN => intadd_0_n8);
   U11484 : NAND2_X1 port map( A1 => intadd_0_B_0_port, A2 => 
                           IRAM_ADDRESS_1_port, ZN => intadd_0_n19);
   U11485 : OR2_X1 port map( A1 => n7748, A2 => n193, ZN => n10369);
   U11486 : NOR2_X1 port map( A1 => intadd_0_B_0_port, A2 => 
                           IRAM_ADDRESS_1_port, ZN => intadd_0_n18);
   U11487 : NOR2_X1 port map( A1 => n7749, A2 => n10160, ZN => 
                           intadd_0_B_0_port);
   U11488 : NOR2_X1 port map( A1 => intadd_0_B_2_port, A2 => 
                           IRAM_ADDRESS_3_port, ZN => intadd_0_n11);
   U11489 : NOR2_X1 port map( A1 => n7748, A2 => n8226, ZN => intadd_0_B_2_port
                           );
   U11490 : NAND2_X1 port map( A1 => n8914, A2 => n8224, ZN => 
                           intadd_0_B_1_port);
   U11491 : NAND2_X1 port map( A1 => n10258, A2 => n10257, ZN => n10298);
   U11492 : NAND2_X1 port map( A1 => n10263, A2 => n8231, ZN => n10257);
   U11493 : NOR2_X1 port map( A1 => n8372, A2 => n8385, ZN => n8371);
   U11494 : INV_X1 port map( A => n10341, ZN => n8372);
   U11495 : AND2_X1 port map( A1 => n10243, A2 => n10334, ZN => n10341);
   U11496 : OR2_X1 port map( A1 => IRAM_ADDRESS_16_port, A2 => n10242, ZN => 
                           n10243);
   U11497 : NAND2_X1 port map( A1 => n10305, A2 => IRAM_ADDRESS_23_port, ZN => 
                           n10256);
   U11498 : NAND2_X1 port map( A1 => n10263, A2 => n10255, ZN => n10305);
   U11499 : OR2_X1 port map( A1 => n7604, A2 => n170, ZN => n10255);
   U11500 : OR2_X1 port map( A1 => n10310, A2 => n8274, ZN => n10304);
   U11501 : AND2_X1 port map( A1 => n8390, A2 => n10314, ZN => n8387);
   U11502 : NAND2_X1 port map( A1 => n10310, A2 => n8274, ZN => n10311);
   U11503 : NAND2_X1 port map( A1 => n10258, A2 => n10254, ZN => n10310);
   U11504 : NAND2_X1 port map( A1 => n10263, A2 => n171, ZN => n10254);
   U11505 : NAND2_X1 port map( A1 => n10316, A2 => n8275, ZN => n10303);
   U11506 : OR2_X1 port map( A1 => n10316, A2 => n8275, ZN => n10314);
   U11507 : NAND2_X1 port map( A1 => n10258, A2 => n10253, ZN => n10316);
   U11508 : NAND2_X1 port map( A1 => n10263, A2 => n8232, ZN => n10253);
   U11509 : NAND2_X1 port map( A1 => n10263, A2 => n7604, ZN => n10258);
   U11510 : NOR2_X1 port map( A1 => n10319, A2 => IRAM_ADDRESS_20_port, ZN => 
                           n8389);
   U11511 : OR2_X1 port map( A1 => n8236, A2 => n10325, ZN => n8202);
   U11512 : XNOR2_X1 port map( A => n10250, B => IRAM_ADDRESS_19_port, ZN => 
                           n10325);
   U11513 : XNOR2_X1 port map( A => n10247, B => IRAM_ADDRESS_17_port, ZN => 
                           n10336);
   U11514 : OR2_X1 port map( A1 => n10250, A2 => IRAM_ADDRESS_19_port, ZN => 
                           n10251);
   U11515 : NAND2_X1 port map( A1 => n10263, A2 => n10246, ZN => n10250);
   U11516 : OR2_X1 port map( A1 => n10261, A2 => n173, ZN => n10246);
   U11517 : NOR2_X1 port map( A1 => n10249, A2 => IRAM_ADDRESS_18_port, ZN => 
                           n10326);
   U11518 : NAND2_X1 port map( A1 => n10249, A2 => IRAM_ADDRESS_18_port, ZN => 
                           n10327);
   U11519 : NAND2_X1 port map( A1 => n10263, A2 => n10245, ZN => n10249);
   U11520 : OR2_X1 port map( A1 => n10261, A2 => n174, ZN => n10245);
   U11521 : OR2_X1 port map( A1 => n10247, A2 => IRAM_ADDRESS_17_port, ZN => 
                           n10248);
   U11522 : NAND2_X1 port map( A1 => n10263, A2 => n10244, ZN => n10247);
   U11523 : OR2_X1 port map( A1 => n10261, A2 => n175, ZN => n10244);
   U11524 : NAND2_X1 port map( A1 => n10263, A2 => n10241, ZN => n10242);
   U11525 : OR2_X1 port map( A1 => n10261, A2 => n176, ZN => n10241);
   U11526 : INV_X1 port map( A => n10238, ZN => n10239);
   U11527 : AOI21_X1 port map( B1 => n10384, B2 => n8360, A => 
                           CU_I_i_FILL_delay, ZN => n8584);
   U11528 : INV_X1 port map( A => n8890, ZN => n8891);
   U11529 : INV_X1 port map( A => n10225, ZN => n10382);
   U11530 : INV_X1 port map( A => n10384, ZN => n10372);
   U11531 : AND2_X1 port map( A1 => n7962, A2 => n8354, ZN => n10384);
   U11532 : NOR2_X1 port map( A1 => n8889, A2 => n8907, ZN => n10385);
   U11533 : NAND2_X1 port map( A1 => n8237, A2 => n163, ZN => n8907);
   U11534 : INV_X1 port map( A => n10393, ZN => n10400);
   U11535 : NAND2_X1 port map( A1 => n8881, A2 => n8880, ZN => n8882);
   U11536 : INV_X1 port map( A => n8876, ZN => n8878);
   U11537 : INV_X1 port map( A => n8875, ZN => n8879);
   U11538 : OAI211_X1 port map( C1 => i_RD1_26_port, C2 => n8870, A => n8869, B
                           => n8868, ZN => n8871);
   U11539 : OAI22_X1 port map( A1 => n8867, A2 => n8866, B1 => n8865, B2 => 
                           n10292, ZN => n8869);
   U11540 : INV_X1 port map( A => n8864, ZN => n8866);
   U11541 : INV_X1 port map( A => n8865, ZN => n8870);
   U11542 : OAI21_X1 port map( B1 => n8875, B2 => n8863, A => n8886, ZN => 
                           n8885);
   U11543 : NAND2_X1 port map( A1 => n8862, A2 => i_RD1_30_port, ZN => n8863);
   U11544 : INV_X1 port map( A => n8861, ZN => n8862);
   U11545 : NAND2_X1 port map( A1 => n8875, A2 => n8860, ZN => n8886);
   U11546 : AND2_X1 port map( A1 => n8902, A2 => n10438, ZN => n8860);
   U11547 : INV_X1 port map( A => CU_I_CW_ID_UNSIGNED_ID_port, ZN => n10438);
   U11548 : OR3_X1 port map( A1 => n10194, A2 => n8900, A3 => n8895, ZN => 
                           n8902);
   U11549 : NAND2_X1 port map( A1 => n8894, A2 => n8859, ZN => n8895);
   U11550 : AND2_X1 port map( A1 => IR_4_port, A2 => IR_3_port, ZN => n8859);
   U11551 : NOR2_X1 port map( A1 => n8858, A2 => IR_6_port, ZN => n8894);
   U11552 : NAND2_X1 port map( A1 => IR_5_port, A2 => n11754, ZN => n8858);
   U11553 : XNOR2_X1 port map( A => IR_2_port, B => IR_1_port, ZN => n8900);
   U11554 : NAND2_X1 port map( A1 => n8857, A2 => n10225, ZN => n8887);
   U11555 : NOR2_X1 port map( A1 => n8848, A2 => n8847, ZN => n8849);
   U11556 : INV_X1 port map( A => n8843, ZN => n8844);
   U11557 : INV_X1 port map( A => n8877, ZN => n8840);
   U11558 : AND2_X1 port map( A1 => n8839, A2 => i_RD1_29_port, ZN => n8877);
   U11559 : NOR2_X1 port map( A1 => n8838, A2 => n8837, ZN => n8841);
   U11560 : OAI21_X1 port map( B1 => n8569, B2 => n8835, A => i_RD1_0_port, ZN 
                           => n8836);
   U11561 : INV_X1 port map( A => n8834, ZN => n8838);
   U11562 : NOR2_X1 port map( A1 => n8833, A2 => n8876, ZN => n8883);
   U11563 : XNOR2_X1 port map( A => n8861, B => n8832, ZN => n8876);
   U11564 : INV_X1 port map( A => i_RD1_30_port, ZN => n8832);
   U11565 : NAND2_X1 port map( A1 => n8831, A2 => n8830, ZN => n8861);
   U11566 : NAND2_X1 port map( A1 => n7768, A2 => i_RD2_30_port, ZN => n8830);
   U11567 : NAND2_X1 port map( A1 => n10165, A2 => n8569, ZN => n8831);
   U11568 : NAND2_X1 port map( A1 => n8829, A2 => n8828, ZN => n10165);
   U11569 : AOI21_X1 port map( B1 => n8424, B2 => IRAM_ADDRESS_30_port, A => 
                           n8827, ZN => n8828);
   U11570 : NOR2_X1 port map( A1 => n7621, A2 => n570, ZN => n8827);
   U11571 : OR2_X1 port map( A1 => n8875, A2 => n8826, ZN => n8833);
   U11572 : OAI22_X1 port map( A1 => i_RD1_28_port, A2 => n8825, B1 => n8839, 
                           B2 => i_RD1_29_port, ZN => n8826);
   U11573 : OAI21_X1 port map( B1 => n10166, B2 => n7768, A => n8824, ZN => 
                           n8839);
   U11574 : NAND2_X1 port map( A1 => n7768, A2 => n8823, ZN => n8824);
   U11575 : INV_X1 port map( A => i_RD2_29_port, ZN => n8823);
   U11576 : NAND2_X1 port map( A1 => n8829, A2 => n8822, ZN => n10166);
   U11577 : NAND2_X1 port map( A1 => n8880, A2 => n8821, ZN => n8875);
   U11578 : NAND2_X1 port map( A1 => n8820, A2 => n8819, ZN => n8821);
   U11579 : INV_X1 port map( A => i_RD1_31_port, ZN => n8819);
   U11580 : INV_X1 port map( A => n8818, ZN => n8820);
   U11581 : NAND2_X1 port map( A1 => n8818, A2 => i_RD1_31_port, ZN => n8880);
   U11582 : AOI21_X1 port map( B1 => n10164, B2 => n8569, A => n8817, ZN => 
                           n8818);
   U11583 : AND2_X1 port map( A1 => n7768, A2 => i_RD2_31_port, ZN => n8817);
   U11584 : NAND2_X1 port map( A1 => n8829, A2 => n8816, ZN => n10164);
   U11585 : NOR2_X1 port map( A1 => n8812, A2 => n8811, ZN => n8813);
   U11586 : NAND4_X1 port map( A1 => n8810, A2 => n8809, A3 => n8808, A4 => 
                           n8807, ZN => n8811);
   U11587 : NOR3_X1 port map( A1 => n8806, A2 => n8805, A3 => n8804, ZN => 
                           n8814);
   U11588 : INV_X1 port map( A => n8803, ZN => n8804);
   U11589 : NAND4_X1 port map( A1 => n8872, A2 => n8802, A3 => n8801, A4 => 
                           n8800, ZN => n8806);
   U11590 : NAND2_X1 port map( A1 => n8825, A2 => i_RD1_28_port, ZN => n8872);
   U11591 : OAI21_X1 port map( B1 => n10167, B2 => n7768, A => n8799, ZN => 
                           n8825);
   U11592 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => n8798, ZN => n8799);
   U11593 : INV_X1 port map( A => i_RD2_28_port, ZN => n8798);
   U11594 : NAND2_X1 port map( A1 => n8829, A2 => n8797, ZN => n10167);
   U11595 : AOI21_X1 port map( B1 => n8421, B2 => IRAM_ADDRESS_28_port, A => 
                           n8796, ZN => n8797);
   U11596 : NOR2_X1 port map( A1 => n7621, A2 => n569, ZN => n8796);
   U11597 : OAI211_X1 port map( C1 => n8791, C2 => i_RD1_24_port, A => n8867, B
                           => n8873, ZN => n8792);
   U11598 : NAND2_X1 port map( A1 => n8790, A2 => i_RD1_27_port, ZN => n8873);
   U11599 : AOI22_X1 port map( A1 => n8789, A2 => i_RD1_25_port, B1 => n8791, 
                           B2 => i_RD1_24_port, ZN => n8867);
   U11600 : AOI21_X1 port map( B1 => n10171, B2 => n8569, A => n8788, ZN => 
                           n8791);
   U11601 : AND2_X1 port map( A1 => n7768, A2 => i_RD2_24_port, ZN => n8788);
   U11602 : NAND2_X1 port map( A1 => n8829, A2 => n8787, ZN => n10171);
   U11603 : NAND2_X1 port map( A1 => n8868, A2 => n8864, ZN => n8793);
   U11604 : NAND2_X1 port map( A1 => n8786, A2 => n8785, ZN => n8864);
   U11605 : INV_X1 port map( A => i_RD1_25_port, ZN => n8785);
   U11606 : INV_X1 port map( A => n8789, ZN => n8786);
   U11607 : AOI21_X1 port map( B1 => n10170, B2 => n8569, A => n8784, ZN => 
                           n8789);
   U11608 : AND2_X1 port map( A1 => n7768, A2 => i_RD2_25_port, ZN => n8784);
   U11609 : NAND2_X1 port map( A1 => n8829, A2 => n8783, ZN => n10170);
   U11610 : AOI21_X1 port map( B1 => n8424, B2 => IRAM_ADDRESS_25_port, A => 
                           n8782, ZN => n8783);
   U11611 : NOR2_X1 port map( A1 => n7621, A2 => n566, ZN => n8782);
   U11612 : OR2_X1 port map( A1 => n8790, A2 => i_RD1_27_port, ZN => n8868);
   U11613 : OAI21_X1 port map( B1 => n10168, B2 => n7768, A => n8781, ZN => 
                           n8790);
   U11614 : NAND2_X1 port map( A1 => n7768, A2 => n8780, ZN => n8781);
   U11615 : INV_X1 port map( A => i_RD2_27_port, ZN => n8780);
   U11616 : NAND2_X1 port map( A1 => n8829, A2 => n8779, ZN => n10168);
   U11617 : AOI21_X1 port map( B1 => n8422, B2 => IRAM_ADDRESS_27_port, A => 
                           n8778, ZN => n8779);
   U11618 : NOR2_X1 port map( A1 => n7621, A2 => n568, ZN => n8778);
   U11619 : XNOR2_X1 port map( A => n8865, B => n10292, ZN => n8794);
   U11620 : INV_X1 port map( A => i_RD1_26_port, ZN => n10292);
   U11621 : NAND2_X1 port map( A1 => n8777, A2 => n8776, ZN => n8865);
   U11622 : NAND2_X1 port map( A1 => n7768, A2 => i_RD2_26_port, ZN => n8776);
   U11623 : NAND2_X1 port map( A1 => n10169, A2 => n8569, ZN => n8777);
   U11624 : NAND2_X1 port map( A1 => n8829, A2 => n8775, ZN => n10169);
   U11625 : OAI22_X1 port map( A1 => n8773, A2 => n8772, B1 => n8771, B2 => 
                           n8770, ZN => n8774);
   U11626 : INV_X1 port map( A => n8769, ZN => n8770);
   U11627 : AND2_X1 port map( A1 => n8768, A2 => n8767, ZN => n8771);
   U11628 : NAND2_X1 port map( A1 => n8766, A2 => i_RD1_22_port, ZN => n8767);
   U11629 : INV_X1 port map( A => n8765, ZN => n8766);
   U11630 : NAND2_X1 port map( A1 => n8764, A2 => n8763, ZN => n8772);
   U11631 : NAND2_X1 port map( A1 => n8762, A2 => n8761, ZN => n8764);
   U11632 : NAND2_X1 port map( A1 => n8760, A2 => i_RD1_20_port, ZN => n8761);
   U11633 : INV_X1 port map( A => n8759, ZN => n8760);
   U11634 : NOR2_X1 port map( A1 => n8773, A2 => n8758, ZN => n8815);
   U11635 : NAND2_X1 port map( A1 => n8756, A2 => n10318, ZN => n8763);
   U11636 : INV_X1 port map( A => i_RD1_21_port, ZN => n10318);
   U11637 : INV_X1 port map( A => n8755, ZN => n8756);
   U11638 : NAND2_X1 port map( A1 => n8755, A2 => i_RD1_21_port, ZN => n8762);
   U11639 : AOI21_X1 port map( B1 => n10174, B2 => n8569, A => n8754, ZN => 
                           n8755);
   U11640 : AND2_X1 port map( A1 => n7768, A2 => i_RD2_21_port, ZN => n8754);
   U11641 : NAND2_X1 port map( A1 => n8829, A2 => n8753, ZN => n10174);
   U11642 : AOI21_X1 port map( B1 => n8421, B2 => IRAM_ADDRESS_21_port, A => 
                           n8752, ZN => n8753);
   U11643 : NOR2_X1 port map( A1 => n7621, A2 => n562, ZN => n8752);
   U11644 : XNOR2_X1 port map( A => n8759, B => i_RD1_20_port, ZN => n8757);
   U11645 : NAND2_X1 port map( A1 => n8751, A2 => n8750, ZN => n8759);
   U11646 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_20_port, ZN => 
                           n8750);
   U11647 : NAND2_X1 port map( A1 => n10219, A2 => n8569, ZN => n8751);
   U11648 : NAND2_X1 port map( A1 => n8829, A2 => n8749, ZN => n10219);
   U11649 : NAND2_X1 port map( A1 => n8747, A2 => i_RD1_23_port, ZN => n8768);
   U11650 : NAND2_X1 port map( A1 => n8746, A2 => n8745, ZN => n8769);
   U11651 : INV_X1 port map( A => i_RD1_23_port, ZN => n8745);
   U11652 : INV_X1 port map( A => n8747, ZN => n8746);
   U11653 : AOI21_X1 port map( B1 => n10172, B2 => n8569, A => n8744, ZN => 
                           n8747);
   U11654 : AND2_X1 port map( A1 => n7768, A2 => i_RD2_23_port, ZN => n8744);
   U11655 : NAND2_X1 port map( A1 => n8829, A2 => n8743, ZN => n10172);
   U11656 : AOI21_X1 port map( B1 => n8421, B2 => IRAM_ADDRESS_23_port, A => 
                           n8742, ZN => n8743);
   U11657 : NOR2_X1 port map( A1 => n7621, A2 => n564, ZN => n8742);
   U11658 : XNOR2_X1 port map( A => n8765, B => i_RD1_22_port, ZN => n8748);
   U11659 : NAND2_X1 port map( A1 => n8741, A2 => n8740, ZN => n8765);
   U11660 : NAND2_X1 port map( A1 => i_SEL_CMPB, A2 => i_RD2_22_port, ZN => 
                           n8740);
   U11661 : NAND2_X1 port map( A1 => n10173, A2 => n8569, ZN => n8741);
   U11662 : NAND2_X1 port map( A1 => n8829, A2 => n8739, ZN => n10173);
   U11663 : OAI211_X1 port map( C1 => n8733, C2 => n8732, A => n8731, B => 
                           n8730, ZN => n8736);
   U11664 : NAND2_X1 port map( A1 => n8729, A2 => i_RD1_17_port, ZN => n8730);
   U11665 : NOR2_X1 port map( A1 => n8729, A2 => i_RD1_17_port, ZN => n8733);
   U11666 : INV_X1 port map( A => n8728, ZN => n8729);
   U11667 : OR2_X1 port map( A1 => n8724, A2 => i_RD1_19_port, ZN => n8735);
   U11668 : NAND2_X1 port map( A1 => n8724, A2 => i_RD1_19_port, ZN => n8738);
   U11669 : OAI21_X1 port map( B1 => n10175, B2 => n7768, A => n8723, ZN => 
                           n8724);
   U11670 : NAND2_X1 port map( A1 => n7768, A2 => n8722, ZN => n8723);
   U11671 : INV_X1 port map( A => i_RD2_19_port, ZN => n8722);
   U11672 : NAND2_X1 port map( A1 => n8829, A2 => n8721, ZN => n10175);
   U11673 : AOI21_X1 port map( B1 => n8421, B2 => IRAM_ADDRESS_19_port, A => 
                           n8720, ZN => n8721);
   U11674 : NOR2_X1 port map( A1 => n7621, A2 => n560, ZN => n8720);
   U11675 : XNOR2_X1 port map( A => n8728, B => i_RD1_17_port, ZN => n8725);
   U11676 : NAND2_X1 port map( A1 => n8719, A2 => n8718, ZN => n8728);
   U11677 : NAND2_X1 port map( A1 => n7768, A2 => i_RD2_17_port, ZN => n8718);
   U11678 : NAND2_X1 port map( A1 => n10177, A2 => n8569, ZN => n8719);
   U11679 : NAND2_X1 port map( A1 => n8829, A2 => n8717, ZN => n10177);
   U11680 : AOI21_X1 port map( B1 => n8421, B2 => IRAM_ADDRESS_17_port, A => 
                           n8716, ZN => n8717);
   U11681 : NOR2_X1 port map( A1 => n7621, A2 => n558, ZN => n8716);
   U11682 : NOR2_X1 port map( A1 => n8715, A2 => n8714, ZN => n8726);
   U11683 : OAI22_X1 port map( A1 => n8713, A2 => i_RD1_16_port, B1 => n8712, 
                           B2 => i_RD1_15_port, ZN => n8714);
   U11684 : OAI21_X1 port map( B1 => n10176, B2 => n7768, A => n8711, ZN => 
                           n8734);
   U11685 : AOI21_X1 port map( B1 => i_SEL_CMPB, B2 => n8710, A => 
                           i_RD1_18_port, ZN => n8711);
   U11686 : INV_X1 port map( A => i_RD2_18_port, ZN => n8710);
   U11687 : NAND2_X1 port map( A1 => n8709, A2 => n8708, ZN => n8731);
   U11688 : AOI21_X1 port map( B1 => i_SEL_CMPB, B2 => i_RD2_18_port, A => 
                           n10333, ZN => n8708);
   U11689 : INV_X1 port map( A => i_RD1_18_port, ZN => n10333);
   U11690 : NAND2_X1 port map( A1 => n10176, A2 => n8569, ZN => n8709);
   U11691 : NAND2_X1 port map( A1 => n8829, A2 => n8707, ZN => n10176);
   U11692 : NAND2_X1 port map( A1 => n8713, A2 => i_RD1_16_port, ZN => n8732);
   U11693 : OAI21_X1 port map( B1 => n10178, B2 => i_SEL_CMPB, A => n8706, ZN 
                           => n8713);
   U11694 : NAND2_X1 port map( A1 => n7768, A2 => n8705, ZN => n8706);
   U11695 : INV_X1 port map( A => i_RD2_16_port, ZN => n8705);
   U11696 : NAND2_X1 port map( A1 => n8829, A2 => n8704, ZN => n10178);
   U11697 : NAND2_X1 port map( A1 => n8712, A2 => i_RD1_15_port, ZN => n8800);
   U11698 : AOI21_X1 port map( B1 => n10179, B2 => n8569, A => n8702, ZN => 
                           n8712);
   U11699 : AND2_X1 port map( A1 => n7768, A2 => i_RD2_15_port, ZN => n8702);
   U11700 : AOI21_X1 port map( B1 => n8424, B2 => IRAM_ADDRESS_15_port, A => 
                           n8700, ZN => n8701);
   U11701 : NOR2_X1 port map( A1 => n7621, A2 => n556, ZN => n8700);
   U11702 : NAND2_X1 port map( A1 => n8699, A2 => i_RD1_14_port, ZN => n8846);
   U11703 : OAI22_X1 port map( A1 => n8699, A2 => i_RD1_14_port, B1 => n8697, 
                           B2 => i_RD1_13_port, ZN => n8698);
   U11704 : AOI21_X1 port map( B1 => n10217, B2 => n8569, A => n8696, ZN => 
                           n8699);
   U11705 : AND2_X1 port map( A1 => n7768, A2 => i_RD2_14_port, ZN => n8696);
   U11706 : NAND2_X1 port map( A1 => n8697, A2 => i_RD1_13_port, ZN => n8801);
   U11707 : OAI21_X1 port map( B1 => n10215, B2 => n7768, A => n8694, ZN => 
                           n8697);
   U11708 : NAND2_X1 port map( A1 => n7768, A2 => n11797, ZN => n8694);
   U11709 : INV_X1 port map( A => i_RD2_13_port, ZN => n11797);
   U11710 : AOI21_X1 port map( B1 => n8422, B2 => IRAM_ADDRESS_13_port, A => 
                           n8692, ZN => n8693);
   U11711 : NOR2_X1 port map( A1 => n7621, A2 => n554, ZN => n8692);
   U11712 : OAI21_X1 port map( B1 => n10213, B2 => n7768, A => n8690, ZN => 
                           n8845);
   U11713 : AOI21_X1 port map( B1 => i_SEL_CMPB, B2 => n8689, A => 
                           i_RD1_12_port, ZN => n8690);
   U11714 : INV_X1 port map( A => i_RD2_12_port, ZN => n8689);
   U11715 : NAND2_X1 port map( A1 => n8688, A2 => n8687, ZN => n8834);
   U11716 : AOI21_X1 port map( B1 => i_SEL_CMPB, B2 => i_RD2_12_port, A => 
                           n8686, ZN => n8687);
   U11717 : NAND2_X1 port map( A1 => n10213, A2 => n8569, ZN => n8688);
   U11718 : AOI21_X1 port map( B1 => n8421, B2 => IRAM_ADDRESS_12_port, A => 
                           n8684, ZN => n8685);
   U11719 : NOR2_X1 port map( A1 => n7621, A2 => n8265, ZN => n8684);
   U11720 : NAND2_X1 port map( A1 => n8683, A2 => i_RD1_11_port, ZN => n8808);
   U11721 : OAI21_X1 port map( B1 => n8683, B2 => i_RD1_11_port, A => n8681, ZN
                           => n8805);
   U11722 : NAND2_X1 port map( A1 => n8680, A2 => n8679, ZN => n8681);
   U11723 : INV_X1 port map( A => n8678, ZN => n8680);
   U11724 : OAI21_X1 port map( B1 => n10180, B2 => n7768, A => n8677, ZN => 
                           n8683);
   U11725 : NAND2_X1 port map( A1 => n7768, A2 => n8676, ZN => n8677);
   U11726 : INV_X1 port map( A => i_RD2_11_port, ZN => n8676);
   U11727 : AOI21_X1 port map( B1 => n8422, B2 => IRAM_ADDRESS_11_port, A => 
                           n8674, ZN => n8675);
   U11728 : NOR2_X1 port map( A1 => n7621, A2 => n552, ZN => n8674);
   U11729 : AOI22_X1 port map( A1 => n8678, A2 => i_RD1_10_port, B1 => n8673, 
                           B2 => i_RD1_9_port, ZN => n8842);
   U11730 : INV_X1 port map( A => n8672, ZN => n8673);
   U11731 : AOI21_X1 port map( B1 => n10211, B2 => n8569, A => n8671, ZN => 
                           n8678);
   U11732 : AND2_X1 port map( A1 => n7768, A2 => i_RD2_10_port, ZN => n8671);
   U11733 : AOI22_X1 port map( A1 => n8667, A2 => n10349, B1 => n8672, B2 => 
                           n8666, ZN => n8803);
   U11734 : INV_X1 port map( A => i_RD1_9_port, ZN => n8666);
   U11735 : NAND2_X1 port map( A1 => n8665, A2 => n8664, ZN => n8672);
   U11736 : NAND2_X1 port map( A1 => n7768, A2 => i_RD2_9_port, ZN => n8664);
   U11737 : NAND2_X1 port map( A1 => n10181, A2 => n8569, ZN => n8665);
   U11738 : AOI21_X1 port map( B1 => n8423, B2 => IRAM_ADDRESS_9_port, A => 
                           n8662, ZN => n8663);
   U11739 : NOR2_X1 port map( A1 => n7621, A2 => n550, ZN => n8662);
   U11740 : INV_X1 port map( A => i_RD1_8_port, ZN => n10349);
   U11741 : INV_X1 port map( A => n8661, ZN => n8667);
   U11742 : OAI211_X1 port map( C1 => n8660, C2 => n8659, A => n8658, B => 
                           n8810, ZN => n8668);
   U11743 : NAND2_X1 port map( A1 => n8661, A2 => i_RD1_8_port, ZN => n8810);
   U11744 : OAI21_X1 port map( B1 => n10182, B2 => n7768, A => n8657, ZN => 
                           n8661);
   U11745 : NAND2_X1 port map( A1 => n7768, A2 => n8656, ZN => n8657);
   U11746 : INV_X1 port map( A => i_RD2_8_port, ZN => n8656);
   U11747 : INV_X1 port map( A => n8654, ZN => n8660);
   U11748 : AOI21_X1 port map( B1 => n8653, B2 => n8652, A => n8812, ZN => 
                           n8669);
   U11749 : NAND4_X1 port map( A1 => n8659, A2 => n8658, A3 => n8654, A4 => 
                           n8651, ZN => n8812);
   U11750 : NAND2_X1 port map( A1 => n8650, A2 => n8649, ZN => n8651);
   U11751 : INV_X1 port map( A => i_RD1_6_port, ZN => n8649);
   U11752 : INV_X1 port map( A => n8648, ZN => n8650);
   U11753 : NAND2_X1 port map( A1 => n8647, A2 => n10354, ZN => n8654);
   U11754 : INV_X1 port map( A => i_RD1_7_port, ZN => n10354);
   U11755 : INV_X1 port map( A => n8646, ZN => n8647);
   U11756 : NAND2_X1 port map( A1 => n8646, A2 => i_RD1_7_port, ZN => n8658);
   U11757 : AOI21_X1 port map( B1 => n10183, B2 => n8569, A => n8645, ZN => 
                           n8646);
   U11758 : AND2_X1 port map( A1 => n7768, A2 => i_RD2_7_port, ZN => n8645);
   U11759 : AOI21_X1 port map( B1 => n8423, B2 => IRAM_ADDRESS_7_port, A => 
                           n8643, ZN => n8644);
   U11760 : NOR2_X1 port map( A1 => n7621, A2 => n548, ZN => n8643);
   U11761 : NAND2_X1 port map( A1 => n8648, A2 => i_RD1_6_port, ZN => n8659);
   U11762 : AOI21_X1 port map( B1 => n10209, B2 => n8569, A => n8642, ZN => 
                           n8648);
   U11763 : AND2_X1 port map( A1 => n7768, A2 => i_RD2_6_port, ZN => n8642);
   U11764 : BUF_X1 port map( A => n8420, Z => n8423);
   U11765 : NAND2_X1 port map( A1 => n8640, A2 => i_RD1_5_port, ZN => n8652);
   U11766 : INV_X1 port map( A => n8639, ZN => n8640);
   U11767 : XNOR2_X1 port map( A => n8639, B => i_RD1_5_port, ZN => n8851);
   U11768 : NAND2_X1 port map( A1 => n8638, A2 => n8637, ZN => n8639);
   U11769 : NAND2_X1 port map( A1 => n7768, A2 => i_RD2_5_port, ZN => n8637);
   U11770 : NAND2_X1 port map( A1 => n10184, A2 => n8569, ZN => n8638);
   U11771 : AOI21_X1 port map( B1 => n8423, B2 => IRAM_ADDRESS_5_port, A => 
                           n8635, ZN => n8636);
   U11772 : NOR2_X1 port map( A1 => n7621, A2 => n546, ZN => n8635);
   U11773 : AND2_X1 port map( A1 => n8634, A2 => i_RD1_4_port, ZN => n8843);
   U11774 : OAI22_X1 port map( A1 => i_RD1_3_port, A2 => n8630, B1 => n8634, B2
                           => i_RD1_4_port, ZN => n8631);
   U11775 : OAI21_X1 port map( B1 => n10207, B2 => n7768, A => n8629, ZN => 
                           n8634);
   U11776 : NAND2_X1 port map( A1 => n7768, A2 => n8628, ZN => n8629);
   U11777 : INV_X1 port map( A => i_RD2_4_port, ZN => n8628);
   U11778 : OAI211_X1 port map( C1 => n7621, C2 => n8266, A => n8627, B => 
                           n8626, ZN => n10207);
   U11779 : NAND2_X1 port map( A1 => n10187, A2 => n8190, ZN => n8625);
   U11780 : INV_X1 port map( A => n10402, ZN => n10194);
   U11781 : NAND2_X1 port map( A1 => n8423, A2 => IRAM_ADDRESS_4_port, ZN => 
                           n8627);
   U11782 : AND2_X1 port map( A1 => n8802, A2 => n8807, ZN => n8632);
   U11783 : NAND2_X1 port map( A1 => n8630, A2 => i_RD1_3_port, ZN => n8807);
   U11784 : AOI21_X1 port map( B1 => n10205, B2 => n8569, A => n8624, ZN => 
                           n8630);
   U11785 : AND2_X1 port map( A1 => n7768, A2 => i_RD2_3_port, ZN => n8624);
   U11786 : AOI21_X1 port map( B1 => n8420, B2 => IRAM_ADDRESS_3_port, A => 
                           n8622, ZN => n8623);
   U11787 : NOR2_X1 port map( A1 => n7621, A2 => n544, ZN => n8622);
   U11788 : NAND2_X1 port map( A1 => n8620, A2 => n8619, ZN => n8633);
   U11789 : NAND2_X1 port map( A1 => n8621, A2 => n7896, ZN => n8619);
   U11790 : NAND2_X1 port map( A1 => n7768, A2 => i_RD2_2_port, ZN => n8617);
   U11791 : NAND2_X1 port map( A1 => n8615, A2 => n8809, ZN => n8620);
   U11792 : NAND2_X1 port map( A1 => n8614, A2 => i_RD1_1_port, ZN => n8809);
   U11793 : OAI21_X1 port map( B1 => n8614, B2 => i_RD1_1_port, A => n8613, ZN 
                           => n8615);
   U11794 : AOI21_X1 port map( B1 => i_SEL_CMPB, B2 => n8835, A => i_RD1_0_port
                           , ZN => n8612);
   U11795 : INV_X1 port map( A => i_RD2_0_port, ZN => n8835);
   U11796 : AOI21_X1 port map( B1 => n8420, B2 => IRAM_ADDRESS_0_port, A => 
                           n8610, ZN => n8611);
   U11797 : NOR2_X1 port map( A1 => n7621, A2 => n541, ZN => n8610);
   U11798 : OAI21_X1 port map( B1 => n10203, B2 => n7768, A => n8609, ZN => 
                           n8614);
   U11799 : NAND2_X1 port map( A1 => n7768, A2 => n8608, ZN => n8609);
   U11800 : INV_X1 port map( A => i_RD2_1_port, ZN => n8608);
   U11801 : AOI21_X1 port map( B1 => n8420, B2 => IRAM_ADDRESS_1_port, A => 
                           n8606, ZN => n8607);
   U11802 : NOR2_X1 port map( A1 => n7621, A2 => n542, ZN => n8606);
   U11803 : NAND2_X1 port map( A1 => n10128, A2 => IR_29_port, ZN => n8903);
   U11804 : OAI21_X1 port map( B1 => IR_26_port, B2 => n8237, A => n8598, ZN =>
                           n8595);
   U11805 : NAND2_X1 port map( A1 => n161, A2 => n163, ZN => n8596);
   U11806 : NAND2_X1 port map( A1 => n10421, A2 => n10187, ZN => 
                           CU_I_CW_MUXA_SEL_port);
   U11807 : NAND2_X1 port map( A1 => n10374, A2 => n10393, ZN => n10187);
   U11808 : NAND2_X1 port map( A1 => n8195, A2 => n8396, ZN => n8890);
   U11809 : NAND2_X1 port map( A1 => n10389, A2 => n8396, ZN => n8599);
   U11810 : NAND2_X1 port map( A1 => n8587, A2 => n8354, ZN => n8600);
   U11811 : AND2_X1 port map( A1 => IR_26_port, A2 => n10149, ZN => n10393);
   U11812 : AND2_X1 port map( A1 => n8230, A2 => n465, ZN => n10436);
   U11813 : NOR2_X1 port map( A1 => n11818, A2 => n8203, ZN => n11996);
   U11814 : NOR2_X1 port map( A1 => n8381, A2 => n10444, ZN => n8364);
   U11815 : OAI211_X1 port map( C1 => n11800, C2 => n10444, A => n8363, B => 
                           n8380, ZN => n8365);
   U11816 : OR2_X1 port map( A1 => n8358, A2 => n10444, ZN => n8363);
   U11817 : NAND2_X1 port map( A1 => n8220, A2 => n8382, ZN => n8375);
   U11818 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n711, B => n9567, ZN => 
                           n9110);
   U11819 : INV_X1 port map( A => n9197, ZN => n9202);
   U11820 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1119, B => n9754, ZN =>
                           n9089);
   U11821 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n1221, B => n9807, ZN =>
                           n9086);
   U11822 : XNOR2_X1 port map( A => n9872, B => DP_OP_751_130_6421_n1425, ZN =>
                           n9079);
   U11823 : OAI21_X1 port map( B1 => n7817, B2 => DP_OP_751_130_6421_n711, A =>
                           n9108, ZN => n9109);
   U11824 : NAND2_X1 port map( A1 => n8219, A2 => DataPath_RF_c_swin_1_port, ZN
                           => n8192);
   U11825 : XNOR2_X1 port map( A => n9823, B => DP_OP_751_130_6421_n1323, ZN =>
                           n9081);
   U11826 : OAI211_X1 port map( C1 => n9271, C2 => DP_OP_751_130_6421_n1425, A 
                           => n9073, B => n9072, ZN => n9074);
   U11827 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n1629, B2 => n9241, A 
                           => n9068, ZN => n9069);
   U11828 : NOR2_X1 port map( A1 => n7985, A2 => n11879, ZN => n9704);
   U11829 : NAND2_X1 port map( A1 => n10096, A2 => n9370, ZN => n9064);
   U11830 : XNOR2_X1 port map( A => n8560, B => n9241, ZN => n9070);
   U11831 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_16_port, A2 => n7617, 
                           ZN => n9753);
   U11832 : XOR2_X1 port map( A => n8141, B => intadd_1_n3, Z => n8204);
   U11833 : XNOR2_X1 port map( A => intadd_0_n8, B => intadd_0_n1, ZN => n8205)
                           ;
   U11834 : INV_X1 port map( A => n10314, ZN => n8386);
   U11835 : XNOR2_X1 port map( A => intadd_1_n13, B => intadd_1_n1, ZN => n8206
                           );
   U11836 : XNOR2_X1 port map( A => intadd_1_n18, B => intadd_1_n2, ZN => n8207
                           );
   U11837 : XOR2_X1 port map( A => intadd_0_n13, B => intadd_0_n2, Z => n8208);
   U11838 : INV_X1 port map( A => n11853, ZN => n8943);
   U11839 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_19_port, A2 => n7618, 
                           ZN => n9692);
   U11840 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n405, B2 => n7816, A =>
                           n9121, ZN => n9123);
   U11841 : NOR2_X1 port map( A1 => n10503, A2 => n10500, ZN => n8218);
   U11842 : NAND2_X1 port map( A1 => DataPath_i_PIPLIN_A_20_port, A2 => n7618, 
                           ZN => n9312);
   U11843 : OAI21_X1 port map( B1 => DP_OP_751_130_6421_n915, B2 => 
                           DP_OP_751_130_6421_n813, A => n9098, ZN => n9099);
   U11844 : INV_X1 port map( A => DP_OP_751_130_6421_n1119, ZN => n8562);
   U11845 : XNOR2_X1 port map( A => DP_OP_751_130_6421_n813, B => n9637, ZN => 
                           n9105);
   U11846 : NOR2_X1 port map( A1 => n8021, A2 => n8146, ZN => n10099);
   U11847 : OR2_X1 port map( A1 => n11879, A2 => n11882, ZN => n8229);
   U11848 : OR2_X1 port map( A1 => n10336, A2 => n10326, ZN => n8236);
   U11849 : BUF_X1 port map( A => n8420, Z => n8424);
   U11850 : AND2_X1 port map( A1 => intadd_1_n14, A2 => n8222, ZN => n8267);
   U11851 : AND4_X1 port map( A1 => n8726, A2 => n8725, A3 => n8738, A4 => 
                           n8735, ZN => n8269);
   U11852 : NOR2_X1 port map( A1 => n10298, A2 => n7611, ZN => n8270);
   U11853 : AND2_X1 port map( A1 => n10304, A2 => n10256, ZN => n8271);
   U11854 : AND2_X1 port map( A1 => n10303, A2 => n10311, ZN => n8273);
   U11855 : AND2_X1 port map( A1 => n10443, A2 => n8572, ZN => n8277);
   U11856 : INV_X1 port map( A => n9692, ZN => n8434);
   U11857 : OR2_X1 port map( A1 => n11556, A2 => n8191, ZN => n8294);
   U11858 : OR2_X1 port map( A1 => n11583, A2 => n8191, ZN => n8295);
   U11859 : AND3_X1 port map( A1 => n8188, A2 => n9602, A3 => n11852, ZN => 
                           n8303);
   U11860 : XOR2_X1 port map( A => n10427, B => n11856, Z => n8304);
   U11861 : INV_X1 port map( A => n10081, ZN => n10095);
   U11862 : INV_X1 port map( A => n10053, ZN => n10054);
   U11863 : INV_X1 port map( A => n9753, ZN => n8438);
   U11864 : INV_X1 port map( A => i_RD1_10_port, ZN => n8679);
   U11865 : INV_X1 port map( A => i_RD1_12_port, ZN => n8686);
   U11866 : NAND3_X1 port map( A1 => n8362, A2 => n8365, A3 => n8366, ZN => 
                           DP_OP_1091J1_126_6973_n75);
   U11867 : OAI22_X2 port map( A1 => n8529, A2 => n11896, B1 => n11897, B2 => 
                           n8191, ZN => n11504);
   U11868 : OAI22_X2 port map( A1 => n8529, A2 => n11523, B1 => n11524, B2 => 
                           n8191, ZN => n11541);
   U11869 : AOI21_X1 port map( B1 => DataPath_RF_c_win_0_port, B2 => n8242, A 
                           => n8348, ZN => n8347);
   U11870 : XNOR2_X1 port map( A => DataPath_RF_c_win_1_port, B => n824, ZN => 
                           n8348);
   U11871 : INV_X1 port map( A => n8350, ZN => n8349);
   U11872 : OAI21_X1 port map( B1 => n8242, B2 => DataPath_RF_c_win_0_port, A 
                           => n8351, ZN => n8350);
   U11873 : NOR2_X1 port map( A1 => n8353, A2 => n8352, ZN => n8351);
   U11874 : NOR2_X1 port map( A1 => DataPath_RF_c_win_2_port, A2 => n825, ZN =>
                           n8352);
   U11875 : XNOR2_X1 port map( A => DataPath_RF_c_win_3_port, B => n826, ZN => 
                           n8353);
   U11876 : NOR2_X1 port map( A1 => n8375, A2 => n8377, ZN => n8355);
   U11877 : NOR2_X1 port map( A1 => IR_26_port, A2 => n8586, ZN => n8356);
   U11878 : NAND2_X1 port map( A1 => n11803, A2 => n8357, ZN => n8361);
   U11879 : INV_X1 port map( A => n9191, ZN => n8359);
   U11880 : OAI21_X1 port map( B1 => n8361, B2 => n8240, A => n8378, ZN => 
                           n8366);
   U11881 : NAND2_X1 port map( A1 => n11998, A2 => n8364, ZN => n8362);
   U11882 : NAND2_X1 port map( A1 => n8368, A2 => n8367, ZN => n10260);
   U11883 : NAND2_X1 port map( A1 => n10340, A2 => n8369, ZN => n8367);
   U11884 : AOI21_X1 port map( B1 => n8369, B2 => n8370, A => n8270, ZN => 
                           n8368);
   U11885 : NAND2_X1 port map( A1 => n8289, A2 => n8374, ZN => n8373);
   U11886 : INV_X1 port map( A => n10305, ZN => n8374);
   U11887 : NOR2_X1 port map( A1 => n8416, A2 => n11993, ZN => n8380);
   U11888 : NAND2_X1 port map( A1 => DP_OP_1091J1_126_6973_n72, A2 => 
                           DRAMRF_READY, ZN => n8381);
   U11889 : XNOR2_X1 port map( A => DataPath_RF_c_swin_4_port, B => 
                           DataPath_RF_c_win_2_port, ZN => n8382);
   U11890 : INV_X1 port map( A => C620_DATA2_31, ZN => n8383);
   U11891 : OAI22_X1 port map( A1 => n11791, A2 => n8136, B1 => n11790, B2 => 
                           n11788, ZN => n7086);
   U11892 : AOI211_X1 port map( C1 => n10441, C2 => n159, A => n10395, B => 
                           n10394, ZN => n10396);
   U11893 : AOI21_X1 port map( B1 => n8904, B2 => n8903, A => n159, ZN => 
                           n10378);
   U11894 : NOR2_X1 port map( A1 => n8596, A2 => n159, ZN => n10230);
   U11895 : NAND2_X1 port map( A1 => IR_29_port, A2 => n159, ZN => n10392);
   U11896 : NOR3_X1 port map( A1 => n8414, A2 => n8415, A3 => n10442, ZN => 
                           n8413);
   U11897 : AOI22_X1 port map( A1 => n10186, A2 => n7758, B1 => n8543, B2 => 
                           DataPath_i_PIPLIN_IN2_0_port, ZN => n2387);
   U11898 : XNOR2_X1 port map( A => n8934, B => n8929, ZN => n8930);
   U11899 : NAND2_X1 port map( A1 => n10282, A2 => n10287, ZN => n10283);
   U11900 : OAI21_X1 port map( B1 => intadd_0_n18, B2 => n7594, A => 
                           intadd_0_n19, ZN => intadd_0_n17);
   U11901 : AOI21_X1 port map( B1 => n10186, B2 => n8569, A => n8836, ZN => 
                           n8837);
   U11902 : OAI21_X1 port map( B1 => n10186, B2 => n7768, A => n8612, ZN => 
                           n8613);
   U11903 : INV_X1 port map( A => n10435, ZN => n8416);
   U11904 : NOR2_X1 port map( A1 => n8230, A2 => n465, ZN => n10435);
   U11905 : XNOR2_X1 port map( A => n8135, B => n10364, ZN => n10366);
   U11906 : NAND2_X1 port map( A1 => n10415, A2 => n10416, ZN => n10268);
   U11907 : OAI21_X1 port map( B1 => intadd_0_n16, B2 => intadd_0_n14, A => 
                           intadd_0_n15, ZN => intadd_0_n13);
   U11908 : NOR2_X1 port map( A1 => intadd_0_n14, A2 => intadd_0_n11, ZN => 
                           intadd_0_n9);
   U11909 : OAI21_X1 port map( B1 => n8669, B2 => n8668, A => n8803, ZN => 
                           n8682);
   U11910 : AND2_X1 port map( A1 => n8005, A2 => n7903, ZN => n10395);
   U11911 : INV_X1 port map( A => n8005, ZN => n10227);
   U11912 : AOI22_X1 port map( A1 => n10203, A2 => n7758, B1 => n8542, B2 => 
                           DataPath_i_PIPLIN_IN2_1_port, ZN => n10204);
   U11913 : NAND2_X1 port map( A1 => n10339, A2 => n10334, ZN => n10335);
   U11914 : OAI21_X1 port map( B1 => n10339, B2 => n10336, A => n10329, ZN => 
                           n10330);
   U11915 : OAI211_X1 port map( C1 => n8005, C2 => n10386, A => n8281, B => 
                           n8195, ZN => n8597);
   U11916 : NAND2_X1 port map( A1 => intadd_0_B_2_port, A2 => 
                           IRAM_ADDRESS_3_port, ZN => intadd_0_n12);
   U11917 : AOI22_X1 port map( A1 => n10185, A2 => n7758, B1 => n8543, B2 => 
                           DataPath_i_PIPLIN_IN2_2_port, ZN => n2384);
   U11918 : NAND2_X1 port map( A1 => n10185, A2 => n8569, ZN => n8618);
   U11919 : INV_X1 port map( A => n7749, ZN => n8914);
   U11920 : OAI211_X1 port map( C1 => n10341, C2 => n10340, A => n10339, B => 
                           n8194, ZN => n10343);
   U11921 : OAI21_X1 port map( B1 => n10274, B2 => n10273, A => n8194, ZN => 
                           n10278);
   U11922 : NOR2_X1 port map( A1 => n10280, A2 => n10279, ZN => n10274);
   U11923 : AOI21_X1 port map( B1 => n8633, B2 => n8632, A => n8631, ZN => 
                           n8850);
   U11924 : OAI21_X1 port map( B1 => intadd_0_n11, B2 => intadd_0_n15, A => 
                           intadd_0_n12, ZN => intadd_0_n10);
   U11925 : AOI21_X1 port map( B1 => intadd_0_CO, B2 => n10361, A => n10362, ZN
                           => n10358);
   U11926 : NAND2_X1 port map( A1 => n10199, A2 => n7758, ZN => n10201);
   U11927 : XNOR2_X1 port map( A => n10321, B => n10320, ZN => n10323);
   U11928 : NAND2_X1 port map( A1 => n10199, A2 => n8005, ZN => n8857);
   U11929 : NAND4_X1 port map( A1 => n8883, A2 => n8851, A3 => n8850, A4 => 
                           n8849, ZN => n8852);
   U11930 : OAI21_X1 port map( B1 => n8850, B2 => n8843, A => n8851, ZN => 
                           n8653);
   U11931 : XNOR2_X1 port map( A => n8139, B => n8937, ZN => n11844);
   U11932 : XNOR2_X1 port map( A => n8928, B => n8925, ZN => n11839);
   U11933 : XNOR2_X1 port map( A => n10358, B => n10357, ZN => n10360);
   U11934 : XNOR2_X1 port map( A => n8138, B => n10352, ZN => n10353);
   U11935 : NAND2_X1 port map( A1 => n10230, A2 => n7752, ZN => n10221);
   U11936 : AND2_X1 port map( A1 => n7752, A2 => n8396, ZN => n10386);
   U11937 : NOR2_X1 port map( A1 => IR_26_port, A2 => n7752, ZN => n10229);
   U11938 : NAND2_X1 port map( A1 => IR_26_port, A2 => n7752, ZN => n10225);
   U11939 : NAND4_X1 port map( A1 => n10422, A2 => n10421, A3 => n10194, A4 => 
                           n8625, ZN => n8626);
   U11940 : XNOR2_X1 port map( A => n10348, B => n10347, ZN => n10350);
   U11941 : XNOR2_X1 port map( A => n10300, B => n10299, ZN => n10301);
   U11942 : OAI21_X1 port map( B1 => n10317, B2 => n10315, A => n10314, ZN => 
                           n10313);
   U11943 : NOR2_X1 port map( A1 => n8912, A2 => n8913, ZN => n8425);
   U11944 : AOI21_X1 port map( B1 => intadd_1_n23, B2 => intadd_1_n27, A => 
                           intadd_1_n20, ZN => intadd_1_n18);
   U11945 : AOI21_X1 port map( B1 => n8141, B2 => intadd_1_n14, A => 
                           intadd_1_n15, ZN => intadd_1_n13);
   U11946 : AOI22_X1 port map( A1 => n7949, A2 => n8210, B1 => n10401, B2 => 
                           n8305, ZN => n10192);
   U11947 : AOI22_X1 port map( A1 => n7949, A2 => n8282, B1 => n10401, B2 => 
                           IR_24_port, ZN => n10193);
   U11948 : AOI22_X1 port map( A1 => n7949, A2 => n8196, B1 => n10401, B2 => 
                           n8302, ZN => n10198);
   U11949 : AOI22_X1 port map( A1 => n7949, A2 => n8280, B1 => n10401, B2 => 
                           IR_21_port, ZN => n10403);
   U11950 : OR2_X1 port map( A1 => n7880, A2 => n178, ZN => n8931);
   U11951 : OR3_X1 port map( A1 => n7880, A2 => n8199, A3 => n8290, ZN => 
                           n10344);
   U11952 : OAI21_X1 port map( B1 => n7880, B2 => n8199, A => n8290, ZN => 
                           n10345);
   U11953 : NOR2_X1 port map( A1 => n7880, A2 => n8238, ZN => n10346);
   U11954 : NOR3_X1 port map( A1 => n8852, A2 => n8853, A3 => n8854, ZN => 
                           n8855);
   U11955 : AOI22_X1 port map( A1 => n8422, A2 => IRAM_ADDRESS_26_port, B1 => 
                           n10401, B2 => DECODEhw_i_tickcounter_26_port, ZN => 
                           n8775);
   U11956 : AOI22_X1 port map( A1 => n8420, A2 => IRAM_ADDRESS_24_port, B1 => 
                           n10401, B2 => DECODEhw_i_tickcounter_24_port, ZN => 
                           n8787);
   U11957 : OAI21_X1 port map( B1 => n7622, B2 => n178, A => n8695, ZN => 
                           n10217);
   U11958 : AOI22_X1 port map( A1 => n8422, A2 => IRAM_ADDRESS_29_port, B1 => 
                           n10401, B2 => DECODEhw_i_tickcounter_29_port, ZN => 
                           n8822);
   U11959 : OAI21_X1 port map( B1 => n7622, B2 => n8199, A => n8693, ZN => 
                           n10215);
   U11960 : AOI22_X1 port map( A1 => n8421, A2 => IRAM_ADDRESS_14_port, B1 => 
                           n10401, B2 => DECODEhw_i_tickcounter_14_port, ZN => 
                           n8695);
   U11961 : AOI22_X1 port map( A1 => n8424, A2 => IRAM_ADDRESS_22_port, B1 => 
                           n10401, B2 => DECODEhw_i_tickcounter_22_port, ZN => 
                           n8739);
   U11962 : AOI22_X1 port map( A1 => n8424, A2 => IRAM_ADDRESS_31_port, B1 => 
                           n10401, B2 => DECODEhw_i_tickcounter_31_port, ZN => 
                           n8816);
   U11963 : OAI21_X1 port map( B1 => n7622, B2 => n177, A => n8701, ZN => 
                           n10179);
   U11964 : OAI21_X1 port map( B1 => n7622, B2 => n179, A => n8685, ZN => 
                           n10213);
   U11965 : OAI21_X1 port map( B1 => n7622, B2 => n180, A => n8675, ZN => 
                           n10180);
   U11966 : AOI22_X1 port map( A1 => n8422, A2 => IRAM_ADDRESS_20_port, B1 => 
                           n10401, B2 => DECODEhw_i_tickcounter_20_port, ZN => 
                           n8749);
   U11967 : AOI22_X1 port map( A1 => n8422, A2 => IRAM_ADDRESS_18_port, B1 => 
                           n10401, B2 => DECODEhw_i_tickcounter_18_port, ZN => 
                           n8707);
   U11968 : AOI22_X1 port map( A1 => n8421, A2 => IRAM_ADDRESS_16_port, B1 => 
                           n10401, B2 => DECODEhw_i_tickcounter_16_port, ZN => 
                           n8704);
   U11969 : OAI21_X1 port map( B1 => n7622, B2 => n8233, A => n8670, ZN => 
                           n10211);
   U11970 : OAI21_X1 port map( B1 => n7622, B2 => n8241, A => n8663, ZN => 
                           n10181);
   U11971 : OAI21_X1 port map( B1 => n7622, B2 => n8238, A => n8655, ZN => 
                           n10182);
   U11972 : AOI22_X1 port map( A1 => n8421, A2 => IRAM_ADDRESS_10_port, B1 => 
                           n10401, B2 => DECODEhw_i_tickcounter_10_port, ZN => 
                           n8670);
   U11973 : AOI22_X1 port map( A1 => n8424, A2 => IRAM_ADDRESS_8_port, B1 => 
                           n10401, B2 => DECODEhw_i_tickcounter_8_port, ZN => 
                           n8655);
   U11974 : OAI21_X1 port map( B1 => n7622, B2 => n8228, A => n8641, ZN => 
                           n10209);
   U11975 : OAI21_X1 port map( B1 => n7622, B2 => n8234, A => n8644, ZN => 
                           n10183);
   U11976 : OAI21_X1 port map( B1 => n7622, B2 => n8198, A => n8636, ZN => 
                           n10184);
   U11977 : OAI21_X1 port map( B1 => n8140, B2 => n8226, A => n8623, ZN => 
                           n10205);
   U11978 : OAI21_X1 port map( B1 => n8703, B2 => n193, A => n8611, ZN => 
                           n10186);
   U11979 : OAI21_X1 port map( B1 => n8703, B2 => n10160, A => n8607, ZN => 
                           n10203);
   U11980 : AOI22_X1 port map( A1 => n8424, A2 => IRAM_ADDRESS_6_port, B1 => 
                           n10401, B2 => DECODEhw_i_tickcounter_6_port, ZN => 
                           n8641);
   U11981 : OAI21_X1 port map( B1 => n8703, B2 => n8224, A => n8616, ZN => 
                           n10185);
   U11982 : AOI22_X1 port map( A1 => n8420, A2 => IRAM_ADDRESS_2_port, B1 => 
                           n10401, B2 => DECODEhw_i_tickcounter_2_port, ZN => 
                           n8616);
   U11983 : INV_X2 port map( A => n8558, ZN => n8555);
   U11984 : INV_X1 port map( A => n9070, ZN => n8448);
   U11985 : INV_X1 port map( A => n8448, ZN => n8450);
   U11986 : INV_X1 port map( A => n8448, ZN => n8451);
   U11987 : INV_X1 port map( A => intadd_0_n17, ZN => intadd_0_n16);
   U11988 : INV_X1 port map( A => intadd_0_n6, ZN => intadd_0_n21);
   U11989 : INV_X1 port map( A => intadd_0_n11, ZN => intadd_0_n22);
   U11990 : INV_X1 port map( A => intadd_0_n14, ZN => intadd_0_n23);
   U11991 : INV_X1 port map( A => intadd_1_n21, ZN => intadd_1_n27);
   U11992 : INV_X1 port map( A => intadd_1_n22, ZN => intadd_1_n20);
   U11993 : INV_X1 port map( A => intadd_1_n16, ZN => intadd_1_n26);
   U11994 : NAND3_X1 port map( A1 => n8417, A2 => n8584, A3 => n10440, ZN => 
                           n8585);
   U11995 : NAND3_X1 port map( A1 => IR_29_port, A2 => n8588, A3 => n8589, ZN 
                           => n8591);
   U11996 : NAND3_X1 port map( A1 => n8604, A2 => n8597, A3 => n10221, ZN => 
                           n10222);
   U11997 : NAND3_X1 port map( A1 => n8223, A2 => n159, A3 => n10376, ZN => 
                           n8602);
   U11998 : NAND3_X1 port map( A1 => n8732, A2 => n8731, A3 => n8734, ZN => 
                           n8715);
   U11999 : NAND3_X1 port map( A1 => n8736, A2 => n8735, A3 => n8734, ZN => 
                           n8737);
   U12000 : NAND3_X1 port map( A1 => n8748, A2 => n8769, A3 => n8768, ZN => 
                           n8773);
   U12001 : NAND3_X1 port map( A1 => n8757, A2 => n8762, A3 => n8763, ZN => 
                           n8758);
   U12002 : NAND3_X1 port map( A1 => n8815, A2 => n8814, A3 => n8813, ZN => 
                           n8853);
   U12003 : NAND3_X1 port map( A1 => n8842, A2 => n8841, A3 => n8840, ZN => 
                           n8848);
   U12004 : NAND3_X1 port map( A1 => n8846, A2 => n8845, A3 => n8844, ZN => 
                           n8847);
   U12005 : NAND3_X1 port map( A1 => n8879, A2 => n8878, A3 => n8877, ZN => 
                           n8881);
   U12006 : MUX2_X1 port map( A => n8886, B => n8885, S => n8884, Z => n10200);
   U12007 : MUX2_X1 port map( A => n8005, B => n10382, S => n10199, Z => n8892)
                           ;
   U12008 : NAND3_X1 port map( A1 => n8892, A2 => n8891, A3 => n8051, ZN => 
                           n8893);
   U12009 : NAND3_X1 port map( A1 => n10146, A2 => IR_1_port, A3 => n8224, ZN 
                           => n11780);
   U12010 : NAND3_X1 port map( A1 => n10138, A2 => n8910, A3 => n8224, ZN => 
                           n11778);
   U12011 : NAND3_X1 port map( A1 => n10146, A2 => n8910, A3 => n11785, ZN => 
                           n11786);
   U12012 : NAND3_X1 port map( A1 => n8948, A2 => n9056, A3 => n8953, ZN => 
                           n9419);
   U12013 : NAND3_X1 port map( A1 => n8983, A2 => n9056, A3 => n8982, ZN => 
                           n9501);
   U12014 : NAND3_X1 port map( A1 => n8997, A2 => n9056, A3 => n8996, ZN => 
                           n9470);
   U12015 : NAND3_X1 port map( A1 => n9032, A2 => n9056, A3 => n9031, ZN => 
                           n9366);
   U12016 : NAND3_X1 port map( A1 => n9040, A2 => n9039, A3 => n9038, ZN => 
                           n9971);
   U12017 : MUX2_X1 port map( A => n9693, B => n7794, S => n9651, Z => n9098);
   U12018 : MUX2_X1 port map( A => n9601, B => n9935, S => n9567, Z => n9108);
   U12019 : MUX2_X1 port map( A => n9914, B => n10083, S => n9398, Z => n9121);
   U12020 : NAND3_X1 port map( A1 => n10033, A2 => n9169, A3 => n9168, ZN => 
                           n9167);
   U12021 : NAND3_X1 port map( A1 => n9780, A2 => n11854, A3 => n8188, ZN => 
                           n9166);
   U12022 : NAND3_X1 port map( A1 => n9200, A2 => n9199, A3 => n9198, ZN => 
                           n9205);
   U12023 : NAND3_X1 port map( A1 => n9212, A2 => n9211, A3 => n9210, ZN => 
                           n9218);
   U12024 : NAND3_X1 port map( A1 => n9228, A2 => n7788, A3 => n11853, ZN => 
                           n9232);
   U12025 : MUX2_X1 port map( A => n10033, B => n10088, S => n9271, Z => n9262)
                           ;
   U12026 : MUX2_X1 port map( A => n10088, B => n10035, S => n9271, Z => n9272)
                           ;
   U12027 : NAND3_X1 port map( A1 => n9323, A2 => n9455, A3 => n9452, ZN => 
                           n9326);
   U12028 : NAND3_X1 port map( A1 => n10103, A2 => n7806, A3 => n9366, ZN => 
                           n9329);
   U12029 : MUX2_X1 port map( A => n9913, B => n9961, S => n8566, Z => n9415);
   U12030 : MUX2_X1 port map( A => n10088, B => n10035, S => n9441, Z => n9413)
                           ;
   U12031 : MUX2_X1 port map( A => n10082, B => n10036, S => n9441, Z => n9443)
                           ;
   U12032 : XOR2_X1 port map( A => n9458, B => n9456, Z => n9467);
   U12033 : MUX2_X1 port map( A => n10082, B => n10036, S => n9727, Z => n9520)
                           ;
   U12034 : MUX2_X1 port map( A => n10036, B => n10084, S => n9727, Z => n9519)
                           ;
   U12035 : MUX2_X1 port map( A => n9520, B => n9519, S => n9518, Z => n9521);
   U12036 : MUX2_X1 port map( A => n10035, B => n10088, S => n9528, Z => n9566)
                           ;
   U12037 : MUX2_X1 port map( A => n10082, B => n10036, S => n7805, Z => n9529)
                           ;
   U12038 : NAND3_X1 port map( A1 => n9599, A2 => n9598, A3 => n9597, ZN => 
                           n9609);
   U12039 : NAND3_X1 port map( A1 => n10033, A2 => n9601, A3 => n9600, ZN => 
                           n9604);
   U12040 : NAND3_X1 port map( A1 => n10035, A2 => n9602, A3 => 
                           DP_OP_751_130_6421_n711, ZN => n9603);
   U12041 : NAND3_X1 port map( A1 => n9624, A2 => n9724, A3 => n9623, ZN => 
                           n9625);
   U12042 : MUX2_X1 port map( A => n10082, B => n10036, S => n7606, Z => n9639)
                           ;
   U12043 : MUX2_X1 port map( A => n10036, B => n10084, S => n7606, Z => n9638)
                           ;
   U12044 : MUX2_X1 port map( A => n9639, B => n9638, S => n9637, Z => n9640);
   U12045 : MUX2_X1 port map( A => n9653, B => n9652, S => n8433, Z => n9654);
   U12046 : NAND3_X1 port map( A1 => n9719, A2 => n9689, A3 => n9688, ZN => 
                           n9690);
   U12047 : NAND3_X1 port map( A1 => n10052, A2 => n9691, A3 => n9690, ZN => 
                           n9698);
   U12048 : MUX2_X1 port map( A => n10082, B => n10036, S => n7777, Z => n9745)
                           ;
   U12049 : MUX2_X1 port map( A => n10036, B => n10084, S => n7777, Z => n9744)
                           ;
   U12050 : MUX2_X1 port map( A => n9745, B => n9744, S => n9743, Z => n9746);
   U12051 : NAND3_X1 port map( A1 => n10033, A2 => n7727, A3 => n8562, ZN => 
                           n9787);
   U12052 : NAND3_X1 port map( A1 => n10035, A2 => n7983, A3 => 
                           DP_OP_751_130_6421_n1119, ZN => n9786);
   U12053 : XOR2_X1 port map( A => n9804, B => n9802, Z => n9812);
   U12054 : XOR2_X1 port map( A => n9804, B => n9803, Z => n9805);
   U12055 : MUX2_X1 port map( A => n10082, B => n10036, S => n7893, Z => n9809)
                           ;
   U12056 : MUX2_X1 port map( A => n10036, B => n10084, S => n7893, Z => n9808)
                           ;
   U12057 : MUX2_X1 port map( A => n9809, B => n9808, S => n9807, Z => n9810);
   U12058 : MUX2_X1 port map( A => n10033, B => n10088, S => n9821, Z => n9825)
                           ;
   U12059 : MUX2_X1 port map( A => n10035, B => n10088, S => n9822, Z => n9824)
                           ;
   U12060 : MUX2_X1 port map( A => n9825, B => n9824, S => n9823, Z => n9826);
   U12061 : MUX2_X1 port map( A => n10082, B => n10036, S => n9871, Z => n9874)
                           ;
   U12062 : MUX2_X1 port map( A => n10036, B => n10084, S => n9871, Z => n9873)
                           ;
   U12063 : MUX2_X1 port map( A => n9874, B => n9873, S => n9872, Z => n9875);
   U12064 : NAND3_X1 port map( A1 => n9893, A2 => n9892, A3 => n9891, ZN => 
                           n9898);
   U12065 : MUX2_X1 port map( A => n10084, B => n10036, S => n8021, Z => n9894)
                           ;
   U12066 : XOR2_X1 port map( A => n9910, B => n9909, Z => n9911);
   U12067 : NAND3_X1 port map( A1 => n10033, A2 => n9935, A3 => n8402, ZN => 
                           n9938);
   U12068 : NAND3_X1 port map( A1 => n10035, A2 => n9936, A3 => n7817, ZN => 
                           n9937);
   U12069 : XOR2_X1 port map( A => n10076, B => n10073, Z => n10080);
   U12070 : XOR2_X1 port map( A => n10081, B => n7816, Z => n10087);
   U12071 : NAND3_X1 port map( A1 => n7558, A2 => IR_1_port, A3 => n10129, ZN 
                           => n10136);
   U12072 : NAND3_X1 port map( A1 => n10144, A2 => IR_1_port, A3 => n10143, ZN 
                           => n10148);
   U12073 : NAND3_X1 port map( A1 => n7903, A2 => IR_29_port, A3 => n10232, ZN 
                           => n10233);
   U12074 : XOR2_X1 port map( A => n10284, B => n10283, Z => n10286);
   U12075 : XOR2_X1 port map( A => n10290, B => n10289, Z => n10291);
   U12076 : XOR2_X1 port map( A => IRAM_ADDRESS_20_port, B => n10319, Z => 
                           n10320);
   U12077 : XOR2_X1 port map( A => n10331, B => n10330, Z => n10332);
   U12078 : XOR2_X1 port map( A => n10336, B => n10335, Z => n10338);
   U12079 : NAND3_X1 port map( A1 => n7594, A2 => IRAM_ADDRESS_0_port, A3 => 
                           n11845, ZN => n10371);
   DataPath_RF_bus_complete_win_data_0_port <= '0';
   U12081 : NOR2_X1 port map( A1 => n7752, A2 => n8396, ZN => n10441);
   U12082 : NOR2_X1 port map( A1 => n11753, A2 => n6692, ZN => 
                           CU_I_CW_IF_WB_EN_port);
   U12083 : AND2_X1 port map( A1 => n10439, A2 => CU_I_CW_MEM_WB_EN_port, ZN =>
                           CU_I_N304);
   U12084 : AND2_X1 port map( A1 => n10439, A2 => CU_I_CW_MEM_WB_MUX_SEL_port, 
                           ZN => CU_I_N305);
   U12085 : NOR2_X1 port map( A1 => RST, A2 => n8412, ZN => CU_I_N317);
   U12086 : NOR2_X1 port map( A1 => n10437, A2 => RST, ZN => CU_I_N318);
   U12087 : NOR2_X1 port map( A1 => DataPath_RF_PUSH_ADDRGEN_curr_state_0_port,
                           A2 => n838, ZN => n10444);
   U12088 : NAND2_X1 port map( A1 => n10444, A2 => DRAMRF_READY, ZN => n11818);
   U12089 : XOR2_X1 port map( A => DataPath_RF_PUSH_ADDRGEN_curr_state_0_port, 
                           B => n838, Z => n11816);
   U12090 : NOR2_X1 port map( A1 => n8417, A2 => n10961, ZN => n10448);
   U12091 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, B2 => 
                           n10449, ZN => n10474);
   U12092 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, B2 => 
                           n10449, ZN => n10471);
   U12093 : NAND2_X1 port map( A1 => n10474, A2 => n10471, ZN => n10447);
   U12094 : AOI22_X1 port map( A1 => n10445, A2 => n11816, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, B2 => 
                           n10449, ZN => n10492);
   U12095 : AOI22_X1 port map( A1 => n11817, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, B2 => 
                           n10449, ZN => n10491);
   U12096 : NAND2_X1 port map( A1 => n10492, A2 => n10491, ZN => n10452);
   U12097 : NOR2_X1 port map( A1 => n10447, A2 => n10452, ZN => n10479);
   U12098 : AOI22_X1 port map( A1 => n11817, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, B2 => 
                           n10449, ZN => n10463);
   U12099 : AOI22_X1 port map( A1 => n11817, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, B2 => 
                           n10449, ZN => n10469);
   U12100 : NAND2_X1 port map( A1 => n10463, A2 => n10469, ZN => n10451);
   U12101 : INV_X1 port map( A => n10451, ZN => n10446);
   U12102 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, B2 => 
                           n10449, ZN => n10453);
   U12103 : AOI22_X1 port map( A1 => n11817, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, B2 => 
                           n10449, ZN => n10467);
   U12104 : AND2_X1 port map( A1 => n10453, A2 => n10467, ZN => n10450);
   U12105 : NAND2_X1 port map( A1 => n10446, A2 => n10450, ZN => n10481);
   U12106 : OAI21_X1 port map( B1 => n11818, B2 => n8310, A => n8203, ZN => 
                           n10456);
   U12107 : NAND2_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, ZN => 
                           n10963);
   U12108 : OAI21_X1 port map( B1 => n10448, B2 => n8310, A => n10963, ZN => 
                           n10458);
   U12109 : NOR2_X1 port map( A1 => n10456, A2 => n10458, ZN => n10475);
   U12110 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, B2 => 
                           n10449, ZN => n10455);
   U12111 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, B2 => 
                           n10449, ZN => n10459);
   U12112 : NAND2_X1 port map( A1 => n10455, A2 => n10459, ZN => n10477);
   U12113 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, B2 => 
                           n10449, ZN => n10457);
   U12114 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, B2 => 
                           n10449, ZN => n10461);
   U12115 : NAND2_X1 port map( A1 => n10457, A2 => n10461, ZN => n10478);
   U12116 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, B2 => 
                           n10449, ZN => n10465);
   U12117 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, B2 => 
                           n10449, ZN => n10454);
   U12118 : NAND2_X1 port map( A1 => n10465, A2 => n10454, ZN => n10476);
   U12119 : INV_X1 port map( A => n10453, ZN => n10470);
   U12120 : INV_X1 port map( A => n10454, ZN => n10466);
   U12121 : INV_X1 port map( A => n10455, ZN => n10462);
   U12122 : INV_X1 port map( A => n10456, ZN => n10965);
   U12123 : OAI21_X1 port map( B1 => n10965, B2 => n10458, A => n10457, ZN => 
                           n10460);
   U12124 : OAI221_X1 port map( B1 => n10462, B2 => n10461, C1 => n10462, C2 =>
                           n10460, A => n10459, ZN => n10464);
   U12125 : OAI221_X1 port map( B1 => n10466, B2 => n10465, C1 => n10466, C2 =>
                           n10464, A => n10463, ZN => n10468);
   U12126 : OAI221_X1 port map( B1 => n10470, B2 => n10469, C1 => n10470, C2 =>
                           n10468, A => n10467, ZN => n10473);
   U12127 : INV_X1 port map( A => n10471, ZN => n10472);
   U12128 : AOI21_X1 port map( B1 => n10474, B2 => n10473, A => n10472, ZN => 
                           n10494);
   U12129 : NAND2_X1 port map( A1 => n10496, A2 => n10494, ZN => n10486);
   U12130 : NOR2_X1 port map( A1 => n10477, A2 => n10476, ZN => n10482);
   U12131 : INV_X1 port map( A => n10482, ZN => n10483);
   U12132 : NAND2_X1 port map( A1 => n10480, A2 => n10501, ZN => n10498);
   U12133 : NOR2_X1 port map( A1 => n10498, A2 => n10486, ZN => n10811);
   U12134 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_224_port, B1 => 
                           n8460, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_96_port, ZN => 
                           n10490);
   U12135 : INV_X1 port map( A => n10496, ZN => n10495);
   U12136 : NOR2_X1 port map( A1 => n10501, A2 => n10485, ZN => n10816);
   U12137 : NOR2_X1 port map( A1 => n10481, A2 => n10480, ZN => n10484);
   U12138 : NAND2_X1 port map( A1 => n10482, A2 => n10484, ZN => n10500);
   U12139 : NOR2_X1 port map( A1 => n10500, A2 => n10485, ZN => n10815);
   U12140 : AOI22_X1 port map( A1 => n8461, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_192_port, B1 => 
                           n8463, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_448_port, ZN => 
                           n10489);
   U12141 : NAND2_X1 port map( A1 => n10484, A2 => n10483, ZN => n10502);
   U12142 : NOR2_X1 port map( A1 => n10498, A2 => n10485, ZN => n10814);
   U12143 : AOI22_X1 port map( A1 => n10813, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_320_port, B1 => 
                           n10814, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_64_port, ZN => 
                           n10488);
   U12144 : NOR2_X1 port map( A1 => n10500, A2 => n10486, ZN => n10812);
   U12145 : NOR2_X1 port map( A1 => n10502, A2 => n10486, ZN => n10810);
   U12146 : AOI22_X1 port map( A1 => n8466, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_480_port, B1 => 
                           n8468, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_352_port, ZN => 
                           n10487);
   U12147 : NAND4_X1 port map( A1 => n10490, A2 => n10489, A3 => n10488, A4 => 
                           n10487, ZN => n10509);
   U12148 : INV_X1 port map( A => n10491, ZN => n10493);
   U12149 : OAI21_X1 port map( B1 => n10494, B2 => n10493, A => n10492, ZN => 
                           n10497);
   U12150 : NAND2_X1 port map( A1 => n10495, A2 => n10497, ZN => n10503);
   U12151 : AOI22_X1 port map( A1 => n8214, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_384_port, B1 => 
                           n8470, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_32_port, ZN => 
                           n10507);
   U12152 : NOR2_X1 port map( A1 => n10499, A2 => n10502, ZN => n10823);
   U12153 : NOR2_X1 port map( A1 => n10503, A2 => n10498, ZN => n10826);
   U12154 : AOI22_X1 port map( A1 => n8213, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_288_port, B1 => 
                           n8472, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_0_port, ZN => 
                           n10506);
   U12155 : NOR2_X1 port map( A1 => n10499, A2 => n10501, ZN => n10822);
   U12156 : NOR2_X1 port map( A1 => n10500, A2 => n10499, ZN => n10827);
   U12157 : AOI22_X1 port map( A1 => n8473, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_160_port, B1 => 
                           n8474, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_416_port, ZN => 
                           n10505);
   U12158 : NOR2_X1 port map( A1 => n10503, A2 => n10502, ZN => n10825);
   U12159 : AOI22_X1 port map( A1 => n10828, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_128_port, B1 => 
                           n10825, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_256_port, ZN => 
                           n10504);
   U12160 : NAND4_X1 port map( A1 => n10507, A2 => n10506, A3 => n10505, A4 => 
                           n10504, ZN => n10508);
   U12161 : OR2_X1 port map( A1 => n10509, A2 => n10508, ZN => 
                           DRAMRF_DATA_OUT(0));
   U12162 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_234_port, B1 => 
                           n10814, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_74_port, ZN => 
                           n10513);
   U12163 : AOI22_X1 port map( A1 => n8461, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_202_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_330_port, ZN => 
                           n10512);
   U12164 : AOI22_X1 port map( A1 => n10815, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_458_port, B1 => 
                           n10812, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_490_port, ZN => 
                           n10511);
   U12165 : AOI22_X1 port map( A1 => n8212, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_106_port, B1 => 
                           n8468, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_362_port, ZN => 
                           n10510);
   U12166 : NAND4_X1 port map( A1 => n10513, A2 => n10512, A3 => n10511, A4 => 
                           n10510, ZN => n10519);
   U12167 : AOI22_X1 port map( A1 => n8473, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_170_port, B1 => 
                           n8474, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_426_port, ZN => 
                           n10517);
   U12168 : AOI22_X1 port map( A1 => n8213, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_298_port, B1 => 
                           n8476, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_138_port, ZN => 
                           n10516);
   U12169 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_42_port, B1 => 
                           n8472, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_10_port, ZN => 
                           n10515);
   U12170 : AOI22_X1 port map( A1 => n8214, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_394_port, B1 => 
                           n10825, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_266_port, ZN => 
                           n10514);
   U12171 : NAND4_X1 port map( A1 => n10517, A2 => n10516, A3 => n10515, A4 => 
                           n10514, ZN => n10518);
   U12172 : OR2_X1 port map( A1 => n10519, A2 => n10518, ZN => 
                           DRAMRF_DATA_OUT(10));
   U12173 : AOI22_X1 port map( A1 => n8212, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_107_port, B1 => 
                           n8468, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_363_port, ZN => 
                           n10523);
   U12174 : AOI22_X1 port map( A1 => n8463, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_459_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_331_port, ZN => 
                           n10522);
   U12175 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_235_port, B1 => 
                           n8462, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_203_port, ZN => 
                           n10521);
   U12176 : AOI22_X1 port map( A1 => n8465, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_75_port, B1 => 
                           n10812, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_491_port, ZN => 
                           n10520);
   U12177 : NAND4_X1 port map( A1 => n10523, A2 => n10522, A3 => n10521, A4 => 
                           n10520, ZN => n10529);
   U12178 : AOI22_X1 port map( A1 => n10826, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_11_port, B1 => 
                           n8473, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_171_port, ZN => 
                           n10527);
   U12179 : AOI22_X1 port map( A1 => n8214, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_395_port, B1 => 
                           n10825, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_267_port, ZN => 
                           n10526);
   U12180 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_43_port, B1 => 
                           n8474, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_427_port, ZN => 
                           n10525);
   U12181 : AOI22_X1 port map( A1 => n8213, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_299_port, B1 => 
                           n8476, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_139_port, ZN => 
                           n10524);
   U12182 : NAND4_X1 port map( A1 => n10527, A2 => n10526, A3 => n10525, A4 => 
                           n10524, ZN => n10528);
   U12183 : OR2_X1 port map( A1 => n10529, A2 => n10528, ZN => 
                           DRAMRF_DATA_OUT(11));
   U12184 : AOI22_X1 port map( A1 => n8461, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_204_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_332_port, ZN => 
                           n10533);
   U12185 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_236_port, B1 => 
                           n8460, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_108_port, ZN => 
                           n10532);
   U12186 : AOI22_X1 port map( A1 => n10815, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_460_port, B1 => 
                           n10814, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_76_port, ZN => 
                           n10531);
   U12187 : AOI22_X1 port map( A1 => n8466, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_492_port, B1 => 
                           n8468, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_364_port, ZN => 
                           n10530);
   U12188 : NAND4_X1 port map( A1 => n10533, A2 => n10532, A3 => n10531, A4 => 
                           n10530, ZN => n10539);
   U12189 : AOI22_X1 port map( A1 => n8214, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_396_port, B1 => 
                           n8471, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_300_port, ZN => 
                           n10537);
   U12190 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_44_port, B1 => 
                           n8472, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_12_port, ZN => 
                           n10536);
   U12191 : AOI22_X1 port map( A1 => n8473, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_172_port, B1 => 
                           n8474, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_428_port, ZN => 
                           n10535);
   U12192 : AOI22_X1 port map( A1 => n8476, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_140_port, B1 => 
                           n10825, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_268_port, ZN => 
                           n10534);
   U12193 : NAND4_X1 port map( A1 => n10537, A2 => n10536, A3 => n10535, A4 => 
                           n10534, ZN => n10538);
   U12194 : OR2_X1 port map( A1 => n10539, A2 => n10538, ZN => 
                           DRAMRF_DATA_OUT(12));
   U12195 : AOI22_X1 port map( A1 => n8461, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_205_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_333_port, ZN => 
                           n10543);
   U12196 : AOI22_X1 port map( A1 => n8465, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_77_port, B1 => 
                           n8469, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_365_port, ZN => 
                           n10542);
   U12197 : AOI22_X1 port map( A1 => n8463, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_461_port, B1 => 
                           n10812, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_493_port, ZN => 
                           n10541);
   U12198 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_237_port, B1 => 
                           n8460, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_109_port, ZN => 
                           n10540);
   U12199 : NAND4_X1 port map( A1 => n10543, A2 => n10542, A3 => n10541, A4 => 
                           n10540, ZN => n10549);
   U12200 : AOI22_X1 port map( A1 => n8477, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_269_port, B1 => 
                           n8473, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_173_port, ZN => 
                           n10547);
   U12201 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_45_port, B1 => 
                           n8471, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_301_port, ZN => 
                           n10546);
   U12202 : AOI22_X1 port map( A1 => n8476, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_141_port, B1 => 
                           n8475, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_429_port, ZN => 
                           n10545);
   U12203 : AOI22_X1 port map( A1 => n8215, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_397_port, B1 => 
                           n8472, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_13_port, ZN => 
                           n10544);
   U12204 : NAND4_X1 port map( A1 => n10547, A2 => n10546, A3 => n10545, A4 => 
                           n10544, ZN => n10548);
   U12205 : OR2_X1 port map( A1 => n10549, A2 => n10548, ZN => 
                           DRAMRF_DATA_OUT(13));
   U12206 : AOI22_X1 port map( A1 => n8212, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_110_port, B1 => 
                           n8463, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_462_port, ZN => 
                           n10553);
   U12207 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_238_port, B1 => 
                           n8462, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_206_port, ZN => 
                           n10552);
   U12208 : AOI22_X1 port map( A1 => n8464, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_334_port, B1 => 
                           n10812, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_494_port, ZN => 
                           n10551);
   U12209 : AOI22_X1 port map( A1 => n8465, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_78_port, B1 => 
                           n8469, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_366_port, ZN => 
                           n10550);
   U12210 : NAND4_X1 port map( A1 => n10553, A2 => n10552, A3 => n10551, A4 => 
                           n10550, ZN => n10559);
   U12211 : AOI22_X1 port map( A1 => n8215, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_398_port, B1 => 
                           n8475, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_430_port, ZN => 
                           n10557);
   U12212 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_46_port, B1 => 
                           n8471, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_302_port, ZN => 
                           n10556);
   U12213 : AOI22_X1 port map( A1 => n8477, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_270_port, B1 => 
                           n8473, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_174_port, ZN => 
                           n10555);
   U12214 : AOI22_X1 port map( A1 => n8472, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_14_port, B1 => 
                           n8476, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_142_port, ZN => 
                           n10554);
   U12215 : NAND4_X1 port map( A1 => n10557, A2 => n10556, A3 => n10555, A4 => 
                           n10554, ZN => n10558);
   U12216 : OR2_X1 port map( A1 => n10559, A2 => n10558, ZN => 
                           DRAMRF_DATA_OUT(14));
   U12217 : AOI22_X1 port map( A1 => n8464, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_335_port, B1 => 
                           n8466, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_495_port, ZN => 
                           n10563);
   U12218 : AOI22_X1 port map( A1 => n8212, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_111_port, B1 => 
                           n8463, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_463_port, ZN => 
                           n10562);
   U12219 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_239_port, B1 => 
                           n8469, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_367_port, ZN => 
                           n10561);
   U12220 : AOI22_X1 port map( A1 => n8461, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_207_port, B1 => 
                           n10814, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_79_port, ZN => 
                           n10560);
   U12221 : NAND4_X1 port map( A1 => n10563, A2 => n10562, A3 => n10561, A4 => 
                           n10560, ZN => n10569);
   U12222 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_47_port, B1 => 
                           n8475, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_431_port, ZN => 
                           n10567);
   U12223 : AOI22_X1 port map( A1 => n8476, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_143_port, B1 => 
                           n8477, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_271_port, ZN => 
                           n10566);
   U12224 : AOI22_X1 port map( A1 => n8213, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_303_port, B1 => 
                           n8472, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_15_port, ZN => 
                           n10565);
   U12225 : AOI22_X1 port map( A1 => n8215, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_399_port, B1 => 
                           n8473, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_175_port, ZN => 
                           n10564);
   U12226 : NAND4_X1 port map( A1 => n10567, A2 => n10566, A3 => n10565, A4 => 
                           n10564, ZN => n10568);
   U12227 : OR2_X1 port map( A1 => n10569, A2 => n10568, ZN => 
                           DRAMRF_DATA_OUT(15));
   U12228 : AOI22_X1 port map( A1 => n8461, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_208_port, B1 => 
                           n8463, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_464_port, ZN => 
                           n10573);
   U12229 : AOI22_X1 port map( A1 => n8466, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_496_port, B1 => 
                           n8469, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_368_port, ZN => 
                           n10572);
   U12230 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_240_port, B1 => 
                           n8460, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_112_port, ZN => 
                           n10571);
   U12231 : AOI22_X1 port map( A1 => n8464, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_336_port, B1 => 
                           n8465, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_80_port, ZN => 
                           n10570);
   U12232 : NAND4_X1 port map( A1 => n10573, A2 => n10572, A3 => n10571, A4 => 
                           n10570, ZN => n10579);
   U12233 : AOI22_X1 port map( A1 => n8215, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_400_port, B1 => 
                           n8470, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_48_port, ZN => 
                           n10577);
   U12234 : AOI22_X1 port map( A1 => n8471, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_304_port, B1 => 
                           n8476, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_144_port, ZN => 
                           n10576);
   U12235 : AOI22_X1 port map( A1 => n10826, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_16_port, B1 => 
                           n8217, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_176_port, ZN => 
                           n10575);
   U12236 : AOI22_X1 port map( A1 => n8477, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_272_port, B1 => 
                           n8475, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_432_port, ZN => 
                           n10574);
   U12237 : NAND4_X1 port map( A1 => n10577, A2 => n10576, A3 => n10575, A4 => 
                           n10574, ZN => n10578);
   U12238 : OR2_X1 port map( A1 => n10579, A2 => n10578, ZN => 
                           DRAMRF_DATA_OUT(16));
   U12239 : AOI22_X1 port map( A1 => n10817, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_241_port, B1 => 
                           n8468, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_369_port, ZN => 
                           n10583);
   U12240 : AOI22_X1 port map( A1 => n8461, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_209_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_337_port, ZN => 
                           n10582);
   U12241 : AOI22_X1 port map( A1 => n8463, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_465_port, B1 => 
                           n8465, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_81_port, ZN => 
                           n10581);
   U12242 : AOI22_X1 port map( A1 => n8212, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_113_port, B1 => 
                           n8466, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_497_port, ZN => 
                           n10580);
   U12243 : NAND4_X1 port map( A1 => n10583, A2 => n10582, A3 => n10581, A4 => 
                           n10580, ZN => n10589);
   U12244 : AOI22_X1 port map( A1 => n8472, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_17_port, B1 => 
                           n8474, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_433_port, ZN => 
                           n10587);
   U12245 : AOI22_X1 port map( A1 => n8214, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_401_port, B1 => 
                           n8476, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_145_port, ZN => 
                           n10586);
   U12246 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_49_port, B1 => 
                           n8217, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_177_port, ZN => 
                           n10585);
   U12247 : AOI22_X1 port map( A1 => n8471, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_305_port, B1 => 
                           n8477, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_273_port, ZN => 
                           n10584);
   U12248 : NAND4_X1 port map( A1 => n10587, A2 => n10586, A3 => n10585, A4 => 
                           n10584, ZN => n10588);
   U12249 : OR2_X1 port map( A1 => n10589, A2 => n10588, ZN => 
                           DRAMRF_DATA_OUT(17));
   U12250 : AOI22_X1 port map( A1 => n8466, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_498_port, B1 => 
                           n8468, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_370_port, ZN => 
                           n10593);
   U12251 : AOI22_X1 port map( A1 => n8212, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_114_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_338_port, ZN => 
                           n10592);
   U12252 : AOI22_X1 port map( A1 => n8463, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_466_port, B1 => 
                           n8465, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_82_port, ZN => 
                           n10591);
   U12253 : AOI22_X1 port map( A1 => n10817, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_242_port, B1 => 
                           n8462, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_210_port, ZN => 
                           n10590);
   U12254 : NAND4_X1 port map( A1 => n10593, A2 => n10592, A3 => n10591, A4 => 
                           n10590, ZN => n10599);
   U12255 : AOI22_X1 port map( A1 => n10824, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_50_port, B1 => 
                           n8472, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_18_port, ZN => 
                           n10597);
   U12256 : AOI22_X1 port map( A1 => n8471, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_306_port, B1 => 
                           n8476, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_146_port, ZN => 
                           n10596);
   U12257 : AOI22_X1 port map( A1 => n8214, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_402_port, B1 => 
                           n8217, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_178_port, ZN => 
                           n10595);
   U12258 : AOI22_X1 port map( A1 => n8477, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_274_port, B1 => 
                           n8474, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_434_port, ZN => 
                           n10594);
   U12259 : NAND4_X1 port map( A1 => n10597, A2 => n10596, A3 => n10595, A4 => 
                           n10594, ZN => n10598);
   U12260 : OR2_X1 port map( A1 => n10599, A2 => n10598, ZN => 
                           DRAMRF_DATA_OUT(18));
   U12261 : AOI22_X1 port map( A1 => n8466, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_499_port, B1 => 
                           n8468, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_371_port, ZN => 
                           n10603);
   U12262 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_243_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_339_port, ZN => 
                           n10602);
   U12263 : AOI22_X1 port map( A1 => n8212, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_115_port, B1 => 
                           n8462, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_211_port, ZN => 
                           n10601);
   U12264 : AOI22_X1 port map( A1 => n8463, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_467_port, B1 => 
                           n8465, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_83_port, ZN => 
                           n10600);
   U12265 : NAND4_X1 port map( A1 => n10603, A2 => n10602, A3 => n10601, A4 => 
                           n10600, ZN => n10609);
   U12266 : AOI22_X1 port map( A1 => n8472, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_19_port, B1 => 
                           n8477, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_275_port, ZN => 
                           n10607);
   U12267 : AOI22_X1 port map( A1 => n8476, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_147_port, B1 => 
                           n8217, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_179_port, ZN => 
                           n10606);
   U12268 : AOI22_X1 port map( A1 => n10824, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_51_port, B1 => 
                           n8471, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_307_port, ZN => 
                           n10605);
   U12269 : AOI22_X1 port map( A1 => n8214, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_403_port, B1 => 
                           n8474, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_435_port, ZN => 
                           n10604);
   U12270 : NAND4_X1 port map( A1 => n10607, A2 => n10606, A3 => n10605, A4 => 
                           n10604, ZN => n10608);
   U12271 : OR2_X1 port map( A1 => n10609, A2 => n10608, ZN => 
                           DRAMRF_DATA_OUT(19));
   U12272 : AOI22_X1 port map( A1 => n8212, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_97_port, B1 => 
                           n8465, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_65_port, ZN => 
                           n10613);
   U12273 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_225_port, B1 => 
                           n10813, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_321_port, ZN => 
                           n10612);
   U12274 : AOI22_X1 port map( A1 => n8462, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_193_port, B1 => 
                           n8468, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_353_port, ZN => 
                           n10611);
   U12275 : AOI22_X1 port map( A1 => n10815, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_449_port, B1 => 
                           n8466, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_481_port, ZN => 
                           n10610);
   U12276 : NAND4_X1 port map( A1 => n10613, A2 => n10612, A3 => n10611, A4 => 
                           n10610, ZN => n10619);
   U12277 : AOI22_X1 port map( A1 => n10824, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_33_port, B1 => 
                           n8474, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_417_port, ZN => 
                           n10617);
   U12278 : AOI22_X1 port map( A1 => n8471, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_289_port, B1 => 
                           n10826, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_1_port, ZN => 
                           n10616);
   U12279 : AOI22_X1 port map( A1 => n8214, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_385_port, B1 => 
                           n8477, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_257_port, ZN => 
                           n10615);
   U12280 : AOI22_X1 port map( A1 => n8476, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_129_port, B1 => 
                           n8473, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_161_port, ZN => 
                           n10614);
   U12281 : NAND4_X1 port map( A1 => n10617, A2 => n10616, A3 => n10615, A4 => 
                           n10614, ZN => n10618);
   U12282 : OR2_X1 port map( A1 => n10619, A2 => n10618, ZN => 
                           DRAMRF_DATA_OUT(1));
   U12283 : AOI22_X1 port map( A1 => n8463, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_468_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_340_port, ZN => 
                           n10623);
   U12284 : AOI22_X1 port map( A1 => n8460, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_116_port, B1 => 
                           n8466, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_500_port, ZN => 
                           n10622);
   U12285 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_244_port, B1 => 
                           n10816, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_212_port, ZN => 
                           n10621);
   U12286 : AOI22_X1 port map( A1 => n8465, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_84_port, B1 => 
                           n10810, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_372_port, ZN => 
                           n10620);
   U12287 : NAND4_X1 port map( A1 => n10623, A2 => n10622, A3 => n10621, A4 => 
                           n10620, ZN => n10629);
   U12288 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_52_port, B1 => 
                           n8477, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_276_port, ZN => 
                           n10627);
   U12289 : AOI22_X1 port map( A1 => n8476, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_148_port, B1 => 
                           n10827, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_436_port, ZN => 
                           n10626);
   U12290 : AOI22_X1 port map( A1 => n8218, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_404_port, B1 => 
                           n8472, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_20_port, ZN => 
                           n10625);
   U12291 : AOI22_X1 port map( A1 => n8213, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_308_port, B1 => 
                           n8473, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_180_port, ZN => 
                           n10624);
   U12292 : NAND4_X1 port map( A1 => n10627, A2 => n10626, A3 => n10625, A4 => 
                           n10624, ZN => n10628);
   U12293 : OR2_X1 port map( A1 => n10629, A2 => n10628, ZN => 
                           DRAMRF_DATA_OUT(20));
   U12294 : AOI22_X1 port map( A1 => n10817, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_245_port, B1 => 
                           n8465, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_85_port, ZN => 
                           n10633);
   U12295 : AOI22_X1 port map( A1 => n8460, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_117_port, B1 => 
                           n8463, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_469_port, ZN => 
                           n10632);
   U12296 : AOI22_X1 port map( A1 => n10813, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_341_port, B1 => 
                           n10810, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_373_port, ZN => 
                           n10631);
   U12297 : AOI22_X1 port map( A1 => n8462, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_213_port, B1 => 
                           n8467, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_501_port, ZN => 
                           n10630);
   U12298 : NAND4_X1 port map( A1 => n10633, A2 => n10632, A3 => n10631, A4 => 
                           n10630, ZN => n10639);
   U12299 : AOI22_X1 port map( A1 => n8218, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_405_port, B1 => 
                           n10823, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_309_port, ZN => 
                           n10637);
   U12300 : AOI22_X1 port map( A1 => n10828, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_149_port, B1 => 
                           n10827, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_437_port, ZN => 
                           n10636);
   U12301 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_53_port, B1 => 
                           n8473, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_181_port, ZN => 
                           n10635);
   U12302 : AOI22_X1 port map( A1 => n8472, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_21_port, B1 => 
                           n8477, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_277_port, ZN => 
                           n10634);
   U12303 : NAND4_X1 port map( A1 => n10637, A2 => n10636, A3 => n10635, A4 => 
                           n10634, ZN => n10638);
   U12304 : OR2_X1 port map( A1 => n10639, A2 => n10638, ZN => 
                           DRAMRF_DATA_OUT(21));
   U12305 : AOI22_X1 port map( A1 => n8462, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_214_port, B1 => 
                           n8216, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_86_port, ZN => 
                           n10643);
   U12306 : AOI22_X1 port map( A1 => n8460, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_118_port, B1 => 
                           n8463, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_470_port, ZN => 
                           n10642);
   U12307 : AOI22_X1 port map( A1 => n8464, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_342_port, B1 => 
                           n10810, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_374_port, ZN => 
                           n10641);
   U12308 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_246_port, B1 => 
                           n8467, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_502_port, ZN => 
                           n10640);
   U12309 : NAND4_X1 port map( A1 => n10643, A2 => n10642, A3 => n10641, A4 => 
                           n10640, ZN => n10649);
   U12310 : AOI22_X1 port map( A1 => n8472, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_22_port, B1 => 
                           n8473, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_182_port, ZN => 
                           n10647);
   U12311 : AOI22_X1 port map( A1 => n8213, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_310_port, B1 => 
                           n8478, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_278_port, ZN => 
                           n10646);
   U12312 : AOI22_X1 port map( A1 => n8218, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_406_port, B1 => 
                           n10827, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_438_port, ZN => 
                           n10645);
   U12313 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_54_port, B1 => 
                           n8476, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_150_port, ZN => 
                           n10644);
   U12314 : NAND4_X1 port map( A1 => n10647, A2 => n10646, A3 => n10645, A4 => 
                           n10644, ZN => n10648);
   U12315 : OR2_X1 port map( A1 => n10649, A2 => n10648, ZN => 
                           DRAMRF_DATA_OUT(22));
   U12316 : AOI22_X1 port map( A1 => n8464, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_343_port, B1 => 
                           n10810, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_375_port, ZN => 
                           n10653);
   U12317 : AOI22_X1 port map( A1 => n8460, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_119_port, B1 => 
                           n10816, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_215_port, ZN => 
                           n10652);
   U12318 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_247_port, B1 => 
                           n10815, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_471_port, ZN => 
                           n10651);
   U12319 : AOI22_X1 port map( A1 => n8465, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_87_port, B1 => 
                           n8466, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_503_port, ZN => 
                           n10650);
   U12320 : NAND4_X1 port map( A1 => n10653, A2 => n10652, A3 => n10651, A4 => 
                           n10650, ZN => n10659);
   U12321 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_55_port, B1 => 
                           n10823, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_311_port, ZN => 
                           n10657);
   U12322 : AOI22_X1 port map( A1 => n8218, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_407_port, B1 => 
                           n10827, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_439_port, ZN => 
                           n10656);
   U12323 : AOI22_X1 port map( A1 => n10826, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_23_port, B1 => 
                           n8477, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_279_port, ZN => 
                           n10655);
   U12324 : AOI22_X1 port map( A1 => n10828, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_151_port, B1 => 
                           n8217, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_183_port, ZN => 
                           n10654);
   U12325 : NAND4_X1 port map( A1 => n10657, A2 => n10656, A3 => n10655, A4 => 
                           n10654, ZN => n10658);
   U12326 : OR2_X1 port map( A1 => n10659, A2 => n10658, ZN => 
                           DRAMRF_DATA_OUT(23));
   U12327 : AOI22_X1 port map( A1 => n8464, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_344_port, B1 => 
                           n8466, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_504_port, ZN => 
                           n10663);
   U12328 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_248_port, B1 => 
                           n8468, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_376_port, ZN => 
                           n10662);
   U12329 : AOI22_X1 port map( A1 => n10815, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_472_port, B1 => 
                           n8465, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_88_port, ZN => 
                           n10661);
   U12330 : AOI22_X1 port map( A1 => n8460, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_120_port, B1 => 
                           n10816, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_216_port, ZN => 
                           n10660);
   U12331 : NAND4_X1 port map( A1 => n10663, A2 => n10662, A3 => n10661, A4 => 
                           n10660, ZN => n10669);
   U12332 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_56_port, B1 => 
                           n10823, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_312_port, ZN => 
                           n10667);
   U12333 : AOI22_X1 port map( A1 => n8214, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_408_port, B1 => 
                           n8472, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_24_port, ZN => 
                           n10666);
   U12334 : AOI22_X1 port map( A1 => n8477, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_280_port, B1 => 
                           n8474, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_440_port, ZN => 
                           n10665);
   U12335 : AOI22_X1 port map( A1 => n10828, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_152_port, B1 => 
                           n8217, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_184_port, ZN => 
                           n10664);
   U12336 : NAND4_X1 port map( A1 => n10667, A2 => n10666, A3 => n10665, A4 => 
                           n10664, ZN => n10668);
   U12337 : OR2_X1 port map( A1 => n10669, A2 => n10668, ZN => 
                           DRAMRF_DATA_OUT(24));
   U12338 : AOI22_X1 port map( A1 => n10817, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_249_port, B1 => 
                           n8216, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_89_port, ZN => 
                           n10673);
   U12339 : AOI22_X1 port map( A1 => n8460, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_121_port, B1 => 
                           n8463, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_473_port, ZN => 
                           n10672);
   U12340 : AOI22_X1 port map( A1 => n8462, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_217_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_345_port, ZN => 
                           n10671);
   U12341 : AOI22_X1 port map( A1 => n8466, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_505_port, B1 => 
                           n8468, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_377_port, ZN => 
                           n10670);
   U12342 : NAND4_X1 port map( A1 => n10673, A2 => n10672, A3 => n10671, A4 => 
                           n10670, ZN => n10679);
   U12343 : AOI22_X1 port map( A1 => n8214, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_409_port, B1 => 
                           n8476, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_153_port, ZN => 
                           n10677);
   U12344 : AOI22_X1 port map( A1 => n8472, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_25_port, B1 => 
                           n8474, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_441_port, ZN => 
                           n10676);
   U12345 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_57_port, B1 => 
                           n8217, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_185_port, ZN => 
                           n10675);
   U12346 : AOI22_X1 port map( A1 => n8213, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_313_port, B1 => 
                           n8478, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_281_port, ZN => 
                           n10674);
   U12347 : NAND4_X1 port map( A1 => n10677, A2 => n10676, A3 => n10675, A4 => 
                           n10674, ZN => n10678);
   U12348 : OR2_X1 port map( A1 => n10679, A2 => n10678, ZN => 
                           DRAMRF_DATA_OUT(25));
   U12349 : AOI22_X1 port map( A1 => n10817, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_250_port, B1 => 
                           n10816, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_218_port, ZN => 
                           n10683);
   U12350 : AOI22_X1 port map( A1 => n8460, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_122_port, B1 => 
                           n8216, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_90_port, ZN => 
                           n10682);
   U12351 : AOI22_X1 port map( A1 => n10813, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_346_port, B1 => 
                           n8468, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_378_port, ZN => 
                           n10681);
   U12352 : AOI22_X1 port map( A1 => n8463, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_474_port, B1 => 
                           n8467, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_506_port, ZN => 
                           n10680);
   U12353 : NAND4_X1 port map( A1 => n10683, A2 => n10682, A3 => n10681, A4 => 
                           n10680, ZN => n10689);
   U12354 : AOI22_X1 port map( A1 => n10824, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_58_port, B1 => 
                           n10823, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_314_port, ZN => 
                           n10687);
   U12355 : AOI22_X1 port map( A1 => n8214, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_410_port, B1 => 
                           n8472, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_26_port, ZN => 
                           n10686);
   U12356 : AOI22_X1 port map( A1 => n8476, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_154_port, B1 => 
                           n8474, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_442_port, ZN => 
                           n10685);
   U12357 : AOI22_X1 port map( A1 => n8478, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_282_port, B1 => 
                           n8217, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_186_port, ZN => 
                           n10684);
   U12358 : NAND4_X1 port map( A1 => n10687, A2 => n10686, A3 => n10685, A4 => 
                           n10684, ZN => n10688);
   U12359 : OR2_X1 port map( A1 => n10689, A2 => n10688, ZN => 
                           DRAMRF_DATA_OUT(26));
   U12360 : AOI22_X1 port map( A1 => n8462, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_219_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_347_port, ZN => 
                           n10693);
   U12361 : AOI22_X1 port map( A1 => n8460, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_123_port, B1 => 
                           n8463, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_475_port, ZN => 
                           n10692);
   U12362 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_251_port, B1 => 
                           n8468, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_379_port, ZN => 
                           n10691);
   U12363 : AOI22_X1 port map( A1 => n8216, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_91_port, B1 => 
                           n8467, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_507_port, ZN => 
                           n10690);
   U12364 : NAND4_X1 port map( A1 => n10693, A2 => n10692, A3 => n10691, A4 => 
                           n10690, ZN => n10699);
   U12365 : AOI22_X1 port map( A1 => n8214, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_411_port, B1 => 
                           n8471, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_315_port, ZN => 
                           n10697);
   U12366 : AOI22_X1 port map( A1 => n8476, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_155_port, B1 => 
                           n8478, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_283_port, ZN => 
                           n10696);
   U12367 : AOI22_X1 port map( A1 => n10824, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_59_port, B1 => 
                           n10822, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_187_port, ZN => 
                           n10695);
   U12368 : AOI22_X1 port map( A1 => n10826, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_27_port, B1 => 
                           n8474, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_443_port, ZN => 
                           n10694);
   U12369 : NAND4_X1 port map( A1 => n10697, A2 => n10696, A3 => n10695, A4 => 
                           n10694, ZN => n10698);
   U12370 : OR2_X1 port map( A1 => n10699, A2 => n10698, ZN => 
                           DRAMRF_DATA_OUT(27));
   U12371 : AOI22_X1 port map( A1 => n10815, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_476_port, B1 => 
                           n8216, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_92_port, ZN => 
                           n10703);
   U12372 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_252_port, B1 => 
                           n10811, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_124_port, ZN => 
                           n10702);
   U12373 : AOI22_X1 port map( A1 => n8467, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_508_port, B1 => 
                           n8469, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_380_port, ZN => 
                           n10701);
   U12374 : AOI22_X1 port map( A1 => n8461, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_220_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_348_port, ZN => 
                           n10700);
   U12375 : NAND4_X1 port map( A1 => n10703, A2 => n10702, A3 => n10701, A4 => 
                           n10700, ZN => n10709);
   U12376 : AOI22_X1 port map( A1 => n8215, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_412_port, B1 => 
                           n10828, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_156_port, ZN => 
                           n10707);
   U12377 : AOI22_X1 port map( A1 => n10824, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_60_port, B1 => 
                           n8472, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_28_port, ZN => 
                           n10706);
   U12378 : AOI22_X1 port map( A1 => n8213, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_316_port, B1 => 
                           n8475, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_444_port, ZN => 
                           n10705);
   U12379 : AOI22_X1 port map( A1 => n8478, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_284_port, B1 => 
                           n10822, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_188_port, ZN => 
                           n10704);
   U12380 : NAND4_X1 port map( A1 => n10707, A2 => n10706, A3 => n10705, A4 => 
                           n10704, ZN => n10708);
   U12381 : OR2_X1 port map( A1 => n10709, A2 => n10708, ZN => 
                           DRAMRF_DATA_OUT(28));
   U12382 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_253_port, B1 => 
                           n10811, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_125_port, ZN => 
                           n10713);
   U12383 : AOI22_X1 port map( A1 => n10813, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_349_port, B1 => 
                           n8469, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_381_port, ZN => 
                           n10712);
   U12384 : AOI22_X1 port map( A1 => n8462, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_221_port, B1 => 
                           n8463, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_477_port, ZN => 
                           n10711);
   U12385 : AOI22_X1 port map( A1 => n8216, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_93_port, B1 => 
                           n8467, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_509_port, ZN => 
                           n10710);
   U12386 : NAND4_X1 port map( A1 => n10713, A2 => n10712, A3 => n10711, A4 => 
                           n10710, ZN => n10719);
   U12387 : AOI22_X1 port map( A1 => n10823, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_317_port, B1 => 
                           n10826, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_29_port, ZN => 
                           n10717);
   U12388 : AOI22_X1 port map( A1 => n8215, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_413_port, B1 => 
                           n8478, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_285_port, ZN => 
                           n10716);
   U12389 : AOI22_X1 port map( A1 => n10828, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_157_port, B1 => 
                           n8475, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_445_port, ZN => 
                           n10715);
   U12390 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_61_port, B1 => 
                           n10822, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_189_port, ZN => 
                           n10714);
   U12391 : NAND4_X1 port map( A1 => n10717, A2 => n10716, A3 => n10715, A4 => 
                           n10714, ZN => n10718);
   U12392 : OR2_X1 port map( A1 => n10719, A2 => n10718, ZN => 
                           DRAMRF_DATA_OUT(29));
   U12393 : AOI22_X1 port map( A1 => n10811, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_98_port, B1 => 
                           n8469, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_354_port, ZN => 
                           n10723);
   U12394 : AOI22_X1 port map( A1 => n10817, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_226_port, B1 => 
                           n8467, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_482_port, ZN => 
                           n10722);
   U12395 : AOI22_X1 port map( A1 => n8463, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_450_port, B1 => 
                           n8216, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_66_port, ZN => 
                           n10721);
   U12396 : AOI22_X1 port map( A1 => n8462, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_194_port, B1 => 
                           n10813, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_322_port, ZN => 
                           n10720);
   U12397 : NAND4_X1 port map( A1 => n10723, A2 => n10722, A3 => n10721, A4 => 
                           n10720, ZN => n10729);
   U12398 : AOI22_X1 port map( A1 => n10823, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_290_port, B1 => 
                           n10822, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_162_port, ZN => 
                           n10727);
   U12399 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_34_port, B1 => 
                           n8475, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_418_port, ZN => 
                           n10726);
   U12400 : AOI22_X1 port map( A1 => n8476, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_130_port, B1 => 
                           n8478, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_258_port, ZN => 
                           n10725);
   U12401 : AOI22_X1 port map( A1 => n8215, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_386_port, B1 => 
                           n8472, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_2_port, ZN => 
                           n10724);
   U12402 : NAND4_X1 port map( A1 => n10727, A2 => n10726, A3 => n10725, A4 => 
                           n10724, ZN => n10728);
   U12403 : OR2_X1 port map( A1 => n10729, A2 => n10728, ZN => 
                           DRAMRF_DATA_OUT(2));
   U12404 : AOI22_X1 port map( A1 => n10811, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_126_port, B1 => 
                           n10812, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_510_port, ZN => 
                           n10733);
   U12405 : AOI22_X1 port map( A1 => n8464, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_350_port, B1 => 
                           n10814, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_94_port, ZN => 
                           n10732);
   U12406 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_254_port, B1 => 
                           n8463, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_478_port, ZN => 
                           n10731);
   U12407 : AOI22_X1 port map( A1 => n10816, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_222_port, B1 => 
                           n8469, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_382_port, ZN => 
                           n10730);
   U12408 : NAND4_X1 port map( A1 => n10733, A2 => n10732, A3 => n10731, A4 => 
                           n10730, ZN => n10739);
   U12409 : AOI22_X1 port map( A1 => n10823, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_318_port, B1 => 
                           n8475, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_446_port, ZN => 
                           n10737);
   U12410 : AOI22_X1 port map( A1 => n8472, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_30_port, B1 => 
                           n8217, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_190_port, ZN => 
                           n10736);
   U12411 : AOI22_X1 port map( A1 => n8215, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_414_port, B1 => 
                           n8476, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_158_port, ZN => 
                           n10735);
   U12412 : AOI22_X1 port map( A1 => n10824, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_62_port, B1 => 
                           n10825, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_286_port, ZN => 
                           n10734);
   U12413 : NAND4_X1 port map( A1 => n10737, A2 => n10736, A3 => n10735, A4 => 
                           n10734, ZN => n10738);
   U12414 : OR2_X1 port map( A1 => n10739, A2 => n10738, ZN => 
                           DRAMRF_DATA_OUT(30));
   U12415 : AOI22_X1 port map( A1 => n10811, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_127_port, B1 => 
                           n10812, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_511_port, ZN => 
                           n10743);
   U12416 : AOI22_X1 port map( A1 => n10816, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_223_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_351_port, ZN => 
                           n10742);
   U12417 : AOI22_X1 port map( A1 => n8463, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_479_port, B1 => 
                           n8469, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_383_port, ZN => 
                           n10741);
   U12418 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_255_port, B1 => 
                           n10814, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_95_port, ZN => 
                           n10740);
   U12419 : NAND4_X1 port map( A1 => n10743, A2 => n10742, A3 => n10741, A4 => 
                           n10740, ZN => n10749);
   U12420 : AOI22_X1 port map( A1 => n8215, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_415_port, B1 => 
                           n10826, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_31_port, ZN => 
                           n10747);
   U12421 : AOI22_X1 port map( A1 => n8478, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_287_port, B1 => 
                           n8475, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_447_port, ZN => 
                           n10746);
   U12422 : AOI22_X1 port map( A1 => n8476, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_159_port, B1 => 
                           n8217, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_191_port, ZN => 
                           n10745);
   U12423 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_63_port, B1 => 
                           n8471, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_319_port, ZN => 
                           n10744);
   U12424 : NAND4_X1 port map( A1 => n10747, A2 => n10746, A3 => n10745, A4 => 
                           n10744, ZN => n10748);
   U12425 : OR2_X1 port map( A1 => n10749, A2 => n10748, ZN => 
                           DRAMRF_DATA_OUT(31));
   U12426 : AOI22_X1 port map( A1 => n10816, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_195_port, B1 => 
                           n10813, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_323_port, ZN => 
                           n10753);
   U12427 : AOI22_X1 port map( A1 => n10811, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_99_port, B1 => 
                           n10815, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_451_port, ZN => 
                           n10752);
   U12428 : AOI22_X1 port map( A1 => n8467, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_483_port, B1 => 
                           n8469, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_355_port, ZN => 
                           n10751);
   U12429 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_227_port, B1 => 
                           n10814, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_67_port, ZN => 
                           n10750);
   U12430 : NAND4_X1 port map( A1 => n10753, A2 => n10752, A3 => n10751, A4 => 
                           n10750, ZN => n10759);
   U12431 : AOI22_X1 port map( A1 => n8476, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_131_port, B1 => 
                           n8217, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_163_port, ZN => 
                           n10757);
   U12432 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_35_port, B1 => 
                           n8471, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_291_port, ZN => 
                           n10756);
   U12433 : AOI22_X1 port map( A1 => n8215, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_387_port, B1 => 
                           n8475, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_419_port, ZN => 
                           n10755);
   U12434 : AOI22_X1 port map( A1 => n10826, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_3_port, B1 => 
                           n10825, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_259_port, ZN => 
                           n10754);
   U12435 : NAND4_X1 port map( A1 => n10757, A2 => n10756, A3 => n10755, A4 => 
                           n10754, ZN => n10758);
   U12436 : OR2_X1 port map( A1 => n10759, A2 => n10758, ZN => 
                           DRAMRF_DATA_OUT(3));
   U12437 : AOI22_X1 port map( A1 => n10815, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_452_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_324_port, ZN => 
                           n10763);
   U12438 : AOI22_X1 port map( A1 => n10816, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_196_port, B1 => 
                           n8469, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_356_port, ZN => 
                           n10762);
   U12439 : AOI22_X1 port map( A1 => n10817, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_228_port, B1 => 
                           n10811, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_100_port, ZN => 
                           n10761);
   U12440 : AOI22_X1 port map( A1 => n8216, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_68_port, B1 => 
                           n10812, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_484_port, ZN => 
                           n10760);
   U12441 : NAND4_X1 port map( A1 => n10763, A2 => n10762, A3 => n10761, A4 => 
                           n10760, ZN => n10769);
   U12442 : AOI22_X1 port map( A1 => n8215, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_388_port, B1 => 
                           n8475, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_420_port, ZN => 
                           n10767);
   U12443 : AOI22_X1 port map( A1 => n10828, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_132_port, B1 => 
                           n10825, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_260_port, ZN => 
                           n10766);
   U12444 : AOI22_X1 port map( A1 => n8470, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_36_port, B1 => 
                           n8472, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_4_port, ZN => 
                           n10765);
   U12445 : AOI22_X1 port map( A1 => n10823, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_292_port, B1 => 
                           n8217, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_164_port, ZN => 
                           n10764);
   U12446 : NAND4_X1 port map( A1 => n10767, A2 => n10766, A3 => n10765, A4 => 
                           n10764, ZN => n10768);
   U12447 : OR2_X1 port map( A1 => n10769, A2 => n10768, ZN => 
                           DRAMRF_DATA_OUT(4));
   U12448 : AOI22_X1 port map( A1 => n8467, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_485_port, B1 => 
                           n8469, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_357_port, ZN => 
                           n10773);
   U12449 : AOI22_X1 port map( A1 => n8461, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_197_port, B1 => 
                           n10813, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_325_port, ZN => 
                           n10772);
   U12450 : AOI22_X1 port map( A1 => n8212, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_101_port, B1 => 
                           n10814, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_69_port, ZN => 
                           n10771);
   U12451 : AOI22_X1 port map( A1 => n10817, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_229_port, B1 => 
                           n8463, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_453_port, ZN => 
                           n10770);
   U12452 : NAND4_X1 port map( A1 => n10773, A2 => n10772, A3 => n10771, A4 => 
                           n10770, ZN => n10779);
   U12453 : AOI22_X1 port map( A1 => n10824, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_37_port, B1 => 
                           n8476, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_133_port, ZN => 
                           n10777);
   U12454 : AOI22_X1 port map( A1 => n8213, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_293_port, B1 => 
                           n10826, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_5_port, ZN => 
                           n10776);
   U12455 : AOI22_X1 port map( A1 => n8215, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_389_port, B1 => 
                           n8475, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_421_port, ZN => 
                           n10775);
   U12456 : AOI22_X1 port map( A1 => n8478, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_261_port, B1 => 
                           n10822, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_165_port, ZN => 
                           n10774);
   U12457 : NAND4_X1 port map( A1 => n10777, A2 => n10776, A3 => n10775, A4 => 
                           n10774, ZN => n10778);
   U12458 : OR2_X1 port map( A1 => n10779, A2 => n10778, ZN => 
                           DRAMRF_DATA_OUT(5));
   U12459 : AOI22_X1 port map( A1 => n8467, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_486_port, B1 => 
                           n10810, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_358_port, ZN => 
                           n10783);
   U12460 : AOI22_X1 port map( A1 => n10813, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_326_port, B1 => 
                           n8216, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_70_port, ZN => 
                           n10782);
   U12461 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_230_port, B1 => 
                           n10811, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_102_port, ZN => 
                           n10781);
   U12462 : AOI22_X1 port map( A1 => n8461, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_198_port, B1 => 
                           n10815, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_454_port, ZN => 
                           n10780);
   U12463 : NAND4_X1 port map( A1 => n10783, A2 => n10782, A3 => n10781, A4 => 
                           n10780, ZN => n10789);
   U12464 : AOI22_X1 port map( A1 => n8218, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_390_port, B1 => 
                           n10822, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_166_port, ZN => 
                           n10787);
   U12465 : AOI22_X1 port map( A1 => n8213, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_294_port, B1 => 
                           n10827, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_422_port, ZN => 
                           n10786);
   U12466 : AOI22_X1 port map( A1 => n10824, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_38_port, B1 => 
                           n8476, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_134_port, ZN => 
                           n10785);
   U12467 : AOI22_X1 port map( A1 => n8472, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_6_port, B1 => 
                           n10825, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_262_port, ZN => 
                           n10784);
   U12468 : NAND4_X1 port map( A1 => n10787, A2 => n10786, A3 => n10785, A4 => 
                           n10784, ZN => n10788);
   U12469 : OR2_X1 port map( A1 => n10789, A2 => n10788, ZN => 
                           DRAMRF_DATA_OUT(6));
   U12470 : AOI22_X1 port map( A1 => n10817, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_231_port, B1 => 
                           n8464, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_327_port, ZN => 
                           n10793);
   U12471 : AOI22_X1 port map( A1 => n8212, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_103_port, B1 => 
                           n8463, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_455_port, ZN => 
                           n10792);
   U12472 : AOI22_X1 port map( A1 => n8216, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_71_port, B1 => 
                           n10812, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_487_port, ZN => 
                           n10791);
   U12473 : AOI22_X1 port map( A1 => n8461, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_199_port, B1 => 
                           n10810, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_359_port, ZN => 
                           n10790);
   U12474 : NAND4_X1 port map( A1 => n10793, A2 => n10792, A3 => n10791, A4 => 
                           n10790, ZN => n10799);
   U12475 : AOI22_X1 port map( A1 => n10824, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_39_port, B1 => 
                           n8471, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_295_port, ZN => 
                           n10797);
   U12476 : AOI22_X1 port map( A1 => n8472, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_7_port, B1 => 
                           n10827, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_423_port, ZN => 
                           n10796);
   U12477 : AOI22_X1 port map( A1 => n8218, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_391_port, B1 => 
                           n10822, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_167_port, ZN => 
                           n10795);
   U12478 : AOI22_X1 port map( A1 => n10828, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_135_port, B1 => 
                           n8478, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_263_port, ZN => 
                           n10794);
   U12479 : NAND4_X1 port map( A1 => n10797, A2 => n10796, A3 => n10795, A4 => 
                           n10794, ZN => n10798);
   U12480 : OR2_X1 port map( A1 => n10799, A2 => n10798, ZN => 
                           DRAMRF_DATA_OUT(7));
   U12481 : AOI22_X1 port map( A1 => n8464, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_328_port, B1 => 
                           n8216, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_72_port, ZN => 
                           n10803);
   U12482 : AOI22_X1 port map( A1 => n8459, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_232_port, B1 => 
                           n10810, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_360_port, ZN => 
                           n10802);
   U12483 : AOI22_X1 port map( A1 => n8461, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_200_port, B1 => 
                           n10815, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_456_port, ZN => 
                           n10801);
   U12484 : AOI22_X1 port map( A1 => n8212, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_104_port, B1 => 
                           n8467, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_488_port, ZN => 
                           n10800);
   U12485 : NAND4_X1 port map( A1 => n10803, A2 => n10802, A3 => n10801, A4 => 
                           n10800, ZN => n10809);
   U12486 : AOI22_X1 port map( A1 => n8473, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_168_port, B1 => 
                           n10827, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_424_port, ZN => 
                           n10807);
   U12487 : AOI22_X1 port map( A1 => n8213, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_296_port, B1 => 
                           n8478, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_264_port, ZN => 
                           n10806);
   U12488 : AOI22_X1 port map( A1 => n10826, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_8_port, B1 => 
                           n10828, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_136_port, ZN => 
                           n10805);
   U12489 : AOI22_X1 port map( A1 => n8218, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_392_port, B1 => 
                           n8470, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_40_port, ZN => 
                           n10804);
   U12490 : NAND4_X1 port map( A1 => n10807, A2 => n10806, A3 => n10805, A4 => 
                           n10804, ZN => n10808);
   U12491 : OR2_X1 port map( A1 => n10809, A2 => n10808, ZN => 
                           DRAMRF_DATA_OUT(8));
   U12492 : AOI22_X1 port map( A1 => n8212, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_105_port, B1 => 
                           n10810, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_361_port, ZN => 
                           n10821);
   U12493 : AOI22_X1 port map( A1 => n10813, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_329_port, B1 => 
                           n8467, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_489_port, ZN => 
                           n10820);
   U12494 : AOI22_X1 port map( A1 => n8463, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_457_port, B1 => 
                           n8216, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_73_port, ZN => 
                           n10819);
   U12495 : AOI22_X1 port map( A1 => n10817, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_233_port, B1 => 
                           n8462, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_201_port, ZN => 
                           n10818);
   U12496 : NAND4_X1 port map( A1 => n10821, A2 => n10820, A3 => n10819, A4 => 
                           n10818, ZN => n10834);
   U12497 : AOI22_X1 port map( A1 => n8213, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_297_port, B1 => 
                           n10822, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_169_port, ZN => 
                           n10832);
   U12498 : AOI22_X1 port map( A1 => n8218, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_393_port, B1 => 
                           n8470, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_41_port, ZN => 
                           n10831);
   U12499 : AOI22_X1 port map( A1 => n8472, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_9_port, B1 => 
                           n8478, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_265_port, ZN => 
                           n10830);
   U12500 : AOI22_X1 port map( A1 => n10828, A2 => 
                           DataPath_RF_bus_sel_savedwin_data_137_port, B1 => 
                           n10827, B2 => 
                           DataPath_RF_bus_sel_savedwin_data_425_port, ZN => 
                           n10829);
   U12501 : NAND4_X1 port map( A1 => n10832, A2 => n10831, A3 => n10830, A4 => 
                           n10829, ZN => n10833);
   U12502 : OR2_X1 port map( A1 => n10834, A2 => n10833, ZN => 
                           DRAMRF_DATA_OUT(9));
   U12503 : OR2_X1 port map( A1 => n11832, A2 => n8291, ZN => n11820);
   U12504 : NAND2_X1 port map( A1 => n11449, A2 => n11820, ZN => n11995);
   U12505 : INV_X1 port map( A => n11995, ZN => DRAMRF_READNOTWRITE);
   U12506 : NOR2_X1 port map( A1 => n494, A2 => n376, ZN => DRAM_ADDRESS_0_port
                           );
   U12507 : AOI21_X1 port map( B1 => n376, B2 => n375, A => n495, ZN => 
                           DRAM_ADDRESS_1_port);
   U12508 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(8), B1 =>
                           DataPath_i_REG_ME_DATA_DATAMEM_8_port, B2 => n8293, 
                           ZN => n10899);
   U12509 : NAND2_X1 port map( A1 => DATA_SIZE_1_port, A2 => n375, ZN => n10846
                           );
   U12510 : OAI221_X1 port map( B1 => DATA_SIZE_0_port, B2 => DATA_SIZE_1_port,
                           C1 => n495, C2 => DATA_SIZE_1_port, A => 
                           i_DATAMEM_RM, ZN => n10835);
   U12511 : NAND4_X1 port map( A1 => n494, A2 => n10945, A3 => n10902, A4 => 
                           n8285, ZN => n10880);
   U12512 : NAND3_X1 port map( A1 => i_DATAMEM_RM, A2 => n495, A3 => n10945, ZN
                           => n10838);
   U12513 : NOR2_X1 port map( A1 => n8278, A2 => n10838, ZN => n10875);
   U12514 : MUX2_X1 port map( A => DRAM_DATA_IN(24), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_24_port, S => n8293, 
                           Z => n10935);
   U12515 : AOI22_X1 port map( A1 => n10875, A2 => n10935, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_0_port, B2 => n8293, 
                           ZN => n10840);
   U12516 : NOR2_X1 port map( A1 => n495, A2 => n10846, ZN => n10836);
   U12517 : AOI21_X1 port map( B1 => n10836, B2 => n8278, A => n10835, ZN => 
                           n10837);
   U12518 : NOR2_X1 port map( A1 => n10837, A2 => n8293, ZN => n10877);
   U12519 : NOR2_X1 port map( A1 => n375, A2 => DATA_SIZE_1_port, ZN => n10871)
                           ;
   U12520 : NAND3_X1 port map( A1 => i_DATAMEM_RM, A2 => n495, A3 => n10871, ZN
                           => n10867);
   U12521 : OAI21_X1 port map( B1 => n494, B2 => n10838, A => n10867, ZN => 
                           n10876);
   U12522 : MUX2_X1 port map( A => DRAM_DATA_IN(16), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_16_port, S => n8293, 
                           Z => n10873);
   U12523 : AOI22_X1 port map( A1 => n10877, A2 => DRAM_DATA_IN(0), B1 => 
                           n10876, B2 => n10873, ZN => n10839);
   U12524 : OAI211_X1 port map( C1 => n10899, C2 => n10880, A => n10840, B => 
                           n10839, ZN => DRAM_DATA_OUT_0_port);
   U12525 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(15), B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_15_port, B2 => 
                           n8293, ZN => n10868);
   U12526 : MUX2_X1 port map( A => DRAM_DATA_IN(31), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_31_port, S => n8293, 
                           Z => n10866);
   U12527 : AOI22_X1 port map( A1 => n10875, A2 => n10866, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_7_port, B2 => n8293, 
                           ZN => n10842);
   U12528 : MUX2_X1 port map( A => DRAM_DATA_IN(23), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_23_port, S => n8293, 
                           Z => n10894);
   U12529 : AOI22_X1 port map( A1 => n10877, A2 => DRAM_DATA_IN(7), B1 => 
                           n10894, B2 => n10876, ZN => n10841);
   U12530 : OAI211_X1 port map( C1 => n10868, C2 => n10880, A => n10842, B => 
                           n10841, ZN => DRAM_DATA_OUT_7_port);
   U12531 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(10), B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_10_port, B2 => 
                           n8293, ZN => n10845);
   U12532 : MUX2_X1 port map( A => DRAM_DATA_IN(26), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_26_port, S => n8293, 
                           Z => n10905);
   U12533 : AOI22_X1 port map( A1 => n10875, A2 => n10905, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_2_port, B2 => n8293, 
                           ZN => n10844);
   U12534 : MUX2_X1 port map( A => DRAM_DATA_IN(18), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_18_port, S => n8293, 
                           Z => n10883);
   U12535 : AOI22_X1 port map( A1 => n10877, A2 => DRAM_DATA_IN(2), B1 => 
                           n10876, B2 => n10883, ZN => n10843);
   U12536 : OAI211_X1 port map( C1 => n10845, C2 => n10880, A => n10844, B => 
                           n10843, ZN => DRAM_DATA_OUT_2_port);
   U12537 : NOR2_X1 port map( A1 => n10902, A2 => n10845, ZN => n10906);
   U12538 : AOI21_X1 port map( B1 => n10940, B2 => n10905, A => n10906, ZN => 
                           n10847);
   U12539 : NAND3_X1 port map( A1 => n10945, A2 => n212, A3 => 
                           DRAM_DATA_OUT_7_port, ZN => n10896);
   U12540 : AOI21_X1 port map( B1 => n10941, B2 => DRAM_DATA_OUT_2_port, A => 
                           n10898, ZN => n10908);
   U12541 : OAI21_X1 port map( B1 => n10945, B2 => n10847, A => n10908, ZN => 
                           DRAM_DATA_OUT_10_port);
   U12542 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(11), B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_11_port, B2 => 
                           n8293, ZN => n10850);
   U12543 : MUX2_X1 port map( A => DRAM_DATA_IN(27), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_27_port, S => n8293, 
                           Z => n10910);
   U12544 : AOI22_X1 port map( A1 => n10875, A2 => n10910, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_3_port, B2 => n8293, 
                           ZN => n10849);
   U12545 : MUX2_X1 port map( A => DRAM_DATA_IN(19), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_19_port, S => n8293, 
                           Z => n10885);
   U12546 : AOI22_X1 port map( A1 => n10877, A2 => DRAM_DATA_IN(3), B1 => 
                           n10876, B2 => n10885, ZN => n10848);
   U12547 : OAI211_X1 port map( C1 => n10850, C2 => n10880, A => n10849, B => 
                           n10848, ZN => DRAM_DATA_OUT_3_port);
   U12548 : NOR2_X1 port map( A1 => n10902, A2 => n10850, ZN => n10909);
   U12549 : AOI21_X1 port map( B1 => n10940, B2 => n10910, A => n10909, ZN => 
                           n10852);
   U12550 : NAND2_X1 port map( A1 => n10941, A2 => DRAM_DATA_OUT_3_port, ZN => 
                           n10851);
   U12551 : INV_X1 port map( A => n10898, ZN => n10942);
   U12552 : OAI211_X1 port map( C1 => n10945, C2 => n10852, A => n10851, B => 
                           n10942, ZN => DRAM_DATA_OUT_11_port);
   U12553 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(12), B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_12_port, B2 => 
                           n8293, ZN => n10855);
   U12554 : MUX2_X1 port map( A => DRAM_DATA_IN(28), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_28_port, S => n8293, 
                           Z => n10913);
   U12555 : AOI22_X1 port map( A1 => n10875, A2 => n10913, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_4_port, B2 => n8293, 
                           ZN => n10854);
   U12556 : MUX2_X1 port map( A => DRAM_DATA_IN(20), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_20_port, S => n8293, 
                           Z => n10887);
   U12557 : AOI22_X1 port map( A1 => n10877, A2 => DRAM_DATA_IN(4), B1 => 
                           n10876, B2 => n10887, ZN => n10853);
   U12558 : OAI211_X1 port map( C1 => n10855, C2 => n10880, A => n10854, B => 
                           n10853, ZN => DRAM_DATA_OUT_4_port);
   U12559 : NOR2_X1 port map( A1 => n10902, A2 => n10855, ZN => n10914);
   U12560 : AOI21_X1 port map( B1 => n10940, B2 => n10913, A => n10914, ZN => 
                           n10856);
   U12561 : AOI21_X1 port map( B1 => n10941, B2 => DRAM_DATA_OUT_4_port, A => 
                           n10898, ZN => n10916);
   U12562 : OAI21_X1 port map( B1 => n10945, B2 => n10856, A => n10916, ZN => 
                           DRAM_DATA_OUT_12_port);
   U12563 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(13), B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_13_port, B2 => 
                           n8293, ZN => n10859);
   U12564 : MUX2_X1 port map( A => DRAM_DATA_IN(29), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_29_port, S => n8293, 
                           Z => n10917);
   U12565 : AOI22_X1 port map( A1 => n10875, A2 => n10917, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_5_port, B2 => n8293, 
                           ZN => n10858);
   U12566 : MUX2_X1 port map( A => DRAM_DATA_IN(21), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_21_port, S => n8293, 
                           Z => n10889);
   U12567 : AOI22_X1 port map( A1 => n10877, A2 => DRAM_DATA_IN(5), B1 => 
                           n10876, B2 => n10889, ZN => n10857);
   U12568 : OAI211_X1 port map( C1 => n10859, C2 => n10880, A => n10858, B => 
                           n10857, ZN => DRAM_DATA_OUT_5_port);
   U12569 : NOR2_X1 port map( A1 => n10902, A2 => n10859, ZN => n10918);
   U12570 : AOI21_X1 port map( B1 => n10940, B2 => n10917, A => n10918, ZN => 
                           n10860);
   U12571 : AOI21_X1 port map( B1 => n10941, B2 => DRAM_DATA_OUT_5_port, A => 
                           n10898, ZN => n10922);
   U12572 : OAI21_X1 port map( B1 => n10945, B2 => n10860, A => n10922, ZN => 
                           DRAM_DATA_OUT_13_port);
   U12573 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(14), B1 
                           => DataPath_i_REG_ME_DATA_DATAMEM_14_port, B2 => 
                           n8293, ZN => n10863);
   U12574 : MUX2_X1 port map( A => DRAM_DATA_IN(30), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_30_port, S => n8293, 
                           Z => n10924);
   U12575 : AOI22_X1 port map( A1 => n10875, A2 => n10924, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_6_port, B2 => n8293, 
                           ZN => n10862);
   U12576 : MUX2_X1 port map( A => DRAM_DATA_IN(22), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_22_port, S => n8293, 
                           Z => n10891);
   U12577 : AOI22_X1 port map( A1 => n10877, A2 => DRAM_DATA_IN(6), B1 => 
                           n10876, B2 => n10891, ZN => n10861);
   U12578 : OAI211_X1 port map( C1 => n10863, C2 => n10880, A => n10862, B => 
                           n10861, ZN => DRAM_DATA_OUT_6_port);
   U12579 : NOR2_X1 port map( A1 => n10902, A2 => n10863, ZN => n10923);
   U12580 : AOI21_X1 port map( B1 => n10940, B2 => n10924, A => n10923, ZN => 
                           n10865);
   U12581 : NAND2_X1 port map( A1 => n10941, A2 => DRAM_DATA_OUT_6_port, ZN => 
                           n10864);
   U12582 : OAI211_X1 port map( C1 => n10945, C2 => n10865, A => n10864, B => 
                           n10942, ZN => DRAM_DATA_OUT_14_port);
   U12583 : INV_X1 port map( A => n10866, ZN => n10933);
   U12584 : OAI22_X1 port map( A1 => n10868, A2 => n10902, B1 => n10933, B2 => 
                           n10867, ZN => n10870);
   U12585 : INV_X1 port map( A => n10870, ZN => n10869);
   U12586 : OAI211_X1 port map( C1 => n212, C2 => n8293, A => n10945, B => 
                           DRAM_DATA_OUT_7_port, ZN => n10931);
   U12587 : OAI21_X1 port map( B1 => n10945, B2 => n10869, A => n10931, ZN => 
                           DRAM_DATA_OUT_15_port);
   U12588 : OAI211_X1 port map( C1 => n212, C2 => n8293, A => n10871, B => 
                           n10870, ZN => n10930);
   U12589 : NOR2_X1 port map( A1 => n8293, A2 => n10930, ZN => n10895);
   U12590 : AOI21_X1 port map( B1 => n376, B2 => n375, A => n8293, ZN => n10872
                           );
   U12591 : NAND2_X1 port map( A1 => n10871, A2 => n8293, ZN => n10927);
   U12592 : INV_X1 port map( A => n10927, ZN => n10919);
   U12593 : AOI22_X1 port map( A1 => n10929, A2 => n10873, B1 => 
                           DRAM_DATA_OUT_0_port, B2 => n10893, ZN => n10874);
   U12594 : NAND2_X1 port map( A1 => n10926, A2 => n10874, ZN => 
                           DRAM_DATA_OUT_16_port);
   U12595 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => DRAM_DATA_IN(9), B1 =>
                           DataPath_i_REG_ME_DATA_DATAMEM_9_port, B2 => n8293, 
                           ZN => n10901);
   U12596 : MUX2_X1 port map( A => DRAM_DATA_IN(25), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_25_port, S => n8293, 
                           Z => n10939);
   U12597 : AOI22_X1 port map( A1 => n10875, A2 => n10939, B1 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_1_port, B2 => n8293, 
                           ZN => n10879);
   U12598 : MUX2_X1 port map( A => DRAM_DATA_IN(17), B => 
                           DataPath_i_REG_ME_DATA_DATAMEM_17_port, S => n8293, 
                           Z => n10881);
   U12599 : AOI22_X1 port map( A1 => n10877, A2 => DRAM_DATA_IN(1), B1 => 
                           n10876, B2 => n10881, ZN => n10878);
   U12600 : OAI211_X1 port map( C1 => n10901, C2 => n10880, A => n10879, B => 
                           n10878, ZN => DRAM_DATA_OUT_1_port);
   U12601 : AOI22_X1 port map( A1 => n10929, A2 => n10881, B1 => n10893, B2 => 
                           DRAM_DATA_OUT_1_port, ZN => n10882);
   U12602 : NAND2_X1 port map( A1 => n10926, A2 => n10882, ZN => 
                           DRAM_DATA_OUT_17_port);
   U12603 : AOI22_X1 port map( A1 => n10929, A2 => n10883, B1 => 
                           DRAM_DATA_OUT_2_port, B2 => n10893, ZN => n10884);
   U12604 : NAND2_X1 port map( A1 => n10926, A2 => n10884, ZN => 
                           DRAM_DATA_OUT_18_port);
   U12605 : AOI22_X1 port map( A1 => n10929, A2 => n10885, B1 => n10893, B2 => 
                           DRAM_DATA_OUT_3_port, ZN => n10886);
   U12606 : NAND2_X1 port map( A1 => n10926, A2 => n10886, ZN => 
                           DRAM_DATA_OUT_19_port);
   U12607 : AOI22_X1 port map( A1 => n10929, A2 => n10887, B1 => 
                           DRAM_DATA_OUT_4_port, B2 => n10893, ZN => n10888);
   U12608 : NAND2_X1 port map( A1 => n10926, A2 => n10888, ZN => 
                           DRAM_DATA_OUT_20_port);
   U12609 : AOI22_X1 port map( A1 => n10929, A2 => n10889, B1 => 
                           DRAM_DATA_OUT_5_port, B2 => n10893, ZN => n10890);
   U12610 : NAND2_X1 port map( A1 => n10926, A2 => n10890, ZN => 
                           DRAM_DATA_OUT_21_port);
   U12611 : AOI22_X1 port map( A1 => n10929, A2 => n10891, B1 => n10893, B2 => 
                           DRAM_DATA_OUT_6_port, ZN => n10892);
   U12612 : NAND2_X1 port map( A1 => n10926, A2 => n10892, ZN => 
                           DRAM_DATA_OUT_22_port);
   U12613 : AOI22_X1 port map( A1 => n10929, A2 => n10894, B1 => 
                           DRAM_DATA_OUT_7_port, B2 => n10893, ZN => n10897);
   U12614 : INV_X1 port map( A => n10895, ZN => n10920);
   U12615 : NAND3_X1 port map( A1 => n10897, A2 => n10896, A3 => n10920, ZN => 
                           DRAM_DATA_OUT_23_port);
   U12616 : AOI21_X1 port map( B1 => n10941, B2 => DRAM_DATA_OUT_0_port, A => 
                           n10898, ZN => n10936);
   U12617 : NOR2_X1 port map( A1 => n10902, A2 => n10899, ZN => n10934);
   U12618 : AOI22_X1 port map( A1 => n10919, A2 => n10934, B1 => n10929, B2 => 
                           n10935, ZN => n10900);
   U12619 : NAND3_X1 port map( A1 => n10936, A2 => n10900, A3 => n10920, ZN => 
                           DRAM_DATA_OUT_24_port);
   U12620 : NOR2_X1 port map( A1 => n10902, A2 => n10901, ZN => n10938);
   U12621 : INV_X1 port map( A => n10938, ZN => n10904);
   U12622 : AOI22_X1 port map( A1 => n10941, A2 => DRAM_DATA_OUT_1_port, B1 => 
                           n10929, B2 => n10939, ZN => n10903);
   U12623 : OAI211_X1 port map( C1 => n10904, C2 => n10927, A => n10926, B => 
                           n10903, ZN => DRAM_DATA_OUT_25_port);
   U12624 : AOI22_X1 port map( A1 => n10919, A2 => n10906, B1 => n10929, B2 => 
                           n10905, ZN => n10907);
   U12625 : NAND3_X1 port map( A1 => n10908, A2 => n10907, A3 => n10920, ZN => 
                           DRAM_DATA_OUT_26_port);
   U12626 : INV_X1 port map( A => n10909, ZN => n10912);
   U12627 : AOI22_X1 port map( A1 => n10941, A2 => DRAM_DATA_OUT_3_port, B1 => 
                           n10929, B2 => n10910, ZN => n10911);
   U12628 : OAI211_X1 port map( C1 => n10912, C2 => n10927, A => n10926, B => 
                           n10911, ZN => DRAM_DATA_OUT_27_port);
   U12629 : AOI22_X1 port map( A1 => n10919, A2 => n10914, B1 => n10929, B2 => 
                           n10913, ZN => n10915);
   U12630 : NAND3_X1 port map( A1 => n10916, A2 => n10915, A3 => n10920, ZN => 
                           DRAM_DATA_OUT_28_port);
   U12631 : AOI22_X1 port map( A1 => n10919, A2 => n10918, B1 => n10929, B2 => 
                           n10917, ZN => n10921);
   U12632 : NAND3_X1 port map( A1 => n10922, A2 => n10921, A3 => n10920, ZN => 
                           DRAM_DATA_OUT_29_port);
   U12633 : INV_X1 port map( A => n10923, ZN => n10928);
   U12634 : AOI22_X1 port map( A1 => n10941, A2 => DRAM_DATA_OUT_6_port, B1 => 
                           n10929, B2 => n10924, ZN => n10925);
   U12635 : OAI211_X1 port map( C1 => n10928, C2 => n10927, A => n10926, B => 
                           n10925, ZN => DRAM_DATA_OUT_30_port);
   U12636 : INV_X1 port map( A => n10929, ZN => n10932);
   U12637 : OAI211_X1 port map( C1 => n10933, C2 => n10932, A => n10931, B => 
                           n10930, ZN => DRAM_DATA_OUT_31_port);
   U12638 : AOI21_X1 port map( B1 => n10940, B2 => n10935, A => n10934, ZN => 
                           n10937);
   U12639 : OAI21_X1 port map( B1 => n10945, B2 => n10937, A => n10936, ZN => 
                           DRAM_DATA_OUT_8_port);
   U12640 : AOI21_X1 port map( B1 => n10940, B2 => n10939, A => n10938, ZN => 
                           n10944);
   U12641 : NAND2_X1 port map( A1 => n10941, A2 => DRAM_DATA_OUT_1_port, ZN => 
                           n10943);
   U12642 : OAI211_X1 port map( C1 => n10945, C2 => n10944, A => n10943, B => 
                           n10942, ZN => DRAM_DATA_OUT_9_port);
   U12643 : OAI211_X1 port map( C1 => n11831, C2 => n8327, A => n8577, B => 
                           n11051, ZN => DataPath_RF_POP_ADDRGEN_N46);
   U12644 : AOI22_X1 port map( A1 => n11831, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_0_port, B1 => 
                           n10947, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_1_port, ZN => 
                           n11056);
   U12645 : NOR2_X1 port map( A1 => RST, A2 => n11056, ZN => 
                           DataPath_RF_POP_ADDRGEN_N47);
   U12646 : AOI22_X1 port map( A1 => n11831, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_1_port, B1 => 
                           n10947, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_2_port, ZN => 
                           n11060);
   U12647 : NOR2_X1 port map( A1 => RST, A2 => n11060, ZN => 
                           DataPath_RF_POP_ADDRGEN_N48);
   U12648 : AOI22_X1 port map( A1 => n11831, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_2_port, B1 => 
                           n10947, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_3_port, ZN => 
                           n11075);
   U12649 : NOR2_X1 port map( A1 => RST, A2 => n11075, ZN => 
                           DataPath_RF_POP_ADDRGEN_N49);
   U12650 : AOI22_X1 port map( A1 => n11831, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_3_port, B1 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_4_port, B2 => 
                           n10947, ZN => n11083);
   U12651 : NOR2_X1 port map( A1 => RST, A2 => n11083, ZN => 
                           DataPath_RF_POP_ADDRGEN_N50);
   U12652 : AOI22_X1 port map( A1 => n11831, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_4_port, B1 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_5_port, B2 => 
                           n10947, ZN => n10968);
   U12653 : NOR2_X1 port map( A1 => RST, A2 => n10968, ZN => 
                           DataPath_RF_POP_ADDRGEN_N51);
   U12654 : INV_X1 port map( A => n11831, ZN => n11052);
   U12655 : OAI221_X1 port map( B1 => n11052, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_5_port, C1 => 
                           n11831, C2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_6_port, A => 
                           n11051, ZN => n10976);
   U12656 : NOR2_X1 port map( A1 => n10976, A2 => RST, ZN => 
                           DataPath_RF_POP_ADDRGEN_N52);
   U12657 : AOI22_X1 port map( A1 => n11831, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_6_port, B1 => 
                           n10947, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_7_port, ZN => 
                           n11004);
   U12658 : NOR2_X1 port map( A1 => RST, A2 => n11004, ZN => 
                           DataPath_RF_POP_ADDRGEN_N53);
   U12659 : AOI22_X1 port map( A1 => n11831, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_7_port, B1 => 
                           n10947, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_8_port, ZN => 
                           n11009);
   U12660 : NOR2_X1 port map( A1 => RST, A2 => n11009, ZN => 
                           DataPath_RF_POP_ADDRGEN_N54);
   U12661 : AOI22_X1 port map( A1 => n11831, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_8_port, B1 => 
                           n10947, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_9_port, ZN => 
                           n11017);
   U12662 : NOR2_X1 port map( A1 => RST, A2 => n11017, ZN => 
                           DataPath_RF_POP_ADDRGEN_N55);
   U12663 : AOI22_X1 port map( A1 => n11831, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_9_port, B1 => 
                           n10947, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_10_port, ZN => 
                           n11021);
   U12664 : NOR2_X1 port map( A1 => RST, A2 => n11021, ZN => 
                           DataPath_RF_POP_ADDRGEN_N56);
   U12665 : AOI22_X1 port map( A1 => n11831, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_10_port, B1 => 
                           n10947, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_11_port, ZN => 
                           n11026);
   U12666 : NOR2_X1 port map( A1 => RST, A2 => n11026, ZN => 
                           DataPath_RF_POP_ADDRGEN_N57);
   U12667 : AOI22_X1 port map( A1 => n11831, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_11_port, B1 => 
                           n10947, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_12_port, ZN => 
                           n11030);
   U12668 : NOR2_X1 port map( A1 => RST, A2 => n11030, ZN => 
                           DataPath_RF_POP_ADDRGEN_N58);
   U12669 : AOI22_X1 port map( A1 => n11831, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_12_port, B1 => 
                           n10947, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_13_port, ZN => 
                           n11034);
   U12670 : NOR2_X1 port map( A1 => RST, A2 => n11034, ZN => 
                           DataPath_RF_POP_ADDRGEN_N59);
   U12671 : AOI22_X1 port map( A1 => n11831, A2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_13_port, B1 => 
                           n10947, B2 => 
                           DataPath_RF_POP_ADDRGEN_curr_addr_14_port, ZN => 
                           n11039);
   U12672 : NOR2_X1 port map( A1 => RST, A2 => n11039, ZN => 
                           DataPath_RF_POP_ADDRGEN_N60);
   U12673 : OAI22_X1 port map( A1 => n11830, A2 => n8291, B1 => n11052, B2 => 
                           n8211, ZN => n11047);
   U12674 : AND2_X1 port map( A1 => n8580, A2 => n11047, ZN => 
                           DataPath_RF_POP_ADDRGEN_N61);
   U12675 : NOR2_X1 port map( A1 => RST, A2 => n11816, ZN => n10964);
   U12676 : OAI21_X1 port map( B1 => n11817, B2 => n8325, A => n10964, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N46);
   U12677 : AOI22_X1 port map( A1 => n11817, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_0_port, B1 => 
                           n10961, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, ZN => 
                           n10948);
   U12678 : NOR2_X1 port map( A1 => RST, A2 => n10948, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N47);
   U12679 : AOI22_X1 port map( A1 => n11817, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_1_port, B1 => 
                           n10961, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, ZN => 
                           n10949);
   U12680 : NOR2_X1 port map( A1 => RST, A2 => n10949, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N48);
   U12681 : AOI22_X1 port map( A1 => n11817, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_2_port, B1 => 
                           n10961, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, ZN => 
                           n10950);
   U12682 : NOR2_X1 port map( A1 => RST, A2 => n10950, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N49);
   U12683 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_3_port, B1 => 
                           n10961, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, ZN => 
                           n10951);
   U12684 : NOR2_X1 port map( A1 => RST, A2 => n10951, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N50);
   U12685 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_4_port, B1 => 
                           n10961, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, ZN => 
                           n10952);
   U12686 : NOR2_X1 port map( A1 => RST, A2 => n10952, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N51);
   U12687 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_5_port, B1 => 
                           n10961, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, ZN => 
                           n10953);
   U12688 : NOR2_X1 port map( A1 => RST, A2 => n10953, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N52);
   U12689 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_6_port, B1 => 
                           n10961, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, ZN => 
                           n10954);
   U12690 : NOR2_X1 port map( A1 => RST, A2 => n10954, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N53);
   U12691 : AOI22_X1 port map( A1 => n11817, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_7_port, B1 => 
                           n10961, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, ZN => 
                           n10955);
   U12692 : NOR2_X1 port map( A1 => RST, A2 => n10955, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N54);
   U12693 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_8_port, B1 => 
                           n10961, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, ZN => 
                           n10956);
   U12694 : NOR2_X1 port map( A1 => RST, A2 => n10956, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N55);
   U12695 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_9_port, B1 => 
                           n10961, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, ZN => 
                           n10957);
   U12696 : NOR2_X1 port map( A1 => RST, A2 => n10957, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N56);
   U12697 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_10_port, B1 => 
                           n10961, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, ZN => 
                           n10958);
   U12698 : NOR2_X1 port map( A1 => RST, A2 => n10958, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N57);
   U12699 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_11_port, B1 => 
                           n10961, B2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, ZN => 
                           n10959);
   U12700 : NOR2_X1 port map( A1 => RST, A2 => n10959, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N58);
   U12701 : AOI22_X1 port map( A1 => n8541, A2 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_12_port, B1 => 
                           DataPath_RF_PUSH_ADDRGEN_curr_addr_13_port, B2 => 
                           n10961, ZN => n10960);
   U12702 : NOR2_X1 port map( A1 => RST, A2 => n10960, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N59);
   U12703 : INV_X1 port map( A => n10961, ZN => n10962);
   U12704 : AOI221_X1 port map( B1 => n8310, B2 => n10963, C1 => n10962, C2 => 
                           n10963, A => RST, ZN => DataPath_RF_PUSH_ADDRGEN_N60
                           );
   U12705 : INV_X1 port map( A => n10964, ZN => n11997);
   U12706 : NOR2_X1 port map( A1 => n10965, A2 => n11997, ZN => 
                           DataPath_RF_PUSH_ADDRGEN_N61);
   U12707 : NOR2_X1 port map( A1 => n10437, A2 => n465, ZN => n11990);
   U12708 : AOI22_X1 port map( A1 => DRAMRF_READY, A2 => n11990, B1 => 
                           DP_OP_1091J1_126_6973_n72, B2 => n11820, ZN => 
                           n10967);
   U12709 : NOR2_X1 port map( A1 => n11996, A2 => n7438, ZN => n11991);
   U12710 : OAI22_X1 port map( A1 => n10436, A2 => n10435, B1 => n11991, B2 => 
                           n11449, ZN => n10966);
   U12711 : AOI21_X1 port map( B1 => n10967, B2 => n10966, A => RST, ZN => 
                           DataPath_WRF_CUhw_N145);
   U12712 : INV_X1 port map( A => n10968, ZN => n10969);
   U12713 : NAND2_X1 port map( A1 => n11082, A2 => n11638, ZN => n11512);
   U12714 : MUX2_X1 port map( A => DRAMRF_DATA_IN(16), B => 
                           DataPath_WRF_CUhw_curr_data_16_port, S => n11993, Z 
                           => n11470);
   U12715 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_16_port, B => 
                           DataPath_i_REG_LDSTR_OUT_16_port, S => n8565, Z => 
                           n11469);
   U12716 : OAI22_X1 port map( A1 => n11923, A2 => n11470, B1 => n11469, B2 => 
                           n7782, ZN => n10992);
   U12717 : OAI22_X1 port map( A1 => n11975, A2 => n11910, B1 => 
                           DataPath_RF_bus_reg_dataout_2384_port, B2 => n8550, 
                           ZN => n6134);
   U12718 : MUX2_X1 port map( A => DRAMRF_DATA_IN(17), B => 
                           DataPath_WRF_CUhw_curr_data_17_port, S => n11993, Z 
                           => n11472);
   U12719 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_17_port, B => 
                           DataPath_i_REG_LDSTR_OUT_17_port, S => n8565, Z => 
                           n11471);
   U12720 : OAI22_X1 port map( A1 => n11923, A2 => n11472, B1 => n11471, B2 => 
                           n7782, ZN => n10993);
   U12721 : OAI22_X1 port map( A1 => n8551, A2 => n11940, B1 => 
                           DataPath_RF_bus_reg_dataout_2385_port, B2 => n8550, 
                           ZN => n6133);
   U12722 : MUX2_X1 port map( A => DRAMRF_DATA_IN(18), B => 
                           DataPath_WRF_CUhw_curr_data_18_port, S => n11993, Z 
                           => n11701);
   U12723 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_18_port, B => 
                           DataPath_i_REG_LDSTR_OUT_18_port, S => n8565, Z => 
                           n10970);
   U12724 : AOI22_X1 port map( A1 => n7782, A2 => n11473, B1 => n11663, B2 => 
                           n11923, ZN => n11941);
   U12725 : OAI22_X1 port map( A1 => n8551, A2 => n11911, B1 => 
                           DataPath_RF_bus_reg_dataout_2386_port, B2 => n8550, 
                           ZN => n6132);
   U12726 : MUX2_X1 port map( A => DRAMRF_DATA_IN(19), B => 
                           DataPath_WRF_CUhw_curr_data_19_port, S => n11993, Z 
                           => n11475);
   U12727 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_19_port, B => 
                           DataPath_i_REG_LDSTR_OUT_19_port, S => n8565, Z => 
                           n11474);
   U12728 : OAI22_X1 port map( A1 => n11923, A2 => n11475, B1 => n11474, B2 => 
                           n7782, ZN => n10994);
   U12729 : OAI22_X1 port map( A1 => n8551, A2 => n11942, B1 => 
                           DataPath_RF_bus_reg_dataout_2387_port, B2 => n8550, 
                           ZN => n6131);
   U12730 : MUX2_X1 port map( A => DRAMRF_DATA_IN(20), B => 
                           DataPath_WRF_CUhw_curr_data_20_port, S => n11993, Z 
                           => n11476);
   U12731 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_20_port, B => 
                           DataPath_i_REG_LDSTR_OUT_20_port, S => n8565, Z => 
                           n10971);
   U12732 : AOI22_X1 port map( A1 => n7782, A2 => n11319, B1 => n11665, B2 => 
                           n11923, ZN => n11902);
   U12733 : OAI22_X1 port map( A1 => n8551, A2 => n11943, B1 => 
                           DataPath_RF_bus_reg_dataout_2388_port, B2 => n8550, 
                           ZN => n6130);
   U12734 : MUX2_X1 port map( A => DRAMRF_DATA_IN(21), B => 
                           DataPath_WRF_CUhw_curr_data_21_port, S => n11993, Z 
                           => n11702);
   U12735 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_21_port, B => 
                           DataPath_i_REG_LDSTR_OUT_21_port, S => n8565, Z => 
                           n10972);
   U12736 : AOI22_X1 port map( A1 => n7782, A2 => n11477, B1 => n11666, B2 => 
                           n11923, ZN => n11903);
   U12737 : OAI22_X1 port map( A1 => n8551, A2 => n11945, B1 => 
                           DataPath_RF_bus_reg_dataout_2389_port, B2 => n8550, 
                           ZN => n6129);
   U12738 : MUX2_X1 port map( A => DRAMRF_DATA_IN(22), B => 
                           DataPath_WRF_CUhw_curr_data_22_port, S => n11993, Z 
                           => n11703);
   U12739 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_22_port, B => 
                           DataPath_i_REG_LDSTR_OUT_22_port, S => n8565, Z => 
                           n10973);
   U12740 : AOI22_X1 port map( A1 => n7782, A2 => n11478, B1 => n11667, B2 => 
                           n11923, ZN => n11946);
   U12741 : OAI22_X1 port map( A1 => n8551, A2 => n11912, B1 => 
                           DataPath_RF_bus_reg_dataout_2390_port, B2 => n8550, 
                           ZN => n6128);
   U12742 : MUX2_X1 port map( A => DRAMRF_DATA_IN(23), B => 
                           DataPath_WRF_CUhw_curr_data_23_port, S => n11993, Z 
                           => n11480);
   U12743 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_23_port, B => 
                           DataPath_i_REG_LDSTR_OUT_23_port, S => n8565, Z => 
                           n11479);
   U12744 : OAI22_X1 port map( A1 => n11923, A2 => n11480, B1 => n11479, B2 => 
                           n7782, ZN => n10995);
   U12745 : OAI22_X1 port map( A1 => n11975, A2 => n11913, B1 => 
                           DataPath_RF_bus_reg_dataout_2391_port, B2 => n8550, 
                           ZN => n6127);
   U12746 : MUX2_X1 port map( A => DRAMRF_DATA_IN(24), B => 
                           DataPath_WRF_CUhw_curr_data_24_port, S => n11993, Z 
                           => n11482);
   U12747 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_24_port, B => 
                           DataPath_i_REG_LDSTR_OUT_24_port, S => n8565, Z => 
                           n11481);
   U12748 : OAI22_X1 port map( A1 => n11923, A2 => n11482, B1 => n11481, B2 => 
                           n7782, ZN => n10996);
   U12749 : OAI22_X1 port map( A1 => n8551, A2 => n11914, B1 => 
                           DataPath_RF_bus_reg_dataout_2392_port, B2 => n8550, 
                           ZN => n6126);
   U12750 : MUX2_X1 port map( A => DRAMRF_DATA_IN(25), B => 
                           DataPath_WRF_CUhw_curr_data_25_port, S => n11993, Z 
                           => n11484);
   U12751 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_25_port, B => 
                           DataPath_i_REG_LDSTR_OUT_25_port, S => n8565, Z => 
                           n11483);
   U12752 : OAI22_X1 port map( A1 => n11923, A2 => n11484, B1 => n11483, B2 => 
                           n7782, ZN => n10997);
   U12753 : OAI22_X1 port map( A1 => n8551, A2 => n11915, B1 => 
                           DataPath_RF_bus_reg_dataout_2393_port, B2 => n8550, 
                           ZN => n6125);
   U12754 : MUX2_X1 port map( A => DRAMRF_DATA_IN(26), B => 
                           DataPath_WRF_CUhw_curr_data_26_port, S => n11993, Z 
                           => n11704);
   U12755 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_26_port, B => 
                           DataPath_i_REG_LDSTR_OUT_26_port, S => n8565, Z => 
                           n10974);
   U12756 : OAI22_X1 port map( A1 => n11923, A2 => n11485, B1 => n11671, B2 => 
                           n7782, ZN => n11950);
   U12757 : OAI22_X1 port map( A1 => n11916, A2 => n8551, B1 => 
                           DataPath_RF_bus_reg_dataout_2394_port, B2 => n8550, 
                           ZN => n6124);
   U12758 : MUX2_X1 port map( A => DRAMRF_DATA_IN(27), B => 
                           DataPath_WRF_CUhw_curr_data_27_port, S => n11993, Z 
                           => n11487);
   U12759 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_27_port, B => 
                           DataPath_i_REG_LDSTR_OUT_27_port, S => i_S3, Z => 
                           n11486);
   U12760 : OAI22_X1 port map( A1 => n11923, A2 => n11487, B1 => n11486, B2 => 
                           n7782, ZN => n10998);
   U12761 : OAI22_X1 port map( A1 => n11975, A2 => n11917, B1 => 
                           DataPath_RF_bus_reg_dataout_2395_port, B2 => n8550, 
                           ZN => n6123);
   U12762 : MUX2_X1 port map( A => DRAMRF_DATA_IN(28), B => 
                           DataPath_WRF_CUhw_curr_data_28_port, S => n11993, Z 
                           => n11489);
   U12763 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_28_port, B => 
                           DataPath_i_REG_LDSTR_OUT_28_port, S => i_S3, Z => 
                           n11488);
   U12764 : OAI22_X1 port map( A1 => n11923, A2 => n11489, B1 => n11488, B2 => 
                           n7782, ZN => n10999);
   U12765 : OAI22_X1 port map( A1 => n8551, A2 => n11918, B1 => 
                           DataPath_RF_bus_reg_dataout_2396_port, B2 => n8550, 
                           ZN => n6122);
   U12766 : MUX2_X1 port map( A => DRAMRF_DATA_IN(29), B => 
                           DataPath_WRF_CUhw_curr_data_29_port, S => n11993, Z 
                           => n11490);
   U12767 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_29_port, B => 
                           DataPath_i_REG_LDSTR_OUT_29_port, S => i_S3, Z => 
                           n10975);
   U12768 : OAI22_X1 port map( A1 => n11923, A2 => n11320, B1 => n11674, B2 => 
                           n7782, ZN => n11953);
   U12769 : OAI22_X1 port map( A1 => n11919, A2 => n8551, B1 => 
                           DataPath_RF_bus_reg_dataout_2397_port, B2 => n8550, 
                           ZN => n6121);
   U12770 : MUX2_X1 port map( A => DRAMRF_DATA_IN(30), B => 
                           DataPath_WRF_CUhw_curr_data_30_port, S => n11993, Z 
                           => n11493);
   U12771 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_30_port, B => 
                           DataPath_i_REG_LDSTR_OUT_30_port, S => i_S3, Z => 
                           n11492);
   U12772 : OAI22_X1 port map( A1 => n11923, A2 => n11493, B1 => n11492, B2 => 
                           n7782, ZN => n11000);
   U12773 : OAI22_X1 port map( A1 => n8551, A2 => n11920, B1 => 
                           DataPath_RF_bus_reg_dataout_2398_port, B2 => n8550, 
                           ZN => n6120);
   U12774 : MUX2_X1 port map( A => DRAMRF_DATA_IN(31), B => 
                           DataPath_WRF_CUhw_curr_data_31_port, S => n11993, Z 
                           => n11495);
   U12775 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_31_port, B => 
                           DataPath_i_REG_LDSTR_OUT_31_port, S => i_S3, Z => 
                           n11494);
   U12776 : OAI22_X1 port map( A1 => n11923, A2 => n11495, B1 => n11494, B2 => 
                           n7782, ZN => n11001);
   U12777 : OAI22_X1 port map( A1 => n11975, A2 => n11921, B1 => 
                           DataPath_RF_bus_reg_dataout_2399_port, B2 => n8550, 
                           ZN => n6119);
   U12778 : INV_X1 port map( A => n10976, ZN => n10977);
   U12779 : NAND2_X1 port map( A1 => n11082, A2 => n11643, ZN => n11517);
   U12780 : OAI22_X1 port map( A1 => n11518, A2 => n11923, B1 => n8219, B2 => 
                           n11517, ZN => n10987);
   U12781 : MUX2_X1 port map( A => DRAMRF_DATA_IN(0), B => 
                           DataPath_WRF_CUhw_curr_data_0_port, S => n11993, Z 
                           => n11688);
   U12782 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_0_port, B => 
                           DataPath_i_REG_LDSTR_OUT_0_port, S => i_S3, Z => 
                           n10978);
   U12783 : AOI22_X1 port map( A1 => n7782, A2 => n11450, B1 => n11645, B2 => 
                           n11923, ZN => n11925);
   U12784 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2336_port, A2 
                           => n11003, B1 => n11002, B2 => n11925, ZN => n6116);
   U12785 : MUX2_X1 port map( A => DRAMRF_DATA_IN(1), B => 
                           DataPath_WRF_CUhw_curr_data_1_port, S => n11993, Z 
                           => n11689);
   U12786 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_1_port, B => 
                           DataPath_i_REG_LDSTR_OUT_1_port, S => i_S3, Z => 
                           n10979);
   U12787 : AOI22_X1 port map( A1 => n7782, A2 => n11451, B1 => n11646, B2 => 
                           n11923, ZN => n11926);
   U12788 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2337_port, A2 
                           => n8479, B1 => n11002, B2 => n11926, ZN => n6115);
   U12789 : MUX2_X1 port map( A => DRAMRF_DATA_IN(2), B => 
                           DataPath_WRF_CUhw_curr_data_2_port, S => n11993, Z 
                           => n11690);
   U12790 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_2_port, B => 
                           DataPath_i_REG_LDSTR_OUT_2_port, S => i_S3, Z => 
                           n10980);
   U12791 : AOI22_X1 port map( A1 => n7782, A2 => n11452, B1 => n11647, B2 => 
                           n11923, ZN => n11927);
   U12792 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2338_port, A2 
                           => n8479, B1 => n11002, B2 => n11927, ZN => n6114);
   U12793 : MUX2_X1 port map( A => DRAMRF_DATA_IN(3), B => 
                           DataPath_WRF_CUhw_curr_data_3_port, S => n11993, Z 
                           => n11691);
   U12794 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_3_port, B => 
                           DataPath_i_REG_LDSTR_OUT_3_port, S => i_S3, Z => 
                           n10981);
   U12795 : AOI22_X1 port map( A1 => n7782, A2 => n11453, B1 => n11648, B2 => 
                           n11923, ZN => n11928);
   U12796 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2339_port, A2 
                           => n8479, B1 => n11002, B2 => n11928, ZN => n6113);
   U12797 : MUX2_X1 port map( A => DRAMRF_DATA_IN(4), B => 
                           DataPath_WRF_CUhw_curr_data_4_port, S => n11993, Z 
                           => n11692);
   U12798 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_4_port, B => 
                           DataPath_i_REG_LDSTR_OUT_4_port, S => i_S3, Z => 
                           n10982);
   U12799 : AOI22_X1 port map( A1 => n7782, A2 => n11454, B1 => n11649, B2 => 
                           n11923, ZN => n11929);
   U12800 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2340_port, A2 
                           => n11003, B1 => n11002, B2 => n11929, ZN => n6112);
   U12801 : MUX2_X1 port map( A => DRAMRF_DATA_IN(5), B => 
                           DataPath_WRF_CUhw_curr_data_5_port, S => n11993, Z 
                           => n11456);
   U12802 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_5_port, B => 
                           DataPath_i_REG_LDSTR_OUT_5_port, S => i_S3, Z => 
                           n11455);
   U12803 : OAI22_X1 port map( A1 => n11923, A2 => n11456, B1 => n11455, B2 => 
                           n7782, ZN => n11012);
   U12804 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2341_port, A2 
                           => n11003, B1 => n11002, B2 => n11930, ZN => n6111);
   U12805 : MUX2_X1 port map( A => DRAMRF_DATA_IN(6), B => 
                           DataPath_WRF_CUhw_curr_data_6_port, S => n11993, Z 
                           => n11693);
   U12806 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_6_port, B => 
                           DataPath_i_REG_LDSTR_OUT_6_port, S => i_S3, Z => 
                           n10983);
   U12807 : AOI22_X1 port map( A1 => n7782, A2 => n11457, B1 => n11651, B2 => 
                           n11923, ZN => n11931);
   U12808 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2342_port, A2 
                           => n8479, B1 => n11002, B2 => n11931, ZN => n6110);
   U12809 : MUX2_X1 port map( A => DRAMRF_DATA_IN(7), B => 
                           DataPath_WRF_CUhw_curr_data_7_port, S => n11993, Z 
                           => n11694);
   U12810 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_7_port, B => 
                           DataPath_i_REG_LDSTR_OUT_7_port, S => i_S3, Z => 
                           n10984);
   U12811 : AOI22_X1 port map( A1 => n7782, A2 => n11458, B1 => n11652, B2 => 
                           n11923, ZN => n11932);
   U12812 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2343_port, A2 
                           => n11003, B1 => n11002, B2 => n11932, ZN => n6109);
   U12813 : MUX2_X1 port map( A => DRAMRF_DATA_IN(8), B => 
                           DataPath_WRF_CUhw_curr_data_8_port, S => n11993, Z 
                           => n11695);
   U12814 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_8_port, B => 
                           DataPath_i_REG_LDSTR_OUT_8_port, S => i_S3, Z => 
                           n10985);
   U12815 : AOI22_X1 port map( A1 => n7782, A2 => n11459, B1 => n11653, B2 => 
                           n11923, ZN => n11898);
   U12816 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2344_port, A2 
                           => n11003, B1 => n11002, B2 => n11898, ZN => n6108);
   U12817 : MUX2_X1 port map( A => DRAMRF_DATA_IN(9), B => 
                           DataPath_WRF_CUhw_curr_data_9_port, S => n11993, Z 
                           => n11461);
   U12818 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_9_port, B => 
                           DataPath_i_REG_LDSTR_OUT_9_port, S => n8565, Z => 
                           n11460);
   U12819 : OAI22_X1 port map( A1 => n11923, A2 => n11461, B1 => n11460, B2 => 
                           n7782, ZN => n11013);
   U12820 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2345_port, A2 
                           => n8479, B1 => n11002, B2 => n11933, ZN => n6107);
   U12821 : MUX2_X1 port map( A => DRAMRF_DATA_IN(10), B => 
                           DataPath_WRF_CUhw_curr_data_10_port, S => n11993, Z 
                           => n11696);
   U12822 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_10_port, B => 
                           DataPath_i_REG_LDSTR_OUT_10_port, S => i_S3, Z => 
                           n10986);
   U12823 : AOI22_X1 port map( A1 => n7782, A2 => n11462, B1 => n11655, B2 => 
                           n11923, ZN => n11934);
   U12824 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2346_port, A2 
                           => n8479, B1 => n11968, B2 => n10987, ZN => n6106);
   U12825 : MUX2_X1 port map( A => DRAMRF_DATA_IN(11), B => 
                           DataPath_WRF_CUhw_curr_data_11_port, S => n11993, Z 
                           => n11697);
   U12826 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_11_port, B => 
                           DataPath_i_REG_LDSTR_OUT_11_port, S => i_S3, Z => 
                           n10988);
   U12827 : AOI22_X1 port map( A1 => n7782, A2 => n11463, B1 => n11656, B2 => 
                           n11923, ZN => n11935);
   U12828 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2347_port, A2 
                           => n8479, B1 => n11002, B2 => n11935, ZN => n6105);
   U12829 : MUX2_X1 port map( A => DRAMRF_DATA_IN(12), B => 
                           DataPath_WRF_CUhw_curr_data_12_port, S => n11993, Z 
                           => n11698);
   U12830 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_12_port, B => 
                           DataPath_i_REG_LDSTR_OUT_12_port, S => i_S3, Z => 
                           n10989);
   U12831 : AOI22_X1 port map( A1 => n7782, A2 => n11464, B1 => n11657, B2 => 
                           n11923, ZN => n11936);
   U12832 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2348_port, A2 
                           => n8479, B1 => n11002, B2 => n11936, ZN => n6104);
   U12833 : MUX2_X1 port map( A => DRAMRF_DATA_IN(13), B => 
                           DataPath_WRF_CUhw_curr_data_13_port, S => n11993, Z 
                           => n11699);
   U12834 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_13_port, B => 
                           DataPath_i_REG_LDSTR_OUT_13_port, S => i_S3, Z => 
                           n10990);
   U12835 : AOI22_X1 port map( A1 => n7782, A2 => n11465, B1 => n11658, B2 => 
                           n11923, ZN => n11937);
   U12836 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2349_port, A2 
                           => n11003, B1 => n11002, B2 => n11937, ZN => n6103);
   U12837 : MUX2_X1 port map( A => DRAMRF_DATA_IN(14), B => 
                           DataPath_WRF_CUhw_curr_data_14_port, S => n11993, Z 
                           => n11700);
   U12838 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_14_port, B => 
                           DataPath_i_REG_LDSTR_OUT_14_port, S => i_S3, Z => 
                           n10991);
   U12839 : AOI22_X1 port map( A1 => n7782, A2 => n11466, B1 => n11659, B2 => 
                           n11923, ZN => n11899);
   U12840 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2350_port, A2 
                           => n11003, B1 => n11002, B2 => n11899, ZN => n6102);
   U12841 : MUX2_X1 port map( A => DRAMRF_DATA_IN(15), B => 
                           DataPath_WRF_CUhw_curr_data_15_port, S => n11993, Z 
                           => n11468);
   U12842 : MUX2_X1 port map( A => DataPath_i_REG_MEM_ALUOUT_15_port, B => 
                           DataPath_i_REG_LDSTR_OUT_15_port, S => i_S3, Z => 
                           n11467);
   U12843 : OAI22_X1 port map( A1 => n11923, A2 => n11468, B1 => n11467, B2 => 
                           n7782, ZN => n11014);
   U12844 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2351_port, A2 
                           => n8479, B1 => n11002, B2 => n11938, ZN => n6101);
   U12845 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2352_port, A2 
                           => n11003, B1 => n11002, B2 => n11939, ZN => n6100);
   U12846 : INV_X1 port map( A => n10993, ZN => n11900);
   U12847 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2353_port, A2 
                           => n8479, B1 => n11002, B2 => n11900, ZN => n6099);
   U12848 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2354_port, A2 
                           => n8479, B1 => n11002, B2 => n11941, ZN => n6098);
   U12849 : INV_X1 port map( A => n10994, ZN => n11901);
   U12850 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2355_port, A2 
                           => n8479, B1 => n11002, B2 => n11901, ZN => n6097);
   U12851 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2356_port, A2 
                           => n8479, B1 => n11002, B2 => n11902, ZN => n6096);
   U12852 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2357_port, A2 
                           => n8479, B1 => n11002, B2 => n11903, ZN => n6095);
   U12853 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2358_port, A2 
                           => n11003, B1 => n11002, B2 => n11946, ZN => n6094);
   U12854 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2359_port, A2 
                           => n11003, B1 => n11002, B2 => n11947, ZN => n6093);
   U12855 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2360_port, A2 
                           => n8479, B1 => n11002, B2 => n11948, ZN => n6092);
   U12856 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2361_port, A2 
                           => n8479, B1 => n11002, B2 => n11949, ZN => n6091);
   U12857 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2362_port, A2 
                           => n8479, B1 => n11002, B2 => n11950, ZN => n6090);
   U12858 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2363_port, A2 
                           => n8479, B1 => n11002, B2 => n11951, ZN => n6089);
   U12859 : INV_X1 port map( A => n10999, ZN => n11952);
   U12860 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2364_port, A2 
                           => n8479, B1 => n11002, B2 => n11952, ZN => n6088);
   U12861 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2365_port, A2 
                           => n8479, B1 => n11002, B2 => n11953, ZN => n6087);
   U12862 : INV_X1 port map( A => n11000, ZN => n11954);
   U12863 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2366_port, A2 
                           => n8479, B1 => n11002, B2 => n11954, ZN => n6086);
   U12864 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2367_port, A2 
                           => n8479, B1 => n11002, B2 => n11955, ZN => n6083);
   U12865 : NAND2_X1 port map( A1 => n11082, A2 => n11046, ZN => n11524);
   U12866 : INV_X1 port map( A => n11004, ZN => n11005);
   U12867 : OAI22_X1 port map( A1 => n8219, A2 => n11524, B1 => n11923, B2 => 
                           n11523, ZN => n11006);
   U12868 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2304_port, A2 
                           => n8480, B1 => n11007, B2 => n11925, ZN => n6080);
   U12869 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2305_port, A2 
                           => n11008, B1 => n11007, B2 => n11926, ZN => n6079);
   U12870 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2306_port, A2 
                           => n8480, B1 => n11007, B2 => n11927, ZN => n6078);
   U12871 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2307_port, A2 
                           => n11008, B1 => n11007, B2 => n11928, ZN => n6077);
   U12872 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2308_port, A2 
                           => n11008, B1 => n11007, B2 => n11929, ZN => n6076);
   U12873 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2309_port, A2 
                           => n8480, B1 => n11007, B2 => n11930, ZN => n6075);
   U12874 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2310_port, A2 
                           => n8480, B1 => n11007, B2 => n11931, ZN => n6074);
   U12875 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2311_port, A2 
                           => n8480, B1 => n11007, B2 => n11932, ZN => n6073);
   U12876 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2312_port, A2 
                           => n11008, B1 => n11007, B2 => n11898, ZN => n6072);
   U12877 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2313_port, A2 
                           => n8480, B1 => n11007, B2 => n11933, ZN => n6071);
   U12878 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2314_port, A2 
                           => n8480, B1 => n11007, B2 => n11934, ZN => n6070);
   U12879 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2315_port, A2 
                           => n11008, B1 => n11007, B2 => n11935, ZN => n6069);
   U12880 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2316_port, A2 
                           => n11008, B1 => n11007, B2 => n11936, ZN => n6068);
   U12881 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2317_port, A2 
                           => n8480, B1 => n11007, B2 => n11937, ZN => n6067);
   U12882 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2318_port, A2 
                           => n8480, B1 => n11007, B2 => n11899, ZN => n6066);
   U12883 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2319_port, A2 
                           => n11008, B1 => n11007, B2 => n11938, ZN => n6065);
   U12884 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2320_port, A2 
                           => n8480, B1 => n11007, B2 => n11939, ZN => n6064);
   U12885 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2321_port, A2 
                           => n8480, B1 => n11007, B2 => n11900, ZN => n6063);
   U12886 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2322_port, A2 
                           => n8480, B1 => n11007, B2 => n11941, ZN => n6062);
   U12887 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2323_port, A2 
                           => n8480, B1 => n11007, B2 => n11901, ZN => n6061);
   U12888 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2324_port, A2 
                           => n11008, B1 => n11007, B2 => n11902, ZN => n6060);
   U12889 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2325_port, A2 
                           => n8480, B1 => n11007, B2 => n11903, ZN => n6059);
   U12890 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2326_port, A2 
                           => n11008, B1 => n11007, B2 => n11946, ZN => n6058);
   U12891 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2327_port, A2 
                           => n8480, B1 => n11007, B2 => n11947, ZN => n6057);
   U12892 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2328_port, A2 
                           => n8480, B1 => n11007, B2 => n11948, ZN => n6056);
   U12893 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2329_port, A2 
                           => n8480, B1 => n11007, B2 => n11949, ZN => n6055);
   U12894 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2330_port, A2 
                           => n11008, B1 => n11007, B2 => n11950, ZN => n6054);
   U12895 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2331_port, A2 
                           => n8480, B1 => n11007, B2 => n11951, ZN => n6053);
   U12896 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2332_port, A2 
                           => n8480, B1 => n11007, B2 => n11952, ZN => n6052);
   U12897 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2333_port, A2 
                           => n8480, B1 => n11007, B2 => n11953, ZN => n6051);
   U12898 : AOI22_X1 port map( A1 => n11920, A2 => n11006, B1 => n8480, B2 => 
                           DataPath_RF_bus_reg_dataout_2334_port, ZN => n6050);
   U12899 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2335_port, A2 
                           => n8480, B1 => n11007, B2 => n11955, ZN => n6047);
   U12900 : NAND2_X1 port map( A1 => n11617, A2 => n11045, ZN => n11543);
   U12901 : NAND2_X1 port map( A1 => n11617, A2 => n11044, ZN => n11544);
   U12902 : OAI22_X1 port map( A1 => n576, A2 => n11543, B1 => n11544, B2 => 
                           n8219, ZN => n11011);
   U12903 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2272_port, B1 => n11958,
                           B2 => n11015, ZN => n6043);
   U12904 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2273_port, B1 => n11959,
                           B2 => n11015, ZN => n6042);
   U12905 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2274_port, B1 => n11960,
                           B2 => n11015, ZN => n6041);
   U12906 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2275_port, B1 => n11961,
                           B2 => n11015, ZN => n6040);
   U12907 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2276_port, B1 => n11962,
                           B2 => n11015, ZN => n6039);
   U12908 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2277_port, B1 => n11963,
                           B2 => n11015, ZN => n6038);
   U12909 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2278_port, B1 => n11964,
                           B2 => n11015, ZN => n6037);
   U12910 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2279_port, B1 => n11965,
                           B2 => n11015, ZN => n6036);
   U12911 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2280_port, B1 => n11966,
                           B2 => n11015, ZN => n6035);
   U12912 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2281_port, B1 => n11967,
                           B2 => n11015, ZN => n6034);
   U12913 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2282_port, B1 => n11968,
                           B2 => n11015, ZN => n6033);
   U12914 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2283_port, B1 => n11969,
                           B2 => n11015, ZN => n6032);
   U12915 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2284_port, B1 => n11970,
                           B2 => n11015, ZN => n6031);
   U12916 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2285_port, B1 => n11971,
                           B2 => n11015, ZN => n6030);
   U12917 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2286_port, B1 => n11972,
                           B2 => n11015, ZN => n6029);
   U12918 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2287_port, B1 => n11974,
                           B2 => n11015, ZN => n6028);
   U12919 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2288_port, B1 => n11910,
                           B2 => n11015, ZN => n6027);
   U12920 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2289_port, B1 => n11940,
                           B2 => n11015, ZN => n6026);
   U12921 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2290_port, B1 => n11911,
                           B2 => n11015, ZN => n6025);
   U12922 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2291_port, B1 => n11942,
                           B2 => n11015, ZN => n6024);
   U12923 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2292_port, B1 => n11943,
                           B2 => n11015, ZN => n6023);
   U12924 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2293_port, B1 => n11945,
                           B2 => n11015, ZN => n6022);
   U12925 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2294_port, B1 => n11912,
                           B2 => n11015, ZN => n6021);
   U12926 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2295_port, B1 => n11913,
                           B2 => n11015, ZN => n6020);
   U12927 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2296_port, B1 => n11914,
                           B2 => n11015, ZN => n6019);
   U12928 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2297_port, B1 => n11915,
                           B2 => n11015, ZN => n6018);
   U12929 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2298_port, B1 => n11916,
                           B2 => n11015, ZN => n6017);
   U12930 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2299_port, B1 => n11917,
                           B2 => n11015, ZN => n6016);
   U12931 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2300_port, B1 => n11918,
                           B2 => n11015, ZN => n6015);
   U12932 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2301_port, B1 => n11919,
                           B2 => n11015, ZN => n6014);
   U12933 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2302_port, B1 => n11920,
                           B2 => n11015, ZN => n6013);
   U12934 : AOI22_X1 port map( A1 => n11016, A2 => 
                           DataPath_RF_bus_reg_dataout_2303_port, B1 => n11921,
                           B2 => n11015, ZN => n6010);
   U12935 : NAND2_X1 port map( A1 => n11045, A2 => n11621, ZN => n11102);
   U12936 : NAND2_X1 port map( A1 => n11044, A2 => n11621, ZN => n11550);
   U12937 : INV_X1 port map( A => n11017, ZN => n11018);
   U12938 : OAI22_X1 port map( A1 => n8219, A2 => n11550, B1 => n11923, B2 => 
                           n11549, ZN => n11019);
   U12939 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2240_port, B1 => n11958,
                           B2 => n8407, ZN => n6007);
   U12940 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2241_port, B1 => n11959,
                           B2 => n8407, ZN => n6006);
   U12941 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2242_port, B1 => n11960,
                           B2 => n8407, ZN => n6005);
   U12942 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2243_port, B1 => n11961,
                           B2 => n8407, ZN => n6004);
   U12943 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2244_port, B1 => n11962,
                           B2 => n8407, ZN => n6003);
   U12944 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2245_port, B1 => n11963,
                           B2 => n8407, ZN => n6002);
   U12945 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2246_port, B1 => n11964,
                           B2 => n8407, ZN => n6001);
   U12946 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2247_port, B1 => n11965,
                           B2 => n8407, ZN => n6000);
   U12947 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2248_port, B1 => n11966,
                           B2 => n8407, ZN => n5999);
   U12948 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2249_port, B1 => n11967,
                           B2 => n8407, ZN => n5998);
   U12949 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2250_port, B1 => n11968,
                           B2 => n8407, ZN => n5997);
   U12950 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2251_port, B1 => n11969,
                           B2 => n8407, ZN => n5996);
   U12951 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2252_port, B1 => n11970,
                           B2 => n8407, ZN => n5995);
   U12952 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2253_port, B1 => n11971,
                           B2 => n8407, ZN => n5994);
   U12953 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2254_port, B1 => n11972,
                           B2 => n8407, ZN => n5993);
   U12954 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2255_port, B1 => n11974,
                           B2 => n8407, ZN => n5992);
   U12955 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2256_port, B1 => n11910,
                           B2 => n8407, ZN => n5991);
   U12956 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2257_port, B1 => n11940,
                           B2 => n8407, ZN => n5990);
   U12957 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2258_port, B1 => n11911,
                           B2 => n8407, ZN => n5989);
   U12958 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2259_port, B1 => n11942,
                           B2 => n8407, ZN => n5988);
   U12959 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2260_port, B1 => n11943,
                           B2 => n8407, ZN => n5987);
   U12960 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2261_port, B1 => n11945,
                           B2 => n8407, ZN => n5986);
   U12961 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2262_port, B1 => n11912,
                           B2 => n8407, ZN => n5985);
   U12962 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2263_port, B1 => n11913,
                           B2 => n8407, ZN => n5984);
   U12963 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2264_port, B1 => n11914,
                           B2 => n8407, ZN => n5983);
   U12964 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2265_port, B1 => n11915,
                           B2 => n8407, ZN => n5982);
   U12965 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2266_port, B1 => n11916,
                           B2 => n8407, ZN => n5981);
   U12966 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2267_port, B1 => n11917,
                           B2 => n8407, ZN => n5980);
   U12967 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2268_port, B1 => n11918,
                           B2 => n8407, ZN => n5979);
   U12968 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2269_port, B1 => n11919,
                           B2 => n8407, ZN => n5978);
   U12969 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2270_port, B1 => n11920,
                           B2 => n8407, ZN => n5977);
   U12970 : AOI22_X1 port map( A1 => n7763, A2 => 
                           DataPath_RF_bus_reg_dataout_2271_port, B1 => n11921,
                           B2 => n8407, ZN => n5974);
   U12971 : NAND2_X1 port map( A1 => n11044, A2 => n11625, ZN => n11137);
   U12972 : NAND2_X1 port map( A1 => n11045, A2 => n11625, ZN => n11556);
   U12973 : INV_X1 port map( A => n11021, ZN => n11022);
   U12974 : AOI22_X1 port map( A1 => n11958, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2208_port, ZN => n5971);
   U12975 : AOI22_X1 port map( A1 => n11959, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2209_port, ZN => n5970);
   U12976 : AOI22_X1 port map( A1 => n11960, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2210_port, ZN => n5969);
   U12977 : AOI22_X1 port map( A1 => n11961, A2 => n11024, B1 => n11023, B2 => 
                           DataPath_RF_bus_reg_dataout_2211_port, ZN => n5968);
   U12978 : AOI22_X1 port map( A1 => n11962, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2212_port, ZN => n5967);
   U12979 : AOI22_X1 port map( A1 => n11963, A2 => n11024, B1 => n11023, B2 => 
                           DataPath_RF_bus_reg_dataout_2213_port, ZN => n5966);
   U12980 : AOI22_X1 port map( A1 => n11964, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2214_port, ZN => n5965);
   U12981 : OAI22_X1 port map( A1 => n11965, A2 => n8481, B1 => 
                           DataPath_RF_bus_reg_dataout_2215_port, B2 => n11024,
                           ZN => n5964);
   U12982 : AOI22_X1 port map( A1 => n11966, A2 => n11024, B1 => n11023, B2 => 
                           DataPath_RF_bus_reg_dataout_2216_port, ZN => n5963);
   U12983 : AOI22_X1 port map( A1 => n11967, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2217_port, ZN => n5962);
   U12984 : AOI22_X1 port map( A1 => n11968, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2218_port, ZN => n5961);
   U12985 : AOI22_X1 port map( A1 => n11969, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2219_port, ZN => n5960);
   U12986 : AOI22_X1 port map( A1 => n11970, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2220_port, ZN => n5959);
   U12987 : AOI22_X1 port map( A1 => n11971, A2 => n11024, B1 => n11023, B2 => 
                           DataPath_RF_bus_reg_dataout_2221_port, ZN => n5958);
   U12988 : AOI22_X1 port map( A1 => n11972, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2222_port, ZN => n5957);
   U12989 : AOI22_X1 port map( A1 => n11974, A2 => n11024, B1 => n11023, B2 => 
                           DataPath_RF_bus_reg_dataout_2223_port, ZN => n5956);
   U12990 : AOI22_X1 port map( A1 => n11910, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2224_port, ZN => n5955);
   U12991 : AOI22_X1 port map( A1 => n11940, A2 => n11024, B1 => n11023, B2 => 
                           DataPath_RF_bus_reg_dataout_2225_port, ZN => n5954);
   U12992 : AOI22_X1 port map( A1 => n11911, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2226_port, ZN => n5953);
   U12993 : AOI22_X1 port map( A1 => n11942, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2227_port, ZN => n5952);
   U12994 : AOI22_X1 port map( A1 => n11943, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2228_port, ZN => n5951);
   U12995 : AOI22_X1 port map( A1 => n11945, A2 => n11024, B1 => n11023, B2 => 
                           DataPath_RF_bus_reg_dataout_2229_port, ZN => n5950);
   U12996 : AOI22_X1 port map( A1 => n11912, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2230_port, ZN => n5949);
   U12997 : AOI22_X1 port map( A1 => n11913, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2231_port, ZN => n5948);
   U12998 : AOI22_X1 port map( A1 => n11914, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2232_port, ZN => n5947);
   U12999 : AOI22_X1 port map( A1 => n11915, A2 => n11024, B1 => n11023, B2 => 
                           DataPath_RF_bus_reg_dataout_2233_port, ZN => n5946);
   U13000 : AOI22_X1 port map( A1 => n11916, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2234_port, ZN => n5945);
   U13001 : AOI22_X1 port map( A1 => n11917, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2235_port, ZN => n5944);
   U13002 : AOI22_X1 port map( A1 => n11918, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2236_port, ZN => n5943);
   U13003 : AOI22_X1 port map( A1 => n11919, A2 => n11024, B1 => n11023, B2 => 
                           DataPath_RF_bus_reg_dataout_2237_port, ZN => n5942);
   U13004 : AOI22_X1 port map( A1 => n11920, A2 => n11024, B1 => n11023, B2 => 
                           DataPath_RF_bus_reg_dataout_2238_port, ZN => n5941);
   U13005 : AOI22_X1 port map( A1 => n11921, A2 => n11024, B1 => n8481, B2 => 
                           DataPath_RF_bus_reg_dataout_2239_port, ZN => n5938);
   U13006 : INV_X1 port map( A => n11045, ZN => n11025);
   U13007 : NAND2_X1 port map( A1 => n11044, A2 => n11629, ZN => n11562);
   U13008 : INV_X1 port map( A => n11026, ZN => n11027);
   U13009 : OAI22_X1 port map( A1 => n8219, A2 => n11562, B1 => n11923, B2 => 
                           n11561, ZN => n11028);
   U13010 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2176_port, B1 => n11958,
                           B2 => n8408, ZN => n5935);
   U13011 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2177_port, B1 => n11959,
                           B2 => n8408, ZN => n5934);
   U13012 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2178_port, B1 => n11960,
                           B2 => n8408, ZN => n5933);
   U13013 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2179_port, B1 => n11961,
                           B2 => n8408, ZN => n5932);
   U13014 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2180_port, B1 => n11962,
                           B2 => n8408, ZN => n5931);
   U13015 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2181_port, B1 => n11963,
                           B2 => n8408, ZN => n5930);
   U13016 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2182_port, B1 => n11964,
                           B2 => n8408, ZN => n5929);
   U13017 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2183_port, B1 => n11965,
                           B2 => n8408, ZN => n5928);
   U13018 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2184_port, B1 => n11966,
                           B2 => n8408, ZN => n5927);
   U13019 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2185_port, B1 => n11967,
                           B2 => n8408, ZN => n5926);
   U13020 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2186_port, B1 => n11968,
                           B2 => n8408, ZN => n5925);
   U13021 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2187_port, B1 => n11969,
                           B2 => n8408, ZN => n5924);
   U13022 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2188_port, B1 => n11970,
                           B2 => n8408, ZN => n5923);
   U13023 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2189_port, B1 => n11971,
                           B2 => n8408, ZN => n5922);
   U13024 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2190_port, B1 => n11972,
                           B2 => n8408, ZN => n5921);
   U13025 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2191_port, B1 => n11974,
                           B2 => n8408, ZN => n5920);
   U13026 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2192_port, B1 => n11910,
                           B2 => n8408, ZN => n5919);
   U13027 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2193_port, B1 => n11940,
                           B2 => n8408, ZN => n5918);
   U13028 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2194_port, B1 => n11911,
                           B2 => n8408, ZN => n5917);
   U13029 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2195_port, B1 => n11942,
                           B2 => n8408, ZN => n5916);
   U13030 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2196_port, B1 => n11943,
                           B2 => n8408, ZN => n5915);
   U13031 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2197_port, B1 => n11945,
                           B2 => n8408, ZN => n5914);
   U13032 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2198_port, B1 => n11912,
                           B2 => n8408, ZN => n5913);
   U13033 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2199_port, B1 => n11913,
                           B2 => n8408, ZN => n5912);
   U13034 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2200_port, B1 => n11914,
                           B2 => n8408, ZN => n5911);
   U13035 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2201_port, B1 => n11915,
                           B2 => n8408, ZN => n5910);
   U13036 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2202_port, B1 => n11916,
                           B2 => n8408, ZN => n5909);
   U13037 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2203_port, B1 => n11917,
                           B2 => n8408, ZN => n5908);
   U13038 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2204_port, B1 => n11918,
                           B2 => n8408, ZN => n5907);
   U13039 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2205_port, B1 => n11919,
                           B2 => n8408, ZN => n5906);
   U13040 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2206_port, B1 => n11920,
                           B2 => n8408, ZN => n5905);
   U13041 : AOI22_X1 port map( A1 => n7760, A2 => 
                           DataPath_RF_bus_reg_dataout_2207_port, B1 => n11921,
                           B2 => n8408, ZN => n5902);
   U13042 : NAND2_X1 port map( A1 => n11045, A2 => n11633, ZN => n11567);
   U13043 : NAND2_X1 port map( A1 => n11044, A2 => n11633, ZN => n11568);
   U13044 : INV_X1 port map( A => n11030, ZN => n11031);
   U13045 : OAI22_X1 port map( A1 => n8219, A2 => n11568, B1 => n11923, B2 => 
                           n11569, ZN => n11032);
   U13046 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2144_port, B1 => n11958,
                           B2 => n8409, ZN => n5899);
   U13047 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2145_port, B1 => n11959,
                           B2 => n8409, ZN => n5898);
   U13048 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2146_port, B1 => n11960,
                           B2 => n8409, ZN => n5897);
   U13049 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2147_port, B1 => n11961,
                           B2 => n8409, ZN => n5896);
   U13050 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2148_port, B1 => n11962,
                           B2 => n8409, ZN => n5895);
   U13051 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2149_port, B1 => n11963,
                           B2 => n8409, ZN => n5894);
   U13052 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2150_port, B1 => n11964,
                           B2 => n8409, ZN => n5893);
   U13053 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2151_port, B1 => n11965,
                           B2 => n8409, ZN => n5892);
   U13054 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2152_port, B1 => n11966,
                           B2 => n8409, ZN => n5891);
   U13055 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2153_port, B1 => n11967,
                           B2 => n8409, ZN => n5890);
   U13056 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2154_port, B1 => n11968,
                           B2 => n8409, ZN => n5889);
   U13057 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2155_port, B1 => n11969,
                           B2 => n8409, ZN => n5888);
   U13058 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2156_port, B1 => n11970,
                           B2 => n8409, ZN => n5887);
   U13059 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2157_port, B1 => n11971,
                           B2 => n8409, ZN => n5886);
   U13060 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2158_port, B1 => n11972,
                           B2 => n8409, ZN => n5885);
   U13061 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2159_port, B1 => n11974,
                           B2 => n8409, ZN => n5884);
   U13062 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2160_port, B1 => n11910,
                           B2 => n8409, ZN => n5883);
   U13063 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2161_port, B1 => n11940,
                           B2 => n8409, ZN => n5882);
   U13064 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2162_port, B1 => n11911,
                           B2 => n8409, ZN => n5881);
   U13065 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2163_port, B1 => n11942,
                           B2 => n8409, ZN => n5880);
   U13066 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2164_port, B1 => n11943,
                           B2 => n8409, ZN => n5879);
   U13067 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2165_port, B1 => n11945,
                           B2 => n8409, ZN => n5878);
   U13068 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2166_port, B1 => n11912,
                           B2 => n8409, ZN => n5877);
   U13069 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2167_port, B1 => n11913,
                           B2 => n8409, ZN => n5876);
   U13070 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2168_port, B1 => n11914,
                           B2 => n8409, ZN => n5875);
   U13071 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2169_port, B1 => n11915,
                           B2 => n8409, ZN => n5874);
   U13072 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2170_port, B1 => n11916,
                           B2 => n8409, ZN => n5873);
   U13073 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2171_port, B1 => n11917,
                           B2 => n8409, ZN => n5872);
   U13074 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2172_port, B1 => n11918,
                           B2 => n8409, ZN => n5871);
   U13075 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2173_port, B1 => n11919,
                           B2 => n8409, ZN => n5870);
   U13076 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2174_port, B1 => n11920,
                           B2 => n8409, ZN => n5869);
   U13077 : AOI22_X1 port map( A1 => n7761, A2 => 
                           DataPath_RF_bus_reg_dataout_2175_port, B1 => n11921,
                           B2 => n8409, ZN => n5866);
   U13078 : INV_X1 port map( A => n11034, ZN => n11035);
   U13079 : NAND2_X1 port map( A1 => n11638, A2 => n11045, ZN => n11572);
   U13080 : NAND2_X1 port map( A1 => n11638, A2 => n11044, ZN => n11573);
   U13081 : OAI22_X1 port map( A1 => n576, A2 => n11572, B1 => n11573, B2 => 
                           n8219, ZN => n11036);
   U13082 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2112_port, B1 => n11958,
                           B2 => n11037, ZN => n5863);
   U13083 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2113_port, B1 => n11959,
                           B2 => n11037, ZN => n5862);
   U13084 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2114_port, B1 => n11960,
                           B2 => n11037, ZN => n5861);
   U13085 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2115_port, B1 => n11961,
                           B2 => n11037, ZN => n5860);
   U13086 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2116_port, B1 => n11962,
                           B2 => n11037, ZN => n5859);
   U13087 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2117_port, B1 => n11963,
                           B2 => n11037, ZN => n5858);
   U13088 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2118_port, B1 => n11964,
                           B2 => n11037, ZN => n5857);
   U13089 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2119_port, B1 => n11965,
                           B2 => n11037, ZN => n5856);
   U13090 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2120_port, B1 => n11966,
                           B2 => n11037, ZN => n5855);
   U13091 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2121_port, B1 => n11967,
                           B2 => n11037, ZN => n5854);
   U13092 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2122_port, B1 => n11968,
                           B2 => n11037, ZN => n5853);
   U13093 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2123_port, B1 => n11969,
                           B2 => n11037, ZN => n5852);
   U13094 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2124_port, B1 => n11970,
                           B2 => n11037, ZN => n5851);
   U13095 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2125_port, B1 => n11971,
                           B2 => n11037, ZN => n5850);
   U13096 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2126_port, B1 => n11972,
                           B2 => n11037, ZN => n5849);
   U13097 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2127_port, B1 => n11974,
                           B2 => n11037, ZN => n5848);
   U13098 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2128_port, B1 => n11910,
                           B2 => n11037, ZN => n5847);
   U13099 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2129_port, B1 => n11940,
                           B2 => n11037, ZN => n5846);
   U13100 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2130_port, B1 => n11911,
                           B2 => n11037, ZN => n5845);
   U13101 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2131_port, B1 => n11942,
                           B2 => n11037, ZN => n5844);
   U13102 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2132_port, B1 => n11943,
                           B2 => n11037, ZN => n5843);
   U13103 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2133_port, B1 => n11945,
                           B2 => n11037, ZN => n5842);
   U13104 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2134_port, B1 => n11912,
                           B2 => n11037, ZN => n5841);
   U13105 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2135_port, B1 => n11913,
                           B2 => n11037, ZN => n5840);
   U13106 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2136_port, B1 => n11914,
                           B2 => n11037, ZN => n5839);
   U13107 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2137_port, B1 => n11915,
                           B2 => n11037, ZN => n5838);
   U13108 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2138_port, B1 => n11916,
                           B2 => n11037, ZN => n5837);
   U13109 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2139_port, B1 => n11917,
                           B2 => n11037, ZN => n5836);
   U13110 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2140_port, B1 => n11918,
                           B2 => n11037, ZN => n5835);
   U13111 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2141_port, B1 => n11919,
                           B2 => n11037, ZN => n5834);
   U13112 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2142_port, B1 => n11920,
                           B2 => n11037, ZN => n5833);
   U13113 : AOI22_X1 port map( A1 => n11038, A2 => 
                           DataPath_RF_bus_reg_dataout_2143_port, B1 => n11921,
                           B2 => n11037, ZN => n5830);
   U13114 : NAND2_X1 port map( A1 => n11643, A2 => n11045, ZN => n11578);
   U13115 : NAND2_X1 port map( A1 => n11643, A2 => n11044, ZN => n11579);
   U13116 : OAI22_X1 port map( A1 => n576, A2 => n11578, B1 => n11579, B2 => 
                           n8219, ZN => n11040);
   U13117 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2080_port, B1 => n11958,
                           B2 => n11042, ZN => n5827);
   U13118 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2081_port, B1 => n11959,
                           B2 => n11042, ZN => n5826);
   U13119 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2082_port, B1 => n11960,
                           B2 => n11042, ZN => n5825);
   U13120 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2083_port, B1 => n11961,
                           B2 => n11042, ZN => n5824);
   U13121 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2084_port, B1 => n11962,
                           B2 => n11042, ZN => n5823);
   U13122 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2085_port, B1 => n11963,
                           B2 => n11042, ZN => n5822);
   U13123 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2086_port, B1 => n11964,
                           B2 => n11042, ZN => n5821);
   U13124 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2087_port, B1 => n11965,
                           B2 => n11042, ZN => n5820);
   U13125 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2088_port, B1 => n11966,
                           B2 => n11042, ZN => n5819);
   U13126 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2089_port, B1 => n11967,
                           B2 => n11042, ZN => n5818);
   U13127 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2090_port, B1 => n11968,
                           B2 => n11042, ZN => n5817);
   U13128 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2091_port, B1 => n11969,
                           B2 => n11042, ZN => n5816);
   U13129 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2092_port, B1 => n11970,
                           B2 => n11042, ZN => n5815);
   U13130 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2093_port, B1 => n11971,
                           B2 => n11042, ZN => n5814);
   U13131 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2094_port, B1 => n11972,
                           B2 => n11042, ZN => n5813);
   U13132 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2095_port, B1 => n11974,
                           B2 => n11042, ZN => n5812);
   U13133 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2096_port, B1 => n11910,
                           B2 => n11042, ZN => n5811);
   U13134 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2097_port, B1 => n11940,
                           B2 => n11042, ZN => n5810);
   U13135 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2098_port, B1 => n11911,
                           B2 => n11042, ZN => n5809);
   U13136 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2099_port, B1 => n11942,
                           B2 => n11042, ZN => n5808);
   U13137 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2100_port, B1 => n11943,
                           B2 => n11042, ZN => n5807);
   U13138 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2101_port, B1 => n11945,
                           B2 => n11042, ZN => n5806);
   U13139 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2102_port, B1 => n11912,
                           B2 => n11042, ZN => n5805);
   U13140 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2103_port, B1 => n11913,
                           B2 => n11042, ZN => n5804);
   U13141 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2104_port, B1 => n11914,
                           B2 => n11042, ZN => n5803);
   U13142 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2105_port, B1 => n11915,
                           B2 => n11042, ZN => n5802);
   U13143 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2106_port, B1 => n11916,
                           B2 => n11042, ZN => n5801);
   U13144 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2107_port, B1 => n11917,
                           B2 => n11042, ZN => n5800);
   U13145 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2108_port, B1 => n11918,
                           B2 => n11042, ZN => n5799);
   U13146 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2109_port, B1 => n11919,
                           B2 => n11042, ZN => n5798);
   U13147 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2110_port, B1 => n11920,
                           B2 => n11042, ZN => n5797);
   U13148 : AOI22_X1 port map( A1 => n11043, A2 => 
                           DataPath_RF_bus_reg_dataout_2111_port, B1 => n11921,
                           B2 => n11042, ZN => n5794);
   U13149 : NAND2_X1 port map( A1 => n11046, A2 => n11044, ZN => n11584);
   U13150 : NAND2_X1 port map( A1 => n11046, A2 => n11045, ZN => n11583);
   U13151 : OAI222_X1 port map( A1 => n11584, A2 => n8219, B1 => n11583, B2 => 
                           n576, C1 => n11585, C2 => n11923, ZN => n11048);
   U13152 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2048_port, A2 
                           => n8482, B1 => n11049, B2 => n11925, ZN => n5788);
   U13153 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2049_port, A2 
                           => n11050, B1 => n11049, B2 => n11926, ZN => n5787);
   U13154 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2050_port, A2 
                           => n11050, B1 => n11049, B2 => n11927, ZN => n5786);
   U13155 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2051_port, A2 
                           => n8482, B1 => n11049, B2 => n11928, ZN => n5785);
   U13156 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2052_port, A2 
                           => n8482, B1 => n11049, B2 => n11929, ZN => n5784);
   U13157 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2053_port, A2 
                           => n8482, B1 => n11049, B2 => n11930, ZN => n5783);
   U13158 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2054_port, A2 
                           => n8482, B1 => n11049, B2 => n11931, ZN => n5782);
   U13159 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2055_port, A2 
                           => n8482, B1 => n11049, B2 => n11932, ZN => n5781);
   U13160 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2056_port, A2 
                           => n8482, B1 => n11049, B2 => n11898, ZN => n5780);
   U13161 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2057_port, A2 
                           => n11050, B1 => n11049, B2 => n11933, ZN => n5779);
   U13162 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2058_port, A2 
                           => n8482, B1 => n11049, B2 => n11934, ZN => n5778);
   U13163 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2059_port, A2 
                           => n11050, B1 => n11049, B2 => n11935, ZN => n5777);
   U13164 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2060_port, A2 
                           => n8482, B1 => n11049, B2 => n11936, ZN => n5776);
   U13165 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2061_port, A2 
                           => n8482, B1 => n11049, B2 => n11937, ZN => n5775);
   U13166 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2062_port, A2 
                           => n11050, B1 => n11049, B2 => n11899, ZN => n5774);
   U13167 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2063_port, A2 
                           => n8482, B1 => n11049, B2 => n11938, ZN => n5773);
   U13168 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2064_port, A2 
                           => n11050, B1 => n11049, B2 => n11939, ZN => n5772);
   U13169 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2065_port, A2 
                           => n8482, B1 => n11049, B2 => n11900, ZN => n5771);
   U13170 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2066_port, A2 
                           => n8482, B1 => n11049, B2 => n11941, ZN => n5770);
   U13171 : AOI22_X1 port map( A1 => n11942, A2 => n11048, B1 => n8482, B2 => 
                           DataPath_RF_bus_reg_dataout_2067_port, ZN => n5769);
   U13172 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2068_port, A2 
                           => n11050, B1 => n11049, B2 => n11902, ZN => n5768);
   U13173 : AOI22_X1 port map( A1 => n11945, A2 => n11048, B1 => n8482, B2 => 
                           DataPath_RF_bus_reg_dataout_2069_port, ZN => n5767);
   U13174 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2070_port, A2 
                           => n11050, B1 => n11049, B2 => n11946, ZN => n5766);
   U13175 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2071_port, A2 
                           => n8482, B1 => n11049, B2 => n11947, ZN => n5765);
   U13176 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2072_port, A2 
                           => n8482, B1 => n11049, B2 => n11948, ZN => n5764);
   U13177 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2073_port, A2 
                           => n8482, B1 => n11049, B2 => n11949, ZN => n5763);
   U13178 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2074_port, A2 
                           => n11050, B1 => n11049, B2 => n11950, ZN => n5762);
   U13179 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2075_port, A2 
                           => n8482, B1 => n11049, B2 => n11951, ZN => n5761);
   U13180 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2076_port, A2 
                           => n8482, B1 => n11049, B2 => n11952, ZN => n5760);
   U13181 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2077_port, A2 
                           => n11050, B1 => n11049, B2 => n11953, ZN => n5759);
   U13182 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2078_port, A2 
                           => n8482, B1 => n11049, B2 => n11954, ZN => n5758);
   U13183 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2079_port, A2 
                           => n8482, B1 => n11049, B2 => n11955, ZN => n5755);
   U13184 : OAI22_X1 port map( A1 => n8483, A2 => n11450, B1 => n11645, B2 => 
                           n11150, ZN => n11103);
   U13185 : NAND2_X1 port map( A1 => n11082, A2 => n11617, ZN => n11887);
   U13186 : NOR2_X1 port map( A1 => n8417, A2 => n11051, ZN => n11053);
   U13187 : AOI22_X1 port map( A1 => n11155, A2 => n8484, B1 => n8485, B2 => 
                           DataPath_RF_bus_reg_dataout_2016_port, ZN => n5751);
   U13188 : OAI22_X1 port map( A1 => n8483, A2 => n11451, B1 => n11646, B2 => 
                           n11150, ZN => n11104);
   U13189 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2017_port, A2 
                           => n8485, B1 => n11156, B2 => n8484, ZN => n5750);
   U13190 : OAI22_X1 port map( A1 => n11153, A2 => n11452, B1 => n11647, B2 => 
                           n11150, ZN => n11105);
   U13191 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2018_port, A2 
                           => n8485, B1 => n11157, B2 => n8484, ZN => n5749);
   U13192 : OAI22_X1 port map( A1 => n8483, A2 => n11453, B1 => n11648, B2 => 
                           n11150, ZN => n11106);
   U13193 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2019_port, A2 
                           => n11055, B1 => n11158, B2 => n11054, ZN => n5748);
   U13194 : OAI22_X1 port map( A1 => n11153, A2 => n11454, B1 => n11649, B2 => 
                           n11150, ZN => n11107);
   U13195 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2020_port, A2 
                           => n8485, B1 => n11159, B2 => n11054, ZN => n5747);
   U13196 : AOI22_X1 port map( A1 => n11150, A2 => n11456, B1 => n11455, B2 => 
                           n11153, ZN => n11062);
   U13197 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2021_port, A2 
                           => n11055, B1 => n11160, B2 => n8484, ZN => n5746);
   U13198 : OAI22_X1 port map( A1 => n11153, A2 => n11457, B1 => n11651, B2 => 
                           n11150, ZN => n11109);
   U13199 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2022_port, A2 
                           => n8485, B1 => n11161, B2 => n8484, ZN => n5745);
   U13200 : OAI22_X1 port map( A1 => n11153, A2 => n11458, B1 => n11652, B2 => 
                           n11150, ZN => n11110);
   U13201 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2023_port, A2 
                           => n11055, B1 => n11162, B2 => n8484, ZN => n5744);
   U13202 : OAI22_X1 port map( A1 => n11153, A2 => n11459, B1 => n11653, B2 => 
                           n11150, ZN => n11111);
   U13203 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2024_port, A2 
                           => n8485, B1 => n11163, B2 => n11054, ZN => n5743);
   U13204 : AOI22_X1 port map( A1 => n11150, A2 => n11461, B1 => n11460, B2 => 
                           n11153, ZN => n11063);
   U13205 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2025_port, A2 
                           => n8485, B1 => n11164, B2 => n8484, ZN => n5742);
   U13206 : OAI22_X1 port map( A1 => n11153, A2 => n11462, B1 => n11655, B2 => 
                           n11150, ZN => n11113);
   U13207 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2026_port, A2 
                           => n8485, B1 => n11165, B2 => n8484, ZN => n5741);
   U13208 : OAI22_X1 port map( A1 => n8483, A2 => n11463, B1 => n11656, B2 => 
                           n11150, ZN => n11114);
   U13209 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2027_port, A2 
                           => n8485, B1 => n11166, B2 => n8484, ZN => n5740);
   U13210 : OAI22_X1 port map( A1 => n8483, A2 => n11464, B1 => n11657, B2 => 
                           n11150, ZN => n11115);
   U13211 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2028_port, A2 
                           => n11055, B1 => n11167, B2 => n11054, ZN => n5739);
   U13212 : OAI22_X1 port map( A1 => n8483, A2 => n11465, B1 => n11658, B2 => 
                           n11150, ZN => n11116);
   U13213 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2029_port, A2 
                           => n8485, B1 => n11168, B2 => n11054, ZN => n5738);
   U13214 : OAI22_X1 port map( A1 => n11153, A2 => n11466, B1 => n11659, B2 => 
                           n11150, ZN => n11117);
   U13215 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2030_port, A2 
                           => n11055, B1 => n11169, B2 => n8484, ZN => n5737);
   U13216 : AOI22_X1 port map( A1 => n11150, A2 => n11468, B1 => n11467, B2 => 
                           n8483, ZN => n11064);
   U13217 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2031_port, A2 
                           => n8485, B1 => n11170, B2 => n8484, ZN => n5736);
   U13218 : AOI22_X1 port map( A1 => n11150, A2 => n11470, B1 => n11469, B2 => 
                           n8483, ZN => n11065);
   U13219 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2032_port, A2 
                           => n11055, B1 => n11171, B2 => n8484, ZN => n5735);
   U13220 : AOI22_X1 port map( A1 => n11150, A2 => n11472, B1 => n11471, B2 => 
                           n8483, ZN => n11066);
   U13221 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2033_port, A2 
                           => n8485, B1 => n11172, B2 => n11054, ZN => n5734);
   U13222 : OAI22_X1 port map( A1 => n11153, A2 => n11473, B1 => n11663, B2 => 
                           n11150, ZN => n11121);
   U13223 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2034_port, A2 
                           => n8485, B1 => n11173, B2 => n8484, ZN => n5733);
   U13224 : AOI22_X1 port map( A1 => n11150, A2 => n11475, B1 => n11474, B2 => 
                           n11153, ZN => n11077);
   U13225 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2035_port, A2 
                           => n8485, B1 => n11174, B2 => n8484, ZN => n5732);
   U13226 : OAI22_X1 port map( A1 => n11153, A2 => n11319, B1 => n11665, B2 => 
                           n11150, ZN => n11123);
   U13227 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2036_port, A2 
                           => n8485, B1 => n11175, B2 => n8484, ZN => n5731);
   U13228 : OAI22_X1 port map( A1 => n11153, A2 => n11477, B1 => n11666, B2 => 
                           n11150, ZN => n11124);
   U13229 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2037_port, A2 
                           => n11055, B1 => n11176, B2 => n11054, ZN => n5730);
   U13230 : OAI22_X1 port map( A1 => n8483, A2 => n11478, B1 => n11667, B2 => 
                           n11150, ZN => n11125);
   U13231 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2038_port, A2 
                           => n8485, B1 => n11177, B2 => n11054, ZN => n5729);
   U13232 : AOI22_X1 port map( A1 => n11150, A2 => n11480, B1 => n11479, B2 => 
                           n11153, ZN => n11078);
   U13233 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2039_port, A2 
                           => n11055, B1 => n11178, B2 => n8484, ZN => n5728);
   U13234 : AOI22_X1 port map( A1 => n11150, A2 => n11482, B1 => n11481, B2 => 
                           n8483, ZN => n11067);
   U13235 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2040_port, A2 
                           => n8485, B1 => n11179, B2 => n8484, ZN => n5727);
   U13236 : AOI22_X1 port map( A1 => n11150, A2 => n11484, B1 => n11483, B2 => 
                           n11153, ZN => n11068);
   U13237 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2041_port, A2 
                           => n8485, B1 => n11180, B2 => n8484, ZN => n5726);
   U13238 : OAI22_X1 port map( A1 => n11153, A2 => n11485, B1 => n11671, B2 => 
                           n11150, ZN => n11129);
   U13239 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2042_port, A2 
                           => n8485, B1 => n11181, B2 => n8484, ZN => n5725);
   U13240 : AOI22_X1 port map( A1 => n11150, A2 => n11487, B1 => n11486, B2 => 
                           n8483, ZN => n11086);
   U13241 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2043_port, A2 
                           => n8485, B1 => n11182, B2 => n8484, ZN => n5724);
   U13242 : AOI22_X1 port map( A1 => n11150, A2 => n11489, B1 => n11488, B2 => 
                           n11153, ZN => n11070);
   U13243 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2044_port, A2 
                           => n8485, B1 => n11183, B2 => n8484, ZN => n5723);
   U13244 : OAI22_X1 port map( A1 => n11153, A2 => n11320, B1 => n11674, B2 => 
                           n11150, ZN => n11132);
   U13245 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2045_port, A2 
                           => n11055, B1 => n11184, B2 => n8484, ZN => n5722);
   U13246 : AOI22_X1 port map( A1 => n11150, A2 => n11493, B1 => n11492, B2 => 
                           n8483, ZN => n11071);
   U13247 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2046_port, A2 
                           => n8485, B1 => n11185, B2 => n8484, ZN => n5721);
   U13248 : AOI22_X1 port map( A1 => n11150, A2 => n11495, B1 => n11494, B2 => 
                           n8483, ZN => n11072);
   U13249 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2047_port, A2 
                           => n11055, B1 => n11186, B2 => n11054, ZN => n5718);
   U13250 : NAND2_X1 port map( A1 => n11082, A2 => n11621, ZN => n11892);
   U13251 : INV_X1 port map( A => n11056, ZN => n11057);
   U13252 : AOI22_X1 port map( A1 => n11155, A2 => n8486, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_1984_port, ZN => n5714);
   U13253 : AOI22_X1 port map( A1 => n11156, A2 => n8486, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_1985_port, ZN => n5713);
   U13254 : AOI22_X1 port map( A1 => n11157, A2 => n8486, B1 => n11058, B2 => 
                           DataPath_RF_bus_reg_dataout_1986_port, ZN => n5712);
   U13255 : AOI22_X1 port map( A1 => n11158, A2 => n8486, B1 => n11058, B2 => 
                           DataPath_RF_bus_reg_dataout_1987_port, ZN => n5711);
   U13256 : AOI22_X1 port map( A1 => n11159, A2 => n8486, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_1988_port, ZN => n5710);
   U13257 : AOI22_X1 port map( A1 => n11160, A2 => n8486, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_1989_port, ZN => n5709);
   U13258 : AOI22_X1 port map( A1 => n11161, A2 => n11059, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_1990_port, ZN => n5708);
   U13259 : OAI22_X1 port map( A1 => n11162, A2 => n11058, B1 => 
                           DataPath_RF_bus_reg_dataout_1991_port, B2 => n8486, 
                           ZN => n5707);
   U13260 : AOI22_X1 port map( A1 => n11163, A2 => n8486, B1 => n11058, B2 => 
                           DataPath_RF_bus_reg_dataout_1992_port, ZN => n5706);
   U13261 : AOI22_X1 port map( A1 => n11164, A2 => n11059, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_1993_port, ZN => n5705);
   U13262 : OAI22_X1 port map( A1 => n11165, A2 => n8487, B1 => 
                           DataPath_RF_bus_reg_dataout_1994_port, B2 => n8486, 
                           ZN => n5704);
   U13263 : AOI22_X1 port map( A1 => n11166, A2 => n8486, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_1995_port, ZN => n5703);
   U13264 : AOI22_X1 port map( A1 => n11167, A2 => n11059, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_1996_port, ZN => n5702);
   U13265 : AOI22_X1 port map( A1 => n11168, A2 => n8486, B1 => n11058, B2 => 
                           DataPath_RF_bus_reg_dataout_1997_port, ZN => n5701);
   U13266 : OAI22_X1 port map( A1 => n11169, A2 => n8487, B1 => 
                           DataPath_RF_bus_reg_dataout_1998_port, B2 => n11059,
                           ZN => n5700);
   U13267 : AOI22_X1 port map( A1 => n11170, A2 => n8486, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_1999_port, ZN => n5699);
   U13268 : AOI22_X1 port map( A1 => n11171, A2 => n8486, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_2000_port, ZN => n5698);
   U13269 : AOI22_X1 port map( A1 => n11172, A2 => n8486, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_2001_port, ZN => n5697);
   U13270 : AOI22_X1 port map( A1 => n11173, A2 => n11059, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_2002_port, ZN => n5696);
   U13271 : AOI22_X1 port map( A1 => n11174, A2 => n8486, B1 => n11058, B2 => 
                           DataPath_RF_bus_reg_dataout_2003_port, ZN => n5695);
   U13272 : AOI22_X1 port map( A1 => n11175, A2 => n11059, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_2004_port, ZN => n5694);
   U13273 : OAI22_X1 port map( A1 => n11176, A2 => n8487, B1 => 
                           DataPath_RF_bus_reg_dataout_2005_port, B2 => n8486, 
                           ZN => n5693);
   U13274 : AOI22_X1 port map( A1 => n11177, A2 => n8486, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_2006_port, ZN => n5692);
   U13275 : OAI22_X1 port map( A1 => n11178, A2 => n8487, B1 => 
                           DataPath_RF_bus_reg_dataout_2007_port, B2 => n8486, 
                           ZN => n5691);
   U13276 : OAI22_X1 port map( A1 => n11179, A2 => n11058, B1 => 
                           DataPath_RF_bus_reg_dataout_2008_port, B2 => n8486, 
                           ZN => n5690);
   U13277 : AOI22_X1 port map( A1 => n11180, A2 => n11059, B1 => n11058, B2 => 
                           DataPath_RF_bus_reg_dataout_2009_port, ZN => n5689);
   U13278 : OAI22_X1 port map( A1 => n11181, A2 => n8487, B1 => 
                           DataPath_RF_bus_reg_dataout_2010_port, B2 => n8486, 
                           ZN => n5688);
   U13279 : AOI22_X1 port map( A1 => n11182, A2 => n8486, B1 => n11058, B2 => 
                           DataPath_RF_bus_reg_dataout_2011_port, ZN => n5687);
   U13280 : AOI22_X1 port map( A1 => n11183, A2 => n8486, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_2012_port, ZN => n5686);
   U13281 : AOI22_X1 port map( A1 => n11184, A2 => n8486, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_2013_port, ZN => n5685);
   U13282 : AOI22_X1 port map( A1 => n11185, A2 => n8486, B1 => n8487, B2 => 
                           DataPath_RF_bus_reg_dataout_2014_port, ZN => n5684);
   U13283 : AOI22_X1 port map( A1 => n11186, A2 => n11059, B1 => n11058, B2 => 
                           DataPath_RF_bus_reg_dataout_2015_port, ZN => n5681);
   U13284 : NAND2_X1 port map( A1 => n11082, A2 => n11625, ZN => n11897);
   U13285 : INV_X1 port map( A => n11060, ZN => n11061);
   U13286 : AOI22_X1 port map( A1 => n11155, A2 => n11069, B1 => n8488, B2 => 
                           DataPath_RF_bus_reg_dataout_1952_port, ZN => n5677);
   U13287 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1953_port, A2 
                           => n8488, B1 => n11073, B2 => n11104, ZN => n5676);
   U13288 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1954_port, A2 
                           => n8488, B1 => n11073, B2 => n11105, ZN => n5675);
   U13289 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1955_port, A2 
                           => n8488, B1 => n11073, B2 => n11106, ZN => n5674);
   U13290 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1956_port, A2 
                           => n8488, B1 => n11073, B2 => n11107, ZN => n5673);
   U13291 : INV_X1 port map( A => n11062, ZN => n11108);
   U13292 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1957_port, A2 
                           => n11074, B1 => n11073, B2 => n11108, ZN => n5672);
   U13293 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1958_port, A2 
                           => n11074, B1 => n11073, B2 => n11109, ZN => n5671);
   U13294 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1959_port, A2 
                           => n11074, B1 => n11073, B2 => n11110, ZN => n5670);
   U13295 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1960_port, A2 
                           => n8488, B1 => n11073, B2 => n11111, ZN => n5669);
   U13296 : INV_X1 port map( A => n11063, ZN => n11112);
   U13297 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1961_port, A2 
                           => n8488, B1 => n11073, B2 => n11112, ZN => n5668);
   U13298 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1962_port, A2 
                           => n8488, B1 => n11073, B2 => n11113, ZN => n5667);
   U13299 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1963_port, A2 
                           => n8488, B1 => n11073, B2 => n11114, ZN => n5666);
   U13300 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1964_port, A2 
                           => n8488, B1 => n11073, B2 => n11115, ZN => n5665);
   U13301 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1965_port, A2 
                           => n8488, B1 => n11073, B2 => n11116, ZN => n5664);
   U13302 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1966_port, A2 
                           => n11074, B1 => n11073, B2 => n11117, ZN => n5663);
   U13303 : INV_X1 port map( A => n11064, ZN => n11118);
   U13304 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1967_port, A2 
                           => n11074, B1 => n11073, B2 => n11118, ZN => n5662);
   U13305 : INV_X1 port map( A => n11065, ZN => n11119);
   U13306 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1968_port, A2 
                           => n8488, B1 => n11073, B2 => n11119, ZN => n5661);
   U13307 : INV_X1 port map( A => n11066, ZN => n11120);
   U13308 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1969_port, A2 
                           => n8488, B1 => n11073, B2 => n11120, ZN => n5660);
   U13309 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1970_port, A2 
                           => n8488, B1 => n11073, B2 => n11121, ZN => n5659);
   U13310 : AOI22_X1 port map( A1 => n11174, A2 => n11069, B1 => n11074, B2 => 
                           DataPath_RF_bus_reg_dataout_1971_port, ZN => n5658);
   U13311 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1972_port, A2 
                           => n8488, B1 => n11073, B2 => n11123, ZN => n5657);
   U13312 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1973_port, A2 
                           => n8488, B1 => n11073, B2 => n11124, ZN => n5656);
   U13313 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1974_port, A2 
                           => n11074, B1 => n11073, B2 => n11125, ZN => n5655);
   U13314 : AOI22_X1 port map( A1 => n11178, A2 => n11069, B1 => n11074, B2 => 
                           DataPath_RF_bus_reg_dataout_1975_port, ZN => n5654);
   U13315 : INV_X1 port map( A => n11067, ZN => n11127);
   U13316 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1976_port, A2 
                           => n11074, B1 => n11073, B2 => n11127, ZN => n5653);
   U13317 : INV_X1 port map( A => n11068, ZN => n11128);
   U13318 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1977_port, A2 
                           => n8488, B1 => n11073, B2 => n11128, ZN => n5652);
   U13319 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1978_port, A2 
                           => n11074, B1 => n11073, B2 => n11129, ZN => n5651);
   U13320 : AOI22_X1 port map( A1 => n11182, A2 => n11069, B1 => n8488, B2 => 
                           DataPath_RF_bus_reg_dataout_1979_port, ZN => n5650);
   U13321 : INV_X1 port map( A => n11070, ZN => n11131);
   U13322 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1980_port, A2 
                           => n8488, B1 => n11073, B2 => n11131, ZN => n5649);
   U13323 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1981_port, A2 
                           => n8488, B1 => n11073, B2 => n11132, ZN => n5648);
   U13324 : INV_X1 port map( A => n11071, ZN => n11133);
   U13325 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1982_port, A2 
                           => n8488, B1 => n11073, B2 => n11133, ZN => n5647);
   U13326 : INV_X1 port map( A => n11072, ZN => n11094);
   U13327 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1983_port, A2 
                           => n8488, B1 => n11073, B2 => n11094, ZN => n5644);
   U13328 : NAND2_X1 port map( A1 => n11082, A2 => n11629, ZN => n11908);
   U13329 : INV_X1 port map( A => n11075, ZN => n11076);
   U13330 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1920_port, A2 
                           => n8489, B1 => n11079, B2 => n11103, ZN => n5640);
   U13331 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1921_port, A2 
                           => n8489, B1 => n11079, B2 => n11104, ZN => n5639);
   U13332 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1922_port, A2 
                           => n8489, B1 => n11079, B2 => n11105, ZN => n5638);
   U13333 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1923_port, A2 
                           => n11080, B1 => n11079, B2 => n11106, ZN => n5637);
   U13334 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1924_port, A2 
                           => n11080, B1 => n11079, B2 => n11107, ZN => n5636);
   U13335 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1925_port, A2 
                           => n11080, B1 => n11079, B2 => n11108, ZN => n5635);
   U13336 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1926_port, A2 
                           => n8489, B1 => n11079, B2 => n11109, ZN => n5634);
   U13337 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1927_port, A2 
                           => n8489, B1 => n11079, B2 => n11110, ZN => n5633);
   U13338 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1928_port, A2 
                           => n8489, B1 => n11079, B2 => n11111, ZN => n5632);
   U13339 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1929_port, A2 
                           => n8489, B1 => n11079, B2 => n11112, ZN => n5631);
   U13340 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1930_port, A2 
                           => n8489, B1 => n11079, B2 => n11113, ZN => n5630);
   U13341 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1931_port, A2 
                           => n8489, B1 => n11079, B2 => n11114, ZN => n5629);
   U13342 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1932_port, A2 
                           => n11080, B1 => n11079, B2 => n11115, ZN => n5628);
   U13343 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1933_port, A2 
                           => n11080, B1 => n11079, B2 => n11116, ZN => n5627);
   U13344 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1934_port, A2 
                           => n11080, B1 => n11079, B2 => n11117, ZN => n5626);
   U13345 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1935_port, A2 
                           => n8489, B1 => n11079, B2 => n11118, ZN => n5625);
   U13346 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1936_port, A2 
                           => n11080, B1 => n11079, B2 => n11119, ZN => n5624);
   U13347 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1937_port, A2 
                           => n8489, B1 => n11079, B2 => n11120, ZN => n5623);
   U13348 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1938_port, A2 
                           => n8489, B1 => n11079, B2 => n11121, ZN => n5622);
   U13349 : INV_X1 port map( A => n11077, ZN => n11122);
   U13350 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1939_port, A2 
                           => n8489, B1 => n11079, B2 => n11122, ZN => n5621);
   U13351 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1940_port, A2 
                           => n8489, B1 => n11079, B2 => n11123, ZN => n5620);
   U13352 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1941_port, A2 
                           => n8489, B1 => n11079, B2 => n11124, ZN => n5619);
   U13353 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1942_port, A2 
                           => n8489, B1 => n11079, B2 => n11125, ZN => n5618);
   U13354 : INV_X1 port map( A => n11078, ZN => n11126);
   U13355 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1943_port, A2 
                           => n11080, B1 => n11079, B2 => n11126, ZN => n5617);
   U13356 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1944_port, A2 
                           => n8489, B1 => n11079, B2 => n11127, ZN => n5616);
   U13357 : AOI22_X1 port map( A1 => n11180, A2 => n11081, B1 => n8489, B2 => 
                           DataPath_RF_bus_reg_dataout_1945_port, ZN => n5615);
   U13358 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1946_port, A2 
                           => n8489, B1 => n11079, B2 => n11129, ZN => n5614);
   U13359 : AOI22_X1 port map( A1 => n11182, A2 => n11081, B1 => n11080, B2 => 
                           DataPath_RF_bus_reg_dataout_1947_port, ZN => n5613);
   U13360 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1948_port, A2 
                           => n8489, B1 => n11079, B2 => n11131, ZN => n5612);
   U13361 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1949_port, A2 
                           => n11080, B1 => n11079, B2 => n11132, ZN => n5611);
   U13362 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1950_port, A2 
                           => n8489, B1 => n11079, B2 => n11133, ZN => n5610);
   U13363 : AOI22_X1 port map( A1 => n11186, A2 => n11081, B1 => n8489, B2 => 
                           DataPath_RF_bus_reg_dataout_1951_port, ZN => n5607);
   U13364 : NAND2_X1 port map( A1 => n11082, A2 => n11633, ZN => n11924);
   U13365 : INV_X1 port map( A => n11083, ZN => n11085);
   U13366 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1888_port, A2 
                           => n8490, B1 => n11088, B2 => n11103, ZN => n5601);
   U13367 : AOI22_X1 port map( A1 => n11156, A2 => n11087, B1 => n8490, B2 => 
                           DataPath_RF_bus_reg_dataout_1889_port, ZN => n5600);
   U13368 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1890_port, A2 
                           => n8490, B1 => n11088, B2 => n11105, ZN => n5599);
   U13369 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1891_port, A2 
                           => n8490, B1 => n11088, B2 => n11106, ZN => n5598);
   U13370 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1892_port, A2 
                           => n8490, B1 => n11088, B2 => n11107, ZN => n5597);
   U13371 : AOI22_X1 port map( A1 => n11160, A2 => n11087, B1 => n8490, B2 => 
                           DataPath_RF_bus_reg_dataout_1893_port, ZN => n5596);
   U13372 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1894_port, A2 
                           => n8490, B1 => n11088, B2 => n11109, ZN => n5595);
   U13373 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1895_port, A2 
                           => n11089, B1 => n11088, B2 => n11110, ZN => n5594);
   U13374 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1896_port, A2 
                           => n8490, B1 => n11088, B2 => n11111, ZN => n5593);
   U13375 : AOI22_X1 port map( A1 => n11164, A2 => n11087, B1 => n8490, B2 => 
                           DataPath_RF_bus_reg_dataout_1897_port, ZN => n5592);
   U13376 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1898_port, A2 
                           => n11089, B1 => n11088, B2 => n11113, ZN => n5591);
   U13377 : AOI22_X1 port map( A1 => n11166, A2 => n11087, B1 => n11089, B2 => 
                           DataPath_RF_bus_reg_dataout_1899_port, ZN => n5590);
   U13378 : AOI22_X1 port map( A1 => n11167, A2 => n11087, B1 => n8490, B2 => 
                           DataPath_RF_bus_reg_dataout_1900_port, ZN => n5589);
   U13379 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1901_port, A2 
                           => n11089, B1 => n11088, B2 => n11116, ZN => n5588);
   U13380 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1902_port, A2 
                           => n8490, B1 => n11088, B2 => n11117, ZN => n5587);
   U13381 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1903_port, A2 
                           => n8490, B1 => n11088, B2 => n11118, ZN => n5586);
   U13382 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1904_port, A2 
                           => n8490, B1 => n11088, B2 => n11119, ZN => n5585);
   U13383 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1905_port, A2 
                           => n11089, B1 => n11088, B2 => n11120, ZN => n5584);
   U13384 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1906_port, A2 
                           => n8490, B1 => n11088, B2 => n11121, ZN => n5583);
   U13385 : AOI22_X1 port map( A1 => n11174, A2 => n11087, B1 => n11089, B2 => 
                           DataPath_RF_bus_reg_dataout_1907_port, ZN => n5582);
   U13386 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1908_port, A2 
                           => n8490, B1 => n11088, B2 => n11123, ZN => n5581);
   U13387 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1909_port, A2 
                           => n8490, B1 => n11088, B2 => n11124, ZN => n5580);
   U13388 : AOI22_X1 port map( A1 => n11177, A2 => n11087, B1 => n8490, B2 => 
                           DataPath_RF_bus_reg_dataout_1910_port, ZN => n5579);
   U13389 : AOI22_X1 port map( A1 => n11178, A2 => n11087, B1 => n11089, B2 => 
                           DataPath_RF_bus_reg_dataout_1911_port, ZN => n5578);
   U13390 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1912_port, A2 
                           => n11089, B1 => n11088, B2 => n11127, ZN => n5577);
   U13391 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1913_port, A2 
                           => n8490, B1 => n11088, B2 => n11128, ZN => n5576);
   U13392 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1914_port, A2 
                           => n11089, B1 => n11088, B2 => n11129, ZN => n5575);
   U13393 : INV_X1 port map( A => n11086, ZN => n11130);
   U13394 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1915_port, A2 
                           => n8490, B1 => n11088, B2 => n11130, ZN => n5574);
   U13395 : AOI22_X1 port map( A1 => n11183, A2 => n11087, B1 => n8490, B2 => 
                           DataPath_RF_bus_reg_dataout_1916_port, ZN => n5573);
   U13396 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1917_port, A2 
                           => n8490, B1 => n11088, B2 => n11132, ZN => n5572);
   U13397 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1918_port, A2 
                           => n11089, B1 => n11088, B2 => n11133, ZN => n5571);
   U13398 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1919_port, A2 
                           => n8490, B1 => n11088, B2 => n11094, ZN => n5568);
   U13399 : OAI22_X1 port map( A1 => n576, A2 => n11512, B1 => n11513, B2 => 
                           n11153, ZN => n11090);
   U13400 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1856_port, A2 
                           => n8491, B1 => n11091, B2 => n11103, ZN => n5566);
   U13401 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1857_port, A2 
                           => n8491, B1 => n11091, B2 => n11104, ZN => n5565);
   U13402 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1858_port, A2 
                           => n8491, B1 => n11091, B2 => n11105, ZN => n5564);
   U13403 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1859_port, A2 
                           => n11092, B1 => n11091, B2 => n11106, ZN => n5563);
   U13404 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1860_port, A2 
                           => n8491, B1 => n11091, B2 => n11107, ZN => n5562);
   U13405 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1861_port, A2 
                           => n8491, B1 => n11091, B2 => n11108, ZN => n5561);
   U13406 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1862_port, A2 
                           => n8491, B1 => n11091, B2 => n11109, ZN => n5560);
   U13407 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1863_port, A2 
                           => n8491, B1 => n11091, B2 => n11110, ZN => n5559);
   U13408 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1864_port, A2 
                           => n11092, B1 => n11091, B2 => n11111, ZN => n5558);
   U13409 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1865_port, A2 
                           => n8491, B1 => n11091, B2 => n11112, ZN => n5557);
   U13410 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1866_port, A2 
                           => n11092, B1 => n11091, B2 => n11113, ZN => n5556);
   U13411 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1867_port, A2 
                           => n8491, B1 => n11091, B2 => n11114, ZN => n5555);
   U13412 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1868_port, A2 
                           => n8491, B1 => n11091, B2 => n11115, ZN => n5554);
   U13413 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1869_port, A2 
                           => n11092, B1 => n11091, B2 => n11116, ZN => n5553);
   U13414 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1870_port, A2 
                           => n8491, B1 => n11091, B2 => n11117, ZN => n5552);
   U13415 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1871_port, A2 
                           => n11092, B1 => n11091, B2 => n11118, ZN => n5551);
   U13416 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1872_port, A2 
                           => n8491, B1 => n11091, B2 => n11119, ZN => n5550);
   U13417 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1873_port, A2 
                           => n8491, B1 => n11091, B2 => n11120, ZN => n5549);
   U13418 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1874_port, A2 
                           => n8491, B1 => n11091, B2 => n11121, ZN => n5548);
   U13419 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1875_port, A2 
                           => n8491, B1 => n11091, B2 => n11122, ZN => n5547);
   U13420 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1876_port, A2 
                           => n11092, B1 => n11091, B2 => n11123, ZN => n5546);
   U13421 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1877_port, A2 
                           => n11092, B1 => n11091, B2 => n11124, ZN => n5545);
   U13422 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1878_port, A2 
                           => n11092, B1 => n11091, B2 => n11125, ZN => n5544);
   U13423 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1879_port, A2 
                           => n8491, B1 => n11091, B2 => n11126, ZN => n5543);
   U13424 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1880_port, A2 
                           => n11092, B1 => n11091, B2 => n11127, ZN => n5542);
   U13425 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1881_port, A2 
                           => n8491, B1 => n11091, B2 => n11128, ZN => n5541);
   U13426 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1882_port, A2 
                           => n11092, B1 => n11091, B2 => n11129, ZN => n5540);
   U13427 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1883_port, A2 
                           => n8491, B1 => n11091, B2 => n11130, ZN => n5539);
   U13428 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1884_port, A2 
                           => n8491, B1 => n11091, B2 => n11131, ZN => n5538);
   U13429 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1885_port, A2 
                           => n8491, B1 => n11091, B2 => n11132, ZN => n5537);
   U13430 : AOI22_X1 port map( A1 => n11185, A2 => n11090, B1 => n8491, B2 => 
                           DataPath_RF_bus_reg_dataout_1886_port, ZN => n5536);
   U13431 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1887_port, A2 
                           => n8491, B1 => n11091, B2 => n11094, ZN => n5533);
   U13432 : OAI22_X1 port map( A1 => n576, A2 => n11517, B1 => n11518, B2 => 
                           n11153, ZN => n11093);
   U13433 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1824_port, A2 
                           => n8492, B1 => n11095, B2 => n11103, ZN => n5531);
   U13434 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1825_port, A2 
                           => n8492, B1 => n11095, B2 => n11104, ZN => n5530);
   U13435 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1826_port, A2 
                           => n8492, B1 => n11095, B2 => n11105, ZN => n5529);
   U13436 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1827_port, A2 
                           => n11096, B1 => n11095, B2 => n11106, ZN => n5528);
   U13437 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1828_port, A2 
                           => n11096, B1 => n11095, B2 => n11107, ZN => n5527);
   U13438 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1829_port, A2 
                           => n11096, B1 => n11095, B2 => n11108, ZN => n5526);
   U13439 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1830_port, A2 
                           => n8492, B1 => n11095, B2 => n11109, ZN => n5525);
   U13440 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1831_port, A2 
                           => n8492, B1 => n11095, B2 => n11110, ZN => n5524);
   U13441 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1832_port, A2 
                           => n11096, B1 => n11095, B2 => n11111, ZN => n5523);
   U13442 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1833_port, A2 
                           => n8492, B1 => n11095, B2 => n11112, ZN => n5522);
   U13443 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1834_port, A2 
                           => n8492, B1 => n11095, B2 => n11113, ZN => n5521);
   U13444 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1835_port, A2 
                           => n8492, B1 => n11095, B2 => n11114, ZN => n5520);
   U13445 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1836_port, A2 
                           => n11096, B1 => n11095, B2 => n11115, ZN => n5519);
   U13446 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1837_port, A2 
                           => n11096, B1 => n11095, B2 => n11116, ZN => n5518);
   U13447 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1838_port, A2 
                           => n8492, B1 => n11095, B2 => n11117, ZN => n5517);
   U13448 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1839_port, A2 
                           => n8492, B1 => n11095, B2 => n11118, ZN => n5516);
   U13449 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1840_port, A2 
                           => n11096, B1 => n11095, B2 => n11119, ZN => n5515);
   U13450 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1841_port, A2 
                           => n8492, B1 => n11095, B2 => n11120, ZN => n5514);
   U13451 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1842_port, A2 
                           => n11096, B1 => n11095, B2 => n11121, ZN => n5513);
   U13452 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1843_port, A2 
                           => n8492, B1 => n11095, B2 => n11122, ZN => n5512);
   U13453 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1844_port, A2 
                           => n8492, B1 => n11095, B2 => n11123, ZN => n5511);
   U13454 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1845_port, A2 
                           => n8492, B1 => n11095, B2 => n11124, ZN => n5510);
   U13455 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1846_port, A2 
                           => n8492, B1 => n11095, B2 => n11125, ZN => n5509);
   U13456 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1847_port, A2 
                           => n11096, B1 => n11095, B2 => n11126, ZN => n5508);
   U13457 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1848_port, A2 
                           => n8492, B1 => n11095, B2 => n11127, ZN => n5507);
   U13458 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1849_port, A2 
                           => n8492, B1 => n11095, B2 => n11128, ZN => n5506);
   U13459 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1850_port, A2 
                           => n11096, B1 => n11095, B2 => n11129, ZN => n5505);
   U13460 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1851_port, A2 
                           => n8492, B1 => n11095, B2 => n11130, ZN => n5504);
   U13461 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1852_port, A2 
                           => n8492, B1 => n11095, B2 => n11131, ZN => n5503);
   U13462 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1853_port, A2 
                           => n8492, B1 => n11095, B2 => n11132, ZN => n5502);
   U13463 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1854_port, A2 
                           => n8492, B1 => n11095, B2 => n11133, ZN => n5501);
   U13464 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1855_port, A2 
                           => n8492, B1 => n11095, B2 => n11094, ZN => n5498);
   U13465 : AOI22_X1 port map( A1 => n11155, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1792_port, ZN => n5496);
   U13466 : AOI22_X1 port map( A1 => n11156, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1793_port, ZN => n5495);
   U13467 : AOI22_X1 port map( A1 => n11157, A2 => n11098, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1794_port, ZN => n5494);
   U13468 : AOI22_X1 port map( A1 => n11158, A2 => n8493, B1 => n11097, B2 => 
                           DataPath_RF_bus_reg_dataout_1795_port, ZN => n5493);
   U13469 : AOI22_X1 port map( A1 => n11159, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1796_port, ZN => n5492);
   U13470 : AOI22_X1 port map( A1 => n11160, A2 => n8493, B1 => n11097, B2 => 
                           DataPath_RF_bus_reg_dataout_1797_port, ZN => n5491);
   U13471 : AOI22_X1 port map( A1 => n11161, A2 => n11098, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1798_port, ZN => n5490);
   U13472 : AOI22_X1 port map( A1 => n11162, A2 => n8493, B1 => n11097, B2 => 
                           DataPath_RF_bus_reg_dataout_1799_port, ZN => n5489);
   U13473 : AOI22_X1 port map( A1 => n11163, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1800_port, ZN => n5488);
   U13474 : AOI22_X1 port map( A1 => n11164, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1801_port, ZN => n5487);
   U13475 : AOI22_X1 port map( A1 => n11165, A2 => n11098, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1802_port, ZN => n5486);
   U13476 : AOI22_X1 port map( A1 => n11166, A2 => n11098, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1803_port, ZN => n5485);
   U13477 : AOI22_X1 port map( A1 => n11167, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1804_port, ZN => n5484);
   U13478 : AOI22_X1 port map( A1 => n11168, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1805_port, ZN => n5483);
   U13479 : AOI22_X1 port map( A1 => n11169, A2 => n8493, B1 => n11097, B2 => 
                           DataPath_RF_bus_reg_dataout_1806_port, ZN => n5482);
   U13480 : AOI22_X1 port map( A1 => n11170, A2 => n11098, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1807_port, ZN => n5481);
   U13481 : AOI22_X1 port map( A1 => n11171, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1808_port, ZN => n5480);
   U13482 : AOI22_X1 port map( A1 => n11172, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1809_port, ZN => n5479);
   U13483 : AOI22_X1 port map( A1 => n11173, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1810_port, ZN => n5478);
   U13484 : AOI22_X1 port map( A1 => n11174, A2 => n11098, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1811_port, ZN => n5477);
   U13485 : AOI22_X1 port map( A1 => n11175, A2 => n11098, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1812_port, ZN => n5476);
   U13486 : AOI22_X1 port map( A1 => n11176, A2 => n8493, B1 => n11097, B2 => 
                           DataPath_RF_bus_reg_dataout_1813_port, ZN => n5475);
   U13487 : AOI22_X1 port map( A1 => n11177, A2 => n8493, B1 => n11097, B2 => 
                           DataPath_RF_bus_reg_dataout_1814_port, ZN => n5474);
   U13488 : AOI22_X1 port map( A1 => n11178, A2 => n8493, B1 => n11097, B2 => 
                           DataPath_RF_bus_reg_dataout_1815_port, ZN => n5473);
   U13489 : AOI22_X1 port map( A1 => n11179, A2 => n11098, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1816_port, ZN => n5472);
   U13490 : AOI22_X1 port map( A1 => n11180, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1817_port, ZN => n5471);
   U13491 : AOI22_X1 port map( A1 => n11181, A2 => n8493, B1 => n11097, B2 => 
                           DataPath_RF_bus_reg_dataout_1818_port, ZN => n5470);
   U13492 : AOI22_X1 port map( A1 => n11182, A2 => n8493, B1 => n11097, B2 => 
                           DataPath_RF_bus_reg_dataout_1819_port, ZN => n5469);
   U13493 : AOI22_X1 port map( A1 => n11183, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1820_port, ZN => n5468);
   U13494 : AOI22_X1 port map( A1 => n11184, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1821_port, ZN => n5467);
   U13495 : AOI22_X1 port map( A1 => n11185, A2 => n8493, B1 => n8494, B2 => 
                           DataPath_RF_bus_reg_dataout_1822_port, ZN => n5466);
   U13496 : AOI22_X1 port map( A1 => n11186, A2 => n8493, B1 => n11097, B2 => 
                           DataPath_RF_bus_reg_dataout_1823_port, ZN => n5463);
   U13497 : OAI22_X1 port map( A1 => n575, A2 => n11543, B1 => n576, B2 => 
                           n11544, ZN => n11099);
   U13498 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1760_port, B1 => n11155,
                           B2 => n11100, ZN => n5461);
   U13499 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1761_port, B1 => n11156,
                           B2 => n11100, ZN => n5460);
   U13500 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1762_port, B1 => n11157,
                           B2 => n11100, ZN => n5459);
   U13501 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1763_port, B1 => n11158,
                           B2 => n11100, ZN => n5458);
   U13502 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1764_port, B1 => n11159,
                           B2 => n11100, ZN => n5457);
   U13503 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1765_port, B1 => n11160,
                           B2 => n11100, ZN => n5456);
   U13504 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1766_port, B1 => n11161,
                           B2 => n11100, ZN => n5455);
   U13505 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1767_port, B1 => n11162,
                           B2 => n11100, ZN => n5454);
   U13506 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1768_port, B1 => n11163,
                           B2 => n11100, ZN => n5453);
   U13507 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1769_port, B1 => n11164,
                           B2 => n11100, ZN => n5452);
   U13508 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1770_port, B1 => n11165,
                           B2 => n11100, ZN => n5451);
   U13509 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1771_port, B1 => n11166,
                           B2 => n11100, ZN => n5450);
   U13510 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1772_port, B1 => n11167,
                           B2 => n11100, ZN => n5449);
   U13511 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1773_port, B1 => n11168,
                           B2 => n11100, ZN => n5448);
   U13512 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1774_port, B1 => n11169,
                           B2 => n11100, ZN => n5447);
   U13513 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1775_port, B1 => n11170,
                           B2 => n11100, ZN => n5446);
   U13514 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1776_port, B1 => n11171,
                           B2 => n11100, ZN => n5445);
   U13515 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1777_port, B1 => n11172,
                           B2 => n11100, ZN => n5444);
   U13516 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1778_port, B1 => n11173,
                           B2 => n11100, ZN => n5443);
   U13517 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1779_port, B1 => n11174,
                           B2 => n11100, ZN => n5442);
   U13518 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1780_port, B1 => n11175,
                           B2 => n11100, ZN => n5441);
   U13519 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1781_port, B1 => n11176,
                           B2 => n11100, ZN => n5440);
   U13520 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1782_port, B1 => n11177,
                           B2 => n11100, ZN => n5439);
   U13521 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1783_port, B1 => n11178,
                           B2 => n11100, ZN => n5438);
   U13522 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1784_port, B1 => n11179,
                           B2 => n11100, ZN => n5437);
   U13523 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1785_port, B1 => n11180,
                           B2 => n11100, ZN => n5436);
   U13524 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1786_port, B1 => n11181,
                           B2 => n11100, ZN => n5435);
   U13525 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1787_port, B1 => n11182,
                           B2 => n11100, ZN => n5434);
   U13526 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1788_port, B1 => n11183,
                           B2 => n11100, ZN => n5433);
   U13527 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1789_port, B1 => n11184,
                           B2 => n11100, ZN => n5432);
   U13528 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1790_port, B1 => n11185,
                           B2 => n11100, ZN => n5431);
   U13529 : AOI22_X1 port map( A1 => n11101, A2 => 
                           DataPath_RF_bus_reg_dataout_1791_port, B1 => n11186,
                           B2 => n11100, ZN => n5428);
   U13530 : OAI222_X1 port map( A1 => n8483, A2 => n11549, B1 => n11102, B2 => 
                           n575, C1 => n11550, C2 => n576, ZN => n11136);
   U13531 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1728_port, A2 
                           => n8495, B1 => n11134, B2 => n11103, ZN => n5426);
   U13532 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1729_port, A2 
                           => n8495, B1 => n11134, B2 => n11104, ZN => n5425);
   U13533 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1730_port, A2 
                           => n11135, B1 => n11134, B2 => n11105, ZN => n5424);
   U13534 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1731_port, A2 
                           => n11135, B1 => n11134, B2 => n11106, ZN => n5423);
   U13535 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1732_port, A2 
                           => n8495, B1 => n11134, B2 => n11107, ZN => n5422);
   U13536 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1733_port, A2 
                           => n8495, B1 => n11134, B2 => n11108, ZN => n5421);
   U13537 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1734_port, A2 
                           => n11135, B1 => n11134, B2 => n11109, ZN => n5420);
   U13538 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1735_port, A2 
                           => n8495, B1 => n11134, B2 => n11110, ZN => n5419);
   U13539 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1736_port, A2 
                           => n11135, B1 => n11134, B2 => n11111, ZN => n5418);
   U13540 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1737_port, A2 
                           => n8495, B1 => n11134, B2 => n11112, ZN => n5417);
   U13541 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1738_port, A2 
                           => n11135, B1 => n11134, B2 => n11113, ZN => n5416);
   U13542 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1739_port, A2 
                           => n11135, B1 => n11134, B2 => n11114, ZN => n5415);
   U13543 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1740_port, A2 
                           => n8495, B1 => n11134, B2 => n11115, ZN => n5414);
   U13544 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1741_port, A2 
                           => n11135, B1 => n11134, B2 => n11116, ZN => n5413);
   U13545 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1742_port, A2 
                           => n8495, B1 => n11134, B2 => n11117, ZN => n5412);
   U13546 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1743_port, A2 
                           => n11135, B1 => n11134, B2 => n11118, ZN => n5411);
   U13547 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1744_port, A2 
                           => n8495, B1 => n11134, B2 => n11119, ZN => n5410);
   U13548 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1745_port, A2 
                           => n8495, B1 => n11134, B2 => n11120, ZN => n5409);
   U13549 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1746_port, A2 
                           => n8495, B1 => n11134, B2 => n11121, ZN => n5408);
   U13550 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1747_port, A2 
                           => n8495, B1 => n11134, B2 => n11122, ZN => n5407);
   U13551 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1748_port, A2 
                           => n8495, B1 => n11134, B2 => n11123, ZN => n5406);
   U13552 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1749_port, A2 
                           => n11135, B1 => n11134, B2 => n11124, ZN => n5405);
   U13553 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1750_port, A2 
                           => n8495, B1 => n11134, B2 => n11125, ZN => n5404);
   U13554 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1751_port, A2 
                           => n8495, B1 => n11134, B2 => n11126, ZN => n5403);
   U13555 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1752_port, A2 
                           => n8495, B1 => n11134, B2 => n11127, ZN => n5402);
   U13556 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1753_port, A2 
                           => n8495, B1 => n11134, B2 => n11128, ZN => n5401);
   U13557 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1754_port, A2 
                           => n11135, B1 => n11134, B2 => n11129, ZN => n5400);
   U13558 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1755_port, A2 
                           => n8495, B1 => n11134, B2 => n11130, ZN => n5399);
   U13559 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1756_port, A2 
                           => n8495, B1 => n11134, B2 => n11131, ZN => n5398);
   U13560 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1757_port, A2 
                           => n8495, B1 => n11134, B2 => n11132, ZN => n5397);
   U13561 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1758_port, A2 
                           => n8495, B1 => n11134, B2 => n11133, ZN => n5396);
   U13562 : AOI22_X1 port map( A1 => n11186, A2 => n11136, B1 => n8495, B2 => 
                           DataPath_RF_bus_reg_dataout_1759_port, ZN => n5393);
   U13563 : OAI22_X1 port map( A1 => n575, A2 => n11556, B1 => n11555, B2 => 
                           n8483, ZN => n11138);
   U13564 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1696_port, B1 => n11155,
                           B2 => n8410, ZN => n5391);
   U13565 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1697_port, B1 => n11156,
                           B2 => n8410, ZN => n5390);
   U13566 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1698_port, B1 => n11157,
                           B2 => n8410, ZN => n5389);
   U13567 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1699_port, B1 => n11158,
                           B2 => n8410, ZN => n5388);
   U13568 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1700_port, B1 => n11159,
                           B2 => n8410, ZN => n5387);
   U13569 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1701_port, B1 => n11160,
                           B2 => n8410, ZN => n5386);
   U13570 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1702_port, B1 => n11161,
                           B2 => n8410, ZN => n5385);
   U13571 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1703_port, B1 => n11162,
                           B2 => n8410, ZN => n5384);
   U13572 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1704_port, B1 => n11163,
                           B2 => n8410, ZN => n5383);
   U13573 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1705_port, B1 => n11164,
                           B2 => n8410, ZN => n5382);
   U13574 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1706_port, B1 => n11165,
                           B2 => n8410, ZN => n5381);
   U13575 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1707_port, B1 => n11166,
                           B2 => n8410, ZN => n5380);
   U13576 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1708_port, B1 => n11167,
                           B2 => n8410, ZN => n5379);
   U13577 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1709_port, B1 => n11168,
                           B2 => n8410, ZN => n5378);
   U13578 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1710_port, B1 => n11169,
                           B2 => n8410, ZN => n5377);
   U13579 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1711_port, B1 => n11170,
                           B2 => n8410, ZN => n5376);
   U13580 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1712_port, B1 => n11171,
                           B2 => n8410, ZN => n5375);
   U13581 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1713_port, B1 => n11172,
                           B2 => n8410, ZN => n5374);
   U13582 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1714_port, B1 => n11173,
                           B2 => n8410, ZN => n5373);
   U13583 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1715_port, B1 => n11174,
                           B2 => n8410, ZN => n5372);
   U13584 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1716_port, B1 => n11175,
                           B2 => n8410, ZN => n5371);
   U13585 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1717_port, B1 => n11176,
                           B2 => n8410, ZN => n5370);
   U13586 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1718_port, B1 => n11177,
                           B2 => n8410, ZN => n5369);
   U13587 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1719_port, B1 => n11178,
                           B2 => n8410, ZN => n5368);
   U13588 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1720_port, B1 => n11179,
                           B2 => n8410, ZN => n5367);
   U13589 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1721_port, B1 => n11180,
                           B2 => n8410, ZN => n5366);
   U13590 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1722_port, B1 => n11181,
                           B2 => n8410, ZN => n5365);
   U13591 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1723_port, B1 => n11182,
                           B2 => n8410, ZN => n5364);
   U13592 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1724_port, B1 => n11183,
                           B2 => n8410, ZN => n5363);
   U13593 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1725_port, B1 => n11184,
                           B2 => n8410, ZN => n5362);
   U13594 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1726_port, B1 => n11185,
                           B2 => n8410, ZN => n5361);
   U13595 : AOI22_X1 port map( A1 => n7759, A2 => 
                           DataPath_RF_bus_reg_dataout_1727_port, B1 => n11186,
                           B2 => n8410, ZN => n5358);
   U13596 : OAI22_X1 port map( A1 => n576, A2 => n11562, B1 => n11561, B2 => 
                           n8483, ZN => n11140);
   U13597 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1664_port, B1 => n11155,
                           B2 => n11141, ZN => n5356);
   U13598 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1665_port, B1 => n11156,
                           B2 => n11141, ZN => n5355);
   U13599 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1666_port, B1 => n11157,
                           B2 => n11141, ZN => n5354);
   U13600 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1667_port, B1 => n11158,
                           B2 => n11141, ZN => n5353);
   U13601 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1668_port, B1 => n11159,
                           B2 => n11141, ZN => n5352);
   U13602 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1669_port, B1 => n11160,
                           B2 => n11141, ZN => n5351);
   U13603 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1670_port, B1 => n11161,
                           B2 => n11141, ZN => n5350);
   U13604 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1671_port, B1 => n11162,
                           B2 => n11141, ZN => n5349);
   U13605 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1672_port, B1 => n11163,
                           B2 => n11141, ZN => n5348);
   U13606 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1673_port, B1 => n11164,
                           B2 => n11141, ZN => n5347);
   U13607 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1674_port, B1 => n11165,
                           B2 => n11141, ZN => n5346);
   U13608 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1675_port, B1 => n11166,
                           B2 => n11141, ZN => n5345);
   U13609 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1676_port, B1 => n11167,
                           B2 => n11141, ZN => n5344);
   U13610 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1677_port, B1 => n11168,
                           B2 => n11141, ZN => n5343);
   U13611 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1678_port, B1 => n11169,
                           B2 => n11141, ZN => n5342);
   U13612 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1679_port, B1 => n11170,
                           B2 => n11141, ZN => n5341);
   U13613 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1680_port, B1 => n11171,
                           B2 => n11141, ZN => n5340);
   U13614 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1681_port, B1 => n11172,
                           B2 => n11141, ZN => n5339);
   U13615 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1682_port, B1 => n11173,
                           B2 => n11141, ZN => n5338);
   U13616 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1683_port, B1 => n11174,
                           B2 => n11141, ZN => n5337);
   U13617 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1684_port, B1 => n11175,
                           B2 => n11141, ZN => n5336);
   U13618 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1685_port, B1 => n11176,
                           B2 => n11141, ZN => n5335);
   U13619 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1686_port, B1 => n11177,
                           B2 => n11141, ZN => n5334);
   U13620 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1687_port, B1 => n11178,
                           B2 => n11141, ZN => n5333);
   U13621 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1688_port, B1 => n11179,
                           B2 => n11141, ZN => n5332);
   U13622 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1689_port, B1 => n11180,
                           B2 => n11141, ZN => n5331);
   U13623 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1690_port, B1 => n11181,
                           B2 => n11141, ZN => n5330);
   U13624 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1691_port, B1 => n11182,
                           B2 => n11141, ZN => n5329);
   U13625 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1692_port, B1 => n11183,
                           B2 => n11141, ZN => n5328);
   U13626 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1693_port, B1 => n11184,
                           B2 => n11141, ZN => n5327);
   U13627 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1694_port, B1 => n11185,
                           B2 => n11141, ZN => n5326);
   U13628 : AOI22_X1 port map( A1 => n11142, A2 => 
                           DataPath_RF_bus_reg_dataout_1695_port, B1 => n11186,
                           B2 => n11141, ZN => n5323);
   U13629 : OAI22_X1 port map( A1 => n576, A2 => n11568, B1 => n11569, B2 => 
                           n8483, ZN => n11143);
   U13630 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1632_port, B1 => n11155,
                           B2 => n11144, ZN => n5321);
   U13631 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1633_port, B1 => n11156,
                           B2 => n11144, ZN => n5320);
   U13632 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1634_port, B1 => n11157,
                           B2 => n11144, ZN => n5319);
   U13633 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1635_port, B1 => n11158,
                           B2 => n11144, ZN => n5318);
   U13634 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1636_port, B1 => n11159,
                           B2 => n11144, ZN => n5317);
   U13635 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1637_port, B1 => n11160,
                           B2 => n11144, ZN => n5316);
   U13636 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1638_port, B1 => n11161,
                           B2 => n11144, ZN => n5315);
   U13637 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1639_port, B1 => n11162,
                           B2 => n11144, ZN => n5314);
   U13638 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1640_port, B1 => n11163,
                           B2 => n11144, ZN => n5313);
   U13639 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1641_port, B1 => n11164,
                           B2 => n11144, ZN => n5312);
   U13640 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1642_port, B1 => n11165,
                           B2 => n11144, ZN => n5311);
   U13641 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1643_port, B1 => n11166,
                           B2 => n11144, ZN => n5310);
   U13642 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1644_port, B1 => n11167,
                           B2 => n11144, ZN => n5309);
   U13643 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1645_port, B1 => n11168,
                           B2 => n11144, ZN => n5308);
   U13644 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1646_port, B1 => n11169,
                           B2 => n11144, ZN => n5307);
   U13645 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1647_port, B1 => n11170,
                           B2 => n11144, ZN => n5306);
   U13646 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1648_port, B1 => n11171,
                           B2 => n11144, ZN => n5305);
   U13647 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1649_port, B1 => n11172,
                           B2 => n11144, ZN => n5304);
   U13648 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1650_port, B1 => n11173,
                           B2 => n11144, ZN => n5303);
   U13649 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1651_port, B1 => n11174,
                           B2 => n11144, ZN => n5302);
   U13650 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1652_port, B1 => n11175,
                           B2 => n11144, ZN => n5301);
   U13651 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1653_port, B1 => n11176,
                           B2 => n11144, ZN => n5300);
   U13652 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1654_port, B1 => n11177,
                           B2 => n11144, ZN => n5299);
   U13653 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1655_port, B1 => n11178,
                           B2 => n11144, ZN => n5298);
   U13654 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1656_port, B1 => n11179,
                           B2 => n11144, ZN => n5297);
   U13655 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1657_port, B1 => n11180,
                           B2 => n11144, ZN => n5296);
   U13656 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1658_port, B1 => n11181,
                           B2 => n11144, ZN => n5295);
   U13657 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1659_port, B1 => n11182,
                           B2 => n11144, ZN => n5294);
   U13658 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1660_port, B1 => n11183,
                           B2 => n11144, ZN => n5293);
   U13659 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1661_port, B1 => n11184,
                           B2 => n11144, ZN => n5292);
   U13660 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1662_port, B1 => n11185,
                           B2 => n11144, ZN => n5291);
   U13661 : AOI22_X1 port map( A1 => n11145, A2 => 
                           DataPath_RF_bus_reg_dataout_1663_port, B1 => n11186,
                           B2 => n11144, ZN => n5288);
   U13662 : OAI22_X1 port map( A1 => n575, A2 => n11572, B1 => n576, B2 => 
                           n11573, ZN => n11146);
   U13663 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1600_port, B1 => n11155,
                           B2 => n11147, ZN => n5286);
   U13664 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1601_port, B1 => n11156,
                           B2 => n11147, ZN => n5285);
   U13665 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1602_port, B1 => n11157,
                           B2 => n11147, ZN => n5284);
   U13666 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1603_port, B1 => n11158,
                           B2 => n11147, ZN => n5283);
   U13667 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1604_port, B1 => n11159,
                           B2 => n11147, ZN => n5282);
   U13668 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1605_port, B1 => n11160,
                           B2 => n11147, ZN => n5281);
   U13669 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1606_port, B1 => n11161,
                           B2 => n11147, ZN => n5280);
   U13670 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1607_port, B1 => n11162,
                           B2 => n11147, ZN => n5279);
   U13671 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1608_port, B1 => n11163,
                           B2 => n11147, ZN => n5278);
   U13672 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1609_port, B1 => n11164,
                           B2 => n11147, ZN => n5277);
   U13673 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1610_port, B1 => n11165,
                           B2 => n11147, ZN => n5276);
   U13674 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1611_port, B1 => n11166,
                           B2 => n11147, ZN => n5275);
   U13675 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1612_port, B1 => n11167,
                           B2 => n11147, ZN => n5274);
   U13676 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1613_port, B1 => n11168,
                           B2 => n11147, ZN => n5273);
   U13677 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1614_port, B1 => n11169,
                           B2 => n11147, ZN => n5272);
   U13678 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1615_port, B1 => n11170,
                           B2 => n11147, ZN => n5271);
   U13679 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1616_port, B1 => n11171,
                           B2 => n11147, ZN => n5270);
   U13680 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1617_port, B1 => n11172,
                           B2 => n11147, ZN => n5269);
   U13681 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1618_port, B1 => n11173,
                           B2 => n11147, ZN => n5268);
   U13682 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1619_port, B1 => n11174,
                           B2 => n11147, ZN => n5267);
   U13683 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1620_port, B1 => n11175,
                           B2 => n11147, ZN => n5266);
   U13684 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1621_port, B1 => n11176,
                           B2 => n11147, ZN => n5265);
   U13685 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1622_port, B1 => n11177,
                           B2 => n11147, ZN => n5264);
   U13686 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1623_port, B1 => n11178,
                           B2 => n11147, ZN => n5263);
   U13687 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1624_port, B1 => n11179,
                           B2 => n11147, ZN => n5262);
   U13688 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1625_port, B1 => n11180,
                           B2 => n11147, ZN => n5261);
   U13689 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1626_port, B1 => n11181,
                           B2 => n11147, ZN => n5260);
   U13690 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1627_port, B1 => n11182,
                           B2 => n11147, ZN => n5259);
   U13691 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1628_port, B1 => n11183,
                           B2 => n11147, ZN => n5258);
   U13692 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1629_port, B1 => n11184,
                           B2 => n11147, ZN => n5257);
   U13693 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1630_port, B1 => n11185,
                           B2 => n11147, ZN => n5256);
   U13694 : AOI22_X1 port map( A1 => n11148, A2 => 
                           DataPath_RF_bus_reg_dataout_1631_port, B1 => n11186,
                           B2 => n11147, ZN => n5253);
   U13695 : OAI22_X1 port map( A1 => n575, A2 => n11578, B1 => n576, B2 => 
                           n11579, ZN => n11149);
   U13696 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1568_port, B1 => n11155,
                           B2 => n11151, ZN => n5250);
   U13697 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1569_port, B1 => n11156,
                           B2 => n11151, ZN => n5249);
   U13698 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1570_port, B1 => n11157,
                           B2 => n11151, ZN => n5248);
   U13699 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1571_port, B1 => n11158,
                           B2 => n11151, ZN => n5247);
   U13700 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1572_port, B1 => n11159,
                           B2 => n11151, ZN => n5246);
   U13701 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1573_port, B1 => n11160,
                           B2 => n11151, ZN => n5245);
   U13702 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1574_port, B1 => n11161,
                           B2 => n11151, ZN => n5244);
   U13703 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1575_port, B1 => n11162,
                           B2 => n11151, ZN => n5243);
   U13704 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1576_port, B1 => n11163,
                           B2 => n11151, ZN => n5242);
   U13705 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1577_port, B1 => n11164,
                           B2 => n11151, ZN => n5241);
   U13706 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1578_port, B1 => n11165,
                           B2 => n11151, ZN => n5240);
   U13707 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1579_port, B1 => n11166,
                           B2 => n11151, ZN => n5239);
   U13708 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1580_port, B1 => n11167,
                           B2 => n11151, ZN => n5238);
   U13709 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1581_port, B1 => n11168,
                           B2 => n11151, ZN => n5237);
   U13710 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1582_port, B1 => n11169,
                           B2 => n11151, ZN => n5236);
   U13711 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1583_port, B1 => n11170,
                           B2 => n11151, ZN => n5235);
   U13712 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1584_port, B1 => n11171,
                           B2 => n11151, ZN => n5234);
   U13713 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1585_port, B1 => n11172,
                           B2 => n11151, ZN => n5233);
   U13714 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1586_port, B1 => n11173,
                           B2 => n11151, ZN => n5232);
   U13715 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1587_port, B1 => n11174,
                           B2 => n11151, ZN => n5231);
   U13716 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1588_port, B1 => n11175,
                           B2 => n11151, ZN => n5230);
   U13717 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1589_port, B1 => n11176,
                           B2 => n11151, ZN => n5229);
   U13718 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1590_port, B1 => n11177,
                           B2 => n11151, ZN => n5228);
   U13719 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1591_port, B1 => n11178,
                           B2 => n11151, ZN => n5227);
   U13720 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1592_port, B1 => n11179,
                           B2 => n11151, ZN => n5226);
   U13721 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1593_port, B1 => n11180,
                           B2 => n11151, ZN => n5225);
   U13722 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1594_port, B1 => n11181,
                           B2 => n11151, ZN => n5224);
   U13723 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1595_port, B1 => n11182,
                           B2 => n11151, ZN => n5223);
   U13724 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1596_port, B1 => n11183,
                           B2 => n11151, ZN => n5222);
   U13725 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1597_port, B1 => n11184,
                           B2 => n11151, ZN => n5221);
   U13726 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1598_port, B1 => n11185,
                           B2 => n11151, ZN => n5220);
   U13727 : AOI22_X1 port map( A1 => n11152, A2 => 
                           DataPath_RF_bus_reg_dataout_1599_port, B1 => n11186,
                           B2 => n11151, ZN => n5217);
   U13728 : OAI22_X1 port map( A1 => n575, A2 => n11583, B1 => n11585, B2 => 
                           n8483, ZN => n11154);
   U13729 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1536_port, B1 => n11155,
                           B2 => n8411, ZN => n5214);
   U13730 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1537_port, B1 => n11156,
                           B2 => n8411, ZN => n5212);
   U13731 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1538_port, B1 => n11157,
                           B2 => n8411, ZN => n5210);
   U13732 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1539_port, B1 => n11158,
                           B2 => n8411, ZN => n5208);
   U13733 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1540_port, B1 => n11159,
                           B2 => n8411, ZN => n5206);
   U13734 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1541_port, B1 => n11160,
                           B2 => n8411, ZN => n5204);
   U13735 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1542_port, B1 => n11161,
                           B2 => n8411, ZN => n5202);
   U13736 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1543_port, B1 => n11162,
                           B2 => n8411, ZN => n5200);
   U13737 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1544_port, B1 => n11163,
                           B2 => n8411, ZN => n5198);
   U13738 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1545_port, B1 => n11164,
                           B2 => n8411, ZN => n5196);
   U13739 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1546_port, B1 => n11165,
                           B2 => n8411, ZN => n5194);
   U13740 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1547_port, B1 => n11166,
                           B2 => n8411, ZN => n5192);
   U13741 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1548_port, B1 => n11167,
                           B2 => n8411, ZN => n5190);
   U13742 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1549_port, B1 => n11168,
                           B2 => n8411, ZN => n5188);
   U13743 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1550_port, B1 => n11169,
                           B2 => n8411, ZN => n5186);
   U13744 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1551_port, B1 => n11170,
                           B2 => n8411, ZN => n5184);
   U13745 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1552_port, B1 => n11171,
                           B2 => n8411, ZN => n5182);
   U13746 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1553_port, B1 => n11172,
                           B2 => n8411, ZN => n5180);
   U13747 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1554_port, B1 => n11173,
                           B2 => n8411, ZN => n5178);
   U13748 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1555_port, B1 => n11174,
                           B2 => n8411, ZN => n5176);
   U13749 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1556_port, B1 => n11175,
                           B2 => n8411, ZN => n5174);
   U13750 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1557_port, B1 => n11176,
                           B2 => n8411, ZN => n5172);
   U13751 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1558_port, B1 => n11177,
                           B2 => n8411, ZN => n5170);
   U13752 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1559_port, B1 => n11178,
                           B2 => n8411, ZN => n5168);
   U13753 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1560_port, B1 => n11179,
                           B2 => n8411, ZN => n5166);
   U13754 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1561_port, B1 => n11180,
                           B2 => n8411, ZN => n5164);
   U13755 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1562_port, B1 => n11181,
                           B2 => n8411, ZN => n5162);
   U13756 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1563_port, B1 => n11182,
                           B2 => n8411, ZN => n5160);
   U13757 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1564_port, B1 => n11183,
                           B2 => n8411, ZN => n5158);
   U13758 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1565_port, B1 => n11184,
                           B2 => n8411, ZN => n5156);
   U13759 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1566_port, B1 => n11185,
                           B2 => n8411, ZN => n5154);
   U13760 : AOI22_X1 port map( A1 => n7762, A2 => 
                           DataPath_RF_bus_reg_dataout_1567_port, B1 => n11186,
                           B2 => n8411, ZN => n5150);
   U13761 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1504_port, A2 
                           => n8496, B1 => n11190, B2 => n7818, ZN => n5148);
   U13762 : AOI22_X1 port map( A1 => n11190, A2 => n7820, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1505_port, ZN => n5147);
   U13763 : AOI22_X1 port map( A1 => n7783, A2 => n11452, B1 => n11647, B2 => 
                           n11281, ZN => n11248);
   U13764 : AOI22_X1 port map( A1 => n11190, A2 => n11248, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1506_port, ZN => n5146);
   U13765 : AOI22_X1 port map( A1 => n11190, A2 => n7814, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1507_port, ZN => n5145);
   U13766 : AOI22_X1 port map( A1 => n11190, A2 => n7819, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1508_port, ZN => n5144);
   U13767 : OAI22_X1 port map( A1 => n11281, A2 => n11456, B1 => n11455, B2 => 
                           n7783, ZN => n11191);
   U13768 : AOI22_X1 port map( A1 => n11190, A2 => n11250, B1 => n11189, B2 => 
                           DataPath_RF_bus_reg_dataout_1509_port, ZN => n5143);
   U13769 : AOI22_X1 port map( A1 => n11190, A2 => n7813, B1 => n11189, B2 => 
                           DataPath_RF_bus_reg_dataout_1510_port, ZN => n5142);
   U13770 : AOI22_X1 port map( A1 => n7783, A2 => n11458, B1 => n11652, B2 => 
                           n11281, ZN => n11252);
   U13771 : AOI22_X1 port map( A1 => n11190, A2 => n11252, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1511_port, ZN => n5141);
   U13772 : AOI22_X1 port map( A1 => n7783, A2 => n11459, B1 => n11653, B2 => 
                           n11281, ZN => n11253);
   U13773 : AOI22_X1 port map( A1 => n11190, A2 => n11253, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1512_port, ZN => n5140);
   U13774 : OAI22_X1 port map( A1 => n11281, A2 => n11461, B1 => n11460, B2 => 
                           n7783, ZN => n11223);
   U13775 : AOI22_X1 port map( A1 => n11190, A2 => n11254, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1513_port, ZN => n5139);
   U13776 : AOI22_X1 port map( A1 => n7783, A2 => n11462, B1 => n11655, B2 => 
                           n11281, ZN => n11255);
   U13777 : AOI22_X1 port map( A1 => n11190, A2 => n11255, B1 => n11189, B2 => 
                           DataPath_RF_bus_reg_dataout_1514_port, ZN => n5138);
   U13778 : OAI22_X1 port map( A1 => n11281, A2 => n11463, B1 => n11656, B2 => 
                           n7783, ZN => n11256);
   U13779 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1515_port, A2 
                           => n8496, B1 => n11294, B2 => n11188, ZN => n5137);
   U13780 : AOI22_X1 port map( A1 => n11190, A2 => n7812, B1 => n11189, B2 => 
                           DataPath_RF_bus_reg_dataout_1516_port, ZN => n5136);
   U13781 : AOI22_X1 port map( A1 => n11190, A2 => n7815, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1517_port, ZN => n5135);
   U13782 : AOI22_X1 port map( A1 => n11190, A2 => n11297, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1518_port, ZN => n5134);
   U13783 : OAI22_X1 port map( A1 => n11281, A2 => n11468, B1 => n11467, B2 => 
                           n7783, ZN => n11205);
   U13784 : AOI22_X1 port map( A1 => n11190, A2 => n11259, B1 => n11189, B2 => 
                           DataPath_RF_bus_reg_dataout_1519_port, ZN => n5133);
   U13785 : OAI22_X1 port map( A1 => n11281, A2 => n11470, B1 => n11469, B2 => 
                           n7783, ZN => n11206);
   U13786 : AOI22_X1 port map( A1 => n11190, A2 => n11260, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1520_port, ZN => n5132);
   U13787 : OAI22_X1 port map( A1 => n11281, A2 => n11472, B1 => n11471, B2 => 
                           n7783, ZN => n11224);
   U13788 : AOI22_X1 port map( A1 => n11190, A2 => n11261, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1521_port, ZN => n5131);
   U13789 : AOI22_X1 port map( A1 => n11190, A2 => n7811, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1522_port, ZN => n5130);
   U13790 : OAI22_X1 port map( A1 => n11281, A2 => n11475, B1 => n11474, B2 => 
                           n7783, ZN => n11207);
   U13791 : AOI22_X1 port map( A1 => n11190, A2 => n11262, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1523_port, ZN => n5129);
   U13792 : AOI22_X1 port map( A1 => n11190, A2 => n11303, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1524_port, ZN => n5128);
   U13793 : AOI22_X1 port map( A1 => n7783, A2 => n11477, B1 => n11666, B2 => 
                           n11281, ZN => n11230);
   U13794 : AOI22_X1 port map( A1 => n11190, A2 => n11230, B1 => n11189, B2 => 
                           DataPath_RF_bus_reg_dataout_1525_port, ZN => n5127);
   U13795 : AOI22_X1 port map( A1 => n7783, A2 => n11478, B1 => n11667, B2 => 
                           n11281, ZN => n11264);
   U13796 : AOI22_X1 port map( A1 => n11190, A2 => n11264, B1 => n11189, B2 => 
                           DataPath_RF_bus_reg_dataout_1526_port, ZN => n5126);
   U13797 : OAI22_X1 port map( A1 => n11281, A2 => n11480, B1 => n11479, B2 => 
                           n7783, ZN => n11208);
   U13798 : AOI22_X1 port map( A1 => n11190, A2 => n11265, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1527_port, ZN => n5125);
   U13799 : OAI22_X1 port map( A1 => n11281, A2 => n11482, B1 => n11481, B2 => 
                           n7783, ZN => n11192);
   U13800 : INV_X1 port map( A => n11192, ZN => n11266);
   U13801 : AOI22_X1 port map( A1 => n11190, A2 => n11266, B1 => n11189, B2 => 
                           DataPath_RF_bus_reg_dataout_1528_port, ZN => n5124);
   U13802 : OAI22_X1 port map( A1 => n11281, A2 => n11484, B1 => n11483, B2 => 
                           n7783, ZN => n11226);
   U13803 : AOI22_X1 port map( A1 => n11190, A2 => n11277, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1529_port, ZN => n5123);
   U13804 : AOI22_X1 port map( A1 => n7783, A2 => n11485, B1 => n11671, B2 => 
                           n11281, ZN => n11267);
   U13805 : AOI22_X1 port map( A1 => n11190, A2 => n11267, B1 => n11189, B2 => 
                           DataPath_RF_bus_reg_dataout_1530_port, ZN => n5122);
   U13806 : AOI22_X1 port map( A1 => n7783, A2 => n11487, B1 => n11486, B2 => 
                           n11281, ZN => n11199);
   U13807 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1531_port, A2 
                           => n8496, B1 => n11311, B2 => n11188, ZN => n5121);
   U13808 : OAI22_X1 port map( A1 => n11281, A2 => n11489, B1 => n11488, B2 => 
                           n7783, ZN => n11218);
   U13809 : AOI22_X1 port map( A1 => n11190, A2 => n11269, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1532_port, ZN => n5120);
   U13810 : AOI22_X1 port map( A1 => n7783, A2 => n11320, B1 => n11674, B2 => 
                           n11281, ZN => n11270);
   U13811 : AOI22_X1 port map( A1 => n11190, A2 => n11270, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1533_port, ZN => n5119);
   U13812 : OAI22_X1 port map( A1 => n11281, A2 => n11493, B1 => n11492, B2 => 
                           n7783, ZN => n11194);
   U13813 : AOI22_X1 port map( A1 => n11190, A2 => n11271, B1 => n11189, B2 => 
                           DataPath_RF_bus_reg_dataout_1534_port, ZN => n5118);
   U13814 : OAI22_X1 port map( A1 => n11281, A2 => n11495, B1 => n11494, B2 => 
                           n7783, ZN => n11195);
   U13815 : INV_X1 port map( A => n11195, ZN => n11272);
   U13816 : AOI22_X1 port map( A1 => n11190, A2 => n11272, B1 => n8496, B2 => 
                           DataPath_RF_bus_reg_dataout_1535_port, ZN => n5115);
   U13817 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1472_port, A2 
                           => n8497, B1 => n11193, B2 => n7818, ZN => n5113);
   U13818 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1473_port, A2 
                           => n11197, B1 => n11193, B2 => n7820, ZN => n5112);
   U13819 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1474_port, A2 
                           => n11197, B1 => n11193, B2 => n11248, ZN => n5111);
   U13820 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1475_port, A2 
                           => n11197, B1 => n11193, B2 => n7814, ZN => n5110);
   U13821 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1476_port, A2 
                           => n8497, B1 => n11193, B2 => n7819, ZN => n5109);
   U13822 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1477_port, A2 
                           => n8497, B1 => n11288, B2 => n11196, ZN => n5108);
   U13823 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1478_port, A2 
                           => n8497, B1 => n11193, B2 => n7813, ZN => n5107);
   U13824 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1479_port, A2 
                           => n8497, B1 => n11193, B2 => n11252, ZN => n5106);
   U13825 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1480_port, A2 
                           => n8497, B1 => n11193, B2 => n11253, ZN => n5105);
   U13826 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1481_port, A2 
                           => n8497, B1 => n11193, B2 => n11254, ZN => n5104);
   U13827 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1482_port, A2 
                           => n8497, B1 => n11193, B2 => n11255, ZN => n5103);
   U13828 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1483_port, A2 
                           => n11197, B1 => n11193, B2 => n11256, ZN => n5102);
   U13829 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1484_port, A2 
                           => n11197, B1 => n11193, B2 => n7812, ZN => n5101);
   U13830 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1485_port, A2 
                           => n8497, B1 => n11193, B2 => n7815, ZN => n5100);
   U13831 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1486_port, A2 
                           => n8497, B1 => n11193, B2 => n11297, ZN => n5099);
   U13832 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1487_port, A2 
                           => n11197, B1 => n11193, B2 => n11259, ZN => n5098);
   U13833 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1488_port, A2 
                           => n8497, B1 => n11193, B2 => n11260, ZN => n5097);
   U13834 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1489_port, A2 
                           => n8497, B1 => n11193, B2 => n11261, ZN => n5096);
   U13835 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1490_port, A2 
                           => n8497, B1 => n11193, B2 => n7811, ZN => n5095);
   U13836 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1491_port, A2 
                           => n8497, B1 => n11193, B2 => n11262, ZN => n5094);
   U13837 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1492_port, A2 
                           => n8497, B1 => n11193, B2 => n11303, ZN => n5093);
   U13838 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1493_port, A2 
                           => n11197, B1 => n11193, B2 => n11230, ZN => n5092);
   U13839 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1494_port, A2 
                           => n11197, B1 => n11306, B2 => n11196, ZN => n5091);
   U13840 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1495_port, A2 
                           => n8497, B1 => n11193, B2 => n11265, ZN => n5090);
   U13841 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1496_port, A2 
                           => n11197, B1 => n11308, B2 => n11196, ZN => n5089);
   U13842 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1497_port, A2 
                           => n8497, B1 => n11193, B2 => n11277, ZN => n5088);
   U13843 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1498_port, A2 
                           => n8497, B1 => n11193, B2 => n11267, ZN => n5087);
   U13844 : AOI22_X1 port map( A1 => n11311, A2 => n11196, B1 => n8497, B2 => 
                           DataPath_RF_bus_reg_dataout_1499_port, ZN => n5086);
   U13845 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1500_port, A2 
                           => n8497, B1 => n11193, B2 => n11269, ZN => n5085);
   U13846 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1501_port, A2 
                           => n8497, B1 => n11193, B2 => n11270, ZN => n5084);
   U13847 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1502_port, A2 
                           => n11197, B1 => n11314, B2 => n11196, ZN => n5083);
   U13848 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1503_port, A2 
                           => n8497, B1 => n11316, B2 => n11196, ZN => n5080);
   U13849 : OAI22_X1 port map( A1 => n575, A2 => n11897, B1 => n11896, B2 => 
                           n11281, ZN => n11198);
   U13850 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1440_port, A2 
                           => n8498, B1 => n11200, B2 => n7818, ZN => n5078);
   U13851 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1441_port, A2 
                           => n11201, B1 => n11200, B2 => n7820, ZN => n5077);
   U13852 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1442_port, A2 
                           => n11201, B1 => n11200, B2 => n11248, ZN => n5076);
   U13853 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1443_port, A2 
                           => n11201, B1 => n11200, B2 => n7814, ZN => n5075);
   U13854 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1444_port, A2 
                           => n8498, B1 => n11200, B2 => n7819, ZN => n5074);
   U13855 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1445_port, A2 
                           => n8498, B1 => n11200, B2 => n11250, ZN => n5073);
   U13856 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1446_port, A2 
                           => n8498, B1 => n11200, B2 => n7813, ZN => n5072);
   U13857 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1447_port, A2 
                           => n8498, B1 => n11200, B2 => n11252, ZN => n5071);
   U13858 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1448_port, A2 
                           => n8498, B1 => n11200, B2 => n11253, ZN => n5070);
   U13859 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1449_port, A2 
                           => n8498, B1 => n11200, B2 => n11254, ZN => n5069);
   U13860 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1450_port, A2 
                           => n8498, B1 => n11200, B2 => n11255, ZN => n5068);
   U13861 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1451_port, A2 
                           => n11201, B1 => n11200, B2 => n11256, ZN => n5067);
   U13862 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1452_port, A2 
                           => n11201, B1 => n11200, B2 => n7812, ZN => n5066);
   U13863 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1453_port, A2 
                           => n8498, B1 => n11200, B2 => n7815, ZN => n5065);
   U13864 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1454_port, A2 
                           => n8498, B1 => n11200, B2 => n11297, ZN => n5064);
   U13865 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1455_port, A2 
                           => n11201, B1 => n11200, B2 => n11259, ZN => n5063);
   U13866 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1456_port, A2 
                           => n8498, B1 => n11200, B2 => n11260, ZN => n5062);
   U13867 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1457_port, A2 
                           => n8498, B1 => n11200, B2 => n11261, ZN => n5061);
   U13868 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1458_port, A2 
                           => n8498, B1 => n11200, B2 => n7811, ZN => n5060);
   U13869 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1459_port, A2 
                           => n8498, B1 => n11200, B2 => n11262, ZN => n5059);
   U13870 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1460_port, A2 
                           => n8498, B1 => n11200, B2 => n11303, ZN => n5058);
   U13871 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1461_port, A2 
                           => n11201, B1 => n11200, B2 => n11230, ZN => n5057);
   U13872 : AOI22_X1 port map( A1 => n11306, A2 => n11198, B1 => n8498, B2 => 
                           DataPath_RF_bus_reg_dataout_1462_port, ZN => n5056);
   U13873 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1463_port, A2 
                           => n11201, B1 => n11200, B2 => n11265, ZN => n5055);
   U13874 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1464_port, A2 
                           => n8498, B1 => n11200, B2 => n11266, ZN => n5054);
   U13875 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1465_port, A2 
                           => n11201, B1 => n11200, B2 => n11277, ZN => n5053);
   U13876 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1466_port, A2 
                           => n8498, B1 => n11200, B2 => n11267, ZN => n5052);
   U13877 : INV_X1 port map( A => n11199, ZN => n11268);
   U13878 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1467_port, A2 
                           => n8498, B1 => n11200, B2 => n11268, ZN => n5051);
   U13879 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1468_port, A2 
                           => n8498, B1 => n11200, B2 => n11269, ZN => n5050);
   U13880 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1469_port, A2 
                           => n8498, B1 => n11200, B2 => n11270, ZN => n5049);
   U13881 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1470_port, A2 
                           => n11201, B1 => n11200, B2 => n11271, ZN => n5048);
   U13882 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1471_port, A2 
                           => n8498, B1 => n11200, B2 => n11272, ZN => n5045);
   U13883 : OAI22_X1 port map( A1 => n575, A2 => n11908, B1 => n11907, B2 => 
                           n11281, ZN => n11202);
   U13884 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1408_port, A2 
                           => n11204, B1 => n11203, B2 => n7818, ZN => n5043);
   U13885 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1409_port, A2 
                           => n8499, B1 => n11203, B2 => n7820, ZN => n5042);
   U13886 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1410_port, A2 
                           => n8499, B1 => n11203, B2 => n11248, ZN => n5041);
   U13887 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1411_port, A2 
                           => n11204, B1 => n11203, B2 => n7814, ZN => n5040);
   U13888 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1412_port, A2 
                           => n11204, B1 => n11203, B2 => n7819, ZN => n5039);
   U13889 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1413_port, A2 
                           => n11204, B1 => n11203, B2 => n11250, ZN => n5038);
   U13890 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1414_port, A2 
                           => n8499, B1 => n11203, B2 => n7813, ZN => n5037);
   U13891 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1415_port, A2 
                           => n11204, B1 => n11203, B2 => n11252, ZN => n5036);
   U13892 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1416_port, A2 
                           => n8499, B1 => n11203, B2 => n11253, ZN => n5035);
   U13893 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1417_port, A2 
                           => n8499, B1 => n11203, B2 => n11254, ZN => n5034);
   U13894 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1418_port, A2 
                           => n8499, B1 => n11203, B2 => n11255, ZN => n5033);
   U13895 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1419_port, A2 
                           => n8499, B1 => n11203, B2 => n11256, ZN => n5032);
   U13896 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1420_port, A2 
                           => n8499, B1 => n11203, B2 => n7812, ZN => n5031);
   U13897 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1421_port, A2 
                           => n8499, B1 => n11203, B2 => n7815, ZN => n5030);
   U13898 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1422_port, A2 
                           => n8499, B1 => n11203, B2 => n11297, ZN => n5029);
   U13899 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1423_port, A2 
                           => n8499, B1 => n11203, B2 => n11259, ZN => n5028);
   U13900 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1424_port, A2 
                           => n11204, B1 => n11203, B2 => n11260, ZN => n5027);
   U13901 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1425_port, A2 
                           => n8499, B1 => n11203, B2 => n11261, ZN => n5026);
   U13902 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1426_port, A2 
                           => n8499, B1 => n11203, B2 => n7811, ZN => n5025);
   U13903 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1427_port, A2 
                           => n8499, B1 => n11203, B2 => n11262, ZN => n5024);
   U13904 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1428_port, A2 
                           => n8499, B1 => n11203, B2 => n11303, ZN => n5023);
   U13905 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1429_port, A2 
                           => n11204, B1 => n11203, B2 => n11230, ZN => n5022);
   U13906 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1430_port, A2 
                           => n8499, B1 => n11203, B2 => n11264, ZN => n5021);
   U13907 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1431_port, A2 
                           => n11204, B1 => n11203, B2 => n11265, ZN => n5020);
   U13908 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1432_port, A2 
                           => n8499, B1 => n11203, B2 => n11266, ZN => n5019);
   U13909 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1433_port, A2 
                           => n11204, B1 => n11203, B2 => n11277, ZN => n5018);
   U13910 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1434_port, A2 
                           => n8499, B1 => n11203, B2 => n11267, ZN => n5017);
   U13911 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1435_port, A2 
                           => n8499, B1 => n11203, B2 => n11268, ZN => n5016);
   U13912 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1436_port, A2 
                           => n8499, B1 => n11203, B2 => n11269, ZN => n5015);
   U13913 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1437_port, A2 
                           => n8499, B1 => n11203, B2 => n11270, ZN => n5014);
   U13914 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1438_port, A2 
                           => n11204, B1 => n11203, B2 => n11271, ZN => n5013);
   U13915 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1439_port, A2 
                           => n8499, B1 => n11203, B2 => n11272, ZN => n5010);
   U13916 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1376_port, A2 
                           => n11210, B1 => n11209, B2 => n7818, ZN => n5008);
   U13917 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1377_port, A2 
                           => n8500, B1 => n11209, B2 => n7820, ZN => n5007);
   U13918 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1378_port, A2 
                           => n8500, B1 => n11209, B2 => n11248, ZN => n5006);
   U13919 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1379_port, A2 
                           => n8500, B1 => n11209, B2 => n7814, ZN => n5005);
   U13920 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1380_port, A2 
                           => n11210, B1 => n11209, B2 => n7819, ZN => n5004);
   U13921 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1381_port, A2 
                           => n11210, B1 => n11209, B2 => n11250, ZN => n5003);
   U13922 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1382_port, A2 
                           => n8500, B1 => n11209, B2 => n7813, ZN => n5002);
   U13923 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1383_port, A2 
                           => n8500, B1 => n11209, B2 => n11252, ZN => n5001);
   U13924 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1384_port, A2 
                           => n8500, B1 => n11209, B2 => n11253, ZN => n5000);
   U13925 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1385_port, A2 
                           => n8500, B1 => n11209, B2 => n11254, ZN => n4999);
   U13926 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1386_port, A2 
                           => n8500, B1 => n11209, B2 => n11255, ZN => n4998);
   U13927 : AOI22_X1 port map( A1 => n11294, A2 => n11211, B1 => n8500, B2 => 
                           DataPath_RF_bus_reg_dataout_1387_port, ZN => n4997);
   U13928 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1388_port, A2 
                           => n8500, B1 => n11295, B2 => n11211, ZN => n4996);
   U13929 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1389_port, A2 
                           => n8500, B1 => n11209, B2 => n7815, ZN => n4995);
   U13930 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1390_port, A2 
                           => n11210, B1 => n11209, B2 => n11297, ZN => n4994);
   U13931 : NOR2_X1 port map( A1 => RST, A2 => n11205, ZN => n11298);
   U13932 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1391_port, A2 
                           => n8500, B1 => n11298, B2 => n11211, ZN => n4993);
   U13933 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1392_port, A2 
                           => n8500, B1 => n11299, B2 => n11211, ZN => n4992);
   U13934 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1393_port, A2 
                           => n11210, B1 => n11209, B2 => n11261, ZN => n4991);
   U13935 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1394_port, A2 
                           => n11210, B1 => n11209, B2 => n7811, ZN => n4990);
   U13936 : NOR2_X1 port map( A1 => RST, A2 => n11207, ZN => n11302);
   U13937 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1395_port, A2 
                           => n8500, B1 => n11302, B2 => n11211, ZN => n4989);
   U13938 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1396_port, A2 
                           => n8500, B1 => n11209, B2 => n11303, ZN => n4988);
   U13939 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1397_port, A2 
                           => n8500, B1 => n11209, B2 => n11230, ZN => n4987);
   U13940 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1398_port, A2 
                           => n11210, B1 => n11209, B2 => n11264, ZN => n4986);
   U13941 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1399_port, A2 
                           => n8500, B1 => n11307, B2 => n11211, ZN => n4985);
   U13942 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1400_port, A2 
                           => n11210, B1 => n11209, B2 => n11266, ZN => n4984);
   U13943 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1401_port, A2 
                           => n8500, B1 => n11209, B2 => n11277, ZN => n4983);
   U13944 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1402_port, A2 
                           => n11210, B1 => n11310, B2 => n11211, ZN => n4982);
   U13945 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1403_port, A2 
                           => n8500, B1 => n11209, B2 => n11268, ZN => n4981);
   U13946 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1404_port, A2 
                           => n8500, B1 => n11209, B2 => n11269, ZN => n4980);
   U13947 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1405_port, A2 
                           => n8500, B1 => n11313, B2 => n11211, ZN => n4979);
   U13948 : AOI22_X1 port map( A1 => n11314, A2 => n11211, B1 => n11210, B2 => 
                           DataPath_RF_bus_reg_dataout_1406_port, ZN => n4978);
   U13949 : AOI22_X1 port map( A1 => n11316, A2 => n11211, B1 => n8500, B2 => 
                           DataPath_RF_bus_reg_dataout_1407_port, ZN => n4975);
   U13950 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1344_port, A2 
                           => n8501, B1 => n11213, B2 => n7818, ZN => n4973);
   U13951 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1345_port, A2 
                           => n11214, B1 => n11213, B2 => n7820, ZN => n4972);
   U13952 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1346_port, A2 
                           => n8501, B1 => n11213, B2 => n11248, ZN => n4971);
   U13953 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1347_port, A2 
                           => n8501, B1 => n11213, B2 => n7814, ZN => n4970);
   U13954 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1348_port, A2 
                           => n8501, B1 => n11213, B2 => n7819, ZN => n4969);
   U13955 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1349_port, A2 
                           => n11214, B1 => n11213, B2 => n11250, ZN => n4968);
   U13956 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1350_port, A2 
                           => n11214, B1 => n11213, B2 => n7813, ZN => n4967);
   U13957 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1351_port, A2 
                           => n8501, B1 => n11213, B2 => n11252, ZN => n4966);
   U13958 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1352_port, A2 
                           => n8501, B1 => n11213, B2 => n11253, ZN => n4965);
   U13959 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1353_port, A2 
                           => n8501, B1 => n11213, B2 => n11254, ZN => n4964);
   U13960 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1354_port, A2 
                           => n8501, B1 => n11213, B2 => n11255, ZN => n4963);
   U13961 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1355_port, A2 
                           => n8501, B1 => n11213, B2 => n11256, ZN => n4962);
   U13962 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1356_port, A2 
                           => n8501, B1 => n11213, B2 => n7812, ZN => n4961);
   U13963 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1357_port, A2 
                           => n8501, B1 => n11213, B2 => n7815, ZN => n4960);
   U13964 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1358_port, A2 
                           => n8501, B1 => n11213, B2 => n11297, ZN => n4959);
   U13965 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1359_port, A2 
                           => n11214, B1 => n11213, B2 => n11259, ZN => n4958);
   U13966 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1360_port, A2 
                           => n8501, B1 => n11213, B2 => n11260, ZN => n4957);
   U13967 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1361_port, A2 
                           => n8501, B1 => n11213, B2 => n11261, ZN => n4956);
   U13968 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1362_port, A2 
                           => n8501, B1 => n11213, B2 => n7811, ZN => n4955);
   U13969 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1363_port, A2 
                           => n8501, B1 => n11213, B2 => n11262, ZN => n4954);
   U13970 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1364_port, A2 
                           => n11214, B1 => n11213, B2 => n11303, ZN => n4953);
   U13971 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1365_port, A2 
                           => n8501, B1 => n11213, B2 => n11230, ZN => n4952);
   U13972 : AOI22_X1 port map( A1 => n11306, A2 => n11212, B1 => n8501, B2 => 
                           DataPath_RF_bus_reg_dataout_1366_port, ZN => n4951);
   U13973 : AOI22_X1 port map( A1 => n11307, A2 => n11212, B1 => n11214, B2 => 
                           DataPath_RF_bus_reg_dataout_1367_port, ZN => n4950);
   U13974 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1368_port, A2 
                           => n11214, B1 => n11213, B2 => n11266, ZN => n4949);
   U13975 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1369_port, A2 
                           => n11214, B1 => n11213, B2 => n11277, ZN => n4948);
   U13976 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1370_port, A2 
                           => n11214, B1 => n11213, B2 => n11267, ZN => n4947);
   U13977 : AOI22_X1 port map( A1 => n11311, A2 => n11212, B1 => n11214, B2 => 
                           DataPath_RF_bus_reg_dataout_1371_port, ZN => n4946);
   U13978 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1372_port, A2 
                           => n8501, B1 => n11213, B2 => n11269, ZN => n4945);
   U13979 : AOI22_X1 port map( A1 => n11313, A2 => n11212, B1 => n8501, B2 => 
                           DataPath_RF_bus_reg_dataout_1373_port, ZN => n4944);
   U13980 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1374_port, A2 
                           => n8501, B1 => n11213, B2 => n11271, ZN => n4943);
   U13981 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1375_port, A2 
                           => n8501, B1 => n11213, B2 => n11272, ZN => n4940);
   U13982 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1312_port, A2 
                           => n8502, B1 => n11215, B2 => n7818, ZN => n4938);
   U13983 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1313_port, A2 
                           => n11216, B1 => n11215, B2 => n7820, ZN => n4937);
   U13984 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1314_port, A2 
                           => n8502, B1 => n11215, B2 => n11248, ZN => n4936);
   U13985 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1315_port, A2 
                           => n8502, B1 => n11215, B2 => n7814, ZN => n4935);
   U13986 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1316_port, A2 
                           => n8502, B1 => n11215, B2 => n7819, ZN => n4934);
   U13987 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1317_port, A2 
                           => n8502, B1 => n11215, B2 => n11250, ZN => n4933);
   U13988 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1318_port, A2 
                           => n8502, B1 => n11215, B2 => n7813, ZN => n4932);
   U13989 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1319_port, A2 
                           => n8502, B1 => n11215, B2 => n11252, ZN => n4931);
   U13990 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1320_port, A2 
                           => n8502, B1 => n11215, B2 => n11253, ZN => n4930);
   U13991 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1321_port, A2 
                           => n8502, B1 => n11215, B2 => n11254, ZN => n4929);
   U13992 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1322_port, A2 
                           => n8502, B1 => n11215, B2 => n11255, ZN => n4928);
   U13993 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1323_port, A2 
                           => n8502, B1 => n11215, B2 => n11256, ZN => n4927);
   U13994 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1324_port, A2 
                           => n8502, B1 => n11215, B2 => n7812, ZN => n4926);
   U13995 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1325_port, A2 
                           => n11216, B1 => n11296, B2 => n11217, ZN => n4925);
   U13996 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1326_port, A2 
                           => n11216, B1 => n11215, B2 => n11297, ZN => n4924);
   U13997 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1327_port, A2 
                           => n8502, B1 => n11215, B2 => n11259, ZN => n4923);
   U13998 : AOI22_X1 port map( A1 => n11299, A2 => n11217, B1 => n11216, B2 => 
                           DataPath_RF_bus_reg_dataout_1328_port, ZN => n4922);
   U13999 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1329_port, A2 
                           => n8502, B1 => n11215, B2 => n11261, ZN => n4921);
   U14000 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1330_port, A2 
                           => n11216, B1 => n11244, B2 => n11217, ZN => n4920);
   U14001 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1331_port, A2 
                           => n8502, B1 => n11215, B2 => n11262, ZN => n4919);
   U14002 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1332_port, A2 
                           => n11216, B1 => n11215, B2 => n11303, ZN => n4918);
   U14003 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1333_port, A2 
                           => n8502, B1 => n11215, B2 => n11230, ZN => n4917);
   U14004 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1334_port, A2 
                           => n11216, B1 => n11215, B2 => n11264, ZN => n4916);
   U14005 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1335_port, A2 
                           => n11216, B1 => n11215, B2 => n11265, ZN => n4915);
   U14006 : AOI22_X1 port map( A1 => n11308, A2 => n11217, B1 => n8502, B2 => 
                           DataPath_RF_bus_reg_dataout_1336_port, ZN => n4914);
   U14007 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1337_port, A2 
                           => n8502, B1 => n11215, B2 => n11277, ZN => n4913);
   U14008 : AOI22_X1 port map( A1 => n11310, A2 => n11217, B1 => n8502, B2 => 
                           DataPath_RF_bus_reg_dataout_1338_port, ZN => n4912);
   U14009 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1339_port, A2 
                           => n8502, B1 => n11215, B2 => n11268, ZN => n4911);
   U14010 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1340_port, A2 
                           => n8502, B1 => n11215, B2 => n11269, ZN => n4910);
   U14011 : AOI22_X1 port map( A1 => n11313, A2 => n11217, B1 => n8502, B2 => 
                           DataPath_RF_bus_reg_dataout_1341_port, ZN => n4909);
   U14012 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1342_port, A2 
                           => n11216, B1 => n11215, B2 => n11271, ZN => n4908);
   U14013 : AOI22_X1 port map( A1 => n11316, A2 => n11217, B1 => n11216, B2 => 
                           DataPath_RF_bus_reg_dataout_1343_port, ZN => n4905);
   U14014 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1280_port, A2 
                           => n11221, B1 => n11220, B2 => n7818, ZN => n4903);
   U14015 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1281_port, A2 
                           => n8503, B1 => n11220, B2 => n7820, ZN => n4902);
   U14016 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1282_port, A2 
                           => n8503, B1 => n11220, B2 => n11248, ZN => n4901);
   U14017 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1283_port, A2 
                           => n11221, B1 => n11220, B2 => n7814, ZN => n4900);
   U14018 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1284_port, A2 
                           => n11221, B1 => n11220, B2 => n7819, ZN => n4899);
   U14019 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1285_port, A2 
                           => n11221, B1 => n11220, B2 => n11250, ZN => n4898);
   U14020 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1286_port, A2 
                           => n8503, B1 => n11220, B2 => n7813, ZN => n4897);
   U14021 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1287_port, A2 
                           => n11221, B1 => n11290, B2 => n11219, ZN => n4896);
   U14022 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1288_port, A2 
                           => n8503, B1 => n11220, B2 => n11253, ZN => n4895);
   U14023 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1289_port, A2 
                           => n8503, B1 => n11220, B2 => n11254, ZN => n4894);
   U14024 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1290_port, A2 
                           => n8503, B1 => n11293, B2 => n11219, ZN => n4893);
   U14025 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1291_port, A2 
                           => n8503, B1 => n11220, B2 => n11256, ZN => n4892);
   U14026 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1292_port, A2 
                           => n8503, B1 => n11220, B2 => n7812, ZN => n4891);
   U14027 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1293_port, A2 
                           => n11221, B1 => n11220, B2 => n7815, ZN => n4890);
   U14028 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1294_port, A2 
                           => n8503, B1 => n11220, B2 => n11297, ZN => n4889);
   U14029 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1295_port, A2 
                           => n8503, B1 => n11220, B2 => n11259, ZN => n4888);
   U14030 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1296_port, A2 
                           => n11221, B1 => n11220, B2 => n11260, ZN => n4887);
   U14031 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1297_port, A2 
                           => n8503, B1 => n11220, B2 => n11261, ZN => n4886);
   U14032 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1298_port, A2 
                           => n8503, B1 => n11220, B2 => n7811, ZN => n4885);
   U14033 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1299_port, A2 
                           => n8503, B1 => n11220, B2 => n11262, ZN => n4884);
   U14034 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1300_port, A2 
                           => n8503, B1 => n11220, B2 => n11303, ZN => n4883);
   U14035 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1301_port, A2 
                           => n8503, B1 => n11220, B2 => n11230, ZN => n4882);
   U14036 : AOI22_X1 port map( A1 => n11306, A2 => n11219, B1 => n8503, B2 => 
                           DataPath_RF_bus_reg_dataout_1302_port, ZN => n4881);
   U14037 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1303_port, A2 
                           => n8503, B1 => n11220, B2 => n11265, ZN => n4880);
   U14038 : AOI22_X1 port map( A1 => n11308, A2 => n11219, B1 => n11221, B2 => 
                           DataPath_RF_bus_reg_dataout_1304_port, ZN => n4879);
   U14039 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1305_port, A2 
                           => n11221, B1 => n11220, B2 => n11277, ZN => n4878);
   U14040 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1306_port, A2 
                           => n8503, B1 => n11220, B2 => n11267, ZN => n4877);
   U14041 : AOI22_X1 port map( A1 => n11311, A2 => n11219, B1 => n8503, B2 => 
                           DataPath_RF_bus_reg_dataout_1307_port, ZN => n4876);
   U14042 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1308_port, A2 
                           => n11221, B1 => n11312, B2 => n11219, ZN => n4875);
   U14043 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1309_port, A2 
                           => n8503, B1 => n11220, B2 => n11270, ZN => n4874);
   U14044 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1310_port, A2 
                           => n8503, B1 => n11220, B2 => n11271, ZN => n4873);
   U14045 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1311_port, A2 
                           => n8503, B1 => n11220, B2 => n11272, ZN => n4870);
   U14046 : OAI22_X1 port map( A1 => n575, A2 => n11544, B1 => n11543, B2 => 
                           n8333, ZN => n11222);
   U14047 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1248_port, A2 
                           => n11228, B1 => n11225, B2 => n7818, ZN => n4868);
   U14048 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1249_port, A2 
                           => n11228, B1 => n11225, B2 => n7820, ZN => n4867);
   U14049 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1250_port, B1 => n11285,
                           B2 => n11227, ZN => n4866);
   U14050 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1251_port, B1 => n11286,
                           B2 => n11227, ZN => n4865);
   U14051 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1252_port, A2 
                           => n11228, B1 => n11225, B2 => n7819, ZN => n4864);
   U14052 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1253_port, B1 => n11288,
                           B2 => n11227, ZN => n4863);
   U14053 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1254_port, B1 => n11289,
                           B2 => n11227, ZN => n4862);
   U14054 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1255_port, B1 => n11290,
                           B2 => n11227, ZN => n4861);
   U14055 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1256_port, B1 => n11291,
                           B2 => n11227, ZN => n4860);
   U14056 : NOR2_X1 port map( A1 => RST, A2 => n11223, ZN => n11292);
   U14057 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1257_port, B1 => n11292,
                           B2 => n11227, ZN => n4859);
   U14058 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1258_port, B1 => n11293,
                           B2 => n11227, ZN => n4858);
   U14059 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1259_port, B1 => n11294,
                           B2 => n11227, ZN => n4857);
   U14060 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1260_port, B1 => n11295,
                           B2 => n11227, ZN => n4856);
   U14061 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1261_port, A2 
                           => n11228, B1 => n11225, B2 => n7815, ZN => n4855);
   U14062 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1262_port, A2 
                           => n11228, B1 => n11225, B2 => n11297, ZN => n4854);
   U14063 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1263_port, A2 
                           => n11228, B1 => n11225, B2 => n11259, ZN => n4853);
   U14064 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1264_port, B1 => n11299,
                           B2 => n11227, ZN => n4852);
   U14065 : NOR2_X1 port map( A1 => RST, A2 => n11224, ZN => n11300);
   U14066 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1265_port, B1 => n11300,
                           B2 => n11227, ZN => n4851);
   U14067 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1266_port, B1 => n11244,
                           B2 => n11227, ZN => n4850);
   U14068 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1267_port, B1 => n11302,
                           B2 => n11227, ZN => n4849);
   U14069 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1268_port, A2 
                           => n11228, B1 => n11225, B2 => n11303, ZN => n4848);
   U14070 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1269_port, A2 
                           => n11228, B1 => n11225, B2 => n11230, ZN => n4847);
   U14071 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1270_port, B1 => n11306,
                           B2 => n11227, ZN => n4846);
   U14072 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1271_port, B1 => n11307,
                           B2 => n11227, ZN => n4845);
   U14073 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1272_port, B1 => n11308,
                           B2 => n11227, ZN => n4844);
   U14074 : NOR2_X1 port map( A1 => RST, A2 => n11226, ZN => n11309);
   U14075 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1273_port, B1 => n11309,
                           B2 => n11227, ZN => n4843);
   U14076 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1274_port, B1 => n11310,
                           B2 => n11227, ZN => n4842);
   U14077 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1275_port, B1 => n11311,
                           B2 => n11227, ZN => n4841);
   U14078 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1276_port, B1 => n11312,
                           B2 => n11227, ZN => n4840);
   U14079 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1277_port, B1 => n11313,
                           B2 => n11227, ZN => n4839);
   U14080 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1278_port, B1 => n11314,
                           B2 => n11227, ZN => n4838);
   U14081 : AOI22_X1 port map( A1 => n11228, A2 => 
                           DataPath_RF_bus_reg_dataout_1279_port, B1 => n11316,
                           B2 => n11227, ZN => n4835);
   U14082 : OAI22_X1 port map( A1 => n575, A2 => n11550, B1 => n11549, B2 => 
                           n11281, ZN => n11229);
   U14083 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1216_port, A2 
                           => n11233, B1 => n11231, B2 => n7818, ZN => n4833);
   U14084 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1217_port, A2 
                           => n11233, B1 => n11231, B2 => n7820, ZN => n4832);
   U14085 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1218_port, B1 => n11285,
                           B2 => n11232, ZN => n4831);
   U14086 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1219_port, B1 => n11286,
                           B2 => n11232, ZN => n4830);
   U14087 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1220_port, A2 
                           => n11233, B1 => n11231, B2 => n7819, ZN => n4829);
   U14088 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1221_port, B1 => n11288,
                           B2 => n11232, ZN => n4828);
   U14089 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1222_port, B1 => n11289,
                           B2 => n11232, ZN => n4827);
   U14090 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1223_port, A2 
                           => n11233, B1 => n11231, B2 => n11252, ZN => n4826);
   U14091 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1224_port, B1 => n11291,
                           B2 => n11232, ZN => n4825);
   U14092 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1225_port, B1 => n11292,
                           B2 => n11232, ZN => n4824);
   U14093 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1226_port, B1 => n11293,
                           B2 => n11232, ZN => n4823);
   U14094 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1227_port, B1 => n11294,
                           B2 => n11232, ZN => n4822);
   U14095 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1228_port, B1 => n11295,
                           B2 => n11232, ZN => n4821);
   U14096 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1229_port, B1 => n11296,
                           B2 => n11232, ZN => n4820);
   U14097 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1230_port, A2 
                           => n11233, B1 => n11231, B2 => n11297, ZN => n4819);
   U14098 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1231_port, B1 => n11298,
                           B2 => n11232, ZN => n4818);
   U14099 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1232_port, B1 => n11299,
                           B2 => n11232, ZN => n4817);
   U14100 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1233_port, A2 
                           => n11233, B1 => n11231, B2 => n11261, ZN => n4816);
   U14101 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1234_port, B1 => n11244,
                           B2 => n11232, ZN => n4815);
   U14102 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1235_port, B1 => n11302,
                           B2 => n11232, ZN => n4814);
   U14103 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1236_port, A2 
                           => n11233, B1 => n11231, B2 => n11303, ZN => n4813);
   U14104 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1237_port, B1 => n11305,
                           B2 => n11232, ZN => n4812);
   U14105 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1238_port, B1 => n11306,
                           B2 => n11232, ZN => n4811);
   U14106 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1239_port, A2 
                           => n11233, B1 => n11231, B2 => n11265, ZN => n4810);
   U14107 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1240_port, B1 => n11308,
                           B2 => n11232, ZN => n4809);
   U14108 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1241_port, A2 
                           => n11233, B1 => n11231, B2 => n11277, ZN => n4808);
   U14109 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1242_port, A2 
                           => n11233, B1 => n11231, B2 => n11267, ZN => n4807);
   U14110 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1243_port, B1 => n11311,
                           B2 => n11232, ZN => n4806);
   U14111 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1244_port, B1 => n11312,
                           B2 => n11232, ZN => n4805);
   U14112 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1245_port, B1 => n11313,
                           B2 => n11232, ZN => n4804);
   U14113 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1246_port, B1 => n11314,
                           B2 => n11232, ZN => n4803);
   U14114 : AOI22_X1 port map( A1 => n11233, A2 => 
                           DataPath_RF_bus_reg_dataout_1247_port, B1 => n11316,
                           B2 => n11232, ZN => n4800);
   U14115 : OAI22_X1 port map( A1 => n8333, A2 => n11556, B1 => n11281, B2 => 
                           n11555, ZN => n11234);
   U14116 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1184_port, A2 
                           => n11237, B1 => n11235, B2 => n7818, ZN => n4798);
   U14117 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1185_port, A2 
                           => n11237, B1 => n11235, B2 => n7820, ZN => n4797);
   U14118 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1186_port, B1 => n11285,
                           B2 => n11236, ZN => n4796);
   U14119 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1187_port, A2 
                           => n11237, B1 => n11235, B2 => n7814, ZN => n4795);
   U14120 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1188_port, A2 
                           => n11237, B1 => n11235, B2 => n7819, ZN => n4794);
   U14121 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1189_port, B1 => n11288,
                           B2 => n11236, ZN => n4793);
   U14122 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1190_port, B1 => n11289,
                           B2 => n11236, ZN => n4792);
   U14123 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1191_port, B1 => n11290,
                           B2 => n11236, ZN => n4791);
   U14124 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1192_port, B1 => n11291,
                           B2 => n11236, ZN => n4790);
   U14125 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1193_port, B1 => n11292,
                           B2 => n11236, ZN => n4789);
   U14126 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1194_port, B1 => n11293,
                           B2 => n11236, ZN => n4788);
   U14127 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1195_port, B1 => n11294,
                           B2 => n11236, ZN => n4787);
   U14128 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1196_port, B1 => n11295,
                           B2 => n11236, ZN => n4786);
   U14129 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1197_port, A2 
                           => n11237, B1 => n11235, B2 => n7815, ZN => n4785);
   U14130 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1198_port, A2 
                           => n11237, B1 => n11235, B2 => n11297, ZN => n4784);
   U14131 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1199_port, A2 
                           => n11237, B1 => n11235, B2 => n11259, ZN => n4783);
   U14132 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1200_port, B1 => n11299,
                           B2 => n11236, ZN => n4782);
   U14133 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1201_port, B1 => n11300,
                           B2 => n11236, ZN => n4781);
   U14134 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1202_port, B1 => n11244,
                           B2 => n11236, ZN => n4780);
   U14135 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1203_port, B1 => n11302,
                           B2 => n11236, ZN => n4779);
   U14136 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1204_port, A2 
                           => n11237, B1 => n11235, B2 => n11303, ZN => n4778);
   U14137 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1205_port, B1 => n11305,
                           B2 => n11236, ZN => n4777);
   U14138 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1206_port, B1 => n11306,
                           B2 => n11236, ZN => n4776);
   U14139 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1207_port, B1 => n11307,
                           B2 => n11236, ZN => n4775);
   U14140 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1208_port, B1 => n11308,
                           B2 => n11236, ZN => n4774);
   U14141 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1209_port, B1 => n11309,
                           B2 => n11236, ZN => n4773);
   U14142 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1210_port, B1 => n11310,
                           B2 => n11236, ZN => n4772);
   U14143 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1211_port, B1 => n11311,
                           B2 => n11236, ZN => n4771);
   U14144 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1212_port, B1 => n11312,
                           B2 => n11236, ZN => n4770);
   U14145 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1213_port, B1 => n11313,
                           B2 => n11236, ZN => n4769);
   U14146 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1214_port, B1 => n11314,
                           B2 => n11236, ZN => n4768);
   U14147 : AOI22_X1 port map( A1 => n11237, A2 => 
                           DataPath_RF_bus_reg_dataout_1215_port, B1 => n11316,
                           B2 => n11236, ZN => n4765);
   U14148 : OAI22_X1 port map( A1 => n575, A2 => n11562, B1 => n11561, B2 => 
                           n11281, ZN => n11238);
   U14149 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1152_port, A2 
                           => n11241, B1 => n11239, B2 => n7818, ZN => n4763);
   U14150 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1153_port, A2 
                           => n11241, B1 => n11239, B2 => n7820, ZN => n4762);
   U14151 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1154_port, B1 => n11285,
                           B2 => n11240, ZN => n4761);
   U14152 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1155_port, B1 => n11286,
                           B2 => n11240, ZN => n4760);
   U14153 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1156_port, A2 
                           => n11241, B1 => n11239, B2 => n7819, ZN => n4759);
   U14154 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1157_port, B1 => n11288,
                           B2 => n11240, ZN => n4758);
   U14155 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1158_port, A2 
                           => n11241, B1 => n11239, B2 => n7813, ZN => n4757);
   U14156 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1159_port, B1 => n11290,
                           B2 => n11240, ZN => n4756);
   U14157 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1160_port, B1 => n11291,
                           B2 => n11240, ZN => n4755);
   U14158 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1161_port, B1 => n11292,
                           B2 => n11240, ZN => n4754);
   U14159 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1162_port, B1 => n11293,
                           B2 => n11240, ZN => n4753);
   U14160 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1163_port, B1 => n11294,
                           B2 => n11240, ZN => n4752);
   U14161 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1164_port, A2 
                           => n11241, B1 => n11239, B2 => n7812, ZN => n4751);
   U14162 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1165_port, A2 
                           => n11241, B1 => n11239, B2 => n7815, ZN => n4750);
   U14163 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1166_port, A2 
                           => n11241, B1 => n11239, B2 => n11297, ZN => n4749);
   U14164 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1167_port, B1 => n11298,
                           B2 => n11240, ZN => n4748);
   U14165 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1168_port, B1 => n11299,
                           B2 => n11240, ZN => n4747);
   U14166 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1169_port, B1 => n11300,
                           B2 => n11240, ZN => n4746);
   U14167 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1170_port, B1 => n11244,
                           B2 => n11240, ZN => n4745);
   U14168 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1171_port, A2 
                           => n11241, B1 => n11239, B2 => n11262, ZN => n4744);
   U14169 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1172_port, A2 
                           => n11241, B1 => n11239, B2 => n11303, ZN => n4743);
   U14170 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1173_port, B1 => n11305,
                           B2 => n11240, ZN => n4742);
   U14171 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1174_port, A2 
                           => n11241, B1 => n11239, B2 => n11264, ZN => n4741);
   U14172 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1175_port, B1 => n11307,
                           B2 => n11240, ZN => n4740);
   U14173 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1176_port, B1 => n11308,
                           B2 => n11240, ZN => n4739);
   U14174 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1177_port, B1 => n11309,
                           B2 => n11240, ZN => n4738);
   U14175 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1178_port, B1 => n11310,
                           B2 => n11240, ZN => n4737);
   U14176 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1179_port, B1 => n11311,
                           B2 => n11240, ZN => n4736);
   U14177 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1180_port, B1 => n11312,
                           B2 => n11240, ZN => n4735);
   U14178 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1181_port, A2 
                           => n11241, B1 => n11239, B2 => n11270, ZN => n4734);
   U14179 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1182_port, B1 => n11314,
                           B2 => n11240, ZN => n4733);
   U14180 : AOI22_X1 port map( A1 => n11241, A2 => 
                           DataPath_RF_bus_reg_dataout_1183_port, B1 => n11316,
                           B2 => n11240, ZN => n4730);
   U14181 : OAI22_X1 port map( A1 => n575, A2 => n11568, B1 => n11569, B2 => 
                           n11281, ZN => n11242);
   U14182 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1120_port, A2 
                           => n11247, B1 => n11245, B2 => n7818, ZN => n4728);
   U14183 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1121_port, A2 
                           => n11247, B1 => n11245, B2 => n7820, ZN => n4727);
   U14184 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1122_port, B1 => n11285,
                           B2 => n11246, ZN => n4726);
   U14185 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1123_port, B1 => n11286,
                           B2 => n11246, ZN => n4725);
   U14186 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1124_port, A2 
                           => n11247, B1 => n11245, B2 => n7819, ZN => n4724);
   U14187 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1125_port, B1 => n11288,
                           B2 => n11246, ZN => n4723);
   U14188 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1126_port, B1 => n11289,
                           B2 => n11246, ZN => n4722);
   U14189 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1127_port, B1 => n11290,
                           B2 => n11246, ZN => n4721);
   U14190 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1128_port, B1 => n11291,
                           B2 => n11246, ZN => n4720);
   U14191 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1129_port, B1 => n11292,
                           B2 => n11246, ZN => n4719);
   U14192 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1130_port, B1 => n11293,
                           B2 => n11246, ZN => n4718);
   U14193 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1131_port, A2 
                           => n11247, B1 => n11245, B2 => n11256, ZN => n4717);
   U14194 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1132_port, A2 
                           => n11247, B1 => n11245, B2 => n7812, ZN => n4716);
   U14195 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1133_port, B1 => n11296,
                           B2 => n11246, ZN => n4715);
   U14196 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1134_port, A2 
                           => n11247, B1 => n11245, B2 => n11297, ZN => n4714);
   U14197 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1135_port, B1 => n11298,
                           B2 => n11246, ZN => n4713);
   U14198 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1136_port, B1 => n11299,
                           B2 => n11246, ZN => n4712);
   U14199 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1137_port, B1 => n11300,
                           B2 => n11246, ZN => n4711);
   U14200 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1138_port, B1 => n11244,
                           B2 => n11246, ZN => n4710);
   U14201 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1139_port, A2 
                           => n11247, B1 => n11245, B2 => n11262, ZN => n4709);
   U14202 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1140_port, A2 
                           => n11247, B1 => n11245, B2 => n11303, ZN => n4708);
   U14203 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1141_port, B1 => n11305,
                           B2 => n11246, ZN => n4707);
   U14204 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1142_port, B1 => n11306,
                           B2 => n11246, ZN => n4706);
   U14205 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1143_port, B1 => n11307,
                           B2 => n11246, ZN => n4705);
   U14206 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1144_port, B1 => n11308,
                           B2 => n11246, ZN => n4704);
   U14207 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1145_port, B1 => n11309,
                           B2 => n11246, ZN => n4703);
   U14208 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1146_port, A2 
                           => n11247, B1 => n11245, B2 => n11267, ZN => n4702);
   U14209 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1147_port, A2 
                           => n11247, B1 => n11245, B2 => n11268, ZN => n4701);
   U14210 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1148_port, B1 => n11312,
                           B2 => n11246, ZN => n4700);
   U14211 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1149_port, B1 => n11313,
                           B2 => n11246, ZN => n4699);
   U14212 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1150_port, B1 => n11314,
                           B2 => n11246, ZN => n4698);
   U14213 : AOI22_X1 port map( A1 => n11247, A2 => 
                           DataPath_RF_bus_reg_dataout_1151_port, B1 => n11316,
                           B2 => n11246, ZN => n4695);
   U14214 : OAI222_X1 port map( A1 => n11373, A2 => n11281, B1 => n11573, B2 =>
                           n575, C1 => n11572, C2 => n8333, ZN => n11263);
   U14215 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1088_port, A2 
                           => n8504, B1 => n11273, B2 => n7818, ZN => n4693);
   U14216 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1089_port, A2 
                           => n11274, B1 => n11273, B2 => n7820, ZN => n4692);
   U14217 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1090_port, A2 
                           => n11274, B1 => n11273, B2 => n11248, ZN => n4691);
   U14218 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1091_port, A2 
                           => n11274, B1 => n11273, B2 => n7814, ZN => n4690);
   U14219 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1092_port, A2 
                           => n8504, B1 => n11273, B2 => n7819, ZN => n4689);
   U14220 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1093_port, A2 
                           => n8504, B1 => n11273, B2 => n11250, ZN => n4688);
   U14221 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1094_port, A2 
                           => n8504, B1 => n11273, B2 => n7813, ZN => n4687);
   U14222 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1095_port, A2 
                           => n8504, B1 => n11273, B2 => n11252, ZN => n4686);
   U14223 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1096_port, A2 
                           => n11274, B1 => n11273, B2 => n11253, ZN => n4685);
   U14224 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1097_port, A2 
                           => n8504, B1 => n11273, B2 => n11254, ZN => n4684);
   U14225 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1098_port, A2 
                           => n8504, B1 => n11273, B2 => n11255, ZN => n4683);
   U14226 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1099_port, A2 
                           => n11274, B1 => n11273, B2 => n11256, ZN => n4682);
   U14227 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1100_port, A2 
                           => n11274, B1 => n11273, B2 => n7812, ZN => n4681);
   U14228 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1101_port, A2 
                           => n8504, B1 => n11273, B2 => n7815, ZN => n4680);
   U14229 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1102_port, A2 
                           => n8504, B1 => n11273, B2 => n11297, ZN => n4679);
   U14230 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1103_port, A2 
                           => n11274, B1 => n11273, B2 => n11259, ZN => n4678);
   U14231 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1104_port, A2 
                           => n8504, B1 => n11273, B2 => n11260, ZN => n4677);
   U14232 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1105_port, A2 
                           => n8504, B1 => n11273, B2 => n11261, ZN => n4676);
   U14233 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1106_port, A2 
                           => n8504, B1 => n11273, B2 => n7811, ZN => n4675);
   U14234 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1107_port, A2 
                           => n8504, B1 => n11273, B2 => n11262, ZN => n4674);
   U14235 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1108_port, A2 
                           => n8504, B1 => n11273, B2 => n11303, ZN => n4673);
   U14236 : AOI22_X1 port map( A1 => n11305, A2 => n11263, B1 => n8504, B2 => 
                           DataPath_RF_bus_reg_dataout_1109_port, ZN => n4672);
   U14237 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1110_port, A2 
                           => n8504, B1 => n11273, B2 => n11264, ZN => n4671);
   U14238 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1111_port, A2 
                           => n11274, B1 => n11273, B2 => n11265, ZN => n4670);
   U14239 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1112_port, A2 
                           => n8504, B1 => n11273, B2 => n11266, ZN => n4669);
   U14240 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1113_port, A2 
                           => n11274, B1 => n11273, B2 => n11277, ZN => n4668);
   U14241 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1114_port, A2 
                           => n8504, B1 => n11273, B2 => n11267, ZN => n4667);
   U14242 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1115_port, A2 
                           => n8504, B1 => n11273, B2 => n11268, ZN => n4666);
   U14243 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1116_port, A2 
                           => n8504, B1 => n11273, B2 => n11269, ZN => n4665);
   U14244 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1117_port, A2 
                           => n8504, B1 => n11273, B2 => n11270, ZN => n4664);
   U14245 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1118_port, A2 
                           => n11274, B1 => n11273, B2 => n11271, ZN => n4663);
   U14246 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1119_port, A2 
                           => n8504, B1 => n11273, B2 => n11272, ZN => n4660);
   U14247 : OAI22_X1 port map( A1 => n575, A2 => n11579, B1 => n11578, B2 => 
                           n8333, ZN => n11275);
   U14248 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1056_port, A2 
                           => n11280, B1 => n11278, B2 => n7818, ZN => n4658);
   U14249 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1057_port, A2 
                           => n11280, B1 => n11278, B2 => n7820, ZN => n4657);
   U14250 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1058_port, B1 => n11285,
                           B2 => n11279, ZN => n4656);
   U14251 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1059_port, B1 => n11286,
                           B2 => n11279, ZN => n4655);
   U14252 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1060_port, A2 
                           => n11280, B1 => n11278, B2 => n7819, ZN => n4654);
   U14253 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1061_port, B1 => n11288,
                           B2 => n11279, ZN => n4653);
   U14254 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1062_port, B1 => n11289,
                           B2 => n11279, ZN => n4652);
   U14255 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1063_port, B1 => n11290,
                           B2 => n11279, ZN => n4651);
   U14256 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1064_port, B1 => n11291,
                           B2 => n11279, ZN => n4650);
   U14257 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1065_port, B1 => n11292,
                           B2 => n11279, ZN => n4649);
   U14258 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1066_port, B1 => n11293,
                           B2 => n11279, ZN => n4648);
   U14259 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1067_port, B1 => n11294,
                           B2 => n11279, ZN => n4647);
   U14260 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1068_port, B1 => n11295,
                           B2 => n11279, ZN => n4646);
   U14261 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1069_port, B1 => n11296,
                           B2 => n11279, ZN => n4645);
   U14262 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1070_port, A2 
                           => n11280, B1 => n11278, B2 => n11297, ZN => n4644);
   U14263 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1071_port, B1 => n11298,
                           B2 => n11279, ZN => n4643);
   U14264 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1072_port, B1 => n11299,
                           B2 => n11279, ZN => n4642);
   U14265 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1073_port, B1 => n11300,
                           B2 => n11279, ZN => n4641);
   U14266 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1074_port, A2 
                           => n11280, B1 => n11278, B2 => n7811, ZN => n4640);
   U14267 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1075_port, B1 => n11302,
                           B2 => n11279, ZN => n4639);
   U14268 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1076_port, A2 
                           => n11280, B1 => n11278, B2 => n11303, ZN => n4638);
   U14269 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1077_port, B1 => n11305,
                           B2 => n11279, ZN => n4637);
   U14270 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1078_port, B1 => n11306,
                           B2 => n11279, ZN => n4636);
   U14271 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1079_port, B1 => n11307,
                           B2 => n11279, ZN => n4635);
   U14272 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1080_port, B1 => n11308,
                           B2 => n11279, ZN => n4634);
   U14273 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1081_port, A2 
                           => n11280, B1 => n11278, B2 => n11277, ZN => n4633);
   U14274 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1082_port, B1 => n11310,
                           B2 => n11279, ZN => n4632);
   U14275 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1083_port, B1 => n11311,
                           B2 => n11279, ZN => n4631);
   U14276 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1084_port, B1 => n11312,
                           B2 => n11279, ZN => n4630);
   U14277 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1085_port, B1 => n11313,
                           B2 => n11279, ZN => n4629);
   U14278 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1086_port, B1 => n11314,
                           B2 => n11279, ZN => n4628);
   U14279 : AOI22_X1 port map( A1 => n11280, A2 => 
                           DataPath_RF_bus_reg_dataout_1087_port, B1 => n11316,
                           B2 => n11279, ZN => n4625);
   U14280 : OAI22_X1 port map( A1 => n8333, A2 => n11583, B1 => n11281, B2 => 
                           n11585, ZN => n11282);
   U14281 : NOR2_X1 port map( A1 => RST, A2 => n11317, ZN => n11304);
   U14282 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1024_port, A2 
                           => n11317, B1 => n11304, B2 => n7818, ZN => n4621);
   U14283 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1025_port, A2 
                           => n11317, B1 => n11304, B2 => n7820, ZN => n4619);
   U14284 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1026_port, B1 => n11285,
                           B2 => n11315, ZN => n4617);
   U14285 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1027_port, B1 => n11286,
                           B2 => n11315, ZN => n4615);
   U14286 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1028_port, A2 
                           => n11317, B1 => n11304, B2 => n7819, ZN => n4613);
   U14287 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1029_port, B1 => n11288,
                           B2 => n11315, ZN => n4611);
   U14288 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1030_port, B1 => n11289,
                           B2 => n11315, ZN => n4609);
   U14289 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1031_port, B1 => n11290,
                           B2 => n11315, ZN => n4607);
   U14290 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1032_port, B1 => n11291,
                           B2 => n11315, ZN => n4605);
   U14291 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1033_port, B1 => n11292,
                           B2 => n11315, ZN => n4603);
   U14292 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1034_port, B1 => n11293,
                           B2 => n11315, ZN => n4601);
   U14293 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1035_port, B1 => n11294,
                           B2 => n11315, ZN => n4599);
   U14294 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1036_port, B1 => n11295,
                           B2 => n11315, ZN => n4597);
   U14295 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1037_port, B1 => n11296,
                           B2 => n11315, ZN => n4595);
   U14296 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1038_port, A2 
                           => n11317, B1 => n11304, B2 => n11297, ZN => n4593);
   U14297 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1039_port, B1 => n11298,
                           B2 => n11315, ZN => n4591);
   U14298 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1040_port, B1 => n11299,
                           B2 => n11315, ZN => n4589);
   U14299 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1041_port, B1 => n11300,
                           B2 => n11315, ZN => n4587);
   U14300 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1042_port, A2 
                           => n11317, B1 => n11304, B2 => n7811, ZN => n4585);
   U14301 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1043_port, B1 => n11302,
                           B2 => n11315, ZN => n4583);
   U14302 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_1044_port, A2 
                           => n11317, B1 => n11304, B2 => n11303, ZN => n4581);
   U14303 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1045_port, B1 => n11305,
                           B2 => n11315, ZN => n4579);
   U14304 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1046_port, B1 => n11306,
                           B2 => n11315, ZN => n4577);
   U14305 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1047_port, B1 => n11307,
                           B2 => n11315, ZN => n4575);
   U14306 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1048_port, B1 => n11308,
                           B2 => n11315, ZN => n4573);
   U14307 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1049_port, B1 => n11309,
                           B2 => n11315, ZN => n4571);
   U14308 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1050_port, B1 => n11310,
                           B2 => n11315, ZN => n4569);
   U14309 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1051_port, B1 => n11311,
                           B2 => n11315, ZN => n4567);
   U14310 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1052_port, B1 => n11312,
                           B2 => n11315, ZN => n4565);
   U14311 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1053_port, B1 => n11313,
                           B2 => n11315, ZN => n4563);
   U14312 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1054_port, B1 => n11314,
                           B2 => n11315, ZN => n4561);
   U14313 : AOI22_X1 port map( A1 => n11317, A2 => 
                           DataPath_RF_bus_reg_dataout_1055_port, B1 => n11316,
                           B2 => n11315, ZN => n4557);
   U14314 : OAI22_X1 port map( A1 => n8333, A2 => n11887, B1 => n11886, B2 => 
                           n11412, ZN => n11318);
   U14315 : AOI22_X1 port map( A1 => n7784, A2 => n11450, B1 => n11645, B2 => 
                           n11412, ZN => n11374);
   U14316 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_992_port, A2 
                           => n8505, B1 => n11322, B2 => n11374, ZN => n4555);
   U14317 : AOI22_X1 port map( A1 => n7784, A2 => n11451, B1 => n11646, B2 => 
                           n11412, ZN => n11375);
   U14318 : AOI22_X1 port map( A1 => n11322, A2 => n11375, B1 => n11321, B2 => 
                           DataPath_RF_bus_reg_dataout_993_port, ZN => n4554);
   U14319 : AOI22_X1 port map( A1 => n7784, A2 => n11452, B1 => n11647, B2 => 
                           n11412, ZN => n11376);
   U14320 : AOI22_X1 port map( A1 => n11322, A2 => n11376, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_994_port, ZN => n4553);
   U14321 : AOI22_X1 port map( A1 => n7784, A2 => n11453, B1 => n11648, B2 => 
                           n11412, ZN => n11377);
   U14322 : AOI22_X1 port map( A1 => n11322, A2 => n11377, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_995_port, ZN => n4552);
   U14323 : AOI22_X1 port map( A1 => n7784, A2 => n11454, B1 => n11649, B2 => 
                           n11412, ZN => n11378);
   U14324 : AOI22_X1 port map( A1 => n11322, A2 => n11378, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_996_port, ZN => n4551);
   U14325 : OAI22_X1 port map( A1 => n11412, A2 => n11456, B1 => n11455, B2 => 
                           n7784, ZN => n11344);
   U14326 : AOI22_X1 port map( A1 => n11322, A2 => n11379, B1 => n11321, B2 => 
                           DataPath_RF_bus_reg_dataout_997_port, ZN => n4550);
   U14327 : AOI22_X1 port map( A1 => n7784, A2 => n11457, B1 => n11651, B2 => 
                           n11412, ZN => n11380);
   U14328 : AOI22_X1 port map( A1 => n11322, A2 => n11380, B1 => n11321, B2 => 
                           DataPath_RF_bus_reg_dataout_998_port, ZN => n4549);
   U14329 : AOI22_X1 port map( A1 => n7784, A2 => n11458, B1 => n11652, B2 => 
                           n11412, ZN => n11381);
   U14330 : AOI22_X1 port map( A1 => n11322, A2 => n11381, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_999_port, ZN => n4548);
   U14331 : AOI22_X1 port map( A1 => n7784, A2 => n11459, B1 => n11653, B2 => 
                           n11412, ZN => n11382);
   U14332 : AOI22_X1 port map( A1 => n11322, A2 => n11382, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1000_port, ZN => n4547);
   U14333 : OAI22_X1 port map( A1 => n11412, A2 => n11461, B1 => n11460, B2 => 
                           n7784, ZN => n11345);
   U14334 : AOI22_X1 port map( A1 => n11322, A2 => n11383, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1001_port, ZN => n4546);
   U14335 : AOI22_X1 port map( A1 => n7784, A2 => n11462, B1 => n11655, B2 => 
                           n11412, ZN => n11384);
   U14336 : AOI22_X1 port map( A1 => n11322, A2 => n11384, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1002_port, ZN => n4545);
   U14337 : AOI22_X1 port map( A1 => n7784, A2 => n11463, B1 => n11656, B2 => 
                           n11412, ZN => n11385);
   U14338 : AOI22_X1 port map( A1 => n11322, A2 => n11385, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1003_port, ZN => n4544);
   U14339 : AOI22_X1 port map( A1 => n7784, A2 => n11464, B1 => n11657, B2 => 
                           n11412, ZN => n11386);
   U14340 : AOI22_X1 port map( A1 => n11322, A2 => n11386, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1004_port, ZN => n4543);
   U14341 : AOI22_X1 port map( A1 => n7784, A2 => n11465, B1 => n11658, B2 => 
                           n11412, ZN => n11387);
   U14342 : AOI22_X1 port map( A1 => n11322, A2 => n11387, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1005_port, ZN => n4542);
   U14343 : AOI22_X1 port map( A1 => n7784, A2 => n11466, B1 => n11659, B2 => 
                           n11412, ZN => n11388);
   U14344 : AOI22_X1 port map( A1 => n11322, A2 => n11388, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1006_port, ZN => n4541);
   U14345 : OAI22_X1 port map( A1 => n11412, A2 => n11468, B1 => n11467, B2 => 
                           n7784, ZN => n11346);
   U14346 : AOI22_X1 port map( A1 => n11322, A2 => n11389, B1 => n11321, B2 => 
                           DataPath_RF_bus_reg_dataout_1007_port, ZN => n4540);
   U14347 : OAI22_X1 port map( A1 => n11412, A2 => n11470, B1 => n11469, B2 => 
                           n7784, ZN => n11347);
   U14348 : AOI22_X1 port map( A1 => n11322, A2 => n11390, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1008_port, ZN => n4539);
   U14349 : OAI22_X1 port map( A1 => n11412, A2 => n11472, B1 => n11471, B2 => 
                           n7784, ZN => n11348);
   U14350 : AOI22_X1 port map( A1 => n11322, A2 => n11391, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1009_port, ZN => n4538);
   U14351 : AOI22_X1 port map( A1 => n7784, A2 => n11473, B1 => n11663, B2 => 
                           n11412, ZN => n11392);
   U14352 : AOI22_X1 port map( A1 => n11322, A2 => n11392, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1010_port, ZN => n4537);
   U14353 : OAI22_X1 port map( A1 => n11412, A2 => n11475, B1 => n11474, B2 => 
                           n7784, ZN => n11349);
   U14354 : AOI22_X1 port map( A1 => n11322, A2 => n11393, B1 => n11321, B2 => 
                           DataPath_RF_bus_reg_dataout_1011_port, ZN => n4536);
   U14355 : AOI22_X1 port map( A1 => n7784, A2 => n11319, B1 => n11665, B2 => 
                           n11412, ZN => n11394);
   U14356 : AOI22_X1 port map( A1 => n11322, A2 => n11394, B1 => n11321, B2 => 
                           DataPath_RF_bus_reg_dataout_1012_port, ZN => n4535);
   U14357 : AOI22_X1 port map( A1 => n7784, A2 => n11477, B1 => n11666, B2 => 
                           n11412, ZN => n11395);
   U14358 : AOI22_X1 port map( A1 => n11322, A2 => n11395, B1 => n11321, B2 => 
                           DataPath_RF_bus_reg_dataout_1013_port, ZN => n4534);
   U14359 : AOI22_X1 port map( A1 => n7784, A2 => n11478, B1 => n11667, B2 => 
                           n11412, ZN => n11396);
   U14360 : AOI22_X1 port map( A1 => n11322, A2 => n11396, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1014_port, ZN => n4533);
   U14361 : OAI22_X1 port map( A1 => n11412, A2 => n11480, B1 => n11479, B2 => 
                           n7784, ZN => n11350);
   U14362 : AOI22_X1 port map( A1 => n11322, A2 => n11397, B1 => n11321, B2 => 
                           DataPath_RF_bus_reg_dataout_1015_port, ZN => n4532);
   U14363 : OAI22_X1 port map( A1 => n11412, A2 => n11482, B1 => n11481, B2 => 
                           n7784, ZN => n11326);
   U14364 : INV_X1 port map( A => n11326, ZN => n11369);
   U14365 : AOI22_X1 port map( A1 => n11322, A2 => n11369, B1 => n11321, B2 => 
                           DataPath_RF_bus_reg_dataout_1016_port, ZN => n4531);
   U14366 : OAI22_X1 port map( A1 => n11412, A2 => n11484, B1 => n11483, B2 => 
                           n7784, ZN => n11327);
   U14367 : AOI22_X1 port map( A1 => n11322, A2 => n11399, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1017_port, ZN => n4530);
   U14368 : AOI22_X1 port map( A1 => n7784, A2 => n11485, B1 => n11671, B2 => 
                           n11412, ZN => n11400);
   U14369 : AOI22_X1 port map( A1 => n11322, A2 => n11400, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1018_port, ZN => n4529);
   U14370 : OAI22_X1 port map( A1 => n11412, A2 => n11487, B1 => n11486, B2 => 
                           n7784, ZN => n11328);
   U14371 : AOI22_X1 port map( A1 => n11322, A2 => n11401, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1019_port, ZN => n4528);
   U14372 : OAI22_X1 port map( A1 => n11412, A2 => n11489, B1 => n11488, B2 => 
                           n7784, ZN => n11329);
   U14373 : AOI22_X1 port map( A1 => n11322, A2 => n11402, B1 => n11321, B2 => 
                           DataPath_RF_bus_reg_dataout_1020_port, ZN => n4527);
   U14374 : AOI22_X1 port map( A1 => n7784, A2 => n11320, B1 => n11674, B2 => 
                           n11412, ZN => n11403);
   U14375 : AOI22_X1 port map( A1 => n11322, A2 => n11403, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1021_port, ZN => n4526);
   U14376 : OAI22_X1 port map( A1 => n11412, A2 => n11493, B1 => n11492, B2 => 
                           n7784, ZN => n11333);
   U14377 : AOI22_X1 port map( A1 => n11322, A2 => n11404, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1022_port, ZN => n4525);
   U14378 : OAI22_X1 port map( A1 => n11412, A2 => n11495, B1 => n11494, B2 => 
                           n7784, ZN => n11351);
   U14379 : AOI22_X1 port map( A1 => n11322, A2 => n11405, B1 => n8505, B2 => 
                           DataPath_RF_bus_reg_dataout_1023_port, ZN => n4522);
   U14380 : OAI22_X1 port map( A1 => n8333, A2 => n11892, B1 => n11412, B2 => 
                           n11891, ZN => n11323);
   U14381 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_960_port, A2 
                           => n11325, B1 => n11324, B2 => n11374, ZN => n4520);
   U14382 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_961_port, A2 
                           => n8506, B1 => n11324, B2 => n11375, ZN => n4519);
   U14383 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_962_port, A2 
                           => n8506, B1 => n11324, B2 => n11376, ZN => n4518);
   U14384 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_963_port, A2 
                           => n11325, B1 => n11324, B2 => n11377, ZN => n4517);
   U14385 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_964_port, A2 
                           => n11325, B1 => n11324, B2 => n11378, ZN => n4516);
   U14386 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_965_port, A2 
                           => n11325, B1 => n11324, B2 => n11379, ZN => n4515);
   U14387 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_966_port, A2 
                           => n8506, B1 => n11324, B2 => n11380, ZN => n4514);
   U14388 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_967_port, A2 
                           => n8506, B1 => n11324, B2 => n11381, ZN => n4513);
   U14389 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_968_port, A2 
                           => n8506, B1 => n11324, B2 => n11382, ZN => n4512);
   U14390 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_969_port, A2 
                           => n8506, B1 => n11324, B2 => n11383, ZN => n4511);
   U14391 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_970_port, A2 
                           => n8506, B1 => n11324, B2 => n11384, ZN => n4510);
   U14392 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_971_port, A2 
                           => n8506, B1 => n11324, B2 => n11385, ZN => n4509);
   U14393 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_972_port, A2 
                           => n8506, B1 => n11324, B2 => n11386, ZN => n4508);
   U14394 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_973_port, A2 
                           => n11325, B1 => n11324, B2 => n11387, ZN => n4507);
   U14395 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_974_port, A2 
                           => n8506, B1 => n11324, B2 => n11388, ZN => n4506);
   U14396 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_975_port, A2 
                           => n8506, B1 => n11324, B2 => n11389, ZN => n4505);
   U14397 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_976_port, A2 
                           => n11325, B1 => n11324, B2 => n11390, ZN => n4504);
   U14398 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_977_port, A2 
                           => n8506, B1 => n11324, B2 => n11391, ZN => n4503);
   U14399 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_978_port, A2 
                           => n11325, B1 => n11324, B2 => n11392, ZN => n4502);
   U14400 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_979_port, A2 
                           => n8506, B1 => n11324, B2 => n11393, ZN => n4501);
   U14401 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_980_port, A2 
                           => n8506, B1 => n11324, B2 => n11394, ZN => n4500);
   U14402 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_981_port, A2 
                           => n8506, B1 => n11324, B2 => n11395, ZN => n4499);
   U14403 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_982_port, A2 
                           => n8506, B1 => n11437, B2 => n11323, ZN => n4498);
   U14404 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_983_port, A2 
                           => n11325, B1 => n11324, B2 => n11397, ZN => n4497);
   U14405 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_984_port, A2 
                           => n8506, B1 => n11324, B2 => n11369, ZN => n4496);
   U14406 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_985_port, A2 
                           => n11325, B1 => n11324, B2 => n11399, ZN => n4495);
   U14407 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_986_port, A2 
                           => n8506, B1 => n11324, B2 => n11400, ZN => n4494);
   U14408 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_987_port, A2 
                           => n8506, B1 => n11324, B2 => n11401, ZN => n4493);
   U14409 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_988_port, A2 
                           => n8506, B1 => n11324, B2 => n11402, ZN => n4492);
   U14410 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_989_port, A2 
                           => n8506, B1 => n11324, B2 => n11403, ZN => n4491);
   U14411 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_990_port, A2 
                           => n11325, B1 => n11324, B2 => n11404, ZN => n4490);
   U14412 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_991_port, A2 
                           => n8506, B1 => n11324, B2 => n11405, ZN => n4487);
   U14413 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_928_port, A2 
                           => n8507, B1 => n11331, B2 => n11374, ZN => n4485);
   U14414 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_929_port, A2 
                           => n8507, B1 => n11331, B2 => n11375, ZN => n4484);
   U14415 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_930_port, A2 
                           => n8507, B1 => n11417, B2 => n11330, ZN => n4483);
   U14416 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_931_port, A2 
                           => n8507, B1 => n11331, B2 => n11377, ZN => n4482);
   U14417 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_932_port, A2 
                           => n8507, B1 => n11331, B2 => n11378, ZN => n4481);
   U14418 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_933_port, A2 
                           => n11332, B1 => n11331, B2 => n11379, ZN => n4480);
   U14419 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_934_port, A2 
                           => n11332, B1 => n11331, B2 => n11380, ZN => n4479);
   U14420 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_935_port, A2 
                           => n8507, B1 => n11331, B2 => n11381, ZN => n4478);
   U14421 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_936_port, A2 
                           => n8507, B1 => n11423, B2 => n11330, ZN => n4477);
   U14422 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_937_port, A2 
                           => n8507, B1 => n11331, B2 => n11383, ZN => n4476);
   U14423 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_938_port, A2 
                           => n11332, B1 => n11331, B2 => n11384, ZN => n4475);
   U14424 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_939_port, A2 
                           => n11332, B1 => n11331, B2 => n11385, ZN => n4474);
   U14425 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_940_port, A2 
                           => n11332, B1 => n11331, B2 => n11386, ZN => n4473);
   U14426 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_941_port, A2 
                           => n8507, B1 => n11331, B2 => n11387, ZN => n4472);
   U14427 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_942_port, A2 
                           => n8507, B1 => n11331, B2 => n11388, ZN => n4471);
   U14428 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_943_port, A2 
                           => n8507, B1 => n11331, B2 => n11389, ZN => n4470);
   U14429 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_944_port, A2 
                           => n11332, B1 => n11331, B2 => n11390, ZN => n4469);
   U14430 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_945_port, A2 
                           => n8507, B1 => n11331, B2 => n11391, ZN => n4468);
   U14431 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_946_port, A2 
                           => n8507, B1 => n11331, B2 => n11392, ZN => n4467);
   U14432 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_947_port, A2 
                           => n8507, B1 => n11331, B2 => n11393, ZN => n4466);
   U14433 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_948_port, A2 
                           => n11332, B1 => n11331, B2 => n11394, ZN => n4465);
   U14434 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_949_port, A2 
                           => n8507, B1 => n11331, B2 => n11395, ZN => n4464);
   U14435 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_950_port, A2 
                           => n8507, B1 => n11331, B2 => n11396, ZN => n4463);
   U14436 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_951_port, A2 
                           => n11332, B1 => n11331, B2 => n11397, ZN => n4462);
   U14437 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_952_port, A2 
                           => n8507, B1 => n11439, B2 => n11330, ZN => n4461);
   U14438 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_953_port, A2 
                           => n11332, B1 => n11440, B2 => n11330, ZN => n4460);
   U14439 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_954_port, A2 
                           => n8507, B1 => n11441, B2 => n11330, ZN => n4459);
   U14440 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_955_port, A2 
                           => n8507, B1 => n11442, B2 => n11330, ZN => n4458);
   U14441 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_956_port, A2 
                           => n8507, B1 => n11443, B2 => n11330, ZN => n4457);
   U14442 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_957_port, A2 
                           => n8507, B1 => n11331, B2 => n11403, ZN => n4456);
   U14443 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_958_port, A2 
                           => n11332, B1 => n11331, B2 => n11404, ZN => n4455);
   U14444 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_959_port, A2 
                           => n8507, B1 => n11331, B2 => n11405, ZN => n4452);
   U14445 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_896_port, A2 
                           => n8508, B1 => n11335, B2 => n11374, ZN => n4450);
   U14446 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_897_port, A2 
                           => n8508, B1 => n11335, B2 => n11375, ZN => n4449);
   U14447 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_898_port, A2 
                           => n8508, B1 => n11335, B2 => n11376, ZN => n4448);
   U14448 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_899_port, A2 
                           => n8508, B1 => n11335, B2 => n11377, ZN => n4447);
   U14449 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_900_port, A2 
                           => n11336, B1 => n11335, B2 => n11378, ZN => n4446);
   U14450 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_901_port, A2 
                           => n8508, B1 => n11335, B2 => n11379, ZN => n4445);
   U14451 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_902_port, A2 
                           => n8508, B1 => n11335, B2 => n11380, ZN => n4444);
   U14452 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_903_port, A2 
                           => n11336, B1 => n11335, B2 => n11381, ZN => n4443);
   U14453 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_904_port, A2 
                           => n11336, B1 => n11335, B2 => n11382, ZN => n4442);
   U14454 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_905_port, A2 
                           => n8508, B1 => n11335, B2 => n11383, ZN => n4441);
   U14455 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_906_port, A2 
                           => n8508, B1 => n11335, B2 => n11384, ZN => n4440);
   U14456 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_907_port, A2 
                           => n11336, B1 => n11335, B2 => n11385, ZN => n4439);
   U14457 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_908_port, A2 
                           => n11336, B1 => n11335, B2 => n11386, ZN => n4438);
   U14458 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_909_port, A2 
                           => n8508, B1 => n11335, B2 => n11387, ZN => n4437);
   U14459 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_910_port, A2 
                           => n8508, B1 => n11335, B2 => n11388, ZN => n4436);
   U14460 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_911_port, A2 
                           => n8508, B1 => n11335, B2 => n11389, ZN => n4435);
   U14461 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_912_port, A2 
                           => n8508, B1 => n11335, B2 => n11390, ZN => n4434);
   U14462 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_913_port, A2 
                           => n11336, B1 => n11335, B2 => n11391, ZN => n4433);
   U14463 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_914_port, A2 
                           => n11336, B1 => n11335, B2 => n11392, ZN => n4432);
   U14464 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_915_port, A2 
                           => n8508, B1 => n11335, B2 => n11393, ZN => n4431);
   U14465 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_916_port, A2 
                           => n11336, B1 => n11335, B2 => n11394, ZN => n4430);
   U14466 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_917_port, A2 
                           => n8508, B1 => n11335, B2 => n11395, ZN => n4429);
   U14467 : AOI22_X1 port map( A1 => n11437, A2 => n11334, B1 => n8508, B2 => 
                           DataPath_RF_bus_reg_dataout_918_port, ZN => n4428);
   U14468 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_919_port, A2 
                           => n11336, B1 => n11335, B2 => n11397, ZN => n4427);
   U14469 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_920_port, A2 
                           => n8508, B1 => n11335, B2 => n11369, ZN => n4426);
   U14470 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_921_port, A2 
                           => n8508, B1 => n11335, B2 => n11399, ZN => n4425);
   U14471 : AOI22_X1 port map( A1 => n11441, A2 => n11334, B1 => n8508, B2 => 
                           DataPath_RF_bus_reg_dataout_922_port, ZN => n4424);
   U14472 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_923_port, A2 
                           => n8508, B1 => n11335, B2 => n11401, ZN => n4423);
   U14473 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_924_port, A2 
                           => n11336, B1 => n11335, B2 => n11402, ZN => n4422);
   U14474 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_925_port, A2 
                           => n8508, B1 => n11444, B2 => n11334, ZN => n4421);
   U14475 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_926_port, A2 
                           => n8508, B1 => n11445, B2 => n11334, ZN => n4420);
   U14476 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_927_port, A2 
                           => n8508, B1 => n11335, B2 => n11405, ZN => n4417);
   U14477 : OAI22_X1 port map( A1 => n8333, A2 => n11924, B1 => n11412, B2 => 
                           n11922, ZN => n11337);
   U14478 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_864_port, A2 
                           => n11339, B1 => n11338, B2 => n11374, ZN => n4415);
   U14479 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_865_port, A2 
                           => n8509, B1 => n11416, B2 => n11337, ZN => n4414);
   U14480 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_866_port, A2 
                           => n8509, B1 => n11338, B2 => n11376, ZN => n4413);
   U14481 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_867_port, A2 
                           => n11339, B1 => n11338, B2 => n11377, ZN => n4412);
   U14482 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_868_port, A2 
                           => n11339, B1 => n11338, B2 => n11378, ZN => n4411);
   U14483 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_869_port, A2 
                           => n11339, B1 => n11338, B2 => n11379, ZN => n4410);
   U14484 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_870_port, A2 
                           => n8509, B1 => n11338, B2 => n11380, ZN => n4409);
   U14485 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_871_port, A2 
                           => n8509, B1 => n11338, B2 => n11381, ZN => n4408);
   U14486 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_872_port, A2 
                           => n8509, B1 => n11338, B2 => n11382, ZN => n4407);
   U14487 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_873_port, A2 
                           => n8509, B1 => n11338, B2 => n11383, ZN => n4406);
   U14488 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_874_port, A2 
                           => n8509, B1 => n11338, B2 => n11384, ZN => n4405);
   U14489 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_875_port, A2 
                           => n8509, B1 => n11338, B2 => n11385, ZN => n4404);
   U14490 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_876_port, A2 
                           => n8509, B1 => n11338, B2 => n11386, ZN => n4403);
   U14491 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_877_port, A2 
                           => n11339, B1 => n11338, B2 => n11387, ZN => n4402);
   U14492 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_878_port, A2 
                           => n8509, B1 => n11338, B2 => n11388, ZN => n4401);
   U14493 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_879_port, A2 
                           => n8509, B1 => n11338, B2 => n11389, ZN => n4400);
   U14494 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_880_port, A2 
                           => n11339, B1 => n11338, B2 => n11390, ZN => n4399);
   U14495 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_881_port, A2 
                           => n8509, B1 => n11338, B2 => n11391, ZN => n4398);
   U14496 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_882_port, A2 
                           => n11339, B1 => n11338, B2 => n11392, ZN => n4397);
   U14497 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_883_port, A2 
                           => n8509, B1 => n11338, B2 => n11393, ZN => n4396);
   U14498 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_884_port, A2 
                           => n8509, B1 => n11338, B2 => n11394, ZN => n4395);
   U14499 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_885_port, A2 
                           => n8509, B1 => n11338, B2 => n11395, ZN => n4394);
   U14500 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_886_port, A2 
                           => n8509, B1 => n11338, B2 => n11396, ZN => n4393);
   U14501 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_887_port, A2 
                           => n11339, B1 => n11338, B2 => n11397, ZN => n4392);
   U14502 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_888_port, A2 
                           => n8509, B1 => n11338, B2 => n11369, ZN => n4391);
   U14503 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_889_port, A2 
                           => n11339, B1 => n11338, B2 => n11399, ZN => n4390);
   U14504 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_890_port, A2 
                           => n8509, B1 => n11338, B2 => n11400, ZN => n4389);
   U14505 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_891_port, A2 
                           => n8509, B1 => n11338, B2 => n11401, ZN => n4388);
   U14506 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_892_port, A2 
                           => n8509, B1 => n11338, B2 => n11402, ZN => n4387);
   U14507 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_893_port, A2 
                           => n8509, B1 => n11338, B2 => n11403, ZN => n4386);
   U14508 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_894_port, A2 
                           => n11339, B1 => n11338, B2 => n11404, ZN => n4385);
   U14509 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_895_port, A2 
                           => n8509, B1 => n11338, B2 => n11405, ZN => n4382);
   U14510 : OAI22_X1 port map( A1 => n11513, A2 => n11412, B1 => n8333, B2 => 
                           n11512, ZN => n11340);
   U14511 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_832_port, A2 
                           => n11342, B1 => n11341, B2 => n11374, ZN => n4380);
   U14512 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_833_port, A2 
                           => n8510, B1 => n11341, B2 => n11375, ZN => n4379);
   U14513 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_834_port, A2 
                           => n8510, B1 => n11341, B2 => n11376, ZN => n4378);
   U14514 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_835_port, A2 
                           => n11342, B1 => n11341, B2 => n11377, ZN => n4377);
   U14515 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_836_port, A2 
                           => n11342, B1 => n11341, B2 => n11378, ZN => n4376);
   U14516 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_837_port, A2 
                           => n11342, B1 => n11341, B2 => n11379, ZN => n4375);
   U14517 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_838_port, A2 
                           => n8510, B1 => n11341, B2 => n11380, ZN => n4374);
   U14518 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_839_port, A2 
                           => n8510, B1 => n11341, B2 => n11381, ZN => n4373);
   U14519 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_840_port, A2 
                           => n8510, B1 => n11341, B2 => n11382, ZN => n4372);
   U14520 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_841_port, A2 
                           => n8510, B1 => n11341, B2 => n11383, ZN => n4371);
   U14521 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_842_port, A2 
                           => n8510, B1 => n11341, B2 => n11384, ZN => n4370);
   U14522 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_843_port, A2 
                           => n8510, B1 => n11341, B2 => n11385, ZN => n4369);
   U14523 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_844_port, A2 
                           => n8510, B1 => n11341, B2 => n11386, ZN => n4368);
   U14524 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_845_port, A2 
                           => n11342, B1 => n11341, B2 => n11387, ZN => n4367);
   U14525 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_846_port, A2 
                           => n8510, B1 => n11341, B2 => n11388, ZN => n4366);
   U14526 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_847_port, A2 
                           => n8510, B1 => n11341, B2 => n11389, ZN => n4365);
   U14527 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_848_port, A2 
                           => n11342, B1 => n11341, B2 => n11390, ZN => n4364);
   U14528 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_849_port, A2 
                           => n8510, B1 => n11341, B2 => n11391, ZN => n4363);
   U14529 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_850_port, A2 
                           => n11342, B1 => n11341, B2 => n11392, ZN => n4362);
   U14530 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_851_port, A2 
                           => n8510, B1 => n11341, B2 => n11393, ZN => n4361);
   U14531 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_852_port, A2 
                           => n8510, B1 => n11341, B2 => n11394, ZN => n4360);
   U14532 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_853_port, A2 
                           => n8510, B1 => n11341, B2 => n11395, ZN => n4359);
   U14533 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_854_port, A2 
                           => n8510, B1 => n11341, B2 => n11396, ZN => n4358);
   U14534 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_855_port, A2 
                           => n11342, B1 => n11341, B2 => n11397, ZN => n4357);
   U14535 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_856_port, A2 
                           => n8510, B1 => n11341, B2 => n11369, ZN => n4356);
   U14536 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_857_port, A2 
                           => n11342, B1 => n11341, B2 => n11399, ZN => n4355);
   U14537 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_858_port, A2 
                           => n8510, B1 => n11341, B2 => n11400, ZN => n4354);
   U14538 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_859_port, A2 
                           => n8510, B1 => n11341, B2 => n11401, ZN => n4353);
   U14539 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_860_port, A2 
                           => n8510, B1 => n11341, B2 => n11402, ZN => n4352);
   U14540 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_861_port, A2 
                           => n8510, B1 => n11341, B2 => n11403, ZN => n4351);
   U14541 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_862_port, A2 
                           => n11342, B1 => n11341, B2 => n11404, ZN => n4350);
   U14542 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_863_port, A2 
                           => n8510, B1 => n11341, B2 => n11405, ZN => n4347);
   U14543 : OAI22_X1 port map( A1 => n11518, A2 => n11412, B1 => n8333, B2 => 
                           n11517, ZN => n11343);
   U14544 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_800_port, B1 => n11415, 
                           B2 => n11352, ZN => n4345);
   U14545 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_801_port, B1 => n11416, 
                           B2 => n11352, ZN => n4344);
   U14546 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_802_port, B1 => n11417, 
                           B2 => n11352, ZN => n4343);
   U14547 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_803_port, B1 => n11418, 
                           B2 => n11352, ZN => n4342);
   U14548 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_804_port, B1 => n11419, 
                           B2 => n11352, ZN => n4341);
   U14549 : NOR2_X1 port map( A1 => RST, A2 => n11344, ZN => n11420);
   U14550 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_805_port, B1 => n11420, 
                           B2 => n11352, ZN => n4340);
   U14551 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_806_port, B1 => n11421, 
                           B2 => n11352, ZN => n4339);
   U14552 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_807_port, B1 => n11422, 
                           B2 => n11352, ZN => n4338);
   U14553 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_808_port, B1 => n11423, 
                           B2 => n11352, ZN => n4337);
   U14554 : NOR2_X1 port map( A1 => RST, A2 => n11345, ZN => n11424);
   U14555 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_809_port, B1 => n11424, 
                           B2 => n11352, ZN => n4336);
   U14556 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_810_port, B1 => n11425, 
                           B2 => n11352, ZN => n4335);
   U14557 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_811_port, B1 => n11426, 
                           B2 => n11352, ZN => n4334);
   U14558 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_812_port, B1 => n11427, 
                           B2 => n11352, ZN => n4333);
   U14559 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_813_port, B1 => n11428, 
                           B2 => n11352, ZN => n4332);
   U14560 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_814_port, B1 => n11429, 
                           B2 => n11352, ZN => n4331);
   U14561 : NOR2_X1 port map( A1 => RST, A2 => n11346, ZN => n11430);
   U14562 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_815_port, B1 => n11430, 
                           B2 => n11352, ZN => n4330);
   U14563 : NOR2_X1 port map( A1 => RST, A2 => n11347, ZN => n11431);
   U14564 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_816_port, B1 => n11431, 
                           B2 => n11352, ZN => n4329);
   U14565 : NOR2_X1 port map( A1 => RST, A2 => n11348, ZN => n11432);
   U14566 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_817_port, B1 => n11432, 
                           B2 => n11352, ZN => n4328);
   U14567 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_818_port, B1 => n11433, 
                           B2 => n11352, ZN => n4327);
   U14568 : NOR2_X1 port map( A1 => RST, A2 => n11349, ZN => n11434);
   U14569 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_819_port, B1 => n11434, 
                           B2 => n11352, ZN => n4326);
   U14570 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_820_port, B1 => n11435, 
                           B2 => n11352, ZN => n4325);
   U14571 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_821_port, B1 => n11436, 
                           B2 => n11352, ZN => n4324);
   U14572 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_822_port, B1 => n11437, 
                           B2 => n11352, ZN => n4323);
   U14573 : NOR2_X1 port map( A1 => RST, A2 => n11350, ZN => n11438);
   U14574 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_823_port, B1 => n11438, 
                           B2 => n11352, ZN => n4322);
   U14575 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_824_port, B1 => n11439, 
                           B2 => n11352, ZN => n4321);
   U14576 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_825_port, B1 => n11440, 
                           B2 => n11352, ZN => n4320);
   U14577 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_826_port, B1 => n11441, 
                           B2 => n11352, ZN => n4319);
   U14578 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_827_port, B1 => n11442, 
                           B2 => n11352, ZN => n4318);
   U14579 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_828_port, B1 => n11443, 
                           B2 => n11352, ZN => n4317);
   U14580 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_829_port, B1 => n11444, 
                           B2 => n11352, ZN => n4316);
   U14581 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_830_port, B1 => n11445, 
                           B2 => n11352, ZN => n4315);
   U14582 : NOR2_X1 port map( A1 => RST, A2 => n11351, ZN => n11447);
   U14583 : AOI22_X1 port map( A1 => n8511, A2 => 
                           DataPath_RF_bus_reg_dataout_831_port, B1 => n11447, 
                           B2 => n11352, ZN => n4312);
   U14584 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_768_port, A2 
                           => n8512, B1 => n11355, B2 => n11374, ZN => n4310);
   U14585 : AOI22_X1 port map( A1 => n11416, A2 => n11354, B1 => n8512, B2 => 
                           DataPath_RF_bus_reg_dataout_769_port, ZN => n4309);
   U14586 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_770_port, A2 
                           => n8512, B1 => n11355, B2 => n11376, ZN => n4308);
   U14587 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_771_port, A2 
                           => n8512, B1 => n11355, B2 => n11377, ZN => n4307);
   U14588 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_772_port, A2 
                           => n11356, B1 => n11355, B2 => n11378, ZN => n4306);
   U14589 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_773_port, A2 
                           => n11356, B1 => n11355, B2 => n11379, ZN => n4305);
   U14590 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_774_port, A2 
                           => n8512, B1 => n11355, B2 => n11380, ZN => n4304);
   U14591 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_775_port, A2 
                           => n8512, B1 => n11355, B2 => n11381, ZN => n4303);
   U14592 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_776_port, A2 
                           => n8512, B1 => n11355, B2 => n11382, ZN => n4302);
   U14593 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_777_port, A2 
                           => n11356, B1 => n11355, B2 => n11383, ZN => n4301);
   U14594 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_778_port, A2 
                           => n11356, B1 => n11355, B2 => n11384, ZN => n4300);
   U14595 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_779_port, A2 
                           => n8512, B1 => n11355, B2 => n11385, ZN => n4299);
   U14596 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_780_port, A2 
                           => n11356, B1 => n11355, B2 => n11386, ZN => n4298);
   U14597 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_781_port, A2 
                           => n8512, B1 => n11355, B2 => n11387, ZN => n4297);
   U14598 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_782_port, A2 
                           => n11356, B1 => n11355, B2 => n11388, ZN => n4296);
   U14599 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_783_port, A2 
                           => n8512, B1 => n11355, B2 => n11389, ZN => n4295);
   U14600 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_784_port, A2 
                           => n8512, B1 => n11355, B2 => n11390, ZN => n4294);
   U14601 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_785_port, A2 
                           => n8512, B1 => n11355, B2 => n11391, ZN => n4293);
   U14602 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_786_port, A2 
                           => n8512, B1 => n11355, B2 => n11392, ZN => n4292);
   U14603 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_787_port, A2 
                           => n8512, B1 => n11355, B2 => n11393, ZN => n4291);
   U14604 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_788_port, A2 
                           => n8512, B1 => n11355, B2 => n11394, ZN => n4290);
   U14605 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_789_port, A2 
                           => n11356, B1 => n11355, B2 => n11395, ZN => n4289);
   U14606 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_790_port, A2 
                           => n11356, B1 => n11355, B2 => n11396, ZN => n4288);
   U14607 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_791_port, A2 
                           => n11356, B1 => n11355, B2 => n11397, ZN => n4287);
   U14608 : AOI22_X1 port map( A1 => n11439, A2 => n11354, B1 => n8512, B2 => 
                           DataPath_RF_bus_reg_dataout_792_port, ZN => n4286);
   U14609 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_793_port, A2 
                           => n8512, B1 => n11355, B2 => n11399, ZN => n4285);
   U14610 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_794_port, A2 
                           => n8512, B1 => n11355, B2 => n11400, ZN => n4284);
   U14611 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_795_port, A2 
                           => n8512, B1 => n11355, B2 => n11401, ZN => n4283);
   U14612 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_796_port, A2 
                           => n11356, B1 => n11355, B2 => n11402, ZN => n4282);
   U14613 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_797_port, A2 
                           => n8512, B1 => n11355, B2 => n11403, ZN => n4281);
   U14614 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_798_port, A2 
                           => n8512, B1 => n11355, B2 => n11404, ZN => n4280);
   U14615 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_799_port, A2 
                           => n8512, B1 => n11355, B2 => n11405, ZN => n4277);
   U14616 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_736_port, B1 => n11415, 
                           B2 => n11358, ZN => n4275);
   U14617 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_737_port, B1 => n11416, 
                           B2 => n11358, ZN => n4274);
   U14618 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_738_port, B1 => n11417, 
                           B2 => n11358, ZN => n4273);
   U14619 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_739_port, B1 => n11418, 
                           B2 => n11358, ZN => n4272);
   U14620 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_740_port, B1 => n11419, 
                           B2 => n11358, ZN => n4271);
   U14621 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_741_port, B1 => n11420, 
                           B2 => n11358, ZN => n4270);
   U14622 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_742_port, B1 => n11421, 
                           B2 => n11358, ZN => n4269);
   U14623 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_743_port, B1 => n11422, 
                           B2 => n11358, ZN => n4268);
   U14624 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_744_port, B1 => n11423, 
                           B2 => n11358, ZN => n4267);
   U14625 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_745_port, B1 => n11424, 
                           B2 => n11358, ZN => n4266);
   U14626 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_746_port, B1 => n11425, 
                           B2 => n11358, ZN => n4265);
   U14627 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_747_port, B1 => n11426, 
                           B2 => n11358, ZN => n4264);
   U14628 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_748_port, B1 => n11427, 
                           B2 => n11358, ZN => n4263);
   U14629 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_749_port, B1 => n11428, 
                           B2 => n11358, ZN => n4262);
   U14630 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_750_port, B1 => n11429, 
                           B2 => n11358, ZN => n4261);
   U14631 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_751_port, B1 => n11430, 
                           B2 => n11358, ZN => n4260);
   U14632 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_752_port, B1 => n11431, 
                           B2 => n11358, ZN => n4259);
   U14633 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_753_port, B1 => n11432, 
                           B2 => n11358, ZN => n4258);
   U14634 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_754_port, B1 => n11433, 
                           B2 => n11358, ZN => n4257);
   U14635 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_755_port, B1 => n11434, 
                           B2 => n11358, ZN => n4256);
   U14636 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_756_port, B1 => n11435, 
                           B2 => n11358, ZN => n4255);
   U14637 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_757_port, B1 => n11436, 
                           B2 => n11358, ZN => n4254);
   U14638 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_758_port, B1 => n11437, 
                           B2 => n11358, ZN => n4253);
   U14639 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_759_port, B1 => n11438, 
                           B2 => n11358, ZN => n4252);
   U14640 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_760_port, B1 => n11439, 
                           B2 => n11358, ZN => n4251);
   U14641 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_761_port, B1 => n11440, 
                           B2 => n11358, ZN => n4250);
   U14642 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_762_port, B1 => n11441, 
                           B2 => n11358, ZN => n4249);
   U14643 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_763_port, B1 => n11442, 
                           B2 => n11358, ZN => n4248);
   U14644 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_764_port, B1 => n11443, 
                           B2 => n11358, ZN => n4247);
   U14645 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_765_port, B1 => n11444, 
                           B2 => n11358, ZN => n4246);
   U14646 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_766_port, B1 => n11445, 
                           B2 => n11358, ZN => n4245);
   U14647 : AOI22_X1 port map( A1 => n11359, A2 => 
                           DataPath_RF_bus_reg_dataout_767_port, B1 => n11447, 
                           B2 => n11358, ZN => n4242);
   U14648 : OAI22_X1 port map( A1 => n8333, A2 => n11550, B1 => n11412, B2 => 
                           n11549, ZN => n11360);
   U14649 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_704_port, B1 => n11415, 
                           B2 => n11361, ZN => n4240);
   U14650 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_705_port, B1 => n11416, 
                           B2 => n11361, ZN => n4239);
   U14651 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_706_port, B1 => n11417, 
                           B2 => n11361, ZN => n4238);
   U14652 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_707_port, B1 => n11418, 
                           B2 => n11361, ZN => n4237);
   U14653 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_708_port, B1 => n11419, 
                           B2 => n11361, ZN => n4236);
   U14654 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_709_port, B1 => n11420, 
                           B2 => n11361, ZN => n4235);
   U14655 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_710_port, B1 => n11421, 
                           B2 => n11361, ZN => n4234);
   U14656 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_711_port, B1 => n11422, 
                           B2 => n11361, ZN => n4233);
   U14657 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_712_port, B1 => n11423, 
                           B2 => n11361, ZN => n4232);
   U14658 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_713_port, B1 => n11424, 
                           B2 => n11361, ZN => n4231);
   U14659 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_714_port, B1 => n11425, 
                           B2 => n11361, ZN => n4230);
   U14660 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_715_port, B1 => n11426, 
                           B2 => n11361, ZN => n4229);
   U14661 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_716_port, B1 => n11427, 
                           B2 => n11361, ZN => n4228);
   U14662 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_717_port, B1 => n11428, 
                           B2 => n11361, ZN => n4227);
   U14663 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_718_port, B1 => n11429, 
                           B2 => n11361, ZN => n4226);
   U14664 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_719_port, B1 => n11430, 
                           B2 => n11361, ZN => n4225);
   U14665 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_720_port, B1 => n11431, 
                           B2 => n11361, ZN => n4224);
   U14666 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_721_port, B1 => n11432, 
                           B2 => n11361, ZN => n4223);
   U14667 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_722_port, B1 => n11433, 
                           B2 => n11361, ZN => n4222);
   U14668 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_723_port, B1 => n11434, 
                           B2 => n11361, ZN => n4221);
   U14669 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_724_port, B1 => n11435, 
                           B2 => n11361, ZN => n4220);
   U14670 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_725_port, B1 => n11436, 
                           B2 => n11361, ZN => n4219);
   U14671 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_726_port, B1 => n11437, 
                           B2 => n11361, ZN => n4218);
   U14672 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_727_port, B1 => n11438, 
                           B2 => n11361, ZN => n4217);
   U14673 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_728_port, B1 => n11439, 
                           B2 => n11361, ZN => n4216);
   U14674 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_729_port, B1 => n11440, 
                           B2 => n11361, ZN => n4215);
   U14675 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_730_port, B1 => n11441, 
                           B2 => n11361, ZN => n4214);
   U14676 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_731_port, B1 => n11442, 
                           B2 => n11361, ZN => n4213);
   U14677 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_732_port, B1 => n11443, 
                           B2 => n11361, ZN => n4212);
   U14678 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_733_port, B1 => n11444, 
                           B2 => n11361, ZN => n4211);
   U14679 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_734_port, B1 => n11445, 
                           B2 => n11361, ZN => n4210);
   U14680 : AOI22_X1 port map( A1 => n11362, A2 => 
                           DataPath_RF_bus_reg_dataout_735_port, B1 => n11447, 
                           B2 => n11361, ZN => n4207);
   U14681 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_672_port, B1 => n11415, 
                           B2 => n11364, ZN => n4205);
   U14682 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_673_port, B1 => n11416, 
                           B2 => n11364, ZN => n4204);
   U14683 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_674_port, B1 => n11417, 
                           B2 => n11364, ZN => n4203);
   U14684 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_675_port, B1 => n11418, 
                           B2 => n11364, ZN => n4202);
   U14685 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_676_port, B1 => n11419, 
                           B2 => n11364, ZN => n4201);
   U14686 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_677_port, B1 => n11420, 
                           B2 => n11364, ZN => n4200);
   U14687 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_678_port, B1 => n11421, 
                           B2 => n11364, ZN => n4199);
   U14688 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_679_port, B1 => n11422, 
                           B2 => n11364, ZN => n4198);
   U14689 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_680_port, B1 => n11423, 
                           B2 => n11364, ZN => n4197);
   U14690 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_681_port, B1 => n11424, 
                           B2 => n11364, ZN => n4196);
   U14691 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_682_port, B1 => n11425, 
                           B2 => n11364, ZN => n4195);
   U14692 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_683_port, B1 => n11426, 
                           B2 => n11364, ZN => n4194);
   U14693 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_684_port, B1 => n11427, 
                           B2 => n11364, ZN => n4193);
   U14694 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_685_port, B1 => n11428, 
                           B2 => n11364, ZN => n4192);
   U14695 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_686_port, B1 => n11429, 
                           B2 => n11364, ZN => n4191);
   U14696 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_687_port, B1 => n11430, 
                           B2 => n11364, ZN => n4190);
   U14697 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_688_port, B1 => n11431, 
                           B2 => n11364, ZN => n4189);
   U14698 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_689_port, B1 => n11432, 
                           B2 => n11364, ZN => n4188);
   U14699 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_690_port, B1 => n11433, 
                           B2 => n11364, ZN => n4187);
   U14700 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_691_port, B1 => n11434, 
                           B2 => n11364, ZN => n4186);
   U14701 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_692_port, B1 => n11435, 
                           B2 => n11364, ZN => n4185);
   U14702 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_693_port, B1 => n11436, 
                           B2 => n11364, ZN => n4184);
   U14703 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_694_port, B1 => n11437, 
                           B2 => n11364, ZN => n4183);
   U14704 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_695_port, B1 => n11438, 
                           B2 => n11364, ZN => n4182);
   U14705 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_696_port, B1 => n11439, 
                           B2 => n11364, ZN => n4181);
   U14706 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_697_port, B1 => n11440, 
                           B2 => n11364, ZN => n4180);
   U14707 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_698_port, B1 => n11441, 
                           B2 => n11364, ZN => n4179);
   U14708 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_699_port, B1 => n11442, 
                           B2 => n11364, ZN => n4178);
   U14709 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_700_port, B1 => n11443, 
                           B2 => n11364, ZN => n4177);
   U14710 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_701_port, B1 => n11444, 
                           B2 => n11364, ZN => n4176);
   U14711 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_702_port, B1 => n11445, 
                           B2 => n11364, ZN => n4175);
   U14712 : AOI22_X1 port map( A1 => n11365, A2 => 
                           DataPath_RF_bus_reg_dataout_703_port, B1 => n11447, 
                           B2 => n11364, ZN => n4172);
   U14713 : OAI22_X1 port map( A1 => n8333, A2 => n11562, B1 => n11412, B2 => 
                           n11561, ZN => n11366);
   U14714 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_640_port, B1 => n11415, 
                           B2 => n11367, ZN => n4170);
   U14715 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_641_port, B1 => n11416, 
                           B2 => n11367, ZN => n4169);
   U14716 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_642_port, B1 => n11417, 
                           B2 => n11367, ZN => n4168);
   U14717 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_643_port, B1 => n11418, 
                           B2 => n11367, ZN => n4167);
   U14718 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_644_port, B1 => n11419, 
                           B2 => n11367, ZN => n4166);
   U14719 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_645_port, B1 => n11420, 
                           B2 => n11367, ZN => n4165);
   U14720 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_646_port, B1 => n11421, 
                           B2 => n11367, ZN => n4164);
   U14721 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_647_port, B1 => n11422, 
                           B2 => n11367, ZN => n4163);
   U14722 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_648_port, B1 => n11423, 
                           B2 => n11367, ZN => n4162);
   U14723 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_649_port, B1 => n11424, 
                           B2 => n11367, ZN => n4161);
   U14724 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_650_port, B1 => n11425, 
                           B2 => n11367, ZN => n4160);
   U14725 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_651_port, B1 => n11426, 
                           B2 => n11367, ZN => n4159);
   U14726 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_652_port, B1 => n11427, 
                           B2 => n11367, ZN => n4158);
   U14727 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_653_port, B1 => n11428, 
                           B2 => n11367, ZN => n4157);
   U14728 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_654_port, B1 => n11429, 
                           B2 => n11367, ZN => n4156);
   U14729 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_655_port, B1 => n11430, 
                           B2 => n11367, ZN => n4155);
   U14730 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_656_port, B1 => n11431, 
                           B2 => n11367, ZN => n4154);
   U14731 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_657_port, B1 => n11432, 
                           B2 => n11367, ZN => n4153);
   U14732 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_658_port, B1 => n11433, 
                           B2 => n11367, ZN => n4152);
   U14733 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_659_port, B1 => n11434, 
                           B2 => n11367, ZN => n4151);
   U14734 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_660_port, B1 => n11435, 
                           B2 => n11367, ZN => n4150);
   U14735 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_661_port, B1 => n11436, 
                           B2 => n11367, ZN => n4149);
   U14736 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_662_port, B1 => n11437, 
                           B2 => n11367, ZN => n4148);
   U14737 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_663_port, B1 => n11438, 
                           B2 => n11367, ZN => n4147);
   U14738 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_664_port, B1 => n11439, 
                           B2 => n11367, ZN => n4146);
   U14739 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_665_port, B1 => n11440, 
                           B2 => n11367, ZN => n4145);
   U14740 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_666_port, B1 => n11441, 
                           B2 => n11367, ZN => n4144);
   U14741 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_667_port, B1 => n11442, 
                           B2 => n11367, ZN => n4143);
   U14742 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_668_port, B1 => n11443, 
                           B2 => n11367, ZN => n4142);
   U14743 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_669_port, B1 => n11444, 
                           B2 => n11367, ZN => n4141);
   U14744 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_670_port, B1 => n11445, 
                           B2 => n11367, ZN => n4140);
   U14745 : AOI22_X1 port map( A1 => n11368, A2 => 
                           DataPath_RF_bus_reg_dataout_671_port, B1 => n11447, 
                           B2 => n11367, ZN => n4137);
   U14746 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_608_port, A2 
                           => n11372, B1 => n11371, B2 => n11374, ZN => n4135);
   U14747 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_609_port, A2 
                           => n8513, B1 => n11371, B2 => n11375, ZN => n4134);
   U14748 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_610_port, A2 
                           => n8513, B1 => n11371, B2 => n11376, ZN => n4133);
   U14749 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_611_port, A2 
                           => n11372, B1 => n11371, B2 => n11377, ZN => n4132);
   U14750 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_612_port, A2 
                           => n11372, B1 => n11371, B2 => n11378, ZN => n4131);
   U14751 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_613_port, A2 
                           => n8513, B1 => n11371, B2 => n11379, ZN => n4130);
   U14752 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_614_port, A2 
                           => n8513, B1 => n11371, B2 => n11380, ZN => n4129);
   U14753 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_615_port, A2 
                           => n8513, B1 => n11371, B2 => n11381, ZN => n4128);
   U14754 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_616_port, A2 
                           => n11372, B1 => n11371, B2 => n11382, ZN => n4127);
   U14755 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_617_port, A2 
                           => n8513, B1 => n11371, B2 => n11383, ZN => n4126);
   U14756 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_618_port, A2 
                           => n8513, B1 => n11371, B2 => n11384, ZN => n4125);
   U14757 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_619_port, A2 
                           => n8513, B1 => n11371, B2 => n11385, ZN => n4124);
   U14758 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_620_port, A2 
                           => n8513, B1 => n11371, B2 => n11386, ZN => n4123);
   U14759 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_621_port, A2 
                           => n11372, B1 => n11371, B2 => n11387, ZN => n4122);
   U14760 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_622_port, A2 
                           => n8513, B1 => n11371, B2 => n11388, ZN => n4121);
   U14761 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_623_port, A2 
                           => n8513, B1 => n11371, B2 => n11389, ZN => n4120);
   U14762 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_624_port, A2 
                           => n11372, B1 => n11371, B2 => n11390, ZN => n4119);
   U14763 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_625_port, A2 
                           => n8513, B1 => n11371, B2 => n11391, ZN => n4118);
   U14764 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_626_port, A2 
                           => n8513, B1 => n11371, B2 => n11392, ZN => n4117);
   U14765 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_627_port, A2 
                           => n8513, B1 => n11371, B2 => n11393, ZN => n4116);
   U14766 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_628_port, A2 
                           => n8513, B1 => n11371, B2 => n11394, ZN => n4115);
   U14767 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_629_port, A2 
                           => n8513, B1 => n11371, B2 => n11395, ZN => n4114);
   U14768 : AOI22_X1 port map( A1 => n11437, A2 => n11370, B1 => n11372, B2 => 
                           DataPath_RF_bus_reg_dataout_630_port, ZN => n4113);
   U14769 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_631_port, A2 
                           => n8513, B1 => n11371, B2 => n11397, ZN => n4112);
   U14770 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_632_port, A2 
                           => n11372, B1 => n11371, B2 => n11369, ZN => n4111);
   U14771 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_633_port, A2 
                           => n8513, B1 => n11371, B2 => n11399, ZN => n4110);
   U14772 : AOI22_X1 port map( A1 => n11441, A2 => n11370, B1 => n11372, B2 => 
                           DataPath_RF_bus_reg_dataout_634_port, ZN => n4109);
   U14773 : AOI22_X1 port map( A1 => n11442, A2 => n11370, B1 => n8513, B2 => 
                           DataPath_RF_bus_reg_dataout_635_port, ZN => n4108);
   U14774 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_636_port, A2 
                           => n11372, B1 => n11371, B2 => n11402, ZN => n4107);
   U14775 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_637_port, A2 
                           => n8513, B1 => n11371, B2 => n11403, ZN => n4106);
   U14776 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_638_port, A2 
                           => n8513, B1 => n11371, B2 => n11404, ZN => n4105);
   U14777 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_639_port, A2 
                           => n8513, B1 => n11371, B2 => n11405, ZN => n4102);
   U14778 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_576_port, A2 
                           => n8514, B1 => n11406, B2 => n11374, ZN => n4100);
   U14779 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_577_port, A2 
                           => n8514, B1 => n11406, B2 => n11375, ZN => n4099);
   U14780 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_578_port, A2 
                           => n11407, B1 => n11406, B2 => n11376, ZN => n4098);
   U14781 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_579_port, A2 
                           => n11407, B1 => n11406, B2 => n11377, ZN => n4097);
   U14782 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_580_port, A2 
                           => n8514, B1 => n11406, B2 => n11378, ZN => n4096);
   U14783 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_581_port, A2 
                           => n8514, B1 => n11406, B2 => n11379, ZN => n4095);
   U14784 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_582_port, A2 
                           => n11407, B1 => n11406, B2 => n11380, ZN => n4094);
   U14785 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_583_port, A2 
                           => n8514, B1 => n11406, B2 => n11381, ZN => n4093);
   U14786 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_584_port, A2 
                           => n8514, B1 => n11406, B2 => n11382, ZN => n4092);
   U14787 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_585_port, A2 
                           => n8514, B1 => n11406, B2 => n11383, ZN => n4091);
   U14788 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_586_port, A2 
                           => n11407, B1 => n11406, B2 => n11384, ZN => n4090);
   U14789 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_587_port, A2 
                           => n8514, B1 => n11406, B2 => n11385, ZN => n4089);
   U14790 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_588_port, A2 
                           => n11407, B1 => n11406, B2 => n11386, ZN => n4088);
   U14791 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_589_port, A2 
                           => n8514, B1 => n11406, B2 => n11387, ZN => n4087);
   U14792 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_590_port, A2 
                           => n8514, B1 => n11406, B2 => n11388, ZN => n4086);
   U14793 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_591_port, A2 
                           => n11407, B1 => n11406, B2 => n11389, ZN => n4085);
   U14794 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_592_port, A2 
                           => n8514, B1 => n11406, B2 => n11390, ZN => n4084);
   U14795 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_593_port, A2 
                           => n8514, B1 => n11406, B2 => n11391, ZN => n4083);
   U14796 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_594_port, A2 
                           => n8514, B1 => n11406, B2 => n11392, ZN => n4082);
   U14797 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_595_port, A2 
                           => n8514, B1 => n11406, B2 => n11393, ZN => n4081);
   U14798 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_596_port, A2 
                           => n8514, B1 => n11406, B2 => n11394, ZN => n4080);
   U14799 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_597_port, A2 
                           => n11407, B1 => n11406, B2 => n11395, ZN => n4079);
   U14800 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_598_port, A2 
                           => n11407, B1 => n11406, B2 => n11396, ZN => n4078);
   U14801 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_599_port, A2 
                           => n8514, B1 => n11406, B2 => n11397, ZN => n4077);
   U14802 : AOI22_X1 port map( A1 => n11439, A2 => n11398, B1 => n8514, B2 => 
                           DataPath_RF_bus_reg_dataout_600_port, ZN => n4076);
   U14803 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_601_port, A2 
                           => n11407, B1 => n11406, B2 => n11399, ZN => n4075);
   U14804 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_602_port, A2 
                           => n8514, B1 => n11406, B2 => n11400, ZN => n4074);
   U14805 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_603_port, A2 
                           => n8514, B1 => n11406, B2 => n11401, ZN => n4073);
   U14806 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_604_port, A2 
                           => n8514, B1 => n11406, B2 => n11402, ZN => n4072);
   U14807 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_605_port, A2 
                           => n8514, B1 => n11406, B2 => n11403, ZN => n4071);
   U14808 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_606_port, A2 
                           => n11407, B1 => n11406, B2 => n11404, ZN => n4070);
   U14809 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_607_port, A2 
                           => n8514, B1 => n11406, B2 => n11405, ZN => n4067);
   U14810 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_544_port, B1 => n11415, 
                           B2 => n11410, ZN => n4065);
   U14811 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_545_port, B1 => n11416, 
                           B2 => n11410, ZN => n4064);
   U14812 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_546_port, B1 => n11417, 
                           B2 => n11410, ZN => n4063);
   U14813 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_547_port, B1 => n11418, 
                           B2 => n11410, ZN => n4062);
   U14814 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_548_port, B1 => n11419, 
                           B2 => n11410, ZN => n4061);
   U14815 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_549_port, B1 => n11420, 
                           B2 => n11410, ZN => n4060);
   U14816 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_550_port, B1 => n11421, 
                           B2 => n11410, ZN => n4059);
   U14817 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_551_port, B1 => n11422, 
                           B2 => n11410, ZN => n4058);
   U14818 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_552_port, B1 => n11423, 
                           B2 => n11410, ZN => n4057);
   U14819 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_553_port, B1 => n11424, 
                           B2 => n11410, ZN => n4056);
   U14820 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_554_port, B1 => n11425, 
                           B2 => n11410, ZN => n4055);
   U14821 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_555_port, B1 => n11426, 
                           B2 => n11410, ZN => n4054);
   U14822 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_556_port, B1 => n11427, 
                           B2 => n11410, ZN => n4053);
   U14823 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_557_port, B1 => n11428, 
                           B2 => n11410, ZN => n4052);
   U14824 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_558_port, B1 => n11429, 
                           B2 => n11410, ZN => n4051);
   U14825 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_559_port, B1 => n11430, 
                           B2 => n11410, ZN => n4050);
   U14826 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_560_port, B1 => n11431, 
                           B2 => n11410, ZN => n4049);
   U14827 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_561_port, B1 => n11432, 
                           B2 => n11410, ZN => n4048);
   U14828 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_562_port, B1 => n11433, 
                           B2 => n11410, ZN => n4047);
   U14829 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_563_port, B1 => n11434, 
                           B2 => n11410, ZN => n4046);
   U14830 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_564_port, B1 => n11435, 
                           B2 => n11410, ZN => n4045);
   U14831 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_565_port, B1 => n11436, 
                           B2 => n11410, ZN => n4044);
   U14832 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_566_port, B1 => n11437, 
                           B2 => n11410, ZN => n4043);
   U14833 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_567_port, B1 => n11438, 
                           B2 => n11410, ZN => n4042);
   U14834 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_568_port, B1 => n11439, 
                           B2 => n11410, ZN => n4041);
   U14835 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_569_port, B1 => n11440, 
                           B2 => n11410, ZN => n4040);
   U14836 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_570_port, B1 => n11441, 
                           B2 => n11410, ZN => n4039);
   U14837 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_571_port, B1 => n11442, 
                           B2 => n11410, ZN => n4038);
   U14838 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_572_port, B1 => n11443, 
                           B2 => n11410, ZN => n4037);
   U14839 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_573_port, B1 => n11444, 
                           B2 => n11410, ZN => n4036);
   U14840 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_574_port, B1 => n11445, 
                           B2 => n11410, ZN => n4035);
   U14841 : AOI22_X1 port map( A1 => n11411, A2 => 
                           DataPath_RF_bus_reg_dataout_575_port, B1 => n11447, 
                           B2 => n11410, ZN => n4032);
   U14842 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_512_port, B1 => n11415, 
                           B2 => n11446, ZN => n4028);
   U14843 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_513_port, B1 => n11416, 
                           B2 => n11446, ZN => n4026);
   U14844 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_514_port, B1 => n11417, 
                           B2 => n11446, ZN => n4024);
   U14845 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_515_port, B1 => n11418, 
                           B2 => n11446, ZN => n4022);
   U14846 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_516_port, B1 => n11419, 
                           B2 => n11446, ZN => n4020);
   U14847 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_517_port, B1 => n11420, 
                           B2 => n11446, ZN => n4018);
   U14848 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_518_port, B1 => n11421, 
                           B2 => n11446, ZN => n4016);
   U14849 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_519_port, B1 => n11422, 
                           B2 => n11446, ZN => n4014);
   U14850 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_520_port, B1 => n11423, 
                           B2 => n11446, ZN => n4012);
   U14851 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_521_port, B1 => n11424, 
                           B2 => n11446, ZN => n4010);
   U14852 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_522_port, B1 => n11425, 
                           B2 => n11446, ZN => n4008);
   U14853 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_523_port, B1 => n11426, 
                           B2 => n11446, ZN => n4006);
   U14854 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_524_port, B1 => n11427, 
                           B2 => n11446, ZN => n4004);
   U14855 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_525_port, B1 => n11428, 
                           B2 => n11446, ZN => n4002);
   U14856 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_526_port, B1 => n11429, 
                           B2 => n11446, ZN => n4000);
   U14857 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_527_port, B1 => n11430, 
                           B2 => n11446, ZN => n3998);
   U14858 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_528_port, B1 => n11431, 
                           B2 => n11446, ZN => n3996);
   U14859 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_529_port, B1 => n11432, 
                           B2 => n11446, ZN => n3994);
   U14860 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_530_port, B1 => n11433, 
                           B2 => n11446, ZN => n3992);
   U14861 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_531_port, B1 => n11434, 
                           B2 => n11446, ZN => n3990);
   U14862 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_532_port, B1 => n11435, 
                           B2 => n11446, ZN => n3988);
   U14863 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_533_port, B1 => n11436, 
                           B2 => n11446, ZN => n3986);
   U14864 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_534_port, B1 => n11437, 
                           B2 => n11446, ZN => n3984);
   U14865 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_535_port, B1 => n11438, 
                           B2 => n11446, ZN => n3982);
   U14866 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_536_port, B1 => n11439, 
                           B2 => n11446, ZN => n3980);
   U14867 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_537_port, B1 => n11440, 
                           B2 => n11446, ZN => n3978);
   U14868 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_538_port, B1 => n11441, 
                           B2 => n11446, ZN => n3976);
   U14869 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_539_port, B1 => n11442, 
                           B2 => n11446, ZN => n3974);
   U14870 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_540_port, B1 => n11443, 
                           B2 => n11446, ZN => n3972);
   U14871 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_541_port, B1 => n11444, 
                           B2 => n11446, ZN => n3970);
   U14872 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_542_port, B1 => n11445, 
                           B2 => n11446, ZN => n3968);
   U14873 : AOI22_X1 port map( A1 => n11448, A2 => 
                           DataPath_RF_bus_reg_dataout_543_port, B1 => n11447, 
                           B2 => n11446, ZN => n3964);
   U14874 : OAI22_X1 port map( A1 => n7766, A2 => n11450, B1 => n11645, B2 => 
                           n8296, ZN => n11525);
   U14875 : AOI22_X1 port map( A1 => n11586, A2 => n11491, B1 => n8516, B2 => 
                           DataPath_RF_bus_reg_dataout_480_port, ZN => n3960);
   U14876 : OAI22_X1 port map( A1 => n8529, A2 => n11451, B1 => n11646, B2 => 
                           n8296, ZN => n11526);
   U14877 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_481_port, A2 
                           => n8516, B1 => n11587, B2 => n8515, ZN => n3958);
   U14878 : OAI22_X1 port map( A1 => n7766, A2 => n11452, B1 => n11647, B2 => 
                           n8296, ZN => n11527);
   U14879 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_482_port, A2 
                           => n8516, B1 => n11588, B2 => n11491, ZN => n3956);
   U14880 : OAI22_X1 port map( A1 => n8529, A2 => n11453, B1 => n11648, B2 => 
                           n8296, ZN => n11528);
   U14881 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_483_port, A2 
                           => n8516, B1 => n11589, B2 => n11491, ZN => n3954);
   U14882 : OAI22_X1 port map( A1 => n7766, A2 => n11454, B1 => n11649, B2 => 
                           n8296, ZN => n11529);
   U14883 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_484_port, A2 
                           => n11498, B1 => n11590, B2 => n8515, ZN => n3952);
   U14884 : NAND2_X1 port map( A1 => n8579, A2 => n11456, ZN => n3232);
   U14885 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_485_port, A2 
                           => n8516, B1 => n11591, B2 => n8515, ZN => n3950);
   U14886 : OAI22_X1 port map( A1 => n7766, A2 => n11457, B1 => n11651, B2 => 
                           n8296, ZN => n11530);
   U14887 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_486_port, A2 
                           => n11498, B1 => n11592, B2 => n11491, ZN => n3948);
   U14888 : OAI22_X1 port map( A1 => n7766, A2 => n11458, B1 => n11652, B2 => 
                           n8296, ZN => n11531);
   U14889 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_487_port, A2 
                           => n8516, B1 => n11593, B2 => n11491, ZN => n3946);
   U14890 : OAI22_X1 port map( A1 => n7766, A2 => n11459, B1 => n11653, B2 => 
                           n8296, ZN => n11532);
   U14891 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_488_port, A2 
                           => n8516, B1 => n11594, B2 => n8515, ZN => n3944);
   U14892 : NAND2_X1 port map( A1 => n8581, A2 => n11461, ZN => n3228);
   U14893 : OAI22_X1 port map( A1 => n8516, A2 => n11595, B1 => 
                           DataPath_RF_bus_reg_dataout_489_port, B2 => n8515, 
                           ZN => n3942);
   U14894 : OAI22_X1 port map( A1 => n8529, A2 => n11462, B1 => n11655, B2 => 
                           n8296, ZN => n11533);
   U14895 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_490_port, A2 
                           => n8516, B1 => n11596, B2 => n8515, ZN => n3940);
   U14896 : OAI22_X1 port map( A1 => n7766, A2 => n11463, B1 => n11656, B2 => 
                           n8296, ZN => n11534);
   U14897 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_491_port, A2 
                           => n8516, B1 => n11597, B2 => n11491, ZN => n3938);
   U14898 : OAI22_X1 port map( A1 => n7766, A2 => n11464, B1 => n11657, B2 => 
                           n8296, ZN => n11535);
   U14899 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_492_port, A2 
                           => n11498, B1 => n11598, B2 => n11491, ZN => n3936);
   U14900 : OAI22_X1 port map( A1 => n7766, A2 => n11465, B1 => n11658, B2 => 
                           n8296, ZN => n11536);
   U14901 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_493_port, A2 
                           => n8516, B1 => n11599, B2 => n8515, ZN => n3934);
   U14902 : OAI22_X1 port map( A1 => n7766, A2 => n11466, B1 => n11659, B2 => 
                           n8296, ZN => n11537);
   U14903 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_494_port, A2 
                           => n11498, B1 => n11600, B2 => n8515, ZN => n3932);
   U14904 : NAND2_X1 port map( A1 => n8582, A2 => n11468, ZN => n3222);
   U14905 : OAI22_X1 port map( A1 => n8516, A2 => n11601, B1 => 
                           DataPath_RF_bus_reg_dataout_495_port, B2 => n8515, 
                           ZN => n3930);
   U14906 : NAND2_X1 port map( A1 => n8574, A2 => n11470, ZN => n3221);
   U14907 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_496_port, B1 => n11602, 
                           B2 => n11497, ZN => n3928);
   U14908 : NAND2_X1 port map( A1 => n8574, A2 => n11472, ZN => n3220);
   U14909 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_497_port, B1 => n11603, 
                           B2 => n11497, ZN => n3926);
   U14910 : OAI22_X1 port map( A1 => n7766, A2 => n11473, B1 => n11663, B2 => 
                           n8296, ZN => n11538);
   U14911 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_498_port, A2 
                           => n11498, B1 => n11604, B2 => n11491, ZN => n3924);
   U14912 : NAND2_X1 port map( A1 => n8574, A2 => n11475, ZN => n3218);
   U14913 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_499_port, B1 => n11605, 
                           B2 => n11497, ZN => n3922);
   U14914 : NAND2_X1 port map( A1 => n8574, A2 => n11476, ZN => n3217);
   U14915 : AOI22_X1 port map( A1 => n11498, A2 => 
                           DataPath_RF_bus_reg_dataout_500_port, B1 => n11606, 
                           B2 => n11497, ZN => n3920);
   U14916 : OAI22_X1 port map( A1 => n7766, A2 => n11477, B1 => n11666, B2 => 
                           n8296, ZN => n11539);
   U14917 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_501_port, A2 
                           => n8516, B1 => n11607, B2 => n11491, ZN => n3918);
   U14918 : OAI22_X1 port map( A1 => n7766, A2 => n11478, B1 => n11667, B2 => 
                           n8296, ZN => n11502);
   U14919 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_502_port, A2 
                           => n11498, B1 => n11608, B2 => n8515, ZN => n3916);
   U14920 : NAND2_X1 port map( A1 => n8574, A2 => n11480, ZN => n3214);
   U14921 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_503_port, A2 
                           => n8516, B1 => n11609, B2 => n8515, ZN => n3914);
   U14922 : NAND2_X1 port map( A1 => n8574, A2 => n11482, ZN => n3213);
   U14923 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_504_port, A2 
                           => n8516, B1 => n11610, B2 => n11491, ZN => n3912);
   U14924 : NAND2_X1 port map( A1 => n8573, A2 => n11484, ZN => n3212);
   U14925 : OAI22_X1 port map( A1 => n11498, A2 => n11611, B1 => 
                           DataPath_RF_bus_reg_dataout_505_port, B2 => n11491, 
                           ZN => n3910);
   U14926 : OAI22_X1 port map( A1 => n7766, A2 => n11485, B1 => n11671, B2 => 
                           n8296, ZN => n11519);
   U14927 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_506_port, A2 
                           => n8516, B1 => n11612, B2 => n8515, ZN => n3908);
   U14928 : NAND2_X1 port map( A1 => n8574, A2 => n11487, ZN => n3210);
   U14929 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_507_port, B1 => n11613, 
                           B2 => n11497, ZN => n3906);
   U14930 : NAND2_X1 port map( A1 => n8574, A2 => n11489, ZN => n3209);
   U14931 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_508_port, B1 => n11614, 
                           B2 => n11497, ZN => n3904);
   U14932 : NAND2_X1 port map( A1 => n8574, A2 => n11490, ZN => n3208);
   U14933 : OAI22_X1 port map( A1 => n8516, A2 => n11615, B1 => 
                           DataPath_RF_bus_reg_dataout_509_port, B2 => n11491, 
                           ZN => n3902);
   U14934 : NAND2_X1 port map( A1 => n8574, A2 => n11493, ZN => n3207);
   U14935 : AOI22_X1 port map( A1 => n8516, A2 => 
                           DataPath_RF_bus_reg_dataout_510_port, B1 => n11616, 
                           B2 => n11497, ZN => n3900);
   U14936 : NAND2_X1 port map( A1 => n8573, A2 => n11495, ZN => n3204);
   U14937 : AOI22_X1 port map( A1 => n11498, A2 => 
                           DataPath_RF_bus_reg_dataout_511_port, B1 => n11751, 
                           B2 => n11497, ZN => n3896);
   U14938 : AOI22_X1 port map( A1 => n11586, A2 => n11499, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_448_port, ZN => n3894);
   U14939 : AOI22_X1 port map( A1 => n11587, A2 => n8517, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_449_port, ZN => n3893);
   U14940 : AOI22_X1 port map( A1 => n11588, A2 => n8517, B1 => n11501, B2 => 
                           DataPath_RF_bus_reg_dataout_450_port, ZN => n3892);
   U14941 : AOI22_X1 port map( A1 => n11589, A2 => n11499, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_451_port, ZN => n3891);
   U14942 : AOI22_X1 port map( A1 => n11590, A2 => n11499, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_452_port, ZN => n3890);
   U14943 : AOI22_X1 port map( A1 => n11591, A2 => n8517, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_453_port, ZN => n3889);
   U14944 : AOI22_X1 port map( A1 => n11592, A2 => n8517, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_454_port, ZN => n3888);
   U14945 : AOI22_X1 port map( A1 => n11593, A2 => n11499, B1 => n11501, B2 => 
                           DataPath_RF_bus_reg_dataout_455_port, ZN => n3887);
   U14946 : AOI22_X1 port map( A1 => n11594, A2 => n11499, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_456_port, ZN => n3886);
   U14947 : OAI22_X1 port map( A1 => n11595, A2 => n8518, B1 => 
                           DataPath_RF_bus_reg_dataout_457_port, B2 => n8517, 
                           ZN => n3885);
   U14948 : AOI22_X1 port map( A1 => n11596, A2 => n8517, B1 => n11501, B2 => 
                           DataPath_RF_bus_reg_dataout_458_port, ZN => n3884);
   U14949 : AOI22_X1 port map( A1 => n11597, A2 => n8517, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_459_port, ZN => n3883);
   U14950 : AOI22_X1 port map( A1 => n11598, A2 => n11499, B1 => n11501, B2 => 
                           DataPath_RF_bus_reg_dataout_460_port, ZN => n3882);
   U14951 : AOI22_X1 port map( A1 => n11599, A2 => n11499, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_461_port, ZN => n3881);
   U14952 : AOI22_X1 port map( A1 => n11600, A2 => n8517, B1 => n11501, B2 => 
                           DataPath_RF_bus_reg_dataout_462_port, ZN => n3880);
   U14953 : OAI22_X1 port map( A1 => n11601, A2 => n11501, B1 => 
                           DataPath_RF_bus_reg_dataout_463_port, B2 => n8517, 
                           ZN => n3879);
   U14954 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_464_port, B1 => n11602, 
                           B2 => n11500, ZN => n3878);
   U14955 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_465_port, B1 => n11603, 
                           B2 => n11500, ZN => n3877);
   U14956 : AOI22_X1 port map( A1 => n11604, A2 => n8517, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_466_port, ZN => n3876);
   U14957 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_467_port, B1 => n11605, 
                           B2 => n11500, ZN => n3875);
   U14958 : AOI22_X1 port map( A1 => n11501, A2 => 
                           DataPath_RF_bus_reg_dataout_468_port, B1 => n11606, 
                           B2 => n11500, ZN => n3874);
   U14959 : AOI22_X1 port map( A1 => n11607, A2 => n11499, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_469_port, ZN => n3873);
   U14960 : AOI22_X1 port map( A1 => n11608, A2 => n11499, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_470_port, ZN => n3872);
   U14961 : AOI22_X1 port map( A1 => n11609, A2 => n8517, B1 => n11501, B2 => 
                           DataPath_RF_bus_reg_dataout_471_port, ZN => n3871);
   U14962 : AOI22_X1 port map( A1 => n11610, A2 => n8517, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_472_port, ZN => n3870);
   U14963 : OAI22_X1 port map( A1 => n11611, A2 => n8518, B1 => 
                           DataPath_RF_bus_reg_dataout_473_port, B2 => n8517, 
                           ZN => n3869);
   U14964 : AOI22_X1 port map( A1 => n11612, A2 => n11499, B1 => n8518, B2 => 
                           DataPath_RF_bus_reg_dataout_474_port, ZN => n3868);
   U14965 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_475_port, B1 => n11613, 
                           B2 => n11500, ZN => n3867);
   U14966 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_476_port, B1 => n11614, 
                           B2 => n11500, ZN => n3866);
   U14967 : OAI22_X1 port map( A1 => n11615, A2 => n8518, B1 => 
                           DataPath_RF_bus_reg_dataout_477_port, B2 => n8517, 
                           ZN => n3865);
   U14968 : AOI22_X1 port map( A1 => n8518, A2 => 
                           DataPath_RF_bus_reg_dataout_478_port, B1 => n11616, 
                           B2 => n11500, ZN => n3864);
   U14969 : AOI22_X1 port map( A1 => n11501, A2 => 
                           DataPath_RF_bus_reg_dataout_479_port, B1 => n11751, 
                           B2 => n11500, ZN => n3861);
   U14970 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_416_port, A2 
                           => n8519, B1 => n11503, B2 => n11525, ZN => n3859);
   U14971 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_417_port, A2 
                           => n8519, B1 => n11503, B2 => n11526, ZN => n3858);
   U14972 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_418_port, A2 
                           => n8519, B1 => n11503, B2 => n11527, ZN => n3857);
   U14973 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_419_port, A2 
                           => n11505, B1 => n11503, B2 => n11528, ZN => n3856);
   U14974 : AOI22_X1 port map( A1 => n11590, A2 => n11504, B1 => n8519, B2 => 
                           DataPath_RF_bus_reg_dataout_420_port, ZN => n3855);
   U14975 : OAI22_X1 port map( A1 => n11591, A2 => n8519, B1 => 
                           DataPath_RF_bus_reg_dataout_421_port, B2 => n11504, 
                           ZN => n3854);
   U14976 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_422_port, A2 
                           => n11505, B1 => n11503, B2 => n11530, ZN => n3853);
   U14977 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_423_port, A2 
                           => n8519, B1 => n11503, B2 => n11531, ZN => n3852);
   U14978 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_424_port, A2 
                           => n8519, B1 => n11503, B2 => n11532, ZN => n3851);
   U14979 : OAI22_X1 port map( A1 => n11595, A2 => n11505, B1 => 
                           DataPath_RF_bus_reg_dataout_425_port, B2 => n11504, 
                           ZN => n3850);
   U14980 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_426_port, A2 
                           => n8519, B1 => n11503, B2 => n11533, ZN => n3849);
   U14981 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_427_port, A2 
                           => n11505, B1 => n11503, B2 => n11534, ZN => n3848);
   U14982 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_428_port, A2 
                           => n8519, B1 => n11503, B2 => n11535, ZN => n3847);
   U14983 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_429_port, A2 
                           => n8519, B1 => n11503, B2 => n11536, ZN => n3846);
   U14984 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_430_port, A2 
                           => n8519, B1 => n11503, B2 => n11537, ZN => n3845);
   U14985 : AOI22_X1 port map( A1 => n11601, A2 => n11504, B1 => n11505, B2 => 
                           DataPath_RF_bus_reg_dataout_431_port, ZN => n3844);
   U14986 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_432_port, A2 
                           => n8519, B1 => n11602, B2 => n11504, ZN => n3843);
   U14987 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_433_port, A2 
                           => n11505, B1 => n11603, B2 => n11504, ZN => n3842);
   U14988 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_434_port, A2 
                           => n8519, B1 => n11503, B2 => n11538, ZN => n3841);
   U14989 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_435_port, A2 
                           => n8519, B1 => n11605, B2 => n11504, ZN => n3840);
   U14990 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_436_port, A2 
                           => n8519, B1 => n11606, B2 => n11504, ZN => n3839);
   U14991 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_437_port, A2 
                           => n11505, B1 => n11503, B2 => n11539, ZN => n3838);
   U14992 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_438_port, A2 
                           => n8519, B1 => n11503, B2 => n11502, ZN => n3837);
   U14993 : OAI22_X1 port map( A1 => n11609, A2 => n11505, B1 => 
                           DataPath_RF_bus_reg_dataout_439_port, B2 => n11504, 
                           ZN => n3836);
   U14994 : OAI22_X1 port map( A1 => n11610, A2 => n11505, B1 => 
                           DataPath_RF_bus_reg_dataout_440_port, B2 => n11504, 
                           ZN => n3835);
   U14995 : AOI22_X1 port map( A1 => n11611, A2 => n11504, B1 => n8519, B2 => 
                           DataPath_RF_bus_reg_dataout_441_port, ZN => n3834);
   U14996 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_442_port, A2 
                           => n8519, B1 => n11503, B2 => n11519, ZN => n3833);
   U14997 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_443_port, A2 
                           => n8519, B1 => n11613, B2 => n11504, ZN => n3832);
   U14998 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_444_port, A2 
                           => n11505, B1 => n11614, B2 => n11504, ZN => n3831);
   U14999 : OAI22_X1 port map( A1 => n11615, A2 => n8519, B1 => 
                           DataPath_RF_bus_reg_dataout_445_port, B2 => n11504, 
                           ZN => n3830);
   U15000 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_446_port, A2 
                           => n8519, B1 => n11616, B2 => n11504, ZN => n3829);
   U15001 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_447_port, A2 
                           => n8519, B1 => n11751, B2 => n11504, ZN => n3826);
   U15002 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_384_port, B1 => n11586, 
                           B2 => n11507, ZN => n3824);
   U15003 : AOI22_X1 port map( A1 => n11587, A2 => n11506, B1 => n8520, B2 => 
                           DataPath_RF_bus_reg_dataout_385_port, ZN => n3823);
   U15004 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_386_port, B1 => n11588, 
                           B2 => n11507, ZN => n3822);
   U15005 : AOI22_X1 port map( A1 => n11589, A2 => n11506, B1 => n8520, B2 => 
                           DataPath_RF_bus_reg_dataout_387_port, ZN => n3821);
   U15006 : AOI22_X1 port map( A1 => n11590, A2 => n11506, B1 => n11508, B2 => 
                           DataPath_RF_bus_reg_dataout_388_port, ZN => n3820);
   U15007 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_389_port, B1 => n11591, 
                           B2 => n11507, ZN => n3819);
   U15008 : AOI22_X1 port map( A1 => n11592, A2 => n11506, B1 => n11508, B2 => 
                           DataPath_RF_bus_reg_dataout_390_port, ZN => n3818);
   U15009 : AOI22_X1 port map( A1 => n11593, A2 => n11506, B1 => n8520, B2 => 
                           DataPath_RF_bus_reg_dataout_391_port, ZN => n3817);
   U15010 : AOI22_X1 port map( A1 => n11508, A2 => 
                           DataPath_RF_bus_reg_dataout_392_port, B1 => n11594, 
                           B2 => n11507, ZN => n3816);
   U15011 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_393_port, B1 => n11595, 
                           B2 => n11507, ZN => n3815);
   U15012 : AOI22_X1 port map( A1 => n11596, A2 => n11506, B1 => n8520, B2 => 
                           DataPath_RF_bus_reg_dataout_394_port, ZN => n3814);
   U15013 : AOI22_X1 port map( A1 => n11597, A2 => n11506, B1 => n8520, B2 => 
                           DataPath_RF_bus_reg_dataout_395_port, ZN => n3813);
   U15014 : AOI22_X1 port map( A1 => n11598, A2 => n11506, B1 => n11508, B2 => 
                           DataPath_RF_bus_reg_dataout_396_port, ZN => n3812);
   U15015 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_397_port, B1 => n11599, 
                           B2 => n11507, ZN => n3811);
   U15016 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_398_port, B1 => n11600, 
                           B2 => n11507, ZN => n3810);
   U15017 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_399_port, B1 => n11601, 
                           B2 => n11507, ZN => n3809);
   U15018 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_400_port, B1 => n11602, 
                           B2 => n11507, ZN => n3808);
   U15019 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_401_port, B1 => n11603, 
                           B2 => n11507, ZN => n3807);
   U15020 : AOI22_X1 port map( A1 => n11508, A2 => 
                           DataPath_RF_bus_reg_dataout_402_port, B1 => n11604, 
                           B2 => n11507, ZN => n3806);
   U15021 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_403_port, B1 => n11605, 
                           B2 => n11507, ZN => n3805);
   U15022 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_404_port, B1 => n11606, 
                           B2 => n11507, ZN => n3804);
   U15023 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_405_port, B1 => n11607, 
                           B2 => n11507, ZN => n3803);
   U15024 : AOI22_X1 port map( A1 => n11508, A2 => 
                           DataPath_RF_bus_reg_dataout_406_port, B1 => n11608, 
                           B2 => n11507, ZN => n3802);
   U15025 : AOI22_X1 port map( A1 => n11508, A2 => 
                           DataPath_RF_bus_reg_dataout_407_port, B1 => n11609, 
                           B2 => n11507, ZN => n3801);
   U15026 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_408_port, B1 => n11610, 
                           B2 => n11507, ZN => n3800);
   U15027 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_409_port, B1 => n11611, 
                           B2 => n11507, ZN => n3799);
   U15028 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_410_port, B1 => n11612, 
                           B2 => n11507, ZN => n3798);
   U15029 : AOI22_X1 port map( A1 => n11508, A2 => 
                           DataPath_RF_bus_reg_dataout_411_port, B1 => n11613, 
                           B2 => n11507, ZN => n3797);
   U15030 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_412_port, B1 => n11614, 
                           B2 => n11507, ZN => n3796);
   U15031 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_413_port, B1 => n11615, 
                           B2 => n11507, ZN => n3795);
   U15032 : AOI22_X1 port map( A1 => n8520, A2 => 
                           DataPath_RF_bus_reg_dataout_414_port, B1 => n11616, 
                           B2 => n11507, ZN => n3794);
   U15033 : AOI22_X1 port map( A1 => n11508, A2 => 
                           DataPath_RF_bus_reg_dataout_415_port, B1 => n11751, 
                           B2 => n11507, ZN => n3791);
   U15034 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_352_port, B1 => n11586, 
                           B2 => n11510, ZN => n3789);
   U15035 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_353_port, B1 => n11587, 
                           B2 => n11510, ZN => n3788);
   U15036 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_354_port, B1 => n11588, 
                           B2 => n11510, ZN => n3787);
   U15037 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_355_port, B1 => n11589, 
                           B2 => n11510, ZN => n3786);
   U15038 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_356_port, B1 => n11590, 
                           B2 => n11510, ZN => n3785);
   U15039 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_357_port, B1 => n11591, 
                           B2 => n11510, ZN => n3784);
   U15040 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_358_port, B1 => n11592, 
                           B2 => n11510, ZN => n3783);
   U15041 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_359_port, B1 => n11593, 
                           B2 => n11510, ZN => n3782);
   U15042 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_360_port, B1 => n11594, 
                           B2 => n11510, ZN => n3781);
   U15043 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_361_port, B1 => n11595, 
                           B2 => n11510, ZN => n3780);
   U15044 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_362_port, B1 => n11596, 
                           B2 => n11510, ZN => n3779);
   U15045 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_363_port, B1 => n11597, 
                           B2 => n11510, ZN => n3778);
   U15046 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_364_port, B1 => n11598, 
                           B2 => n11510, ZN => n3777);
   U15047 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_365_port, B1 => n11599, 
                           B2 => n11510, ZN => n3776);
   U15048 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_366_port, B1 => n11600, 
                           B2 => n11510, ZN => n3775);
   U15049 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_367_port, B1 => n11601, 
                           B2 => n11510, ZN => n3774);
   U15050 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_368_port, B1 => n11602, 
                           B2 => n11510, ZN => n3773);
   U15051 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_369_port, B1 => n11603, 
                           B2 => n11510, ZN => n3772);
   U15052 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_370_port, B1 => n11604, 
                           B2 => n11510, ZN => n3771);
   U15053 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_371_port, B1 => n11605, 
                           B2 => n11510, ZN => n3770);
   U15054 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_372_port, B1 => n11606, 
                           B2 => n11510, ZN => n3769);
   U15055 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_373_port, B1 => n11607, 
                           B2 => n11510, ZN => n3768);
   U15056 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_374_port, B1 => n11608, 
                           B2 => n11510, ZN => n3767);
   U15057 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_375_port, B1 => n11609, 
                           B2 => n11510, ZN => n3766);
   U15058 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_376_port, B1 => n11610, 
                           B2 => n11510, ZN => n3765);
   U15059 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_377_port, B1 => n11611, 
                           B2 => n11510, ZN => n3764);
   U15060 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_378_port, B1 => n11612, 
                           B2 => n11510, ZN => n3763);
   U15061 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_379_port, B1 => n11613, 
                           B2 => n11510, ZN => n3762);
   U15062 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_380_port, B1 => n11614, 
                           B2 => n11510, ZN => n3761);
   U15063 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_381_port, B1 => n11615, 
                           B2 => n11510, ZN => n3760);
   U15064 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_382_port, B1 => n11616, 
                           B2 => n11510, ZN => n3759);
   U15065 : AOI22_X1 port map( A1 => n8521, A2 => 
                           DataPath_RF_bus_reg_dataout_383_port, B1 => n11751, 
                           B2 => n11510, ZN => n3756);
   U15066 : AOI22_X1 port map( A1 => n11586, A2 => n11514, B1 => n11516, B2 => 
                           DataPath_RF_bus_reg_dataout_320_port, ZN => n3752);
   U15067 : OAI22_X1 port map( A1 => n11587, A2 => n8523, B1 => 
                           DataPath_RF_bus_reg_dataout_321_port, B2 => n8522, 
                           ZN => n3751);
   U15068 : AOI22_X1 port map( A1 => n11588, A2 => n8522, B1 => n8523, B2 => 
                           DataPath_RF_bus_reg_dataout_322_port, ZN => n3750);
   U15069 : AOI22_X1 port map( A1 => n11589, A2 => n8522, B1 => n11516, B2 => 
                           DataPath_RF_bus_reg_dataout_323_port, ZN => n3749);
   U15070 : OAI22_X1 port map( A1 => n11590, A2 => n8523, B1 => 
                           DataPath_RF_bus_reg_dataout_324_port, B2 => n11514, 
                           ZN => n3748);
   U15071 : AOI22_X1 port map( A1 => n11591, A2 => n11514, B1 => n11516, B2 => 
                           DataPath_RF_bus_reg_dataout_325_port, ZN => n3747);
   U15072 : AOI22_X1 port map( A1 => n11592, A2 => n11514, B1 => n11516, B2 => 
                           DataPath_RF_bus_reg_dataout_326_port, ZN => n3746);
   U15073 : AOI22_X1 port map( A1 => n11593, A2 => n8522, B1 => n8523, B2 => 
                           DataPath_RF_bus_reg_dataout_327_port, ZN => n3745);
   U15074 : AOI22_X1 port map( A1 => n11594, A2 => n8522, B1 => n8523, B2 => 
                           DataPath_RF_bus_reg_dataout_328_port, ZN => n3744);
   U15075 : OAI22_X1 port map( A1 => n11595, A2 => n8523, B1 => 
                           DataPath_RF_bus_reg_dataout_329_port, B2 => n11514, 
                           ZN => n3743);
   U15076 : OAI22_X1 port map( A1 => n11596, A2 => n11516, B1 => 
                           DataPath_RF_bus_reg_dataout_330_port, B2 => n8522, 
                           ZN => n3742);
   U15077 : OAI22_X1 port map( A1 => n11597, A2 => n8523, B1 => 
                           DataPath_RF_bus_reg_dataout_331_port, B2 => n8522, 
                           ZN => n3741);
   U15078 : OAI22_X1 port map( A1 => n11598, A2 => n8523, B1 => 
                           DataPath_RF_bus_reg_dataout_332_port, B2 => n11514, 
                           ZN => n3740);
   U15079 : OAI22_X1 port map( A1 => n11599, A2 => n8523, B1 => 
                           DataPath_RF_bus_reg_dataout_333_port, B2 => n11514, 
                           ZN => n3739);
   U15080 : OAI22_X1 port map( A1 => n11600, A2 => n8523, B1 => 
                           DataPath_RF_bus_reg_dataout_334_port, B2 => n8522, 
                           ZN => n3738);
   U15081 : OAI22_X1 port map( A1 => n11601, A2 => n11516, B1 => 
                           DataPath_RF_bus_reg_dataout_335_port, B2 => n8522, 
                           ZN => n3737);
   U15082 : AOI22_X1 port map( A1 => n8523, A2 => 
                           DataPath_RF_bus_reg_dataout_336_port, B1 => n11602, 
                           B2 => n11515, ZN => n3736);
   U15083 : AOI22_X1 port map( A1 => n8523, A2 => 
                           DataPath_RF_bus_reg_dataout_337_port, B1 => n11603, 
                           B2 => n11515, ZN => n3735);
   U15084 : AOI22_X1 port map( A1 => n11604, A2 => n11514, B1 => n8523, B2 => 
                           DataPath_RF_bus_reg_dataout_338_port, ZN => n3734);
   U15085 : AOI22_X1 port map( A1 => n8523, A2 => 
                           DataPath_RF_bus_reg_dataout_339_port, B1 => n11605, 
                           B2 => n11515, ZN => n3733);
   U15086 : AOI22_X1 port map( A1 => n11516, A2 => 
                           DataPath_RF_bus_reg_dataout_340_port, B1 => n11606, 
                           B2 => n11515, ZN => n3732);
   U15087 : AOI22_X1 port map( A1 => n11607, A2 => n11514, B1 => n8523, B2 => 
                           DataPath_RF_bus_reg_dataout_341_port, ZN => n3731);
   U15088 : AOI22_X1 port map( A1 => n11608, A2 => n8522, B1 => n11516, B2 => 
                           DataPath_RF_bus_reg_dataout_342_port, ZN => n3730);
   U15089 : AOI22_X1 port map( A1 => n11609, A2 => n8522, B1 => n8523, B2 => 
                           DataPath_RF_bus_reg_dataout_343_port, ZN => n3729);
   U15090 : AOI22_X1 port map( A1 => n11610, A2 => n11514, B1 => n8523, B2 => 
                           DataPath_RF_bus_reg_dataout_344_port, ZN => n3728);
   U15091 : OAI22_X1 port map( A1 => n11611, A2 => n8523, B1 => 
                           DataPath_RF_bus_reg_dataout_345_port, B2 => n11514, 
                           ZN => n3727);
   U15092 : AOI22_X1 port map( A1 => n11612, A2 => n11514, B1 => n8523, B2 => 
                           DataPath_RF_bus_reg_dataout_346_port, ZN => n3726);
   U15093 : AOI22_X1 port map( A1 => n8523, A2 => 
                           DataPath_RF_bus_reg_dataout_347_port, B1 => n11613, 
                           B2 => n11515, ZN => n3725);
   U15094 : AOI22_X1 port map( A1 => n8523, A2 => 
                           DataPath_RF_bus_reg_dataout_348_port, B1 => n11614, 
                           B2 => n11515, ZN => n3724);
   U15095 : OAI22_X1 port map( A1 => n11615, A2 => n8523, B1 => 
                           DataPath_RF_bus_reg_dataout_349_port, B2 => n8522, 
                           ZN => n3723);
   U15096 : AOI22_X1 port map( A1 => n8523, A2 => 
                           DataPath_RF_bus_reg_dataout_350_port, B1 => n11616, 
                           B2 => n11515, ZN => n3722);
   U15097 : AOI22_X1 port map( A1 => n11516, A2 => 
                           DataPath_RF_bus_reg_dataout_351_port, B1 => n11751, 
                           B2 => n11515, ZN => n3719);
   U15098 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_288_port, A2 
                           => n8525, B1 => n11520, B2 => n11525, ZN => n3715);
   U15099 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_289_port, A2 
                           => n8525, B1 => n11520, B2 => n11526, ZN => n3714);
   U15100 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_290_port, A2 
                           => n8525, B1 => n11520, B2 => n11527, ZN => n3713);
   U15101 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_291_port, A2 
                           => n11522, B1 => n11520, B2 => n11528, ZN => n3712);
   U15102 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_292_port, A2 
                           => n11522, B1 => n11520, B2 => n11529, ZN => n3711);
   U15103 : OAI22_X1 port map( A1 => n11591, A2 => n8525, B1 => 
                           DataPath_RF_bus_reg_dataout_293_port, B2 => n8524, 
                           ZN => n3710);
   U15104 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_294_port, A2 
                           => n8525, B1 => n11520, B2 => n11530, ZN => n3709);
   U15105 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_295_port, A2 
                           => n8525, B1 => n11520, B2 => n11531, ZN => n3708);
   U15106 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_296_port, A2 
                           => n8525, B1 => n11520, B2 => n11532, ZN => n3707);
   U15107 : AOI22_X1 port map( A1 => n11595, A2 => n11521, B1 => n8525, B2 => 
                           DataPath_RF_bus_reg_dataout_297_port, ZN => n3706);
   U15108 : AOI22_X1 port map( A1 => n11596, A2 => n11521, B1 => n8525, B2 => 
                           DataPath_RF_bus_reg_dataout_298_port, ZN => n3705);
   U15109 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_299_port, A2 
                           => n11522, B1 => n11520, B2 => n11534, ZN => n3704);
   U15110 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_300_port, A2 
                           => n8525, B1 => n11520, B2 => n11535, ZN => n3703);
   U15111 : AOI22_X1 port map( A1 => n11599, A2 => n8524, B1 => n11522, B2 => 
                           DataPath_RF_bus_reg_dataout_301_port, ZN => n3702);
   U15112 : AOI22_X1 port map( A1 => n11600, A2 => n8524, B1 => n11522, B2 => 
                           DataPath_RF_bus_reg_dataout_302_port, ZN => n3701);
   U15113 : OAI22_X1 port map( A1 => n11601, A2 => n8525, B1 => 
                           DataPath_RF_bus_reg_dataout_303_port, B2 => n11521, 
                           ZN => n3700);
   U15114 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_304_port, A2 
                           => n8525, B1 => n11602, B2 => n11521, ZN => n3699);
   U15115 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_305_port, A2 
                           => n8525, B1 => n11603, B2 => n8524, ZN => n3698);
   U15116 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_306_port, A2 
                           => n11522, B1 => n11520, B2 => n11538, ZN => n3697);
   U15117 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_307_port, A2 
                           => n11522, B1 => n11605, B2 => n8524, ZN => n3696);
   U15118 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_308_port, A2 
                           => n8525, B1 => n11606, B2 => n11521, ZN => n3695);
   U15119 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_309_port, A2 
                           => n8525, B1 => n11520, B2 => n11539, ZN => n3694);
   U15120 : AOI22_X1 port map( A1 => n11608, A2 => n11521, B1 => n8525, B2 => 
                           DataPath_RF_bus_reg_dataout_310_port, ZN => n3693);
   U15121 : OAI22_X1 port map( A1 => n11609, A2 => n8525, B1 => 
                           DataPath_RF_bus_reg_dataout_311_port, B2 => n11521, 
                           ZN => n3692);
   U15122 : OAI22_X1 port map( A1 => n11610, A2 => n11522, B1 => 
                           DataPath_RF_bus_reg_dataout_312_port, B2 => n8524, 
                           ZN => n3691);
   U15123 : OAI22_X1 port map( A1 => n11611, A2 => n8525, B1 => 
                           DataPath_RF_bus_reg_dataout_313_port, B2 => n8524, 
                           ZN => n3690);
   U15124 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_314_port, A2 
                           => n8525, B1 => n11520, B2 => n11519, ZN => n3689);
   U15125 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_315_port, A2 
                           => n8525, B1 => n11613, B2 => n11521, ZN => n3688);
   U15126 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_316_port, A2 
                           => n11522, B1 => n11614, B2 => n8524, ZN => n3687);
   U15127 : AOI22_X1 port map( A1 => n11615, A2 => n11521, B1 => n8525, B2 => 
                           DataPath_RF_bus_reg_dataout_317_port, ZN => n3686);
   U15128 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_318_port, A2 
                           => n8525, B1 => n11616, B2 => n8524, ZN => n3685);
   U15129 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_319_port, A2 
                           => n11522, B1 => n11751, B2 => n8524, ZN => n3682);
   U15130 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_256_port, A2 
                           => n8526, B1 => n11540, B2 => n11525, ZN => n3678);
   U15131 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_257_port, A2 
                           => n8526, B1 => n11540, B2 => n11526, ZN => n3677);
   U15132 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_258_port, A2 
                           => n8526, B1 => n11540, B2 => n11527, ZN => n3676);
   U15133 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_259_port, A2 
                           => n11542, B1 => n11540, B2 => n11528, ZN => n3675);
   U15134 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_260_port, A2 
                           => n8526, B1 => n11540, B2 => n11529, ZN => n3674);
   U15135 : OAI22_X1 port map( A1 => n11591, A2 => n11542, B1 => 
                           DataPath_RF_bus_reg_dataout_261_port, B2 => n11541, 
                           ZN => n3673);
   U15136 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_262_port, A2 
                           => n8526, B1 => n11540, B2 => n11530, ZN => n3672);
   U15137 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_263_port, A2 
                           => n8526, B1 => n11540, B2 => n11531, ZN => n3671);
   U15138 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_264_port, A2 
                           => n11542, B1 => n11540, B2 => n11532, ZN => n3670);
   U15139 : OAI22_X1 port map( A1 => n11595, A2 => n8526, B1 => 
                           DataPath_RF_bus_reg_dataout_265_port, B2 => n11541, 
                           ZN => n3669);
   U15140 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_266_port, A2 
                           => n8526, B1 => n11540, B2 => n11533, ZN => n3668);
   U15141 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_267_port, A2 
                           => n8526, B1 => n11540, B2 => n11534, ZN => n3667);
   U15142 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_268_port, A2 
                           => n8526, B1 => n11540, B2 => n11535, ZN => n3666);
   U15143 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_269_port, A2 
                           => n8526, B1 => n11540, B2 => n11536, ZN => n3665);
   U15144 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_270_port, A2 
                           => n11542, B1 => n11540, B2 => n11537, ZN => n3664);
   U15145 : AOI22_X1 port map( A1 => n11601, A2 => n11541, B1 => n8526, B2 => 
                           DataPath_RF_bus_reg_dataout_271_port, ZN => n3663);
   U15146 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_272_port, A2 
                           => n11542, B1 => n11602, B2 => n11541, ZN => n3662);
   U15147 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_273_port, A2 
                           => n8526, B1 => n11603, B2 => n11541, ZN => n3661);
   U15148 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_274_port, A2 
                           => n8526, B1 => n11540, B2 => n11538, ZN => n3660);
   U15149 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_275_port, A2 
                           => n8526, B1 => n11605, B2 => n11541, ZN => n3659);
   U15150 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_276_port, A2 
                           => n11542, B1 => n11606, B2 => n11541, ZN => n3658);
   U15151 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_277_port, A2 
                           => n11542, B1 => n11540, B2 => n11539, ZN => n3657);
   U15152 : AOI22_X1 port map( A1 => n11608, A2 => n11541, B1 => n8526, B2 => 
                           DataPath_RF_bus_reg_dataout_278_port, ZN => n3656);
   U15153 : OAI22_X1 port map( A1 => n11609, A2 => n8526, B1 => 
                           DataPath_RF_bus_reg_dataout_279_port, B2 => n11541, 
                           ZN => n3655);
   U15154 : AOI22_X1 port map( A1 => n11610, A2 => n11541, B1 => n11542, B2 => 
                           DataPath_RF_bus_reg_dataout_280_port, ZN => n3654);
   U15155 : AOI22_X1 port map( A1 => n11611, A2 => n11541, B1 => n11542, B2 => 
                           DataPath_RF_bus_reg_dataout_281_port, ZN => n3653);
   U15156 : AOI22_X1 port map( A1 => n11612, A2 => n11541, B1 => n8526, B2 => 
                           DataPath_RF_bus_reg_dataout_282_port, ZN => n3652);
   U15157 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_283_port, A2 
                           => n8526, B1 => n11613, B2 => n11541, ZN => n3651);
   U15158 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_284_port, A2 
                           => n8526, B1 => n11614, B2 => n11541, ZN => n3650);
   U15159 : AOI22_X1 port map( A1 => n11615, A2 => n11541, B1 => n8526, B2 => 
                           DataPath_RF_bus_reg_dataout_285_port, ZN => n3649);
   U15160 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_286_port, A2 
                           => n8526, B1 => n11616, B2 => n11541, ZN => n3648);
   U15161 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_287_port, A2 
                           => n11542, B1 => n11751, B2 => n11541, ZN => n3645);
   U15162 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_224_port, B1 => n11586, 
                           B2 => n11547, ZN => n3640);
   U15163 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_225_port, B1 => n11587, 
                           B2 => n11547, ZN => n3639);
   U15164 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_226_port, B1 => n11588, 
                           B2 => n11547, ZN => n3638);
   U15165 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_227_port, B1 => n11589, 
                           B2 => n11547, ZN => n3637);
   U15166 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_228_port, B1 => n11590, 
                           B2 => n11547, ZN => n3636);
   U15167 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_229_port, B1 => n11591, 
                           B2 => n11547, ZN => n3635);
   U15168 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_230_port, B1 => n11592, 
                           B2 => n11547, ZN => n3634);
   U15169 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_231_port, B1 => n11593, 
                           B2 => n11547, ZN => n3633);
   U15170 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_232_port, B1 => n11594, 
                           B2 => n11547, ZN => n3632);
   U15171 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_233_port, B1 => n11595, 
                           B2 => n11547, ZN => n3631);
   U15172 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_234_port, B1 => n11596, 
                           B2 => n11547, ZN => n3630);
   U15173 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_235_port, B1 => n11597, 
                           B2 => n11547, ZN => n3629);
   U15174 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_236_port, B1 => n11598, 
                           B2 => n11547, ZN => n3628);
   U15175 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_237_port, B1 => n11599, 
                           B2 => n11547, ZN => n3627);
   U15176 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_238_port, B1 => n11600, 
                           B2 => n11547, ZN => n3626);
   U15177 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_239_port, B1 => n11601, 
                           B2 => n11547, ZN => n3625);
   U15178 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_240_port, B1 => n11602, 
                           B2 => n11547, ZN => n3624);
   U15179 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_241_port, B1 => n11603, 
                           B2 => n11547, ZN => n3623);
   U15180 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_242_port, B1 => n11604, 
                           B2 => n11547, ZN => n3622);
   U15181 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_243_port, B1 => n11605, 
                           B2 => n11547, ZN => n3621);
   U15182 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_244_port, B1 => n11606, 
                           B2 => n11547, ZN => n3620);
   U15183 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_245_port, B1 => n11607, 
                           B2 => n11547, ZN => n3619);
   U15184 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_246_port, B1 => n11608, 
                           B2 => n11547, ZN => n3618);
   U15185 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_247_port, B1 => n11609, 
                           B2 => n11547, ZN => n3617);
   U15186 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_248_port, B1 => n11610, 
                           B2 => n11547, ZN => n3616);
   U15187 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_249_port, B1 => n11611, 
                           B2 => n11547, ZN => n3615);
   U15188 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_250_port, B1 => n11612, 
                           B2 => n11547, ZN => n3614);
   U15189 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_251_port, B1 => n11613, 
                           B2 => n11547, ZN => n3613);
   U15190 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_252_port, B1 => n11614, 
                           B2 => n11547, ZN => n3612);
   U15191 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_253_port, B1 => n11615, 
                           B2 => n11547, ZN => n3611);
   U15192 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_254_port, B1 => n11616, 
                           B2 => n11547, ZN => n3610);
   U15193 : AOI22_X1 port map( A1 => n11548, A2 => 
                           DataPath_RF_bus_reg_dataout_255_port, B1 => n11751, 
                           B2 => n11547, ZN => n3607);
   U15194 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_192_port, B1 => n11586, 
                           B2 => n11553, ZN => n3602);
   U15195 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_193_port, B1 => n11587, 
                           B2 => n11553, ZN => n3601);
   U15196 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_194_port, B1 => n11588, 
                           B2 => n11553, ZN => n3600);
   U15197 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_195_port, B1 => n11589, 
                           B2 => n11553, ZN => n3599);
   U15198 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_196_port, B1 => n11590, 
                           B2 => n11553, ZN => n3598);
   U15199 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_197_port, B1 => n11591, 
                           B2 => n11553, ZN => n3597);
   U15200 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_198_port, B1 => n11592, 
                           B2 => n11553, ZN => n3596);
   U15201 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_199_port, B1 => n11593, 
                           B2 => n11553, ZN => n3595);
   U15202 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_200_port, B1 => n11594, 
                           B2 => n11553, ZN => n3594);
   U15203 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_201_port, B1 => n11595, 
                           B2 => n11553, ZN => n3593);
   U15204 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_202_port, B1 => n11596, 
                           B2 => n11553, ZN => n3592);
   U15205 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_203_port, B1 => n11597, 
                           B2 => n11553, ZN => n3591);
   U15206 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_204_port, B1 => n11598, 
                           B2 => n11553, ZN => n3590);
   U15207 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_205_port, B1 => n11599, 
                           B2 => n11553, ZN => n3589);
   U15208 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_206_port, B1 => n11600, 
                           B2 => n11553, ZN => n3588);
   U15209 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_207_port, B1 => n11601, 
                           B2 => n11553, ZN => n3587);
   U15210 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_208_port, B1 => n11602, 
                           B2 => n11553, ZN => n3586);
   U15211 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_209_port, B1 => n11603, 
                           B2 => n11553, ZN => n3585);
   U15212 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_210_port, B1 => n11604, 
                           B2 => n11553, ZN => n3584);
   U15213 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_211_port, B1 => n11605, 
                           B2 => n11553, ZN => n3583);
   U15214 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_212_port, B1 => n11606, 
                           B2 => n11553, ZN => n3582);
   U15215 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_213_port, B1 => n11607, 
                           B2 => n11553, ZN => n3581);
   U15216 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_214_port, B1 => n11608, 
                           B2 => n11553, ZN => n3580);
   U15217 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_215_port, B1 => n11609, 
                           B2 => n11553, ZN => n3579);
   U15218 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_216_port, B1 => n11610, 
                           B2 => n11553, ZN => n3578);
   U15219 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_217_port, B1 => n11611, 
                           B2 => n11553, ZN => n3577);
   U15220 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_218_port, B1 => n11612, 
                           B2 => n11553, ZN => n3576);
   U15221 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_219_port, B1 => n11613, 
                           B2 => n11553, ZN => n3575);
   U15222 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_220_port, B1 => n11614, 
                           B2 => n11553, ZN => n3574);
   U15223 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_221_port, B1 => n11615, 
                           B2 => n11553, ZN => n3573);
   U15224 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_222_port, B1 => n11616, 
                           B2 => n11553, ZN => n3572);
   U15225 : AOI22_X1 port map( A1 => n11554, A2 => 
                           DataPath_RF_bus_reg_dataout_223_port, B1 => n11751, 
                           B2 => n11553, ZN => n3569);
   U15226 : OAI22_X1 port map( A1 => n8219, A2 => n11556, B1 => n8529, B2 => 
                           n11555, ZN => n11557);
   U15227 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_160_port, B1 => n11586, 
                           B2 => n11559, ZN => n3564);
   U15228 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_161_port, B1 => n11587, 
                           B2 => n11559, ZN => n3563);
   U15229 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_162_port, B1 => n11588, 
                           B2 => n11559, ZN => n3562);
   U15230 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_163_port, B1 => n11589, 
                           B2 => n11559, ZN => n3561);
   U15231 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_164_port, B1 => n11590, 
                           B2 => n11559, ZN => n3560);
   U15232 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_165_port, B1 => n11591, 
                           B2 => n11559, ZN => n3559);
   U15233 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_166_port, B1 => n11592, 
                           B2 => n11559, ZN => n3558);
   U15234 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_167_port, B1 => n11593, 
                           B2 => n11559, ZN => n3557);
   U15235 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_168_port, B1 => n11594, 
                           B2 => n11559, ZN => n3556);
   U15236 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_169_port, B1 => n11595, 
                           B2 => n11559, ZN => n3555);
   U15237 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_170_port, B1 => n11596, 
                           B2 => n11559, ZN => n3554);
   U15238 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_171_port, B1 => n11597, 
                           B2 => n11559, ZN => n3553);
   U15239 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_172_port, B1 => n11598, 
                           B2 => n11559, ZN => n3552);
   U15240 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_173_port, B1 => n11599, 
                           B2 => n11559, ZN => n3551);
   U15241 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_174_port, B1 => n11600, 
                           B2 => n11559, ZN => n3550);
   U15242 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_175_port, B1 => n11601, 
                           B2 => n11559, ZN => n3549);
   U15243 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_176_port, B1 => n11602, 
                           B2 => n11559, ZN => n3548);
   U15244 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_177_port, B1 => n11603, 
                           B2 => n11559, ZN => n3547);
   U15245 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_178_port, B1 => n11604, 
                           B2 => n11559, ZN => n3546);
   U15246 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_179_port, B1 => n11605, 
                           B2 => n11559, ZN => n3545);
   U15247 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_180_port, B1 => n11606, 
                           B2 => n11559, ZN => n3544);
   U15248 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_181_port, B1 => n11607, 
                           B2 => n11559, ZN => n3543);
   U15249 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_182_port, B1 => n11608, 
                           B2 => n11559, ZN => n3542);
   U15250 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_183_port, B1 => n11609, 
                           B2 => n11559, ZN => n3541);
   U15251 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_184_port, B1 => n11610, 
                           B2 => n11559, ZN => n3540);
   U15252 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_185_port, B1 => n11611, 
                           B2 => n11559, ZN => n3539);
   U15253 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_186_port, B1 => n11612, 
                           B2 => n11559, ZN => n3538);
   U15254 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_187_port, B1 => n11613, 
                           B2 => n11559, ZN => n3537);
   U15255 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_188_port, B1 => n11614, 
                           B2 => n11559, ZN => n3536);
   U15256 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_189_port, B1 => n11615, 
                           B2 => n11559, ZN => n3535);
   U15257 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_190_port, B1 => n11616, 
                           B2 => n11559, ZN => n3534);
   U15258 : AOI22_X1 port map( A1 => n11560, A2 => 
                           DataPath_RF_bus_reg_dataout_191_port, B1 => n11751, 
                           B2 => n11559, ZN => n3531);
   U15259 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_128_port, B1 => n11586, 
                           B2 => n11565, ZN => n3526);
   U15260 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_129_port, B1 => n11587, 
                           B2 => n11565, ZN => n3525);
   U15261 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_130_port, B1 => n11588, 
                           B2 => n11565, ZN => n3524);
   U15262 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_131_port, B1 => n11589, 
                           B2 => n11565, ZN => n3523);
   U15263 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_132_port, B1 => n11590, 
                           B2 => n11565, ZN => n3522);
   U15264 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_133_port, B1 => n11591, 
                           B2 => n11565, ZN => n3521);
   U15265 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_134_port, B1 => n11592, 
                           B2 => n11565, ZN => n3520);
   U15266 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_135_port, B1 => n11593, 
                           B2 => n11565, ZN => n3519);
   U15267 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_136_port, B1 => n11594, 
                           B2 => n11565, ZN => n3518);
   U15268 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_137_port, B1 => n11595, 
                           B2 => n11565, ZN => n3517);
   U15269 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_138_port, B1 => n11596, 
                           B2 => n11565, ZN => n3516);
   U15270 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_139_port, B1 => n11597, 
                           B2 => n11565, ZN => n3515);
   U15271 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_140_port, B1 => n11598, 
                           B2 => n11565, ZN => n3514);
   U15272 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_141_port, B1 => n11599, 
                           B2 => n11565, ZN => n3513);
   U15273 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_142_port, B1 => n11600, 
                           B2 => n11565, ZN => n3512);
   U15274 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_143_port, B1 => n11601, 
                           B2 => n11565, ZN => n3511);
   U15275 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_144_port, B1 => n11602, 
                           B2 => n11565, ZN => n3510);
   U15276 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_145_port, B1 => n11603, 
                           B2 => n11565, ZN => n3509);
   U15277 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_146_port, B1 => n11604, 
                           B2 => n11565, ZN => n3508);
   U15278 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_147_port, B1 => n11605, 
                           B2 => n11565, ZN => n3507);
   U15279 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_148_port, B1 => n11606, 
                           B2 => n11565, ZN => n3506);
   U15280 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_149_port, B1 => n11607, 
                           B2 => n11565, ZN => n3505);
   U15281 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_150_port, B1 => n11608, 
                           B2 => n11565, ZN => n3504);
   U15282 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_151_port, B1 => n11609, 
                           B2 => n11565, ZN => n3503);
   U15283 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_152_port, B1 => n11610, 
                           B2 => n11565, ZN => n3502);
   U15284 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_153_port, B1 => n11611, 
                           B2 => n11565, ZN => n3501);
   U15285 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_154_port, B1 => n11612, 
                           B2 => n11565, ZN => n3500);
   U15286 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_155_port, B1 => n11613, 
                           B2 => n11565, ZN => n3499);
   U15287 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_156_port, B1 => n11614, 
                           B2 => n11565, ZN => n3498);
   U15288 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_157_port, B1 => n11615, 
                           B2 => n11565, ZN => n3497);
   U15289 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_158_port, B1 => n11616, 
                           B2 => n11565, ZN => n3496);
   U15290 : AOI22_X1 port map( A1 => n11566, A2 => 
                           DataPath_RF_bus_reg_dataout_159_port, B1 => n11751, 
                           B2 => n11565, ZN => n3493);
   U15291 : OAI22_X1 port map( A1 => n11586, A2 => n8527, B1 => 
                           DataPath_RF_bus_reg_dataout_96_port, B2 => n11570, 
                           ZN => n3488);
   U15292 : AOI22_X1 port map( A1 => n11587, A2 => n11570, B1 => n8527, B2 => 
                           DataPath_RF_bus_reg_dataout_97_port, ZN => n3487);
   U15293 : OAI22_X1 port map( A1 => n11588, A2 => n8527, B1 => 
                           DataPath_RF_bus_reg_dataout_98_port, B2 => n11570, 
                           ZN => n3486);
   U15294 : AOI22_X1 port map( A1 => n11589, A2 => n11570, B1 => n8527, B2 => 
                           DataPath_RF_bus_reg_dataout_99_port, ZN => n3485);
   U15295 : AOI22_X1 port map( A1 => n11590, A2 => n11570, B1 => n11571, B2 => 
                           DataPath_RF_bus_reg_dataout_100_port, ZN => n3484);
   U15296 : OAI22_X1 port map( A1 => n11591, A2 => n11571, B1 => 
                           DataPath_RF_bus_reg_dataout_101_port, B2 => n11570, 
                           ZN => n3483);
   U15297 : AOI22_X1 port map( A1 => n11592, A2 => n11570, B1 => n8527, B2 => 
                           DataPath_RF_bus_reg_dataout_102_port, ZN => n3482);
   U15298 : OAI22_X1 port map( A1 => n11593, A2 => n11571, B1 => 
                           DataPath_RF_bus_reg_dataout_103_port, B2 => n11570, 
                           ZN => n3481);
   U15299 : OAI22_X1 port map( A1 => n11594, A2 => n8527, B1 => 
                           DataPath_RF_bus_reg_dataout_104_port, B2 => n11570, 
                           ZN => n3480);
   U15300 : AOI22_X1 port map( A1 => n11595, A2 => n11570, B1 => n11571, B2 => 
                           DataPath_RF_bus_reg_dataout_105_port, ZN => n3479);
   U15301 : OAI22_X1 port map( A1 => n11596, A2 => n8527, B1 => 
                           DataPath_RF_bus_reg_dataout_106_port, B2 => n11570, 
                           ZN => n3478);
   U15302 : AOI22_X1 port map( A1 => n11597, A2 => n11570, B1 => n8527, B2 => 
                           DataPath_RF_bus_reg_dataout_107_port, ZN => n3477);
   U15303 : AOI22_X1 port map( A1 => n11598, A2 => n11570, B1 => n8527, B2 => 
                           DataPath_RF_bus_reg_dataout_108_port, ZN => n3476);
   U15304 : AOI22_X1 port map( A1 => n11599, A2 => n11570, B1 => n8527, B2 => 
                           DataPath_RF_bus_reg_dataout_109_port, ZN => n3475);
   U15305 : OAI22_X1 port map( A1 => n11600, A2 => n8527, B1 => 
                           DataPath_RF_bus_reg_dataout_110_port, B2 => n11570, 
                           ZN => n3474);
   U15306 : AOI22_X1 port map( A1 => n11601, A2 => n11570, B1 => n8527, B2 => 
                           DataPath_RF_bus_reg_dataout_111_port, ZN => n3473);
   U15307 : OAI22_X1 port map( A1 => n11571, A2 => n11602, B1 => 
                           DataPath_RF_bus_reg_dataout_112_port, B2 => n11570, 
                           ZN => n3472);
   U15308 : OAI22_X1 port map( A1 => n8527, A2 => n11603, B1 => 
                           DataPath_RF_bus_reg_dataout_113_port, B2 => n11570, 
                           ZN => n3471);
   U15309 : OAI22_X1 port map( A1 => n11604, A2 => n8527, B1 => 
                           DataPath_RF_bus_reg_dataout_114_port, B2 => n11570, 
                           ZN => n3470);
   U15310 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_115_port, A2 
                           => n8527, B1 => n11605, B2 => n11570, ZN => n3469);
   U15311 : OAI22_X1 port map( A1 => n11571, A2 => n11606, B1 => 
                           DataPath_RF_bus_reg_dataout_116_port, B2 => n11570, 
                           ZN => n3468);
   U15312 : OAI22_X1 port map( A1 => n11607, A2 => n8527, B1 => 
                           DataPath_RF_bus_reg_dataout_117_port, B2 => n11570, 
                           ZN => n3467);
   U15313 : AOI22_X1 port map( A1 => n11608, A2 => n11570, B1 => n11571, B2 => 
                           DataPath_RF_bus_reg_dataout_118_port, ZN => n3466);
   U15314 : OAI22_X1 port map( A1 => n11609, A2 => n8527, B1 => 
                           DataPath_RF_bus_reg_dataout_119_port, B2 => n11570, 
                           ZN => n3465);
   U15315 : AOI22_X1 port map( A1 => n11610, A2 => n11570, B1 => n8527, B2 => 
                           DataPath_RF_bus_reg_dataout_120_port, ZN => n3464);
   U15316 : AOI22_X1 port map( A1 => n11611, A2 => n11570, B1 => n11571, B2 => 
                           DataPath_RF_bus_reg_dataout_121_port, ZN => n3463);
   U15317 : AOI22_X1 port map( A1 => n11612, A2 => n11570, B1 => n8527, B2 => 
                           DataPath_RF_bus_reg_dataout_122_port, ZN => n3462);
   U15318 : OAI22_X1 port map( A1 => n8527, A2 => n11613, B1 => 
                           DataPath_RF_bus_reg_dataout_123_port, B2 => n11570, 
                           ZN => n3461);
   U15319 : OAI22_X1 port map( A1 => n11571, A2 => n11614, B1 => 
                           DataPath_RF_bus_reg_dataout_124_port, B2 => n11570, 
                           ZN => n3460);
   U15320 : AOI22_X1 port map( A1 => n11615, A2 => n11570, B1 => n11571, B2 => 
                           DataPath_RF_bus_reg_dataout_125_port, ZN => n3459);
   U15321 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_126_port, A2 
                           => n8527, B1 => n11616, B2 => n11570, ZN => n3458);
   U15322 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_127_port, A2 
                           => n8527, B1 => n11751, B2 => n11570, ZN => n3455);
   U15323 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_64_port, B1 => n11586, 
                           B2 => n11576, ZN => n3450);
   U15324 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_65_port, B1 => n11587, 
                           B2 => n11576, ZN => n3449);
   U15325 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_66_port, B1 => n11588, 
                           B2 => n11576, ZN => n3448);
   U15326 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_67_port, B1 => n11589, 
                           B2 => n11576, ZN => n3447);
   U15327 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_68_port, B1 => n11590, 
                           B2 => n11576, ZN => n3446);
   U15328 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_69_port, B1 => n11591, 
                           B2 => n11576, ZN => n3445);
   U15329 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_70_port, B1 => n11592, 
                           B2 => n11576, ZN => n3444);
   U15330 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_71_port, B1 => n11593, 
                           B2 => n11576, ZN => n3443);
   U15331 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_72_port, B1 => n11594, 
                           B2 => n11576, ZN => n3442);
   U15332 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_73_port, B1 => n11595, 
                           B2 => n11576, ZN => n3441);
   U15333 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_74_port, B1 => n11596, 
                           B2 => n11576, ZN => n3440);
   U15334 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_75_port, B1 => n11597, 
                           B2 => n11576, ZN => n3439);
   U15335 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_76_port, B1 => n11598, 
                           B2 => n11576, ZN => n3438);
   U15336 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_77_port, B1 => n11599, 
                           B2 => n11576, ZN => n3437);
   U15337 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_78_port, B1 => n11600, 
                           B2 => n11576, ZN => n3436);
   U15338 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_79_port, B1 => n11601, 
                           B2 => n11576, ZN => n3435);
   U15339 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_80_port, B1 => n11602, 
                           B2 => n11576, ZN => n3434);
   U15340 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_81_port, B1 => n11603, 
                           B2 => n11576, ZN => n3433);
   U15341 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_82_port, B1 => n11604, 
                           B2 => n11576, ZN => n3432);
   U15342 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_83_port, B1 => n11605, 
                           B2 => n11576, ZN => n3431);
   U15343 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_84_port, B1 => n11606, 
                           B2 => n11576, ZN => n3430);
   U15344 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_85_port, B1 => n11607, 
                           B2 => n11576, ZN => n3429);
   U15345 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_86_port, B1 => n11608, 
                           B2 => n11576, ZN => n3428);
   U15346 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_87_port, B1 => n11609, 
                           B2 => n11576, ZN => n3427);
   U15347 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_88_port, B1 => n11610, 
                           B2 => n11576, ZN => n3426);
   U15348 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_89_port, B1 => n11611, 
                           B2 => n11576, ZN => n3425);
   U15349 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_90_port, B1 => n11612, 
                           B2 => n11576, ZN => n3424);
   U15350 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_91_port, B1 => n11613, 
                           B2 => n11576, ZN => n3423);
   U15351 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_92_port, B1 => n11614, 
                           B2 => n11576, ZN => n3422);
   U15352 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_93_port, B1 => n11615, 
                           B2 => n11576, ZN => n3421);
   U15353 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_94_port, B1 => n11616, 
                           B2 => n11576, ZN => n3420);
   U15354 : AOI22_X1 port map( A1 => n11577, A2 => 
                           DataPath_RF_bus_reg_dataout_95_port, B1 => n11751, 
                           B2 => n11576, ZN => n3417);
   U15355 : AOI211_X1 port map( C1 => n8296, C2 => n11581, A => RST, B => 
                           n11580, ZN => n11582);
   U15356 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_32_port, B1 => n11586, 
                           B2 => n8528, ZN => n3412);
   U15357 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_33_port, B1 => n11587, 
                           B2 => n8528, ZN => n3411);
   U15358 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_34_port, B1 => n11588, 
                           B2 => n8528, ZN => n3410);
   U15359 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_35_port, B1 => n11589, 
                           B2 => n8528, ZN => n3409);
   U15360 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_36_port, B1 => n11590, 
                           B2 => n8528, ZN => n3408);
   U15361 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_37_port, B1 => n11591, 
                           B2 => n8528, ZN => n3407);
   U15362 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_38_port, B1 => n11592, 
                           B2 => n8528, ZN => n3406);
   U15363 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_39_port, B1 => n11593, 
                           B2 => n8528, ZN => n3405);
   U15364 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_40_port, B1 => n11594, 
                           B2 => n8528, ZN => n3404);
   U15365 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_41_port, B1 => n11595, 
                           B2 => n8528, ZN => n3403);
   U15366 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_42_port, B1 => n11596, 
                           B2 => n8528, ZN => n3402);
   U15367 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_43_port, B1 => n11597, 
                           B2 => n8528, ZN => n3401);
   U15368 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_44_port, B1 => n11598, 
                           B2 => n8528, ZN => n3400);
   U15369 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_45_port, B1 => n11599, 
                           B2 => n8528, ZN => n3399);
   U15370 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_46_port, B1 => n11600, 
                           B2 => n8528, ZN => n3398);
   U15371 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_47_port, B1 => n11601, 
                           B2 => n8528, ZN => n3397);
   U15372 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_48_port, B1 => n11602, 
                           B2 => n8528, ZN => n3396);
   U15373 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_49_port, B1 => n11603, 
                           B2 => n8528, ZN => n3395);
   U15374 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_50_port, B1 => n11604, 
                           B2 => n8528, ZN => n3394);
   U15375 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_51_port, B1 => n11605, 
                           B2 => n8528, ZN => n3393);
   U15376 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_52_port, B1 => n11606, 
                           B2 => n8528, ZN => n3392);
   U15377 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_53_port, B1 => n11607, 
                           B2 => n8528, ZN => n3391);
   U15378 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_54_port, B1 => n11608, 
                           B2 => n8528, ZN => n3390);
   U15379 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_55_port, B1 => n11609, 
                           B2 => n8528, ZN => n3389);
   U15380 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_56_port, B1 => n11610, 
                           B2 => n8528, ZN => n3388);
   U15381 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_57_port, B1 => n11611, 
                           B2 => n8528, ZN => n3387);
   U15382 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_58_port, B1 => n11612, 
                           B2 => n8528, ZN => n3386);
   U15383 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_59_port, B1 => n11613, 
                           B2 => n8528, ZN => n3385);
   U15384 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_60_port, B1 => n11614, 
                           B2 => n8528, ZN => n3384);
   U15385 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_61_port, B1 => n11615, 
                           B2 => n8528, ZN => n3383);
   U15386 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_62_port, B1 => n11616, 
                           B2 => n8528, ZN => n3382);
   U15387 : AOI22_X1 port map( A1 => n7764, A2 => 
                           DataPath_RF_bus_reg_dataout_63_port, B1 => n11751, 
                           B2 => n8528, ZN => n3379);
   U15388 : OAI22_X1 port map( A1 => n11586, A2 => n8540, B1 => 
                           DataPath_RF_bus_reg_dataout_0_port, B2 => n7765, ZN 
                           => n3372);
   U15389 : OAI22_X1 port map( A1 => n11587, A2 => n8540, B1 => 
                           DataPath_RF_bus_reg_dataout_1_port, B2 => n7765, ZN 
                           => n3370);
   U15390 : OAI22_X1 port map( A1 => n11588, A2 => n8540, B1 => 
                           DataPath_RF_bus_reg_dataout_2_port, B2 => n7765, ZN 
                           => n3368);
   U15391 : OAI22_X1 port map( A1 => n11589, A2 => n8540, B1 => 
                           DataPath_RF_bus_reg_dataout_3_port, B2 => n7765, ZN 
                           => n3366);
   U15392 : AOI22_X1 port map( A1 => n11590, A2 => n7765, B1 => n8540, B2 => 
                           DataPath_RF_bus_reg_dataout_4_port, ZN => n3364);
   U15393 : AOI22_X1 port map( A1 => n11591, A2 => n7765, B1 => n8540, B2 => 
                           DataPath_RF_bus_reg_dataout_5_port, ZN => n3362);
   U15394 : AOI22_X1 port map( A1 => n11592, A2 => n7765, B1 => n11752, B2 => 
                           DataPath_RF_bus_reg_dataout_6_port, ZN => n3360);
   U15395 : OAI22_X1 port map( A1 => n11593, A2 => n8540, B1 => 
                           DataPath_RF_bus_reg_dataout_7_port, B2 => n7765, ZN 
                           => n3358);
   U15396 : OAI22_X1 port map( A1 => n11594, A2 => n8540, B1 => 
                           DataPath_RF_bus_reg_dataout_8_port, B2 => n7765, ZN 
                           => n3356);
   U15397 : AOI22_X1 port map( A1 => n11595, A2 => n7765, B1 => n8540, B2 => 
                           DataPath_RF_bus_reg_dataout_9_port, ZN => n3354);
   U15398 : OAI22_X1 port map( A1 => n11596, A2 => n8540, B1 => 
                           DataPath_RF_bus_reg_dataout_10_port, B2 => n7765, ZN
                           => n3352);
   U15399 : OAI22_X1 port map( A1 => n11597, A2 => n8540, B1 => 
                           DataPath_RF_bus_reg_dataout_11_port, B2 => n7765, ZN
                           => n3350);
   U15400 : AOI22_X1 port map( A1 => n11598, A2 => n7765, B1 => n11752, B2 => 
                           DataPath_RF_bus_reg_dataout_12_port, ZN => n3348);
   U15401 : AOI22_X1 port map( A1 => n11599, A2 => n7765, B1 => n11752, B2 => 
                           DataPath_RF_bus_reg_dataout_13_port, ZN => n3346);
   U15402 : AOI22_X1 port map( A1 => n11600, A2 => n7765, B1 => n11752, B2 => 
                           DataPath_RF_bus_reg_dataout_14_port, ZN => n3344);
   U15403 : AOI22_X1 port map( A1 => n11601, A2 => n7765, B1 => n8540, B2 => 
                           DataPath_RF_bus_reg_dataout_15_port, ZN => n3342);
   U15404 : OAI22_X1 port map( A1 => n8540, A2 => n11602, B1 => 
                           DataPath_RF_bus_reg_dataout_16_port, B2 => n7765, ZN
                           => n3340);
   U15405 : OAI22_X1 port map( A1 => n8540, A2 => n11603, B1 => 
                           DataPath_RF_bus_reg_dataout_17_port, B2 => n7765, ZN
                           => n3338);
   U15406 : AOI22_X1 port map( A1 => n11604, A2 => n7765, B1 => n11752, B2 => 
                           DataPath_RF_bus_reg_dataout_18_port, ZN => n3336);
   U15407 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_19_port, A2 =>
                           n11752, B1 => n11605, B2 => n7765, ZN => n3334);
   U15408 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_20_port, A2 =>
                           n8540, B1 => n11606, B2 => n7765, ZN => n3332);
   U15409 : OAI22_X1 port map( A1 => n11607, A2 => n8540, B1 => 
                           DataPath_RF_bus_reg_dataout_21_port, B2 => n7765, ZN
                           => n3330);
   U15410 : OAI22_X1 port map( A1 => n11608, A2 => n8540, B1 => 
                           DataPath_RF_bus_reg_dataout_22_port, B2 => n7765, ZN
                           => n3328);
   U15411 : AOI22_X1 port map( A1 => n11609, A2 => n7765, B1 => n8540, B2 => 
                           DataPath_RF_bus_reg_dataout_23_port, ZN => n3326);
   U15412 : OAI22_X1 port map( A1 => n11610, A2 => n8540, B1 => 
                           DataPath_RF_bus_reg_dataout_24_port, B2 => n7765, ZN
                           => n3324);
   U15413 : OAI22_X1 port map( A1 => n11611, A2 => n8540, B1 => 
                           DataPath_RF_bus_reg_dataout_25_port, B2 => n7765, ZN
                           => n3322);
   U15414 : AOI22_X1 port map( A1 => n11612, A2 => n7765, B1 => n8540, B2 => 
                           DataPath_RF_bus_reg_dataout_26_port, ZN => n3320);
   U15415 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_27_port, A2 =>
                           n11752, B1 => n11613, B2 => n7765, ZN => n3318);
   U15416 : OAI22_X1 port map( A1 => n8540, A2 => n11614, B1 => 
                           DataPath_RF_bus_reg_dataout_28_port, B2 => n7765, ZN
                           => n3316);
   U15417 : OAI22_X1 port map( A1 => n11615, A2 => n11752, B1 => 
                           DataPath_RF_bus_reg_dataout_29_port, B2 => n7765, ZN
                           => n3314);
   U15418 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_30_port, A2 =>
                           n11752, B1 => n11616, B2 => n7765, ZN => n3312);
   U15419 : NAND2_X1 port map( A1 => n11617, A2 => n11642, ZN => n11618);
   U15420 : OAI22_X1 port map( A1 => n11645, A2 => n11620, B1 => n791, B2 => 
                           n11619, ZN => n6991);
   U15421 : OAI22_X1 port map( A1 => n11646, A2 => n11620, B1 => n792, B2 => 
                           n11619, ZN => n6990);
   U15422 : OAI22_X1 port map( A1 => n11647, A2 => n11620, B1 => n793, B2 => 
                           n11619, ZN => n6989);
   U15423 : OAI22_X1 port map( A1 => n11648, A2 => n11620, B1 => n794, B2 => 
                           n11619, ZN => n6988);
   U15424 : OAI22_X1 port map( A1 => n11649, A2 => n11620, B1 => n795, B2 => 
                           n11619, ZN => n6987);
   U15425 : OAI22_X1 port map( A1 => n11650, A2 => n11620, B1 => n796, B2 => 
                           n11619, ZN => n6986);
   U15426 : OAI22_X1 port map( A1 => n11651, A2 => n11620, B1 => n797, B2 => 
                           n11619, ZN => n6985);
   U15427 : OAI22_X1 port map( A1 => n11652, A2 => n11620, B1 => n798, B2 => 
                           n11619, ZN => n6984);
   U15428 : OAI22_X1 port map( A1 => n11653, A2 => n11620, B1 => n799, B2 => 
                           n11619, ZN => n6983);
   U15429 : OAI22_X1 port map( A1 => n11654, A2 => n11620, B1 => n800, B2 => 
                           n11619, ZN => n6982);
   U15430 : OAI22_X1 port map( A1 => n11655, A2 => n8530, B1 => n801, B2 => 
                           n11619, ZN => n6981);
   U15431 : OAI22_X1 port map( A1 => n11656, A2 => n8530, B1 => n802, B2 => 
                           n11619, ZN => n6980);
   U15432 : OAI22_X1 port map( A1 => n11657, A2 => n8530, B1 => n803, B2 => 
                           n11619, ZN => n6979);
   U15433 : OAI22_X1 port map( A1 => n11658, A2 => n8530, B1 => n804, B2 => 
                           n11619, ZN => n6978);
   U15434 : OAI22_X1 port map( A1 => n11659, A2 => n8530, B1 => n805, B2 => 
                           n11619, ZN => n6977);
   U15435 : OAI22_X1 port map( A1 => n11660, A2 => n8530, B1 => n806, B2 => 
                           n11619, ZN => n6976);
   U15436 : OAI22_X1 port map( A1 => n11661, A2 => n8530, B1 => n807, B2 => 
                           n11619, ZN => n6975);
   U15437 : OAI22_X1 port map( A1 => n11662, A2 => n8530, B1 => n808, B2 => 
                           n11619, ZN => n6974);
   U15438 : OAI22_X1 port map( A1 => n11663, A2 => n8530, B1 => n809, B2 => 
                           n11619, ZN => n6973);
   U15439 : OAI22_X1 port map( A1 => n11664, A2 => n8530, B1 => n810, B2 => 
                           n11619, ZN => n6972);
   U15440 : OAI22_X1 port map( A1 => n11665, A2 => n8530, B1 => n811, B2 => 
                           n11619, ZN => n6971);
   U15441 : OAI22_X1 port map( A1 => n11666, A2 => n8530, B1 => n812, B2 => 
                           n11619, ZN => n6970);
   U15442 : OAI22_X1 port map( A1 => n11667, A2 => n11620, B1 => n813, B2 => 
                           n11619, ZN => n6969);
   U15443 : OAI22_X1 port map( A1 => n11668, A2 => n11620, B1 => n814, B2 => 
                           n11619, ZN => n6968);
   U15444 : OAI22_X1 port map( A1 => n11669, A2 => n11620, B1 => n815, B2 => 
                           n11619, ZN => n6967);
   U15445 : OAI22_X1 port map( A1 => n11670, A2 => n11620, B1 => n816, B2 => 
                           n11619, ZN => n6966);
   U15446 : OAI22_X1 port map( A1 => n11671, A2 => n11620, B1 => n817, B2 => 
                           n11619, ZN => n6965);
   U15447 : OAI22_X1 port map( A1 => n11672, A2 => n8530, B1 => n818, B2 => 
                           n11619, ZN => n6964);
   U15448 : OAI22_X1 port map( A1 => n11673, A2 => n8530, B1 => n819, B2 => 
                           n11619, ZN => n6963);
   U15449 : OAI22_X1 port map( A1 => n11674, A2 => n8530, B1 => n820, B2 => 
                           n11619, ZN => n6962);
   U15450 : OAI22_X1 port map( A1 => n11675, A2 => n8530, B1 => n821, B2 => 
                           n11619, ZN => n6961);
   U15451 : OAI22_X1 port map( A1 => n11678, A2 => n8530, B1 => n822, B2 => 
                           n11619, ZN => n6960);
   U15452 : INV_X1 port map( A => n11621, ZN => n11622);
   U15453 : INV_X1 port map( A => n11642, ZN => n11634);
   U15454 : OAI22_X1 port map( A1 => n11645, A2 => n11624, B1 => n759, B2 => 
                           n8531, ZN => n6959);
   U15455 : OAI22_X1 port map( A1 => n11646, A2 => n11624, B1 => n760, B2 => 
                           n8531, ZN => n6958);
   U15456 : OAI22_X1 port map( A1 => n11647, A2 => n11624, B1 => n761, B2 => 
                           n8531, ZN => n6957);
   U15457 : OAI22_X1 port map( A1 => n11648, A2 => n11624, B1 => n762, B2 => 
                           n8531, ZN => n6956);
   U15458 : OAI22_X1 port map( A1 => n11649, A2 => n11624, B1 => n763, B2 => 
                           n11623, ZN => n6955);
   U15459 : OAI22_X1 port map( A1 => n11650, A2 => n11624, B1 => n764, B2 => 
                           n11623, ZN => n6954);
   U15460 : OAI22_X1 port map( A1 => n11651, A2 => n11624, B1 => n765, B2 => 
                           n11623, ZN => n6953);
   U15461 : OAI22_X1 port map( A1 => n11652, A2 => n11624, B1 => n766, B2 => 
                           n11623, ZN => n6952);
   U15462 : OAI22_X1 port map( A1 => n11653, A2 => n11624, B1 => n767, B2 => 
                           n11623, ZN => n6951);
   U15463 : OAI22_X1 port map( A1 => n11654, A2 => n11624, B1 => n768, B2 => 
                           n8531, ZN => n6950);
   U15464 : OAI22_X1 port map( A1 => n11655, A2 => n8532, B1 => n769, B2 => 
                           n8531, ZN => n6949);
   U15465 : OAI22_X1 port map( A1 => n11656, A2 => n8532, B1 => n770, B2 => 
                           n8531, ZN => n6948);
   U15466 : OAI22_X1 port map( A1 => n11657, A2 => n8532, B1 => n771, B2 => 
                           n8531, ZN => n6947);
   U15467 : OAI22_X1 port map( A1 => n11658, A2 => n8532, B1 => n772, B2 => 
                           n8531, ZN => n6946);
   U15468 : OAI22_X1 port map( A1 => n11659, A2 => n8532, B1 => n773, B2 => 
                           n8531, ZN => n6945);
   U15469 : OAI22_X1 port map( A1 => n11660, A2 => n8532, B1 => n774, B2 => 
                           n8531, ZN => n6944);
   U15470 : OAI22_X1 port map( A1 => n11661, A2 => n8532, B1 => n775, B2 => 
                           n8531, ZN => n6943);
   U15471 : OAI22_X1 port map( A1 => n11662, A2 => n8532, B1 => n776, B2 => 
                           n8531, ZN => n6942);
   U15472 : OAI22_X1 port map( A1 => n11663, A2 => n8532, B1 => n777, B2 => 
                           n8531, ZN => n6941);
   U15473 : OAI22_X1 port map( A1 => n11664, A2 => n8532, B1 => n778, B2 => 
                           n8531, ZN => n6940);
   U15474 : OAI22_X1 port map( A1 => n11665, A2 => n8532, B1 => n779, B2 => 
                           n8531, ZN => n6939);
   U15475 : OAI22_X1 port map( A1 => n11666, A2 => n8532, B1 => n780, B2 => 
                           n8531, ZN => n6938);
   U15476 : OAI22_X1 port map( A1 => n11667, A2 => n11624, B1 => n781, B2 => 
                           n8531, ZN => n6937);
   U15477 : OAI22_X1 port map( A1 => n11668, A2 => n11624, B1 => n782, B2 => 
                           n11623, ZN => n6936);
   U15478 : OAI22_X1 port map( A1 => n11669, A2 => n11624, B1 => n783, B2 => 
                           n8531, ZN => n6935);
   U15479 : OAI22_X1 port map( A1 => n11670, A2 => n11624, B1 => n784, B2 => 
                           n8531, ZN => n6934);
   U15480 : OAI22_X1 port map( A1 => n11671, A2 => n11624, B1 => n785, B2 => 
                           n8531, ZN => n6933);
   U15481 : OAI22_X1 port map( A1 => n11672, A2 => n8532, B1 => n786, B2 => 
                           n11623, ZN => n6932);
   U15482 : OAI22_X1 port map( A1 => n11673, A2 => n8532, B1 => n787, B2 => 
                           n11623, ZN => n6931);
   U15483 : OAI22_X1 port map( A1 => n11674, A2 => n8532, B1 => n788, B2 => 
                           n11623, ZN => n6930);
   U15484 : OAI22_X1 port map( A1 => n11675, A2 => n8532, B1 => n789, B2 => 
                           n8531, ZN => n6929);
   U15485 : OAI22_X1 port map( A1 => n11678, A2 => n8532, B1 => n790, B2 => 
                           n11623, ZN => n6928);
   U15486 : NAND2_X1 port map( A1 => n11625, A2 => n11642, ZN => n11626);
   U15487 : OAI22_X1 port map( A1 => n11645, A2 => n11628, B1 => n727, B2 => 
                           n11627, ZN => n6927);
   U15488 : OAI22_X1 port map( A1 => n11646, A2 => n11628, B1 => n728, B2 => 
                           n11627, ZN => n6926);
   U15489 : OAI22_X1 port map( A1 => n11647, A2 => n11628, B1 => n729, B2 => 
                           n11627, ZN => n6925);
   U15490 : OAI22_X1 port map( A1 => n11648, A2 => n11628, B1 => n730, B2 => 
                           n11627, ZN => n6924);
   U15491 : OAI22_X1 port map( A1 => n11649, A2 => n11628, B1 => n731, B2 => 
                           n11627, ZN => n6923);
   U15492 : OAI22_X1 port map( A1 => n11650, A2 => n11628, B1 => n732, B2 => 
                           n11627, ZN => n6922);
   U15493 : OAI22_X1 port map( A1 => n11651, A2 => n11628, B1 => n733, B2 => 
                           n11627, ZN => n6921);
   U15494 : OAI22_X1 port map( A1 => n11652, A2 => n11628, B1 => n734, B2 => 
                           n11627, ZN => n6920);
   U15495 : OAI22_X1 port map( A1 => n11653, A2 => n11628, B1 => n735, B2 => 
                           n11627, ZN => n6919);
   U15496 : OAI22_X1 port map( A1 => n11654, A2 => n11628, B1 => n736, B2 => 
                           n11627, ZN => n6918);
   U15497 : OAI22_X1 port map( A1 => n11655, A2 => n11628, B1 => n737, B2 => 
                           n11627, ZN => n6917);
   U15498 : OAI22_X1 port map( A1 => n11656, A2 => n8533, B1 => n738, B2 => 
                           n11627, ZN => n6916);
   U15499 : OAI22_X1 port map( A1 => n11657, A2 => n8533, B1 => n739, B2 => 
                           n11627, ZN => n6915);
   U15500 : OAI22_X1 port map( A1 => n11658, A2 => n8533, B1 => n740, B2 => 
                           n11627, ZN => n6914);
   U15501 : OAI22_X1 port map( A1 => n11659, A2 => n8533, B1 => n741, B2 => 
                           n11627, ZN => n6913);
   U15502 : OAI22_X1 port map( A1 => n11660, A2 => n8533, B1 => n742, B2 => 
                           n11627, ZN => n6912);
   U15503 : OAI22_X1 port map( A1 => n11661, A2 => n8533, B1 => n743, B2 => 
                           n11627, ZN => n6911);
   U15504 : OAI22_X1 port map( A1 => n11662, A2 => n8533, B1 => n744, B2 => 
                           n11627, ZN => n6910);
   U15505 : OAI22_X1 port map( A1 => n11663, A2 => n8533, B1 => n745, B2 => 
                           n11627, ZN => n6909);
   U15506 : OAI22_X1 port map( A1 => n11664, A2 => n8533, B1 => n746, B2 => 
                           n11627, ZN => n6908);
   U15507 : OAI22_X1 port map( A1 => n11665, A2 => n8533, B1 => n747, B2 => 
                           n11627, ZN => n6907);
   U15508 : OAI22_X1 port map( A1 => n11666, A2 => n8533, B1 => n748, B2 => 
                           n11627, ZN => n6906);
   U15509 : OAI22_X1 port map( A1 => n11667, A2 => n11628, B1 => n749, B2 => 
                           n11627, ZN => n6905);
   U15510 : OAI22_X1 port map( A1 => n11668, A2 => n11628, B1 => n750, B2 => 
                           n11627, ZN => n6904);
   U15511 : OAI22_X1 port map( A1 => n11669, A2 => n11628, B1 => n751, B2 => 
                           n11627, ZN => n6903);
   U15512 : OAI22_X1 port map( A1 => n11670, A2 => n11628, B1 => n752, B2 => 
                           n11627, ZN => n6902);
   U15513 : OAI22_X1 port map( A1 => n11671, A2 => n11628, B1 => n753, B2 => 
                           n11627, ZN => n6901);
   U15514 : OAI22_X1 port map( A1 => n11672, A2 => n8533, B1 => n754, B2 => 
                           n11627, ZN => n6900);
   U15515 : OAI22_X1 port map( A1 => n11673, A2 => n8533, B1 => n755, B2 => 
                           n11627, ZN => n6899);
   U15516 : OAI22_X1 port map( A1 => n11674, A2 => n8533, B1 => n756, B2 => 
                           n11627, ZN => n6898);
   U15517 : OAI22_X1 port map( A1 => n11675, A2 => n8533, B1 => n757, B2 => 
                           n11627, ZN => n6897);
   U15518 : OAI22_X1 port map( A1 => n11678, A2 => n8533, B1 => n758, B2 => 
                           n11627, ZN => n6896);
   U15519 : OAI22_X1 port map( A1 => n11645, A2 => n11632, B1 => n695, B2 => 
                           n8534, ZN => n6895);
   U15520 : OAI22_X1 port map( A1 => n11646, A2 => n11632, B1 => n696, B2 => 
                           n8534, ZN => n6894);
   U15521 : OAI22_X1 port map( A1 => n11647, A2 => n11632, B1 => n697, B2 => 
                           n8534, ZN => n6893);
   U15522 : OAI22_X1 port map( A1 => n11648, A2 => n11632, B1 => n698, B2 => 
                           n8534, ZN => n6892);
   U15523 : OAI22_X1 port map( A1 => n11649, A2 => n11632, B1 => n699, B2 => 
                           n8534, ZN => n6891);
   U15524 : OAI22_X1 port map( A1 => n11650, A2 => n11632, B1 => n700, B2 => 
                           n8534, ZN => n6890);
   U15525 : OAI22_X1 port map( A1 => n11651, A2 => n11632, B1 => n701, B2 => 
                           n8534, ZN => n6889);
   U15526 : OAI22_X1 port map( A1 => n11652, A2 => n11632, B1 => n702, B2 => 
                           n8534, ZN => n6888);
   U15527 : OAI22_X1 port map( A1 => n11653, A2 => n11632, B1 => n703, B2 => 
                           n8534, ZN => n6887);
   U15528 : OAI22_X1 port map( A1 => n11654, A2 => n11632, B1 => n704, B2 => 
                           n8534, ZN => n6886);
   U15529 : OAI22_X1 port map( A1 => n11655, A2 => n11632, B1 => n705, B2 => 
                           n8534, ZN => n6885);
   U15530 : OAI22_X1 port map( A1 => n11656, A2 => n8535, B1 => n706, B2 => 
                           n8534, ZN => n6884);
   U15531 : OAI22_X1 port map( A1 => n11657, A2 => n8535, B1 => n707, B2 => 
                           n8534, ZN => n6883);
   U15532 : OAI22_X1 port map( A1 => n11658, A2 => n8535, B1 => n708, B2 => 
                           n8534, ZN => n6882);
   U15533 : OAI22_X1 port map( A1 => n11659, A2 => n8535, B1 => n709, B2 => 
                           n8534, ZN => n6881);
   U15534 : OAI22_X1 port map( A1 => n11660, A2 => n8535, B1 => n710, B2 => 
                           n8534, ZN => n6880);
   U15535 : OAI22_X1 port map( A1 => n11661, A2 => n8535, B1 => n711, B2 => 
                           n11631, ZN => n6879);
   U15536 : OAI22_X1 port map( A1 => n11662, A2 => n8535, B1 => n712, B2 => 
                           n11631, ZN => n6878);
   U15537 : OAI22_X1 port map( A1 => n11663, A2 => n8535, B1 => n713, B2 => 
                           n11631, ZN => n6877);
   U15538 : OAI22_X1 port map( A1 => n11664, A2 => n8535, B1 => n714, B2 => 
                           n11631, ZN => n6876);
   U15539 : OAI22_X1 port map( A1 => n11665, A2 => n8535, B1 => n715, B2 => 
                           n11631, ZN => n6875);
   U15540 : OAI22_X1 port map( A1 => n11666, A2 => n8535, B1 => n716, B2 => 
                           n8534, ZN => n6874);
   U15541 : OAI22_X1 port map( A1 => n11667, A2 => n11632, B1 => n717, B2 => 
                           n11631, ZN => n6873);
   U15542 : OAI22_X1 port map( A1 => n11668, A2 => n11632, B1 => n718, B2 => 
                           n8534, ZN => n6872);
   U15543 : OAI22_X1 port map( A1 => n11669, A2 => n11632, B1 => n719, B2 => 
                           n11631, ZN => n6871);
   U15544 : OAI22_X1 port map( A1 => n11670, A2 => n11632, B1 => n720, B2 => 
                           n8534, ZN => n6870);
   U15545 : OAI22_X1 port map( A1 => n11671, A2 => n11632, B1 => n721, B2 => 
                           n8534, ZN => n6869);
   U15546 : OAI22_X1 port map( A1 => n11672, A2 => n8535, B1 => n722, B2 => 
                           n11631, ZN => n6868);
   U15547 : OAI22_X1 port map( A1 => n11673, A2 => n8535, B1 => n723, B2 => 
                           n11631, ZN => n6867);
   U15548 : OAI22_X1 port map( A1 => n11674, A2 => n8535, B1 => n724, B2 => 
                           n8534, ZN => n6866);
   U15549 : OAI22_X1 port map( A1 => n11675, A2 => n8535, B1 => n725, B2 => 
                           n11631, ZN => n6865);
   U15550 : OAI22_X1 port map( A1 => n11678, A2 => n8535, B1 => n726, B2 => 
                           n8534, ZN => n6864);
   U15551 : INV_X1 port map( A => n11633, ZN => n11635);
   U15552 : OAI22_X1 port map( A1 => n11645, A2 => n11637, B1 => n663, B2 => 
                           n8536, ZN => n6863);
   U15553 : OAI22_X1 port map( A1 => n11646, A2 => n11637, B1 => n664, B2 => 
                           n8536, ZN => n6862);
   U15554 : OAI22_X1 port map( A1 => n11647, A2 => n11637, B1 => n665, B2 => 
                           n8536, ZN => n6861);
   U15555 : OAI22_X1 port map( A1 => n11648, A2 => n11637, B1 => n666, B2 => 
                           n8536, ZN => n6860);
   U15556 : OAI22_X1 port map( A1 => n11649, A2 => n11637, B1 => n667, B2 => 
                           n11636, ZN => n6859);
   U15557 : OAI22_X1 port map( A1 => n11650, A2 => n11637, B1 => n668, B2 => 
                           n11636, ZN => n6858);
   U15558 : OAI22_X1 port map( A1 => n11651, A2 => n11637, B1 => n669, B2 => 
                           n11636, ZN => n6857);
   U15559 : OAI22_X1 port map( A1 => n11652, A2 => n11637, B1 => n670, B2 => 
                           n11636, ZN => n6856);
   U15560 : OAI22_X1 port map( A1 => n11653, A2 => n11637, B1 => n671, B2 => 
                           n11636, ZN => n6855);
   U15561 : OAI22_X1 port map( A1 => n11654, A2 => n11637, B1 => n672, B2 => 
                           n8536, ZN => n6854);
   U15562 : OAI22_X1 port map( A1 => n11655, A2 => n8537, B1 => n673, B2 => 
                           n8536, ZN => n6853);
   U15563 : OAI22_X1 port map( A1 => n11656, A2 => n8537, B1 => n674, B2 => 
                           n8536, ZN => n6852);
   U15564 : OAI22_X1 port map( A1 => n11657, A2 => n8537, B1 => n675, B2 => 
                           n8536, ZN => n6851);
   U15565 : OAI22_X1 port map( A1 => n11658, A2 => n8537, B1 => n676, B2 => 
                           n8536, ZN => n6850);
   U15566 : OAI22_X1 port map( A1 => n11659, A2 => n8537, B1 => n677, B2 => 
                           n8536, ZN => n6849);
   U15567 : OAI22_X1 port map( A1 => n11660, A2 => n8537, B1 => n678, B2 => 
                           n8536, ZN => n6848);
   U15568 : OAI22_X1 port map( A1 => n11661, A2 => n8537, B1 => n679, B2 => 
                           n8536, ZN => n6847);
   U15569 : OAI22_X1 port map( A1 => n11662, A2 => n8537, B1 => n680, B2 => 
                           n8536, ZN => n6846);
   U15570 : OAI22_X1 port map( A1 => n11663, A2 => n8537, B1 => n681, B2 => 
                           n8536, ZN => n6845);
   U15571 : OAI22_X1 port map( A1 => n11664, A2 => n8537, B1 => n682, B2 => 
                           n8536, ZN => n6844);
   U15572 : OAI22_X1 port map( A1 => n11665, A2 => n8537, B1 => n683, B2 => 
                           n8536, ZN => n6843);
   U15573 : OAI22_X1 port map( A1 => n11666, A2 => n8537, B1 => n684, B2 => 
                           n8536, ZN => n6842);
   U15574 : OAI22_X1 port map( A1 => n11667, A2 => n11637, B1 => n685, B2 => 
                           n8536, ZN => n6841);
   U15575 : OAI22_X1 port map( A1 => n11668, A2 => n11637, B1 => n686, B2 => 
                           n11636, ZN => n6840);
   U15576 : OAI22_X1 port map( A1 => n11669, A2 => n11637, B1 => n687, B2 => 
                           n8536, ZN => n6839);
   U15577 : OAI22_X1 port map( A1 => n11670, A2 => n11637, B1 => n688, B2 => 
                           n8536, ZN => n6838);
   U15578 : OAI22_X1 port map( A1 => n11671, A2 => n11637, B1 => n689, B2 => 
                           n8536, ZN => n6837);
   U15579 : OAI22_X1 port map( A1 => n11672, A2 => n8537, B1 => n690, B2 => 
                           n11636, ZN => n6836);
   U15580 : OAI22_X1 port map( A1 => n11673, A2 => n8537, B1 => n691, B2 => 
                           n11636, ZN => n6835);
   U15581 : OAI22_X1 port map( A1 => n11674, A2 => n8537, B1 => n692, B2 => 
                           n11636, ZN => n6834);
   U15582 : OAI22_X1 port map( A1 => n11675, A2 => n8537, B1 => n693, B2 => 
                           n8536, ZN => n6833);
   U15583 : OAI22_X1 port map( A1 => n11678, A2 => n8537, B1 => n694, B2 => 
                           n11636, ZN => n6832);
   U15584 : NAND2_X1 port map( A1 => n11638, A2 => n11642, ZN => n11639);
   U15585 : OAI22_X1 port map( A1 => n11645, A2 => n11641, B1 => n631, B2 => 
                           n11640, ZN => n6831);
   U15586 : OAI22_X1 port map( A1 => n11646, A2 => n11641, B1 => n632, B2 => 
                           n11640, ZN => n6830);
   U15587 : OAI22_X1 port map( A1 => n11647, A2 => n11641, B1 => n633, B2 => 
                           n11640, ZN => n6829);
   U15588 : OAI22_X1 port map( A1 => n11648, A2 => n11641, B1 => n634, B2 => 
                           n11640, ZN => n6828);
   U15589 : OAI22_X1 port map( A1 => n11649, A2 => n11641, B1 => n635, B2 => 
                           n11640, ZN => n6827);
   U15590 : OAI22_X1 port map( A1 => n11650, A2 => n11641, B1 => n636, B2 => 
                           n11640, ZN => n6826);
   U15591 : OAI22_X1 port map( A1 => n11651, A2 => n11641, B1 => n637, B2 => 
                           n11640, ZN => n6825);
   U15592 : OAI22_X1 port map( A1 => n11652, A2 => n11641, B1 => n638, B2 => 
                           n11640, ZN => n6824);
   U15593 : OAI22_X1 port map( A1 => n11653, A2 => n11641, B1 => n639, B2 => 
                           n11640, ZN => n6823);
   U15594 : OAI22_X1 port map( A1 => n11654, A2 => n11641, B1 => n640, B2 => 
                           n11640, ZN => n6822);
   U15595 : OAI22_X1 port map( A1 => n11655, A2 => n8538, B1 => n641, B2 => 
                           n11640, ZN => n6821);
   U15596 : OAI22_X1 port map( A1 => n11656, A2 => n8538, B1 => n642, B2 => 
                           n11640, ZN => n6820);
   U15597 : OAI22_X1 port map( A1 => n11657, A2 => n8538, B1 => n643, B2 => 
                           n11640, ZN => n6819);
   U15598 : OAI22_X1 port map( A1 => n11658, A2 => n8538, B1 => n644, B2 => 
                           n11640, ZN => n6818);
   U15599 : OAI22_X1 port map( A1 => n11659, A2 => n8538, B1 => n645, B2 => 
                           n11640, ZN => n6817);
   U15600 : OAI22_X1 port map( A1 => n11660, A2 => n8538, B1 => n646, B2 => 
                           n11640, ZN => n6816);
   U15601 : OAI22_X1 port map( A1 => n11661, A2 => n8538, B1 => n647, B2 => 
                           n11640, ZN => n6815);
   U15602 : OAI22_X1 port map( A1 => n11662, A2 => n8538, B1 => n648, B2 => 
                           n11640, ZN => n6814);
   U15603 : OAI22_X1 port map( A1 => n11663, A2 => n8538, B1 => n649, B2 => 
                           n11640, ZN => n6813);
   U15604 : OAI22_X1 port map( A1 => n11664, A2 => n8538, B1 => n650, B2 => 
                           n11640, ZN => n6812);
   U15605 : OAI22_X1 port map( A1 => n11665, A2 => n8538, B1 => n651, B2 => 
                           n11640, ZN => n6811);
   U15606 : OAI22_X1 port map( A1 => n11666, A2 => n8538, B1 => n652, B2 => 
                           n11640, ZN => n6810);
   U15607 : OAI22_X1 port map( A1 => n11667, A2 => n11641, B1 => n653, B2 => 
                           n11640, ZN => n6809);
   U15608 : OAI22_X1 port map( A1 => n11668, A2 => n11641, B1 => n654, B2 => 
                           n11640, ZN => n6808);
   U15609 : OAI22_X1 port map( A1 => n11669, A2 => n11641, B1 => n655, B2 => 
                           n11640, ZN => n6807);
   U15610 : OAI22_X1 port map( A1 => n11670, A2 => n11641, B1 => n656, B2 => 
                           n11640, ZN => n6806);
   U15611 : OAI22_X1 port map( A1 => n11671, A2 => n11641, B1 => n657, B2 => 
                           n11640, ZN => n6805);
   U15612 : OAI22_X1 port map( A1 => n11672, A2 => n8538, B1 => n658, B2 => 
                           n11640, ZN => n6804);
   U15613 : OAI22_X1 port map( A1 => n11673, A2 => n8538, B1 => n659, B2 => 
                           n11640, ZN => n6803);
   U15614 : OAI22_X1 port map( A1 => n11674, A2 => n8538, B1 => n660, B2 => 
                           n11640, ZN => n6802);
   U15615 : OAI22_X1 port map( A1 => n11675, A2 => n8538, B1 => n661, B2 => 
                           n11640, ZN => n6801);
   U15616 : OAI22_X1 port map( A1 => n11678, A2 => n8538, B1 => n662, B2 => 
                           n11640, ZN => n6800);
   U15617 : NAND2_X1 port map( A1 => n11643, A2 => n11642, ZN => n11644);
   U15618 : OAI22_X1 port map( A1 => n11645, A2 => n11677, B1 => n599, B2 => 
                           n11676, ZN => n6799);
   U15619 : OAI22_X1 port map( A1 => n11646, A2 => n11677, B1 => n600, B2 => 
                           n11676, ZN => n6798);
   U15620 : OAI22_X1 port map( A1 => n11647, A2 => n11677, B1 => n601, B2 => 
                           n11676, ZN => n6797);
   U15621 : OAI22_X1 port map( A1 => n11648, A2 => n11677, B1 => n602, B2 => 
                           n11676, ZN => n6796);
   U15622 : OAI22_X1 port map( A1 => n11649, A2 => n11677, B1 => n603, B2 => 
                           n11676, ZN => n6795);
   U15623 : OAI22_X1 port map( A1 => n11650, A2 => n11677, B1 => n604, B2 => 
                           n11676, ZN => n6794);
   U15624 : OAI22_X1 port map( A1 => n11651, A2 => n11677, B1 => n605, B2 => 
                           n11676, ZN => n6793);
   U15625 : OAI22_X1 port map( A1 => n11652, A2 => n11677, B1 => n606, B2 => 
                           n11676, ZN => n6792);
   U15626 : OAI22_X1 port map( A1 => n11653, A2 => n11677, B1 => n607, B2 => 
                           n11676, ZN => n6791);
   U15627 : OAI22_X1 port map( A1 => n11654, A2 => n11677, B1 => n608, B2 => 
                           n11676, ZN => n6790);
   U15628 : OAI22_X1 port map( A1 => n11655, A2 => n11677, B1 => n609, B2 => 
                           n11676, ZN => n6789);
   U15629 : OAI22_X1 port map( A1 => n11656, A2 => n8539, B1 => n610, B2 => 
                           n11676, ZN => n6788);
   U15630 : OAI22_X1 port map( A1 => n11657, A2 => n8539, B1 => n611, B2 => 
                           n11676, ZN => n6787);
   U15631 : OAI22_X1 port map( A1 => n11658, A2 => n8539, B1 => n612, B2 => 
                           n11676, ZN => n6786);
   U15632 : OAI22_X1 port map( A1 => n11659, A2 => n8539, B1 => n613, B2 => 
                           n11676, ZN => n6785);
   U15633 : OAI22_X1 port map( A1 => n11660, A2 => n8539, B1 => n614, B2 => 
                           n11676, ZN => n6784);
   U15634 : OAI22_X1 port map( A1 => n11661, A2 => n8539, B1 => n615, B2 => 
                           n11676, ZN => n6783);
   U15635 : OAI22_X1 port map( A1 => n11662, A2 => n8539, B1 => n616, B2 => 
                           n11676, ZN => n6782);
   U15636 : OAI22_X1 port map( A1 => n11663, A2 => n8539, B1 => n617, B2 => 
                           n11676, ZN => n6781);
   U15637 : OAI22_X1 port map( A1 => n11664, A2 => n8539, B1 => n618, B2 => 
                           n11676, ZN => n6780);
   U15638 : OAI22_X1 port map( A1 => n11665, A2 => n8539, B1 => n619, B2 => 
                           n11676, ZN => n6779);
   U15639 : OAI22_X1 port map( A1 => n11666, A2 => n8539, B1 => n620, B2 => 
                           n11676, ZN => n6778);
   U15640 : OAI22_X1 port map( A1 => n11667, A2 => n11677, B1 => n621, B2 => 
                           n11676, ZN => n6777);
   U15641 : OAI22_X1 port map( A1 => n11668, A2 => n11677, B1 => n622, B2 => 
                           n11676, ZN => n6776);
   U15642 : OAI22_X1 port map( A1 => n11669, A2 => n11677, B1 => n623, B2 => 
                           n11676, ZN => n6775);
   U15643 : OAI22_X1 port map( A1 => n11670, A2 => n11677, B1 => n624, B2 => 
                           n11676, ZN => n6774);
   U15644 : OAI22_X1 port map( A1 => n11671, A2 => n11677, B1 => n625, B2 => 
                           n11676, ZN => n6773);
   U15645 : OAI22_X1 port map( A1 => n11672, A2 => n8539, B1 => n626, B2 => 
                           n11676, ZN => n6772);
   U15646 : OAI22_X1 port map( A1 => n11673, A2 => n8539, B1 => n627, B2 => 
                           n11676, ZN => n6771);
   U15647 : OAI22_X1 port map( A1 => n11674, A2 => n8539, B1 => n628, B2 => 
                           n11676, ZN => n6770);
   U15648 : OAI22_X1 port map( A1 => n11675, A2 => n8539, B1 => n629, B2 => 
                           n11676, ZN => n6769);
   U15649 : OAI22_X1 port map( A1 => n11678, A2 => n8539, B1 => n630, B2 => 
                           n11676, ZN => n6768);
   U15650 : AOI22_X1 port map( A1 => i_RD1_0_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_0_port, B2 => n8543, ZN => n3261
                           );
   U15651 : AOI22_X1 port map( A1 => i_RD1_1_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_1_port, B2 => n8544, ZN => 
                           n11680);
   U15652 : INV_X1 port map( A => n11680, ZN => n6735);
   U15653 : AOI22_X1 port map( A1 => i_RD1_2_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_2_port, B2 => n8543, ZN => n3260
                           );
   U15654 : AOI22_X1 port map( A1 => i_RD1_3_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_3_port, B2 => n8544, ZN => 
                           n11681);
   U15655 : INV_X1 port map( A => n11681, ZN => n6734);
   U15656 : AOI22_X1 port map( A1 => i_RD1_4_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_4_port, B2 => n8544, ZN => n3259
                           );
   U15657 : AOI22_X1 port map( A1 => i_RD1_5_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_5_port, B2 => n8544, ZN => n3258
                           );
   U15658 : AOI22_X1 port map( A1 => i_RD1_6_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_6_port, B2 => n8544, ZN => n3257
                           );
   U15659 : AOI22_X1 port map( A1 => i_RD1_7_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_7_port, B2 => n8544, ZN => n3256
                           );
   U15660 : AOI22_X1 port map( A1 => i_RD1_8_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_8_port, B2 => n8544, ZN => 
                           n11682);
   U15661 : INV_X1 port map( A => n11682, ZN => n6733);
   U15662 : AOI22_X1 port map( A1 => i_RD1_9_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_9_port, B2 => n8544, ZN => n3255
                           );
   U15663 : AOI22_X1 port map( A1 => i_RD1_10_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_10_port, B2 => n8544, ZN => 
                           n11683);
   U15664 : INV_X1 port map( A => n11683, ZN => n6732);
   U15665 : AOI22_X1 port map( A1 => i_RD1_11_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_11_port, B2 => n8544, ZN => 
                           n3254);
   U15666 : AOI22_X1 port map( A1 => i_RD1_12_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_12_port, B2 => n8544, ZN => 
                           n11684);
   U15667 : INV_X1 port map( A => n11684, ZN => n6731);
   U15668 : AOI22_X1 port map( A1 => i_RD1_13_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_13_port, B2 => n8544, ZN => 
                           n11685);
   U15669 : INV_X1 port map( A => n11685, ZN => n6730);
   U15670 : AOI22_X1 port map( A1 => i_RD1_14_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_14_port, B2 => n8544, ZN => 
                           n11686);
   U15671 : INV_X1 port map( A => n11686, ZN => n6729);
   U15672 : AOI22_X1 port map( A1 => i_RD1_15_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_15_port, B2 => n8544, ZN => 
                           n3253);
   U15673 : AOI22_X1 port map( A1 => i_RD1_16_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_16_port, B2 => n8544, ZN => 
                           n3252);
   U15674 : AOI22_X1 port map( A1 => i_RD1_17_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_17_port, B2 => n8543, ZN => 
                           n3251);
   U15675 : AOI22_X1 port map( A1 => i_RD1_18_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_18_port, B2 => n8544, ZN => 
                           n3250);
   U15676 : AOI22_X1 port map( A1 => i_RD1_19_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_19_port, B2 => n8544, ZN => 
                           n3249);
   U15677 : AOI22_X1 port map( A1 => i_RD1_20_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_20_port, B2 => n8544, ZN => 
                           n11687);
   U15678 : INV_X1 port map( A => n11687, ZN => n6728);
   U15679 : AOI22_X1 port map( A1 => i_RD1_21_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_21_port, B2 => n8544, ZN => 
                           n3248);
   U15680 : AOI22_X1 port map( A1 => i_RD1_22_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_22_port, B2 => n8544, ZN => 
                           n3247);
   U15681 : AOI22_X1 port map( A1 => i_RD1_23_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_A_23_port, B2 => n8544, ZN => 
                           n3246);
   U15682 : AOI22_X1 port map( A1 => i_RD1_24_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_A_24_port, B2 => n8544, ZN => 
                           n3245);
   U15683 : AOI22_X1 port map( A1 => i_RD1_25_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_A_25_port, B2 => n8544, ZN => 
                           n3244);
   U15684 : AOI22_X1 port map( A1 => i_RD1_26_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_A_26_port, B2 => n8544, ZN => 
                           n3243);
   U15685 : AOI22_X1 port map( A1 => i_RD1_27_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_A_27_port, B2 => n8544, ZN => 
                           n3242);
   U15686 : AOI22_X1 port map( A1 => i_RD1_28_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_A_28_port, B2 => n8544, ZN => 
                           n3241);
   U15687 : AOI22_X1 port map( A1 => i_RD1_29_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_A_29_port, B2 => n8544, ZN => 
                           n3240);
   U15688 : AOI22_X1 port map( A1 => i_RD1_30_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_A_30_port, B2 => n8544, ZN => 
                           n3239);
   U15689 : AOI22_X1 port map( A1 => i_RD1_31_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_A_31_port, B2 => n8544, ZN => 
                           n3238);
   U15690 : NAND2_X1 port map( A1 => n8573, A2 => n11688, ZN => n3237);
   U15691 : NAND2_X1 port map( A1 => n8572, A2 => n11689, ZN => n3236);
   U15692 : NAND2_X1 port map( A1 => n8573, A2 => n11690, ZN => n3235);
   U15693 : NAND2_X1 port map( A1 => n8573, A2 => n11691, ZN => n3234);
   U15694 : NAND2_X1 port map( A1 => n8573, A2 => n11692, ZN => n3233);
   U15695 : NAND2_X1 port map( A1 => n8572, A2 => n11693, ZN => n3231);
   U15696 : NAND2_X1 port map( A1 => n8573, A2 => n11694, ZN => n3230);
   U15697 : NAND2_X1 port map( A1 => n8572, A2 => n11695, ZN => n3229);
   U15698 : NAND2_X1 port map( A1 => n8572, A2 => n11696, ZN => n3227);
   U15699 : NAND2_X1 port map( A1 => n8572, A2 => n11697, ZN => n3226);
   U15700 : NAND2_X1 port map( A1 => n8572, A2 => n11698, ZN => n3225);
   U15701 : NAND2_X1 port map( A1 => n8572, A2 => n11699, ZN => n3224);
   U15702 : NAND2_X1 port map( A1 => n8572, A2 => n11700, ZN => n3223);
   U15703 : NAND2_X1 port map( A1 => n8572, A2 => n11701, ZN => n3219);
   U15704 : NAND2_X1 port map( A1 => n8572, A2 => n11702, ZN => n3216);
   U15705 : NAND2_X1 port map( A1 => n8572, A2 => n11703, ZN => n3215);
   U15706 : NAND2_X1 port map( A1 => n8573, A2 => n11704, ZN => n3211);
   U15707 : NOR2_X1 port map( A1 => n541, A2 => n542, ZN => n11706);
   U15708 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_2_port, A2 => 
                           n11706, ZN => n11708);
   U15709 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_4_port, A2 => 
                           n11709, ZN => n11711);
   U15710 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_6_port, A2 => 
                           n11712, ZN => n11714);
   U15711 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_8_port, A2 => 
                           n11715, ZN => n11717);
   U15712 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_10_port, A2 => 
                           n11718, ZN => n11720);
   U15713 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_12_port, A2 => 
                           n11721, ZN => n11723);
   U15714 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_14_port, A2 => 
                           n11724, ZN => n11726);
   U15715 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_16_port, A2 => 
                           n11727, ZN => n11729);
   U15716 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_18_port, A2 => 
                           n11730, ZN => n11732);
   U15717 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_20_port, A2 => 
                           n11733, ZN => n11735);
   U15718 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_22_port, A2 => 
                           n11736, ZN => n11738);
   U15719 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_24_port, A2 => 
                           n11739, ZN => n11741);
   U15720 : NOR2_X1 port map( A1 => n566, A2 => n11741, ZN => n11742);
   U15721 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_26_port, A2 => 
                           n11742, ZN => n11745);
   U15722 : NOR2_X1 port map( A1 => n568, A2 => n11745, ZN => n11744);
   U15723 : INV_X1 port map( A => n11744, ZN => n11746);
   U15724 : NOR2_X1 port map( A1 => n569, A2 => n11746, ZN => n11747);
   U15725 : NAND2_X1 port map( A1 => DECODEhw_i_tickcounter_29_port, A2 => 
                           n11747, ZN => n11749);
   U15726 : NOR2_X1 port map( A1 => n570, A2 => n11749, ZN => n11748);
   U15727 : OAI21_X1 port map( B1 => DECODEhw_i_tickcounter_31_port, B2 => 
                           n11748, A => n8579, ZN => n11705);
   U15728 : AOI21_X1 port map( B1 => DECODEhw_i_tickcounter_31_port, B2 => 
                           n11748, A => n11705, ZN => n7166);
   U15729 : AND2_X1 port map( A1 => n8570, A2 => n541, ZN => n7165);
   U15730 : AOI211_X1 port map( C1 => n542, C2 => n541, A => RST, B => n11706, 
                           ZN => n7164);
   U15731 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_2_port, C2 => 
                           n11706, A => n11708, B => n8577, ZN => n11707);
   U15732 : AOI211_X1 port map( C1 => n544, C2 => n11708, A => RST, B => n11709
                           , ZN => n7162);
   U15733 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_4_port, C2 => 
                           n11709, A => n11711, B => n8571, ZN => n11710);
   U15734 : AOI211_X1 port map( C1 => n546, C2 => n11711, A => RST, B => n11712
                           , ZN => n7160);
   U15735 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_6_port, C2 => 
                           n11712, A => n11714, B => n8578, ZN => n11713);
   U15736 : INV_X1 port map( A => n11713, ZN => n7159);
   U15737 : AOI211_X1 port map( C1 => n548, C2 => n11714, A => RST, B => n11715
                           , ZN => n7158);
   U15738 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_8_port, C2 => 
                           n11715, A => n11717, B => n8572, ZN => n11716);
   U15739 : INV_X1 port map( A => n11716, ZN => n7157);
   U15740 : AOI211_X1 port map( C1 => n550, C2 => n11717, A => RST, B => n11718
                           , ZN => n7156);
   U15741 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_10_port, C2 => 
                           n11718, A => n11720, B => n8577, ZN => n11719);
   U15742 : INV_X1 port map( A => n11719, ZN => n7155);
   U15743 : AOI211_X1 port map( C1 => n552, C2 => n11720, A => RST, B => n11721
                           , ZN => n7154);
   U15744 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_12_port, C2 => 
                           n11721, A => n11723, B => n8574, ZN => n11722);
   U15745 : INV_X1 port map( A => n11722, ZN => n7153);
   U15746 : AOI211_X1 port map( C1 => n554, C2 => n11723, A => RST, B => n11724
                           , ZN => n7152);
   U15747 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_14_port, C2 => 
                           n11724, A => n11726, B => n8571, ZN => n11725);
   U15748 : INV_X1 port map( A => n11725, ZN => n7151);
   U15749 : AOI211_X1 port map( C1 => n556, C2 => n11726, A => RST, B => n11727
                           , ZN => n7150);
   U15750 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_16_port, C2 => 
                           n11727, A => n11729, B => n8570, ZN => n11728);
   U15751 : INV_X1 port map( A => n11728, ZN => n7149);
   U15752 : AOI211_X1 port map( C1 => n558, C2 => n11729, A => RST, B => n11730
                           , ZN => n7148);
   U15753 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_18_port, C2 => 
                           n11730, A => n11732, B => n8581, ZN => n11731);
   U15754 : INV_X1 port map( A => n11731, ZN => n7147);
   U15755 : AOI211_X1 port map( C1 => n560, C2 => n11732, A => RST, B => n11733
                           , ZN => n7146);
   U15756 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_20_port, C2 => 
                           n11733, A => n11735, B => n8582, ZN => n11734);
   U15757 : INV_X1 port map( A => n11734, ZN => n7145);
   U15758 : AOI211_X1 port map( C1 => n562, C2 => n11735, A => RST, B => n11736
                           , ZN => n7144);
   U15759 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_22_port, C2 => 
                           n11736, A => n11738, B => n8573, ZN => n11737);
   U15760 : INV_X1 port map( A => n11737, ZN => n7143);
   U15761 : AOI211_X1 port map( C1 => n564, C2 => n11738, A => RST, B => n11739
                           , ZN => n7142);
   U15762 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_24_port, C2 => 
                           n11739, A => n11741, B => n8576, ZN => n11740);
   U15763 : INV_X1 port map( A => n11740, ZN => n7141);
   U15764 : AOI211_X1 port map( C1 => n566, C2 => n11741, A => RST, B => n11742
                           , ZN => n7140);
   U15765 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_26_port, C2 => 
                           n11742, A => n11745, B => n8575, ZN => n11743);
   U15766 : INV_X1 port map( A => n11743, ZN => n7139);
   U15767 : AOI211_X1 port map( C1 => n568, C2 => n11745, A => RST, B => n11744
                           , ZN => n7138);
   U15768 : AOI211_X1 port map( C1 => n569, C2 => n11746, A => RST, B => n11747
                           , ZN => n7137);
   U15769 : OAI211_X1 port map( C1 => DECODEhw_i_tickcounter_29_port, C2 => 
                           n11747, A => n11749, B => n8572, ZN => n3160);
   U15770 : AOI211_X1 port map( C1 => n570, C2 => n11749, A => RST, B => n11748
                           , ZN => n7136);
   U15771 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_31_port, A2 =>
                           n11752, B1 => n11751, B2 => n7765, ZN => n3154);
   U15772 : NOR4_X1 port map( A1 => IR_8_port, A2 => IR_7_port, A3 => IR_9_port
                           , A4 => IR_10_port, ZN => n11754);
   U15773 : OAI21_X1 port map( B1 => n8238, B2 => n8418, A => n11755, ZN => 
                           n7135);
   U15774 : OAI21_X1 port map( B1 => n8418, B2 => n178, A => n11756, ZN => 
                           n7133);
   U15775 : OAI21_X1 port map( B1 => n8418, B2 => n177, A => n11757, ZN => 
                           n7132);
   U15776 : OAI21_X1 port map( B1 => n8418, B2 => n176, A => n11758, ZN => 
                           n7131);
   U15777 : OAI21_X1 port map( B1 => n8418, B2 => n175, A => n11759, ZN => 
                           n7130);
   U15778 : OAI21_X1 port map( B1 => n8418, B2 => n174, A => n11760, ZN => 
                           n7129);
   U15779 : OAI21_X1 port map( B1 => n10434, B2 => n173, A => n11761, ZN => 
                           n7128);
   U15780 : OAI21_X1 port map( B1 => n8418, B2 => n172, A => n11762, ZN => 
                           n7127);
   U15781 : OAI21_X1 port map( B1 => n8418, B2 => n171, A => n11763, ZN => 
                           n7126);
   U15782 : OAI21_X1 port map( B1 => n8418, B2 => n170, A => n11764, ZN => 
                           n7125);
   U15783 : OAI21_X1 port map( B1 => n8418, B2 => n169, A => n11765, ZN => 
                           n7124);
   U15784 : INV_X1 port map( A => IRAM_DATA(26), ZN => n11766);
   U15785 : INV_X1 port map( A => IRAM_DATA(28), ZN => n11768);
   U15786 : INV_X1 port map( A => IRAM_DATA(30), ZN => n11769);
   U15787 : AOI22_X1 port map( A1 => i_DATAMEM_WM, A2 => n11981, B1 => n10439, 
                           B2 => CU_I_CW_EX_DRAM_WE_port, ZN => n11770);
   U15788 : INV_X1 port map( A => n11770, ZN => n7118);
   U15789 : AOI22_X1 port map( A1 => n10439, A2 => CU_I_CW_ID_WB_EN_port, B1 =>
                           n11981, B2 => CU_I_CW_EX_WB_EN_port, ZN => n2839);
   U15790 : AOI22_X1 port map( A1 => n10439, A2 => CU_I_CW_ID_WB_MUX_SEL_port, 
                           B1 => n11981, B2 => CU_I_CW_EX_WB_MUX_SEL_port, ZN 
                           => n2838);
   U15791 : AOI22_X1 port map( A1 => n10439, A2 => CU_I_CW_EX_WB_EN_port, B1 =>
                           n11981, B2 => CU_I_CW_MEM_WB_EN_port, ZN => n2833);
   U15792 : AOI22_X1 port map( A1 => n10439, A2 => CU_I_CW_EX_WB_MUX_SEL_port, 
                           B1 => n11981, B2 => CU_I_CW_MEM_WB_MUX_SEL_port, ZN 
                           => n2832);
   U15793 : OAI21_X1 port map( B1 => n8458, B2 => CU_I_CW_EX_MEM_EN_port, A => 
                           n8575, ZN => n11771);
   U15794 : INV_X1 port map( A => n11771, ZN => n7099);
   U15795 : AOI22_X1 port map( A1 => DATA_SIZE_0_port, A2 => n11981, B1 => 
                           n10439, B2 => CU_I_CW_EX_DATA_SIZE_0_port, ZN => 
                           n11772);
   U15796 : INV_X1 port map( A => n11772, ZN => n7098);
   U15797 : AOI22_X1 port map( A1 => DATA_SIZE_1_port, A2 => n11981, B1 => 
                           n10439, B2 => CU_I_CW_EX_DATA_SIZE_1_port, ZN => 
                           n11773);
   U15798 : INV_X1 port map( A => n11773, ZN => n7097);
   U15799 : AOI22_X1 port map( A1 => i_DATAMEM_RM, A2 => n11981, B1 => n10439, 
                           B2 => CU_I_CW_EX_DRAM_RE_port, ZN => n11774);
   U15800 : INV_X1 port map( A => n11774, ZN => n7096);
   U15801 : NAND2_X1 port map( A1 => IR_2_port, A2 => IR_1_port, ZN => n11785);
   U15802 : NOR3_X1 port map( A1 => n11785, A2 => n11782, A3 => n11775, ZN => 
                           n11776);
   U15803 : AOI21_X1 port map( B1 => n11981, B2 => i_ALU_OP_0_port, A => n11776
                           , ZN => n11777);
   U15804 : OAI211_X1 port map( C1 => n11781, C2 => n11780, A => n11779, B => 
                           n11778, ZN => n7090);
   U15805 : OAI222_X1 port map( A1 => n11784, A2 => n11782, B1 => n11783, B2 =>
                           IR_26_port, C1 => n11791, C2 => n8283, ZN => n7089);
   U15806 : OAI211_X1 port map( C1 => n217, C2 => n11791, A => n11787, B => 
                           n11786, ZN => n7087);
   U15807 : INV_X1 port map( A => CU_I_CW_ID_MUXB_SEL_port, ZN => n11788);
   U15808 : NAND2_X1 port map( A1 => n10439, A2 => CU_I_CW_ID_MUXA_SEL_port, ZN
                           => n11789);
   U15809 : OAI21_X1 port map( B1 => n11791, B2 => n8557, A => n11789, ZN => 
                           n7085);
   U15810 : AOI22_X1 port map( A1 => n10439, A2 => CU_I_CW_ID_EX_EN_port, B1 =>
                           CU_I_CW_EX_EX_EN_port, B2 => n11981, ZN => n2767);
   U15811 : AOI22_X1 port map( A1 => n10433, A2 => 
                           DataPath_i_PIPLIN_WRB1_0_port, B1 => n7791, B2 => 
                           DataPath_i_PIPLIN_WRB2_0_port, ZN => n2766);
   U15812 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_WRB1_1_port
                           , B1 => n7791, B2 => DataPath_i_PIPLIN_WRB2_1_port, 
                           ZN => n2765);
   U15813 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_WRB1_2_port
                           , B1 => n7791, B2 => DataPath_i_PIPLIN_WRB2_2_port, 
                           ZN => n2764);
   U15814 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_WRB1_3_port
                           , B1 => n7791, B2 => DataPath_i_PIPLIN_WRB2_3_port, 
                           ZN => n2763);
   U15815 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_WRB1_4_port
                           , B1 => n7791, B2 => DataPath_i_PIPLIN_WRB2_4_port, 
                           ZN => n2762);
   U15816 : OAI22_X1 port map( A1 => n213, A2 => n11791, B1 => n10438, B2 => 
                           n11790, ZN => n7084);
   U15817 : OAI22_X1 port map( A1 => n212, A2 => n11791, B1 => n213, B2 => 
                           n11790, ZN => n7083);
   U15818 : AOI22_X1 port map( A1 => i_RD2_0_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_0_port, B2 => n8544, ZN => n2755
                           );
   U15819 : AOI22_X1 port map( A1 => i_RD2_1_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_1_port, B2 => n8544, ZN => n2754
                           );
   U15820 : AOI22_X1 port map( A1 => i_RD2_2_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_2_port, B2 => n8544, ZN => n2753
                           );
   U15821 : AOI22_X1 port map( A1 => i_RD2_3_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_3_port, B2 => n8544, ZN => 
                           n11792);
   U15822 : INV_X1 port map( A => n11792, ZN => n7082);
   U15823 : AOI22_X1 port map( A1 => i_RD2_4_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_B_4_port, B2 => n8544, ZN => 
                           n11793);
   U15824 : INV_X1 port map( A => n11793, ZN => n7081);
   U15825 : AOI22_X1 port map( A1 => i_RD2_5_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_5_port, B2 => n8544, ZN => n2752
                           );
   U15826 : INV_X1 port map( A => i_RD2_6_port, ZN => n11794);
   U15827 : OAI22_X1 port map( A1 => n477, A2 => n11847, B1 => n11794, B2 => 
                           n11846, ZN => n7080);
   U15828 : AOI22_X1 port map( A1 => i_RD2_7_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_7_port, B2 => n8544, ZN => n2751
                           );
   U15829 : AOI22_X1 port map( A1 => i_RD2_8_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_8_port, B2 => n8543, ZN => n2750
                           );
   U15830 : AOI22_X1 port map( A1 => i_RD2_9_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_9_port, B2 => n8543, ZN => n2749
                           );
   U15831 : AOI22_X1 port map( A1 => i_RD2_10_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_10_port, B2 => n8543, ZN => 
                           n11795);
   U15832 : INV_X1 port map( A => n11795, ZN => n7079);
   U15833 : AOI22_X1 port map( A1 => i_RD2_11_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_11_port, B2 => n8543, ZN => 
                           n2748);
   U15834 : AOI22_X1 port map( A1 => i_RD2_12_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_12_port, B2 => n8543, ZN => 
                           n11796);
   U15835 : INV_X1 port map( A => n11796, ZN => n7078);
   U15836 : OAI22_X1 port map( A1 => n11797, A2 => n11846, B1 => n8324, B2 => 
                           n11847, ZN => n7077);
   U15837 : AOI22_X1 port map( A1 => i_RD2_14_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_14_port, B2 => n8543, ZN => 
                           n11798);
   U15838 : INV_X1 port map( A => n11798, ZN => n7076);
   U15839 : AOI22_X1 port map( A1 => i_RD2_15_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_15_port, B2 => n8543, ZN => 
                           n2747);
   U15840 : AOI22_X1 port map( A1 => i_RD2_16_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_16_port, B2 => n8543, ZN => 
                           n2746);
   U15841 : AOI22_X1 port map( A1 => i_RD2_17_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_17_port, B2 => n8543, ZN => 
                           n2745);
   U15842 : AOI22_X1 port map( A1 => i_RD2_18_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_18_port, B2 => n8543, ZN => 
                           n2744);
   U15843 : AOI22_X1 port map( A1 => i_RD2_19_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_B_19_port, B2 => n8543, ZN => 
                           n2743);
   U15844 : AOI22_X1 port map( A1 => i_RD2_20_port, A2 => n7758, B1 => 
                           DataPath_i_PIPLIN_B_20_port, B2 => n8543, ZN => 
                           n11799);
   U15845 : INV_X1 port map( A => n11799, ZN => n7075);
   U15846 : AOI22_X1 port map( A1 => i_RD2_21_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_B_21_port, B2 => n8543, ZN => 
                           n2742);
   U15847 : AOI22_X1 port map( A1 => i_RD2_22_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_B_22_port, B2 => n8543, ZN => 
                           n2741);
   U15848 : AOI22_X1 port map( A1 => i_RD2_23_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_B_23_port, B2 => n8543, ZN => 
                           n2740);
   U15849 : AOI22_X1 port map( A1 => i_RD2_24_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_B_24_port, B2 => n8543, ZN => 
                           n2739);
   U15850 : AOI22_X1 port map( A1 => i_RD2_25_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_B_25_port, B2 => n8543, ZN => 
                           n2738);
   U15851 : AOI22_X1 port map( A1 => i_RD2_26_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_B_26_port, B2 => n8543, ZN => 
                           n2737);
   U15852 : AOI22_X1 port map( A1 => i_RD2_27_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_B_27_port, B2 => n8543, ZN => 
                           n2736);
   U15853 : AOI22_X1 port map( A1 => i_RD2_28_port, A2 => n11848, B1 => 
                           DataPath_i_PIPLIN_B_28_port, B2 => n8543, ZN => 
                           n2735);
   U15854 : AOI22_X1 port map( A1 => i_RD2_29_port, A2 => n11848, B1 => n8543, 
                           B2 => DataPath_i_PIPLIN_B_29_port, ZN => n2734);
   U15855 : AOI22_X1 port map( A1 => i_RD2_30_port, A2 => n7758, B1 => n8544, 
                           B2 => DataPath_i_PIPLIN_B_30_port, ZN => n2733);
   U15856 : AOI22_X1 port map( A1 => i_RD2_31_port, A2 => n7758, B1 => n8543, 
                           B2 => DataPath_i_PIPLIN_B_31_port, ZN => n2732);
   U15857 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_0_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_0_port, ZN => n2731);
   U15858 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_1_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_1_port, ZN => n2730);
   U15859 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_2_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_2_port, ZN => n2729);
   U15860 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_3_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_3_port, ZN => n2728);
   U15861 : AOI22_X1 port map( A1 => n10433, A2 => DataPath_i_PIPLIN_B_4_port, 
                           B1 => n10432, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_4_port, ZN => n2727);
   U15862 : AOI22_X1 port map( A1 => n10433, A2 => DataPath_i_PIPLIN_B_5_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_5_port, ZN => n2726);
   U15863 : AOI22_X1 port map( A1 => n10433, A2 => n8320, B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_6_port, ZN => n2725);
   U15864 : AOI22_X1 port map( A1 => n10433, A2 => DataPath_i_PIPLIN_B_7_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_7_port, ZN => n2724);
   U15865 : AOI22_X1 port map( A1 => n10433, A2 => DataPath_i_PIPLIN_B_8_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_8_port, ZN => n2723);
   U15866 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_9_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_9_port, ZN => n2722);
   U15867 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_10_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_10_port, ZN => n2721)
                           ;
   U15868 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_11_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_11_port, ZN => n2720)
                           ;
   U15869 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_12_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_12_port, ZN => n2719)
                           ;
   U15870 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_13_port, 
                           B1 => n10432, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_13_port, ZN => n2718)
                           ;
   U15871 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_14_port, 
                           B1 => n10432, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_14_port, ZN => n2717)
                           ;
   U15872 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_15_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_15_port, ZN => n2716)
                           ;
   U15873 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_16_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_16_port, ZN => n2715)
                           ;
   U15874 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_17_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_17_port, ZN => n2714)
                           ;
   U15875 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_18_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_18_port, ZN => n2713)
                           ;
   U15876 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_19_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_19_port, ZN => n2712)
                           ;
   U15877 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_20_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_20_port, ZN => n2711)
                           ;
   U15878 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_21_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_21_port, ZN => n2710)
                           ;
   U15879 : AOI22_X1 port map( A1 => n10433, A2 => DataPath_i_PIPLIN_B_22_port,
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_22_port, ZN => n2709)
                           ;
   U15880 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_23_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_23_port, ZN => n2708)
                           ;
   U15881 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_24_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_24_port, ZN => n2707)
                           ;
   U15882 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_25_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_25_port, ZN => n2706)
                           ;
   U15883 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_26_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_26_port, ZN => n2705)
                           ;
   U15884 : AOI22_X1 port map( A1 => n10433, A2 => DataPath_i_PIPLIN_B_27_port,
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_27_port, ZN => n2704)
                           ;
   U15885 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_28_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_28_port, ZN => n2703)
                           ;
   U15886 : AOI22_X1 port map( A1 => n10433, A2 => DataPath_i_PIPLIN_B_29_port,
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_29_port, ZN => n2702)
                           ;
   U15887 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_30_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_30_port, ZN => n2701)
                           ;
   U15888 : AOI22_X1 port map( A1 => n7796, A2 => DataPath_i_PIPLIN_B_31_port, 
                           B1 => n7791, B2 => 
                           DataPath_i_REG_ME_DATA_DATAMEM_31_port, ZN => n2700)
                           ;
   U15889 : INV_X1 port map( A => n11800, ZN => n11801);
   U15890 : OAI21_X1 port map( B1 => n8413, B2 => n11802, A => n11820, ZN => 
                           n11804);
   U15891 : NAND2_X1 port map( A1 => n11805, A2 => n11804, ZN => n11807);
   U15892 : NOR2_X1 port map( A1 => n11805, A2 => n11804, ZN => n11813);
   U15893 : NOR2_X1 port map( A1 => n11813, A2 => n11811, ZN => n11812);
   U15894 : AOI22_X1 port map( A1 => DataPath_RF_c_win_0_port, A2 => n11812, B1
                           => DataPath_RF_c_win_4_port, B2 => n11813, ZN => 
                           n11806);
   U15895 : OAI211_X1 port map( C1 => n8333, C2 => n11807, A => n11806, B => 
                           n8580, ZN => n7074);
   U15896 : AOI222_X1 port map( A1 => n8554, A2 => n11811, B1 => 
                           DataPath_RF_c_win_1_port, B2 => n11812, C1 => 
                           DataPath_RF_c_win_0_port, C2 => n11813, ZN => n11808
                           );
   U15897 : NOR2_X1 port map( A1 => RST, A2 => n11808, ZN => n7073);
   U15898 : AOI222_X1 port map( A1 => n11814, A2 => n11811, B1 => n11813, B2 =>
                           DataPath_RF_c_win_1_port, C1 => n8554, C2 => n11812,
                           ZN => n11809);
   U15899 : NOR2_X1 port map( A1 => RST, A2 => n11809, ZN => n7072);
   U15900 : AOI222_X1 port map( A1 => n11814, A2 => n11812, B1 => 
                           DataPath_RF_c_win_4_port, B2 => n11811, C1 => n8554,
                           C2 => n11813, ZN => n11810);
   U15901 : NOR2_X1 port map( A1 => RST, A2 => n11810, ZN => n7071);
   U15902 : NOR2_X1 port map( A1 => RST, A2 => n11815, ZN => n7070);
   U15903 : AOI21_X1 port map( B1 => DataPath_RF_PUSH_ADDRGEN_curr_state_0_port
                           , B2 => n7724, A => n11816, ZN => n11819);
   U15904 : AOI211_X1 port map( C1 => n11819, C2 => n11818, A => RST, B => 
                           n11817, ZN => n7069);
   U15905 : NAND2_X1 port map( A1 => n11996, A2 => n11820, ZN => n11822);
   U15906 : NOR2_X1 port map( A1 => n11996, A2 => n11820, ZN => n11826);
   U15907 : INV_X1 port map( A => n11822, ZN => n11828);
   U15908 : NOR2_X1 port map( A1 => n11826, A2 => n11828, ZN => n11827);
   U15909 : AOI22_X1 port map( A1 => DataPath_RF_c_swin_0_port, A2 => n11827, 
                           B1 => n11826, B2 => DataPath_RF_c_swin_1_port, ZN =>
                           n11821);
   U15910 : OAI211_X1 port map( C1 => n8334, C2 => n11822, A => n11821, B => 
                           n8575, ZN => n7068);
   U15911 : AOI222_X1 port map( A1 => DataPath_RF_c_swin_2_port, A2 => n11826, 
                           B1 => DataPath_RF_c_swin_0_port, B2 => n11828, C1 =>
                           DataPath_RF_c_swin_1_port, C2 => n11827, ZN => 
                           n11823);
   U15912 : NOR2_X1 port map( A1 => RST, A2 => n11823, ZN => n7067);
   U15913 : AOI222_X1 port map( A1 => DataPath_RF_c_swin_3_port, A2 => n11826, 
                           B1 => DataPath_RF_c_swin_2_port, B2 => n11827, C1 =>
                           DataPath_RF_c_swin_1_port, C2 => n11828, ZN => 
                           n11824);
   U15914 : NOR2_X1 port map( A1 => RST, A2 => n11824, ZN => n7066);
   U15915 : AOI222_X1 port map( A1 => DataPath_RF_c_swin_2_port, A2 => n11828, 
                           B1 => DataPath_RF_c_swin_4_port, B2 => n11826, C1 =>
                           DataPath_RF_c_swin_3_port, C2 => n11827, ZN => 
                           n11825);
   U15916 : NOR2_X1 port map( A1 => RST, A2 => n11825, ZN => n7065);
   U15917 : AOI222_X1 port map( A1 => DataPath_RF_c_swin_3_port, A2 => n11828, 
                           B1 => DataPath_RF_c_swin_4_port, B2 => n11827, C1 =>
                           DataPath_RF_c_swin_0_port, C2 => n11826, ZN => 
                           n11829);
   U15918 : NOR2_X1 port map( A1 => RST, A2 => n11829, ZN => n7064);
   U15919 : NOR2_X1 port map( A1 => n8412, A2 => n11830, ZN => n11833);
   U15920 : AOI211_X1 port map( C1 => n11833, C2 => n11832, A => RST, B => 
                           n11831, ZN => n7063);
   U15921 : AND2_X1 port map( A1 => n11833, A2 => n8572, ZN => n7062);
   U15922 : INV_X1 port map( A => i_RD1_0_port, ZN => n11835);
   U15923 : INV_X1 port map( A => i_RD1_3_port, ZN => n11836);
   U15924 : INV_X1 port map( A => i_RD1_4_port, ZN => n11837);
   U15925 : OAI21_X1 port map( B1 => n7757, B2 => n11839, A => n11838, ZN => 
                           n7052);
   U15926 : INV_X1 port map( A => i_RD1_11_port, ZN => n11840);
   U15927 : INV_X1 port map( A => i_RD1_14_port, ZN => n11842);
   U15928 : OAI21_X1 port map( B1 => n11842, B2 => n11845, A => n11841, ZN => 
                           n7047);
   U15929 : OAI21_X1 port map( B1 => n7757, B2 => n11844, A => n11843, ZN => 
                           n7046);
   U15930 : NOR2_X1 port map( A1 => n8189, A2 => n8197, ZN => n11864);
   U15931 : INV_X1 port map( A => n11864, ZN => n11852);
   U15932 : NAND2_X1 port map( A1 => n8188, A2 => n11879, ZN => n11860);
   U15933 : INV_X1 port map( A => n11860, ZN => n11861);
   U15934 : NOR2_X1 port map( A1 => n8188, A2 => n8189, ZN => n11851);
   U15935 : NAND3_X1 port map( A1 => n8188, A2 => n8197, A3 => i_ALU_OP_4_port,
                           ZN => n11873);
   U15936 : NOR2_X1 port map( A1 => n8197, A2 => n11883, ZN => n11850);
   U15937 : INV_X1 port map( A => n11851, ZN => n11849);
   U15938 : NAND2_X1 port map( A1 => n11852, A2 => n11849, ZN => n11853);
   U15939 : INV_X1 port map( A => n11873, ZN => n11868);
   U15940 : NAND2_X1 port map( A1 => n10431, A2 => n11852, ZN => n11865);
   U15941 : NAND2_X1 port map( A1 => n8188, A2 => n8189, ZN => n11870);
   U15942 : NOR2_X1 port map( A1 => n8566, A2 => n11878, ZN => n11858);
   U15943 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_0_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_0_port, ZN => 
                           n2209);
   U15944 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_1_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_1_port, ZN => 
                           n2208);
   U15945 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_2_port, B1 => 
                           n8553, B2 => DataPath_i_REG_LDSTR_OUT_2_port, ZN => 
                           n2207);
   U15946 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_3_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_3_port, ZN => 
                           n2206);
   U15947 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_4_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_4_port, ZN => 
                           n2205);
   U15948 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_5_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_5_port, ZN => 
                           n2204);
   U15949 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_6_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_6_port, ZN => 
                           n2203);
   U15950 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_7_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_7_port, ZN => 
                           n2202);
   U15951 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_8_port, B1 => 
                           n11988, B2 => DataPath_i_REG_LDSTR_OUT_8_port, ZN =>
                           n2201);
   U15952 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_9_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_9_port, ZN => 
                           n2200);
   U15953 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_10_port, B1 =>
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_10_port, ZN =>
                           n2199);
   U15954 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_11_port, B1 =>
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_11_port, ZN =>
                           n2198);
   U15955 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_12_port, B1 =>
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_12_port, ZN =>
                           n2197);
   U15956 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_13_port, B1 =>
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_13_port, ZN =>
                           n2196);
   U15957 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_14_port, B1 =>
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_14_port, ZN =>
                           n2195);
   U15958 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_15_port, B1 =>
                           n11988, B2 => DataPath_i_REG_LDSTR_OUT_15_port, ZN 
                           => n2194);
   U15959 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_16_port, B1 =>
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_16_port, ZN =>
                           n2193);
   U15960 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_17_port, B1 =>
                           n11988, B2 => DataPath_i_REG_LDSTR_OUT_17_port, ZN 
                           => n2192);
   U15961 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_18_port, B1 =>
                           n11988, B2 => DataPath_i_REG_LDSTR_OUT_18_port, ZN 
                           => n2191);
   U15962 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_19_port, B1 =>
                           n11988, B2 => DataPath_i_REG_LDSTR_OUT_19_port, ZN 
                           => n2190);
   U15963 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_20_port, B1 =>
                           n11988, B2 => DataPath_i_REG_LDSTR_OUT_20_port, ZN 
                           => n2189);
   U15964 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_21_port, B1 =>
                           n11988, B2 => DataPath_i_REG_LDSTR_OUT_21_port, ZN 
                           => n2188);
   U15965 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_22_port, B1 =>
                           n11988, B2 => DataPath_i_REG_LDSTR_OUT_22_port, ZN 
                           => n2187);
   U15966 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_23_port, B1 =>
                           n11988, B2 => DataPath_i_REG_LDSTR_OUT_23_port, ZN 
                           => n2186);
   U15967 : AOI22_X1 port map( A1 => n8552, A2 => DRAM_DATA_OUT_24_port, B1 => 
                           n8553, B2 => DataPath_i_REG_LDSTR_OUT_24_port, ZN =>
                           n2185);
   U15968 : AOI22_X1 port map( A1 => n8552, A2 => DRAM_DATA_OUT_25_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_25_port, ZN =>
                           n2184);
   U15969 : AOI22_X1 port map( A1 => n8552, A2 => DRAM_DATA_OUT_26_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_26_port, ZN =>
                           n2183);
   U15970 : AOI22_X1 port map( A1 => n11987, A2 => DRAM_DATA_OUT_27_port, B1 =>
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_27_port, ZN =>
                           n2182);
   U15971 : AOI22_X1 port map( A1 => n8552, A2 => DRAM_DATA_OUT_28_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_28_port, ZN =>
                           n2181);
   U15972 : AOI22_X1 port map( A1 => n8552, A2 => DRAM_DATA_OUT_29_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_29_port, ZN =>
                           n2180);
   U15973 : AOI22_X1 port map( A1 => n8552, A2 => DRAM_DATA_OUT_30_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_30_port, ZN =>
                           n2179);
   U15974 : AOI22_X1 port map( A1 => n8552, A2 => DRAM_DATA_OUT_31_port, B1 => 
                           n7786, B2 => DataPath_i_REG_LDSTR_OUT_31_port, ZN =>
                           n2178);
   U15975 : XNOR2_X1 port map( A => n10427, B => n11857, ZN => n11854);
   U15976 : AOI22_X1 port map( A1 => n10429, A2 => n11855, B1 => n7791, B2 => 
                           DRAM_ADDRESS_2_port, ZN => n2151);
   U15977 : NOR2_X1 port map( A1 => n11870, A2 => n8197, ZN => n11874);
   U15978 : OAI22_X1 port map( A1 => n498, A2 => n11884, B1 => n11863, B2 => 
                           n11885, ZN => n7015);
   U15979 : INV_X1 port map( A => n11874, ZN => n11867);
   U15980 : INV_X1 port map( A => n11870, ZN => n11869);
   U15981 : NOR2_X1 port map( A1 => n11871, A2 => n7773, ZN => n11872);
   U15982 : NOR3_X1 port map( A1 => n11876, A2 => n10425, A3 => n11875, ZN => 
                           n11877);
   U15983 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_0_port, A2 => 
                           n7786, B1 => n11987, B2 => n8278, ZN => n1149);
   U15984 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_1_port, A2 => 
                           n7786, B1 => n11987, B2 => n8285, ZN => n1148);
   U15985 : AOI22_X1 port map( A1 => DRAM_ADDRESS_2_port, A2 => n8552, B1 => 
                           n7786, B2 => DataPath_i_REG_MEM_ALUOUT_2_port, ZN =>
                           n1147);
   U15986 : AOI22_X1 port map( A1 => DRAM_ADDRESS_3_port, A2 => n8552, B1 => 
                           n7786, B2 => DataPath_i_REG_MEM_ALUOUT_3_port, ZN =>
                           n1146);
   U15987 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_4_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_4_port, ZN 
                           => n1145);
   U15988 : AOI22_X1 port map( A1 => DRAM_ADDRESS_5_port, A2 => n8552, B1 => 
                           n7786, B2 => DataPath_i_REG_MEM_ALUOUT_5_port, ZN =>
                           n1144);
   U15989 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_6_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_6_port, ZN 
                           => n1143);
   U15990 : AOI22_X1 port map( A1 => DRAM_ADDRESS_7_port, A2 => n8552, B1 => 
                           n7786, B2 => DataPath_i_REG_MEM_ALUOUT_7_port, ZN =>
                           n1142);
   U15991 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_8_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_8_port, ZN 
                           => n1141);
   U15992 : AOI22_X1 port map( A1 => DRAM_ADDRESS_9_port, A2 => n8552, B1 => 
                           n7786, B2 => DataPath_i_REG_MEM_ALUOUT_9_port, ZN =>
                           n1140);
   U15993 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_10_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_10_port, ZN 
                           => n1139);
   U15994 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_11_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_11_port, ZN 
                           => n1138);
   U15995 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_12_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_12_port, ZN 
                           => n1137);
   U15996 : AOI22_X1 port map( A1 => DRAM_ADDRESS_13_port, A2 => n8552, B1 => 
                           n7786, B2 => DataPath_i_REG_MEM_ALUOUT_13_port, ZN 
                           => n1136);
   U15997 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_14_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_14_port, ZN 
                           => n1135);
   U15998 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_15_port, A2 => 
                           n7786, B1 => n11987, B2 => DRAM_ADDRESS_15_port, ZN 
                           => n1134);
   U15999 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_16_port, A2 => 
                           n7786, B1 => n8552, B2 => DRAM_ADDRESS_16_port, ZN 
                           => n1133);
   U16000 : AOI22_X1 port map( A1 => DRAM_ADDRESS_17_port, A2 => n8552, B1 => 
                           n7786, B2 => DataPath_i_REG_MEM_ALUOUT_17_port, ZN 
                           => n1132);
   U16001 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_18_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_18_port, ZN 
                           => n1131);
   U16002 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_19_port, A2 => 
                           n7786, B1 => n11987, B2 => DRAM_ADDRESS_19_port, ZN 
                           => n1130);
   U16003 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_20_port, A2 => 
                           n7786, B1 => n11987, B2 => DRAM_ADDRESS_20_port, ZN 
                           => n1129);
   U16004 : AOI22_X1 port map( A1 => DRAM_ADDRESS_21_port, A2 => n8552, B1 => 
                           n7786, B2 => DataPath_i_REG_MEM_ALUOUT_21_port, ZN 
                           => n1128);
   U16005 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_22_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_22_port, ZN 
                           => n1127);
   U16006 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_23_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_23_port, ZN 
                           => n1126);
   U16007 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_24_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_24_port, ZN 
                           => n1125);
   U16008 : AOI22_X1 port map( A1 => DRAM_ADDRESS_25_port, A2 => n8552, B1 => 
                           n7786, B2 => DataPath_i_REG_MEM_ALUOUT_25_port, ZN 
                           => n1124);
   U16009 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_26_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_26_port, ZN 
                           => n1123);
   U16010 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_27_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_27_port, ZN 
                           => n1122);
   U16011 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_28_port, A2 => 
                           n8553, B1 => n8552, B2 => DRAM_ADDRESS_28_port, ZN 
                           => n1121);
   U16012 : AOI22_X1 port map( A1 => DRAM_ADDRESS_29_port, A2 => n8552, B1 => 
                           n7786, B2 => DataPath_i_REG_MEM_ALUOUT_29_port, ZN 
                           => n1120);
   U16013 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_30_port, A2 => 
                           n8553, B1 => n11987, B2 => DRAM_ADDRESS_30_port, ZN 
                           => n1119);
   U16014 : AOI22_X1 port map( A1 => DataPath_i_REG_MEM_ALUOUT_31_port, A2 => 
                           n8553, B1 => n8552, B2 => DRAM_ADDRESS_31_port, ZN 
                           => n1116);
   U16015 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2528_port, B1 => n11889,
                           B2 => n11925, ZN => n1112);
   U16016 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2529_port, B1 => n11889,
                           B2 => n11926, ZN => n1111);
   U16017 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2530_port, B1 => n11889,
                           B2 => n11927, ZN => n1110);
   U16018 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2531_port, B1 => n11889,
                           B2 => n11928, ZN => n1109);
   U16019 : AOI22_X1 port map( A1 => n11890, A2 => 
                           DataPath_RF_bus_reg_dataout_2532_port, B1 => n11889,
                           B2 => n11929, ZN => n1108);
   U16020 : AOI22_X1 port map( A1 => n11890, A2 => 
                           DataPath_RF_bus_reg_dataout_2533_port, B1 => n11889,
                           B2 => n11930, ZN => n1107);
   U16021 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2534_port, B1 => n11889,
                           B2 => n11931, ZN => n1106);
   U16022 : AOI22_X1 port map( A1 => n11890, A2 => 
                           DataPath_RF_bus_reg_dataout_2535_port, B1 => n11889,
                           B2 => n11932, ZN => n1105);
   U16023 : AOI22_X1 port map( A1 => n11890, A2 => 
                           DataPath_RF_bus_reg_dataout_2536_port, B1 => n11889,
                           B2 => n11898, ZN => n1104);
   U16024 : AOI22_X1 port map( A1 => n11890, A2 => 
                           DataPath_RF_bus_reg_dataout_2537_port, B1 => n11889,
                           B2 => n11933, ZN => n1103);
   U16025 : AOI22_X1 port map( A1 => n11890, A2 => 
                           DataPath_RF_bus_reg_dataout_2538_port, B1 => n11889,
                           B2 => n11934, ZN => n1102);
   U16026 : AOI22_X1 port map( A1 => n11890, A2 => 
                           DataPath_RF_bus_reg_dataout_2539_port, B1 => n11889,
                           B2 => n11935, ZN => n1101);
   U16027 : AOI22_X1 port map( A1 => n11890, A2 => 
                           DataPath_RF_bus_reg_dataout_2540_port, B1 => n11889,
                           B2 => n11936, ZN => n1100);
   U16028 : AOI22_X1 port map( A1 => n11890, A2 => 
                           DataPath_RF_bus_reg_dataout_2541_port, B1 => n11889,
                           B2 => n11937, ZN => n1099);
   U16029 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2542_port, B1 => n11889,
                           B2 => n11899, ZN => n1098);
   U16030 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2543_port, B1 => n11889,
                           B2 => n11938, ZN => n1097);
   U16031 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2544_port, B1 => n11889,
                           B2 => n11939, ZN => n1096);
   U16032 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2545_port, B1 => n11889,
                           B2 => n11900, ZN => n1095);
   U16033 : AOI22_X1 port map( A1 => n11890, A2 => 
                           DataPath_RF_bus_reg_dataout_2546_port, B1 => n11889,
                           B2 => n11941, ZN => n1094);
   U16034 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2547_port, B1 => n11889,
                           B2 => n11901, ZN => n1093);
   U16035 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2548_port, B1 => n11889,
                           B2 => n11902, ZN => n1092);
   U16036 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2549_port, B1 => n11889,
                           B2 => n11903, ZN => n1091);
   U16037 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2550_port, B1 => n11889,
                           B2 => n11946, ZN => n1090);
   U16038 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2551_port, B1 => n11889,
                           B2 => n11947, ZN => n1089);
   U16039 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2552_port, B1 => n11889,
                           B2 => n11948, ZN => n1088);
   U16040 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2553_port, B1 => n11889,
                           B2 => n11949, ZN => n1087);
   U16041 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2554_port, A2 
                           => n8545, B1 => n11916, B2 => n11888, ZN => n1086);
   U16042 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2555_port, B1 => n11889,
                           B2 => n11951, ZN => n1085);
   U16043 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2556_port, B1 => n11889,
                           B2 => n11952, ZN => n1084);
   U16044 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2557_port, A2 
                           => n8545, B1 => n11919, B2 => n11888, ZN => n1083);
   U16045 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2558_port, B1 => n11889,
                           B2 => n11954, ZN => n1082);
   U16046 : AOI22_X1 port map( A1 => n8545, A2 => 
                           DataPath_RF_bus_reg_dataout_2559_port, B1 => n11889,
                           B2 => n11955, ZN => n1079);
   U16047 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2496_port, A2 
                           => n11895, B1 => n11894, B2 => n11925, ZN => n1075);
   U16048 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2497_port, A2 
                           => n11895, B1 => n11894, B2 => n11926, ZN => n1074);
   U16049 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2498_port, A2 
                           => n11895, B1 => n11894, B2 => n11927, ZN => n1073);
   U16050 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2499_port, A2 
                           => n11895, B1 => n11894, B2 => n11928, ZN => n1072);
   U16051 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2500_port, A2 
                           => n11895, B1 => n11894, B2 => n11929, ZN => n1071);
   U16052 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2501_port, A2 
                           => n11895, B1 => n11894, B2 => n11930, ZN => n1070);
   U16053 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2502_port, A2 
                           => n11895, B1 => n11894, B2 => n11931, ZN => n1069);
   U16054 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2503_port, A2 
                           => n11895, B1 => n11894, B2 => n11932, ZN => n1068);
   U16055 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2504_port, A2 
                           => n8546, B1 => n11894, B2 => n11898, ZN => n1067);
   U16056 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2505_port, A2 
                           => n8546, B1 => n11894, B2 => n11933, ZN => n1066);
   U16057 : AOI22_X1 port map( A1 => n11968, A2 => n11893, B1 => n11895, B2 => 
                           DataPath_RF_bus_reg_dataout_2506_port, ZN => n1065);
   U16058 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2507_port, A2 
                           => n8546, B1 => n11894, B2 => n11935, ZN => n1064);
   U16059 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2508_port, A2 
                           => n8546, B1 => n11894, B2 => n11936, ZN => n1063);
   U16060 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2509_port, A2 
                           => n8546, B1 => n11894, B2 => n11937, ZN => n1062);
   U16061 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2510_port, A2 
                           => n8546, B1 => n11894, B2 => n11899, ZN => n1061);
   U16062 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2511_port, A2 
                           => n8546, B1 => n11894, B2 => n11938, ZN => n1060);
   U16063 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2512_port, A2 
                           => n8546, B1 => n11894, B2 => n11939, ZN => n1059);
   U16064 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2513_port, A2 
                           => n8546, B1 => n11894, B2 => n11900, ZN => n1058);
   U16065 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2514_port, A2 
                           => n8546, B1 => n11894, B2 => n11941, ZN => n1057);
   U16066 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2515_port, A2 
                           => n8546, B1 => n11894, B2 => n11901, ZN => n1056);
   U16067 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2516_port, A2 
                           => n8546, B1 => n11894, B2 => n11902, ZN => n1055);
   U16068 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2517_port, A2 
                           => n8546, B1 => n11894, B2 => n11903, ZN => n1054);
   U16069 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2518_port, A2 
                           => n11895, B1 => n11894, B2 => n11946, ZN => n1053);
   U16070 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2519_port, A2 
                           => n8546, B1 => n11894, B2 => n11947, ZN => n1052);
   U16071 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2520_port, A2 
                           => n8546, B1 => n11894, B2 => n11948, ZN => n1051);
   U16072 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2521_port, A2 
                           => n8546, B1 => n11894, B2 => n11949, ZN => n1050);
   U16073 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2522_port, A2 
                           => n8546, B1 => n11894, B2 => n11950, ZN => n1049);
   U16074 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2523_port, A2 
                           => n8546, B1 => n11894, B2 => n11951, ZN => n1048);
   U16075 : AOI22_X1 port map( A1 => n11918, A2 => n11893, B1 => n8546, B2 => 
                           DataPath_RF_bus_reg_dataout_2524_port, ZN => n1047);
   U16076 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2525_port, A2 
                           => n8546, B1 => n11894, B2 => n11953, ZN => n1046);
   U16077 : AOI22_X1 port map( A1 => n11920, A2 => n11893, B1 => n8546, B2 => 
                           DataPath_RF_bus_reg_dataout_2526_port, ZN => n1045);
   U16078 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2527_port, A2 
                           => n8546, B1 => n11894, B2 => n11955, ZN => n1042);
   U16079 : OAI22_X1 port map( A1 => n8219, A2 => n11897, B1 => n11923, B2 => 
                           n11896, ZN => n11904);
   U16080 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2464_port, A2 
                           => n8547, B1 => n11905, B2 => n11925, ZN => n1038);
   U16081 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2465_port, A2 
                           => n8547, B1 => n11905, B2 => n11926, ZN => n1037);
   U16082 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2466_port, A2 
                           => n8547, B1 => n11905, B2 => n11927, ZN => n1036);
   U16083 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2467_port, A2 
                           => n8547, B1 => n11905, B2 => n11928, ZN => n1035);
   U16084 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2468_port, A2 
                           => n8547, B1 => n11905, B2 => n11929, ZN => n1034);
   U16085 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2469_port, A2 
                           => n8547, B1 => n11905, B2 => n11930, ZN => n1033);
   U16086 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2470_port, A2 
                           => n8547, B1 => n11905, B2 => n11931, ZN => n1032);
   U16087 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2471_port, A2 
                           => n8547, B1 => n11905, B2 => n11932, ZN => n1031);
   U16088 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2472_port, A2 
                           => n8547, B1 => n11905, B2 => n11898, ZN => n1030);
   U16089 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2473_port, A2 
                           => n8547, B1 => n11905, B2 => n11933, ZN => n1029);
   U16090 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2474_port, A2 
                           => n11906, B1 => n11905, B2 => n11934, ZN => n1028);
   U16091 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2475_port, A2 
                           => n11906, B1 => n11905, B2 => n11935, ZN => n1027);
   U16092 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2476_port, A2 
                           => n11906, B1 => n11905, B2 => n11936, ZN => n1026);
   U16093 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2477_port, A2 
                           => n8547, B1 => n11905, B2 => n11937, ZN => n1025);
   U16094 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2478_port, A2 
                           => n11906, B1 => n11905, B2 => n11899, ZN => n1024);
   U16095 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2479_port, A2 
                           => n8547, B1 => n11905, B2 => n11938, ZN => n1023);
   U16096 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2480_port, A2 
                           => n8547, B1 => n11905, B2 => n11939, ZN => n1022);
   U16097 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2481_port, A2 
                           => n8547, B1 => n11905, B2 => n11900, ZN => n1021);
   U16098 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2482_port, A2 
                           => n11906, B1 => n11905, B2 => n11941, ZN => n1020);
   U16099 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2483_port, A2 
                           => n8547, B1 => n11905, B2 => n11901, ZN => n1019);
   U16100 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2484_port, A2 
                           => n8547, B1 => n11905, B2 => n11902, ZN => n1018);
   U16101 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2485_port, A2 
                           => n11906, B1 => n11905, B2 => n11903, ZN => n1017);
   U16102 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2486_port, A2 
                           => n8547, B1 => n11905, B2 => n11946, ZN => n1016);
   U16103 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2487_port, A2 
                           => n8547, B1 => n11905, B2 => n11947, ZN => n1015);
   U16104 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2488_port, A2 
                           => n8547, B1 => n11905, B2 => n11948, ZN => n1014);
   U16105 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2489_port, A2 
                           => n11906, B1 => n11905, B2 => n11949, ZN => n1013);
   U16106 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2490_port, A2 
                           => n11906, B1 => n11905, B2 => n11950, ZN => n1012);
   U16107 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2491_port, A2 
                           => n11906, B1 => n11905, B2 => n11951, ZN => n1011);
   U16108 : AOI22_X1 port map( A1 => n11918, A2 => n11904, B1 => n8547, B2 => 
                           DataPath_RF_bus_reg_dataout_2492_port, ZN => n1010);
   U16109 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2493_port, A2 
                           => n8547, B1 => n11905, B2 => n11953, ZN => n1009);
   U16110 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2494_port, A2 
                           => n11906, B1 => n11905, B2 => n11954, ZN => n1008);
   U16111 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2495_port, A2 
                           => n8547, B1 => n11905, B2 => n11955, ZN => n1005);
   U16112 : OAI22_X1 port map( A1 => n8219, A2 => n11908, B1 => n11923, B2 => 
                           n11907, ZN => n11909);
   U16113 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2432_port, B1 => n11958,
                           B2 => n8286, ZN => n1001);
   U16114 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2433_port, B1 => n11959,
                           B2 => n8286, ZN => n1000);
   U16115 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2434_port, B1 => n11960,
                           B2 => n8286, ZN => n999);
   U16116 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2435_port, B1 => n11961,
                           B2 => n8286, ZN => n998);
   U16117 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2436_port, B1 => n11962,
                           B2 => n8286, ZN => n997);
   U16118 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2437_port, B1 => n11963,
                           B2 => n8286, ZN => n996);
   U16119 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2438_port, B1 => n11964,
                           B2 => n8286, ZN => n995);
   U16120 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2439_port, B1 => n11965,
                           B2 => n8286, ZN => n994);
   U16121 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2440_port, B1 => n11966,
                           B2 => n8286, ZN => n993);
   U16122 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2441_port, B1 => n11967,
                           B2 => n8286, ZN => n992);
   U16123 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2442_port, B1 => n11968,
                           B2 => n8286, ZN => n991);
   U16124 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_2443_port, B1 => n11969,
                           B2 => n8286, ZN => n990);
   U16125 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_2444_port, B1 => n11970,
                           B2 => n8286, ZN => n989);
   U16126 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_2445_port, B1 => n11971,
                           B2 => n8286, ZN => n988);
   U16127 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_2446_port, B1 => n11972,
                           B2 => n8286, ZN => n987);
   U16128 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_2447_port, B1 => n11974,
                           B2 => n8286, ZN => n986);
   U16129 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_2448_port, B1 => n11910,
                           B2 => n8286, ZN => n985);
   U16130 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_2449_port, B1 => n11940,
                           B2 => n8286, ZN => n984);
   U16131 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_2450_port, B1 => n11911,
                           B2 => n8286, ZN => n983);
   U16132 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_2451_port, B1 => n11942,
                           B2 => n8286, ZN => n982);
   U16133 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_2452_port, B1 => n11943,
                           B2 => n8286, ZN => n981);
   U16134 : AOI22_X1 port map( A1 => n8548, A2 => 
                           DataPath_RF_bus_reg_dataout_2453_port, B1 => n11945,
                           B2 => n8286, ZN => n980);
   U16135 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2454_port, B1 => n11912,
                           B2 => n8286, ZN => n979);
   U16136 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2455_port, B1 => n11913,
                           B2 => n8286, ZN => n978);
   U16137 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2456_port, B1 => n11914,
                           B2 => n8286, ZN => n977);
   U16138 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2457_port, B1 => n11915,
                           B2 => n8286, ZN => n976);
   U16139 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2458_port, B1 => n11916,
                           B2 => n8286, ZN => n975);
   U16140 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2459_port, B1 => n11917,
                           B2 => n8286, ZN => n974);
   U16141 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2460_port, B1 => n11918,
                           B2 => n8286, ZN => n973);
   U16142 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2461_port, B1 => n11919,
                           B2 => n8286, ZN => n972);
   U16143 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2462_port, B1 => n11920,
                           B2 => n8286, ZN => n971);
   U16144 : AOI22_X1 port map( A1 => n7781, A2 => 
                           DataPath_RF_bus_reg_dataout_2463_port, B1 => n11921,
                           B2 => n8286, ZN => n968);
   U16145 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2400_port, A2 
                           => n11957, B1 => n11956, B2 => n11925, ZN => n963);
   U16146 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2401_port, A2 
                           => n11957, B1 => n11956, B2 => n11926, ZN => n962);
   U16147 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2402_port, A2 
                           => n11957, B1 => n11956, B2 => n11927, ZN => n961);
   U16148 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2403_port, A2 
                           => n11957, B1 => n11956, B2 => n11928, ZN => n960);
   U16149 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2404_port, A2 
                           => n8549, B1 => n11956, B2 => n11929, ZN => n959);
   U16150 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2405_port, A2 
                           => n11957, B1 => n11956, B2 => n11930, ZN => n958);
   U16151 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2406_port, A2 
                           => n8549, B1 => n11956, B2 => n11931, ZN => n957);
   U16152 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2407_port, A2 
                           => n8549, B1 => n11956, B2 => n11932, ZN => n956);
   U16153 : AOI22_X1 port map( A1 => n11966, A2 => n11944, B1 => n8549, B2 => 
                           DataPath_RF_bus_reg_dataout_2408_port, ZN => n955);
   U16154 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2409_port, A2 
                           => n8549, B1 => n11956, B2 => n11933, ZN => n954);
   U16155 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2410_port, A2 
                           => n8549, B1 => n11956, B2 => n11934, ZN => n953);
   U16156 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2411_port, A2 
                           => n8549, B1 => n11956, B2 => n11935, ZN => n952);
   U16157 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2412_port, A2 
                           => n8549, B1 => n11956, B2 => n11936, ZN => n951);
   U16158 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2413_port, A2 
                           => n8549, B1 => n11956, B2 => n11937, ZN => n950);
   U16159 : AOI22_X1 port map( A1 => n11972, A2 => n11944, B1 => n11957, B2 => 
                           DataPath_RF_bus_reg_dataout_2414_port, ZN => n949);
   U16160 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2415_port, A2 
                           => n8549, B1 => n11956, B2 => n11938, ZN => n948);
   U16161 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2416_port, A2 
                           => n8549, B1 => n11956, B2 => n11939, ZN => n946);
   U16162 : AOI22_X1 port map( A1 => n11940, A2 => n11944, B1 => n11957, B2 => 
                           DataPath_RF_bus_reg_dataout_2417_port, ZN => n944);
   U16163 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2418_port, A2 
                           => n11957, B1 => n11956, B2 => n11941, ZN => n942);
   U16164 : AOI22_X1 port map( A1 => n11942, A2 => n11944, B1 => n8549, B2 => 
                           DataPath_RF_bus_reg_dataout_2419_port, ZN => n940);
   U16165 : AOI22_X1 port map( A1 => n11943, A2 => n11944, B1 => n8549, B2 => 
                           DataPath_RF_bus_reg_dataout_2420_port, ZN => n938);
   U16166 : AOI22_X1 port map( A1 => n11945, A2 => n11944, B1 => n8549, B2 => 
                           DataPath_RF_bus_reg_dataout_2421_port, ZN => n936);
   U16167 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2422_port, A2 
                           => n11957, B1 => n11956, B2 => n11946, ZN => n934);
   U16168 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2423_port, A2 
                           => n8549, B1 => n11956, B2 => n11947, ZN => n932);
   U16169 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2424_port, A2 
                           => n8549, B1 => n11956, B2 => n11948, ZN => n930);
   U16170 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2425_port, A2 
                           => n8549, B1 => n11956, B2 => n11949, ZN => n928);
   U16171 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2426_port, A2 
                           => n11957, B1 => n11956, B2 => n11950, ZN => n926);
   U16172 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2427_port, A2 
                           => n8549, B1 => n11956, B2 => n11951, ZN => n924);
   U16173 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2428_port, A2 
                           => n8549, B1 => n11956, B2 => n11952, ZN => n922);
   U16174 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2429_port, A2 
                           => n8549, B1 => n11956, B2 => n11953, ZN => n920);
   U16175 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2430_port, A2 
                           => n8549, B1 => n11956, B2 => n11954, ZN => n918);
   U16176 : AOI22_X1 port map( A1 => DataPath_RF_bus_reg_dataout_2431_port, A2 
                           => n8549, B1 => n11956, B2 => n11955, ZN => n914);
   U16177 : OAI22_X1 port map( A1 => n8551, A2 => n11958, B1 => 
                           DataPath_RF_bus_reg_dataout_2368_port, B2 => n8550, 
                           ZN => n912);
   U16178 : OAI22_X1 port map( A1 => n8551, A2 => n11959, B1 => 
                           DataPath_RF_bus_reg_dataout_2369_port, B2 => n8550, 
                           ZN => n910);
   U16179 : OAI22_X1 port map( A1 => n8551, A2 => n11960, B1 => 
                           DataPath_RF_bus_reg_dataout_2370_port, B2 => n8550, 
                           ZN => n908);
   U16180 : OAI22_X1 port map( A1 => n8551, A2 => n11961, B1 => 
                           DataPath_RF_bus_reg_dataout_2371_port, B2 => n8550, 
                           ZN => n906);
   U16181 : OAI22_X1 port map( A1 => n8551, A2 => n11962, B1 => 
                           DataPath_RF_bus_reg_dataout_2372_port, B2 => n11973,
                           ZN => n904);
   U16182 : OAI22_X1 port map( A1 => n8551, A2 => n11963, B1 => 
                           DataPath_RF_bus_reg_dataout_2373_port, B2 => n11973,
                           ZN => n902);
   U16183 : OAI22_X1 port map( A1 => n8551, A2 => n11964, B1 => 
                           DataPath_RF_bus_reg_dataout_2374_port, B2 => n11973,
                           ZN => n900);
   U16184 : OAI22_X1 port map( A1 => n11975, A2 => n11965, B1 => 
                           DataPath_RF_bus_reg_dataout_2375_port, B2 => n11973,
                           ZN => n898);
   U16185 : OAI22_X1 port map( A1 => n8551, A2 => n11966, B1 => 
                           DataPath_RF_bus_reg_dataout_2376_port, B2 => n11973,
                           ZN => n896);
   U16186 : OAI22_X1 port map( A1 => n11975, A2 => n11967, B1 => 
                           DataPath_RF_bus_reg_dataout_2377_port, B2 => n11973,
                           ZN => n894);
   U16187 : OAI22_X1 port map( A1 => n11975, A2 => n11968, B1 => 
                           DataPath_RF_bus_reg_dataout_2378_port, B2 => n11973,
                           ZN => n892);
   U16188 : OAI22_X1 port map( A1 => n11975, A2 => n11969, B1 => 
                           DataPath_RF_bus_reg_dataout_2379_port, B2 => n11973,
                           ZN => n890);
   U16189 : OAI22_X1 port map( A1 => n8551, A2 => n11970, B1 => 
                           DataPath_RF_bus_reg_dataout_2380_port, B2 => n11973,
                           ZN => n888);
   U16190 : OAI22_X1 port map( A1 => n8551, A2 => n11971, B1 => 
                           DataPath_RF_bus_reg_dataout_2381_port, B2 => n8550, 
                           ZN => n886);
   U16191 : OAI22_X1 port map( A1 => n11975, A2 => n11972, B1 => 
                           DataPath_RF_bus_reg_dataout_2382_port, B2 => n8550, 
                           ZN => n884);
   U16192 : OAI22_X1 port map( A1 => n11975, A2 => n11974, B1 => 
                           DataPath_RF_bus_reg_dataout_2383_port, B2 => n8550, 
                           ZN => n880);
   U16193 : INV_X1 port map( A => n11976, ZN => DRAM_ISSUE);
   U16194 : AOI22_X1 port map( A1 => n10439, A2 => CU_I_CW_ID_DRAM_RE_port, B1 
                           => n11981, B2 => CU_I_CW_EX_DRAM_RE_port, ZN => 
                           n11977);
   U16195 : INV_X1 port map( A => n11977, ZN => n368);
   U16196 : AOI22_X1 port map( A1 => n10439, A2 => CU_I_CW_ID_DATA_SIZE_1_port,
                           B1 => n11981, B2 => CU_I_CW_EX_DATA_SIZE_1_port, ZN 
                           => n11978);
   U16197 : INV_X1 port map( A => n11978, ZN => n367);
   U16198 : AOI22_X1 port map( A1 => n10439, A2 => CU_I_CW_ID_DATA_SIZE_0_port,
                           B1 => n11981, B2 => CU_I_CW_EX_DATA_SIZE_0_port, ZN 
                           => n11979);
   U16199 : INV_X1 port map( A => n11979, ZN => n366);
   U16200 : AOI22_X1 port map( A1 => n10439, A2 => CU_I_CW_ID_MEM_EN_port, B1 
                           => n11981, B2 => CU_I_CW_EX_MEM_EN_port, ZN => 
                           n11980);
   U16201 : INV_X1 port map( A => n11980, ZN => n365);
   U16202 : AOI22_X1 port map( A1 => n10439, A2 => CU_I_CW_ID_DRAM_WE_port, B1 
                           => n11981, B2 => CU_I_CW_EX_DRAM_WE_port, ZN => 
                           n11982);
   U16203 : INV_X1 port map( A => n11982, ZN => n364);
   U16204 : AOI22_X1 port map( A1 => n8552, A2 => DataPath_i_PIPLIN_WRB2_4_port
                           , B1 => n7786, B2 => i_ADD_WB_4_port, ZN => n11983);
   U16205 : INV_X1 port map( A => n11983, ZN => n359);
   U16206 : AOI22_X1 port map( A1 => n8552, A2 => DataPath_i_PIPLIN_WRB2_3_port
                           , B1 => n7786, B2 => i_ADD_WB_3_port, ZN => n11984);
   U16207 : INV_X1 port map( A => n11984, ZN => n358);
   U16208 : AOI22_X1 port map( A1 => i_ADD_WB_2_port, A2 => n8553, B1 => n8552,
                           B2 => DataPath_i_PIPLIN_WRB2_2_port, ZN => n11985);
   U16209 : INV_X1 port map( A => n11985, ZN => n357);
   U16210 : AOI22_X1 port map( A1 => n8552, A2 => DataPath_i_PIPLIN_WRB2_1_port
                           , B1 => n7786, B2 => i_ADD_WB_1_port, ZN => n11986);
   U16211 : INV_X1 port map( A => n11986, ZN => n356);
   U16212 : AOI22_X1 port map( A1 => i_ADD_WB_0_port, A2 => n8553, B1 => n11987
                           , B2 => DataPath_i_PIPLIN_WRB2_0_port, ZN => n11989)
                           ;
   U16213 : INV_X1 port map( A => n11989, ZN => n355);
   U16214 : AOI21_X1 port map( B1 => n11991, B2 => n8412, A => n11990, ZN => 
                           n11992);
   U16215 : AOI21_X1 port map( B1 => n466, B2 => n11993, A => n11992, ZN => 
                           n11994);
   U16216 : NOR2_X1 port map( A1 => RST, A2 => n11994, ZN => n99);
   U16217 : OAI21_X1 port map( B1 => n8417, B2 => n11996, A => n11995, ZN => 
                           DRAMRF_ISSUE);
   U16218 : AOI21_X1 port map( B1 => DataPath_RF_PUSH_ADDRGEN_curr_state_0_port
                           , B2 => n7724, A => n11997, ZN => n90);
   U16219 : OAI21_X1 port map( B1 => n8418, B2 => n179, A => n11999, ZN => n43)
                           ;
   U16220 : OAI21_X1 port map( B1 => n8418, B2 => n180, A => n12000, ZN => n42)
                           ;
   U16221 : OAI21_X1 port map( B1 => n8224, B2 => n8418, A => n12001, ZN => n36
                           );
   U16222 : OAI21_X1 port map( B1 => n8418, B2 => n193, A => n12002, ZN => n34)
                           ;
   IRAM_ISSUE <= '1';

end SYN_dlx_rtl;
